module W_half_extend