
module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_con_RegWr, i_addr_Rd, 
        i_data_Rd, o_data_Rs, o_data_Rt, i_addr_Rt_4_, i_addr_Rt_3_, 
        i_addr_Rt_2_, i_addr_Rt_1_, i_addr_Rt_0_ );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr, i_addr_Rt_4_, i_addr_Rt_3_, i_addr_Rt_2_,
         i_addr_Rt_1_, i_addr_Rt_0_;
  wire   n5, n6, n9, n11, n13, n15, n16, n17, n18, n20, n21, n22, n23, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n1, n2, n3, n4, n7, n8, n10, n12, n14, n19, n24,
         n33, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591;
  wire   [1023:0] regs;

  DFEC1 regs_reg_31__30_ ( .D(i_data_Rd[30]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(i_data_Rd[29]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(i_data_Rd[28]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(i_data_Rd[27]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(i_data_Rd[26]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(i_data_Rd[25]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(i_data_Rd[24]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(i_data_Rd[23]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(i_data_Rd[22]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(i_data_Rd[21]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(i_data_Rd[20]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(i_data_Rd[18]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(i_data_Rd[17]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(i_data_Rd[16]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(i_data_Rd[15]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(i_data_Rd[14]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(i_data_Rd[13]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(i_data_Rd[12]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(i_data_Rd[11]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(i_data_Rd[10]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(i_data_Rd[9]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(i_data_Rd[8]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(i_data_Rd[7]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(i_data_Rd[5]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(i_data_Rd[4]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(i_data_Rd[3]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(i_data_Rd[2]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(i_data_Rd[0]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[992]) );
  DFEC1 regs_reg_30__31_ ( .D(i_data_Rd[31]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(i_data_Rd[30]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(i_data_Rd[29]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(i_data_Rd[28]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(i_data_Rd[27]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(i_data_Rd[26]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(i_data_Rd[25]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(i_data_Rd[24]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(i_data_Rd[23]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(i_data_Rd[22]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(i_data_Rd[21]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(i_data_Rd[20]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(i_data_Rd[18]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(i_data_Rd[17]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(i_data_Rd[16]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(i_data_Rd[15]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(i_data_Rd[14]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(i_data_Rd[13]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(i_data_Rd[12]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(i_data_Rd[11]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(i_data_Rd[10]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(i_data_Rd[9]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(i_data_Rd[8]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(i_data_Rd[7]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(i_data_Rd[5]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(i_data_Rd[4]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(i_data_Rd[3]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(i_data_Rd[2]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(i_data_Rd[0]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[960]) );
  DFEC1 regs_reg_29__31_ ( .D(i_data_Rd[31]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(i_data_Rd[30]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(i_data_Rd[29]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(i_data_Rd[28]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[956]) );
  DFEC1 regs_reg_29__27_ ( .D(i_data_Rd[27]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(i_data_Rd[26]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(i_data_Rd[25]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(i_data_Rd[24]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(i_data_Rd[23]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(i_data_Rd[22]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(i_data_Rd[21]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(i_data_Rd[20]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(i_data_Rd[18]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(i_data_Rd[17]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(i_data_Rd[16]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(i_data_Rd[15]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(i_data_Rd[14]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(i_data_Rd[13]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(i_data_Rd[12]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(i_data_Rd[11]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(i_data_Rd[10]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(i_data_Rd[9]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(i_data_Rd[8]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(i_data_Rd[7]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(i_data_Rd[5]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(i_data_Rd[4]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(i_data_Rd[3]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(i_data_Rd[2]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(i_data_Rd[0]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[928]) );
  DFEC1 regs_reg_28__31_ ( .D(i_data_Rd[31]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(i_data_Rd[30]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(i_data_Rd[29]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(i_data_Rd[28]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(i_data_Rd[27]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(i_data_Rd[26]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(i_data_Rd[25]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(i_data_Rd[24]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(i_data_Rd[23]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(i_data_Rd[22]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(i_data_Rd[21]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(i_data_Rd[20]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(i_data_Rd[18]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(i_data_Rd[17]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(i_data_Rd[16]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(i_data_Rd[15]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(i_data_Rd[14]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(i_data_Rd[13]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(i_data_Rd[12]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(i_data_Rd[11]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(i_data_Rd[10]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(i_data_Rd[9]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(i_data_Rd[8]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(i_data_Rd[7]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(i_data_Rd[5]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(i_data_Rd[4]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(i_data_Rd[3]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(i_data_Rd[2]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(i_data_Rd[0]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(i_data_Rd[31]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(i_data_Rd[30]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(i_data_Rd[29]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(i_data_Rd[28]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(i_data_Rd[27]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(i_data_Rd[26]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(i_data_Rd[25]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(i_data_Rd[24]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(i_data_Rd[23]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(i_data_Rd[22]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(i_data_Rd[21]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(i_data_Rd[20]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(i_data_Rd[18]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(i_data_Rd[17]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(i_data_Rd[16]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(i_data_Rd[15]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(i_data_Rd[14]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(i_data_Rd[13]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(i_data_Rd[12]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(i_data_Rd[11]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(i_data_Rd[10]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(i_data_Rd[9]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(i_data_Rd[8]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(i_data_Rd[7]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(i_data_Rd[5]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(i_data_Rd[4]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(i_data_Rd[3]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(i_data_Rd[2]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(i_data_Rd[1]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(i_data_Rd[0]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[864]) );
  DFEC1 regs_reg_26__31_ ( .D(i_data_Rd[31]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(i_data_Rd[30]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(i_data_Rd[29]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(i_data_Rd[28]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(i_data_Rd[27]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(i_data_Rd[26]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(i_data_Rd[25]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(i_data_Rd[24]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(i_data_Rd[23]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(i_data_Rd[22]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(i_data_Rd[21]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(i_data_Rd[20]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(i_data_Rd[18]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(i_data_Rd[17]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(i_data_Rd[16]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(i_data_Rd[15]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(i_data_Rd[14]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(i_data_Rd[13]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(i_data_Rd[12]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(i_data_Rd[11]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(i_data_Rd[10]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(i_data_Rd[9]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(i_data_Rd[8]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(i_data_Rd[7]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(i_data_Rd[5]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(i_data_Rd[4]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(i_data_Rd[3]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(i_data_Rd[2]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(i_data_Rd[0]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[832]) );
  DFEC1 regs_reg_25__31_ ( .D(i_data_Rd[31]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(i_data_Rd[30]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(i_data_Rd[29]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(i_data_Rd[28]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(i_data_Rd[27]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(i_data_Rd[26]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(i_data_Rd[25]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(i_data_Rd[24]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(i_data_Rd[23]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(i_data_Rd[22]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(i_data_Rd[21]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(i_data_Rd[20]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(i_data_Rd[19]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(i_data_Rd[18]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(i_data_Rd[17]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(i_data_Rd[16]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(i_data_Rd[15]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(i_data_Rd[14]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(i_data_Rd[13]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(i_data_Rd[12]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(i_data_Rd[11]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(i_data_Rd[10]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(i_data_Rd[9]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(i_data_Rd[8]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(i_data_Rd[7]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(i_data_Rd[6]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(i_data_Rd[5]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(i_data_Rd[4]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(i_data_Rd[3]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(i_data_Rd[2]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(i_data_Rd[1]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(i_data_Rd[0]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[800]) );
  DFEC1 regs_reg_24__31_ ( .D(i_data_Rd[31]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(i_data_Rd[30]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(i_data_Rd[29]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(i_data_Rd[28]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(i_data_Rd[27]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(i_data_Rd[26]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(i_data_Rd[25]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(i_data_Rd[24]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(i_data_Rd[23]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(i_data_Rd[22]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(i_data_Rd[21]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(i_data_Rd[20]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(i_data_Rd[19]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(i_data_Rd[18]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(i_data_Rd[17]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(i_data_Rd[16]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(i_data_Rd[15]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(i_data_Rd[14]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(i_data_Rd[13]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(i_data_Rd[12]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(i_data_Rd[11]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(i_data_Rd[10]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(i_data_Rd[9]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(i_data_Rd[8]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(i_data_Rd[7]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(i_data_Rd[6]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(i_data_Rd[5]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(i_data_Rd[4]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(i_data_Rd[3]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(i_data_Rd[2]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(i_data_Rd[1]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(i_data_Rd[0]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(i_data_Rd[31]), .E(n22), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(i_data_Rd[30]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(i_data_Rd[29]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(i_data_Rd[28]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(i_data_Rd[27]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(i_data_Rd[26]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(i_data_Rd[25]), .E(n22), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(i_data_Rd[24]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(i_data_Rd[23]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(i_data_Rd[22]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(i_data_Rd[21]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(i_data_Rd[20]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(i_data_Rd[19]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(i_data_Rd[18]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(i_data_Rd[17]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(i_data_Rd[16]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(i_data_Rd[15]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(i_data_Rd[14]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(i_data_Rd[13]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(i_data_Rd[12]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(i_data_Rd[11]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(i_data_Rd[10]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(i_data_Rd[9]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(i_data_Rd[8]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(i_data_Rd[7]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(i_data_Rd[6]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(i_data_Rd[5]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(i_data_Rd[4]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(i_data_Rd[3]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(i_data_Rd[2]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(i_data_Rd[1]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(i_data_Rd[0]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[736]) );
  DFEC1 regs_reg_22__31_ ( .D(i_data_Rd[31]), .E(n21), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(i_data_Rd[30]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(i_data_Rd[29]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(i_data_Rd[28]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(i_data_Rd[27]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(i_data_Rd[26]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(i_data_Rd[25]), .E(n21), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(i_data_Rd[24]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(i_data_Rd[23]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(i_data_Rd[22]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(i_data_Rd[21]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(i_data_Rd[20]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(i_data_Rd[19]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(i_data_Rd[18]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(i_data_Rd[17]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(i_data_Rd[16]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(i_data_Rd[15]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(i_data_Rd[14]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(i_data_Rd[13]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(i_data_Rd[12]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(i_data_Rd[11]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(i_data_Rd[10]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(i_data_Rd[9]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(i_data_Rd[8]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(i_data_Rd[7]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(i_data_Rd[6]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(i_data_Rd[5]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(i_data_Rd[4]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(i_data_Rd[3]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(i_data_Rd[2]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(i_data_Rd[1]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(i_data_Rd[0]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[704]) );
  DFEC1 regs_reg_21__31_ ( .D(i_data_Rd[31]), .E(n20), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(i_data_Rd[30]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(i_data_Rd[29]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(i_data_Rd[28]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(i_data_Rd[27]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(i_data_Rd[26]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(i_data_Rd[25]), .E(n20), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(i_data_Rd[24]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(i_data_Rd[23]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(i_data_Rd[22]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(i_data_Rd[21]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(i_data_Rd[20]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(i_data_Rd[19]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(i_data_Rd[18]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(i_data_Rd[17]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(i_data_Rd[16]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(i_data_Rd[15]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(i_data_Rd[14]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(i_data_Rd[13]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(i_data_Rd[12]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(i_data_Rd[11]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(i_data_Rd[10]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(i_data_Rd[9]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(i_data_Rd[8]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(i_data_Rd[7]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(i_data_Rd[6]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(i_data_Rd[5]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(i_data_Rd[4]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(i_data_Rd[3]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(i_data_Rd[2]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(i_data_Rd[1]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(i_data_Rd[0]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[672]) );
  DFEC1 regs_reg_20__31_ ( .D(i_data_Rd[31]), .E(n18), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(i_data_Rd[30]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(i_data_Rd[29]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(i_data_Rd[28]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(i_data_Rd[27]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(i_data_Rd[26]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(i_data_Rd[25]), .E(n18), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(i_data_Rd[24]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(i_data_Rd[23]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(i_data_Rd[22]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(i_data_Rd[21]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(i_data_Rd[20]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(i_data_Rd[19]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(i_data_Rd[18]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(i_data_Rd[17]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(i_data_Rd[16]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(i_data_Rd[15]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(i_data_Rd[14]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(i_data_Rd[13]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(i_data_Rd[12]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(i_data_Rd[11]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(i_data_Rd[10]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(i_data_Rd[9]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(i_data_Rd[8]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(i_data_Rd[7]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(i_data_Rd[6]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(i_data_Rd[5]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(i_data_Rd[4]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(i_data_Rd[3]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(i_data_Rd[2]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(i_data_Rd[1]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(i_data_Rd[0]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(i_data_Rd[31]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(i_data_Rd[30]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(i_data_Rd[29]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(i_data_Rd[28]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(i_data_Rd[27]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(i_data_Rd[26]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(i_data_Rd[25]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(i_data_Rd[24]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(i_data_Rd[23]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(i_data_Rd[22]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(i_data_Rd[21]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(i_data_Rd[20]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(i_data_Rd[19]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(i_data_Rd[18]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(i_data_Rd[17]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(i_data_Rd[16]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(i_data_Rd[15]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(i_data_Rd[14]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(i_data_Rd[13]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(i_data_Rd[12]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(i_data_Rd[11]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(i_data_Rd[10]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(i_data_Rd[9]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(i_data_Rd[8]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(i_data_Rd[7]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(i_data_Rd[6]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(i_data_Rd[5]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(i_data_Rd[4]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(i_data_Rd[3]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(i_data_Rd[2]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(i_data_Rd[1]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(i_data_Rd[0]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[608]) );
  DFEC1 regs_reg_18__31_ ( .D(i_data_Rd[31]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(i_data_Rd[30]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(i_data_Rd[29]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(i_data_Rd[28]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(i_data_Rd[27]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(i_data_Rd[26]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(i_data_Rd[25]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(i_data_Rd[24]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(i_data_Rd[23]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(i_data_Rd[22]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(i_data_Rd[21]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(i_data_Rd[20]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(i_data_Rd[19]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(i_data_Rd[18]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(i_data_Rd[17]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(i_data_Rd[16]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(i_data_Rd[15]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(i_data_Rd[14]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(i_data_Rd[13]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(i_data_Rd[12]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(i_data_Rd[11]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(i_data_Rd[10]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(i_data_Rd[9]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(i_data_Rd[8]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(i_data_Rd[7]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(i_data_Rd[6]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(i_data_Rd[5]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(i_data_Rd[4]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(i_data_Rd[3]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(i_data_Rd[2]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(i_data_Rd[1]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(i_data_Rd[0]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[576]) );
  DFEC1 regs_reg_17__31_ ( .D(i_data_Rd[31]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(i_data_Rd[30]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(i_data_Rd[29]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(i_data_Rd[28]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(i_data_Rd[27]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(i_data_Rd[26]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(i_data_Rd[25]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(i_data_Rd[24]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(i_data_Rd[23]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(i_data_Rd[22]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(i_data_Rd[21]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(i_data_Rd[20]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(i_data_Rd[19]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(i_data_Rd[18]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(i_data_Rd[17]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(i_data_Rd[16]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(i_data_Rd[15]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(i_data_Rd[14]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(i_data_Rd[13]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(i_data_Rd[12]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(i_data_Rd[11]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(i_data_Rd[10]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(i_data_Rd[9]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(i_data_Rd[8]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(i_data_Rd[7]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(i_data_Rd[6]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(i_data_Rd[5]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(i_data_Rd[4]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(i_data_Rd[3]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(i_data_Rd[2]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(i_data_Rd[1]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(i_data_Rd[0]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(i_data_Rd[31]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(i_data_Rd[30]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(i_data_Rd[29]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(i_data_Rd[28]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(i_data_Rd[27]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(i_data_Rd[26]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(i_data_Rd[25]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(i_data_Rd[24]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(i_data_Rd[23]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(i_data_Rd[22]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(i_data_Rd[21]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(i_data_Rd[20]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(i_data_Rd[19]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(i_data_Rd[18]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(i_data_Rd[17]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(i_data_Rd[16]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(i_data_Rd[15]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(i_data_Rd[14]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(i_data_Rd[13]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(i_data_Rd[12]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(i_data_Rd[11]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(i_data_Rd[10]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(i_data_Rd[9]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(i_data_Rd[8]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(i_data_Rd[7]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(i_data_Rd[6]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(i_data_Rd[5]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(i_data_Rd[4]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(i_data_Rd[3]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(i_data_Rd[2]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(i_data_Rd[1]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(i_data_Rd[0]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[512]) );
  DFEC1 regs_reg_15__31_ ( .D(i_data_Rd[31]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(i_data_Rd[30]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(i_data_Rd[29]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(i_data_Rd[28]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(i_data_Rd[27]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(i_data_Rd[26]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(i_data_Rd[25]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(i_data_Rd[24]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(i_data_Rd[23]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(i_data_Rd[22]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(i_data_Rd[21]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(i_data_Rd[20]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(i_data_Rd[19]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(i_data_Rd[18]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(i_data_Rd[17]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(i_data_Rd[16]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(i_data_Rd[15]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(i_data_Rd[13]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(i_data_Rd[12]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(i_data_Rd[11]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(i_data_Rd[9]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(i_data_Rd[8]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(i_data_Rd[7]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(i_data_Rd[6]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(i_data_Rd[5]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(i_data_Rd[4]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(i_data_Rd[3]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(i_data_Rd[2]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(i_data_Rd[1]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(i_data_Rd[0]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[480]) );
  DFEC1 regs_reg_14__31_ ( .D(i_data_Rd[31]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(i_data_Rd[30]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(i_data_Rd[29]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(i_data_Rd[28]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(i_data_Rd[27]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(i_data_Rd[26]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(i_data_Rd[25]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(i_data_Rd[24]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(i_data_Rd[23]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(i_data_Rd[22]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(i_data_Rd[21]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(i_data_Rd[20]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(i_data_Rd[19]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(i_data_Rd[18]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(i_data_Rd[17]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(i_data_Rd[16]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(i_data_Rd[15]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(i_data_Rd[13]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(i_data_Rd[12]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(i_data_Rd[11]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(i_data_Rd[9]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(i_data_Rd[8]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(i_data_Rd[7]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(i_data_Rd[6]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(i_data_Rd[5]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(i_data_Rd[4]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(i_data_Rd[3]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(i_data_Rd[2]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(i_data_Rd[1]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(i_data_Rd[0]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[448]) );
  DFEC1 regs_reg_13__31_ ( .D(i_data_Rd[31]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(i_data_Rd[30]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(i_data_Rd[29]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(i_data_Rd[28]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[444]) );
  DFEC1 regs_reg_13__27_ ( .D(i_data_Rd[27]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(i_data_Rd[26]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(i_data_Rd[25]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(i_data_Rd[24]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(i_data_Rd[23]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(i_data_Rd[22]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(i_data_Rd[21]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(i_data_Rd[20]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(i_data_Rd[19]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(i_data_Rd[18]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(i_data_Rd[17]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(i_data_Rd[16]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(i_data_Rd[15]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(i_data_Rd[13]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(i_data_Rd[12]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(i_data_Rd[11]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(i_data_Rd[9]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(i_data_Rd[8]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(i_data_Rd[7]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(i_data_Rd[6]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(i_data_Rd[5]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(i_data_Rd[4]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(i_data_Rd[3]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(i_data_Rd[2]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(i_data_Rd[1]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(i_data_Rd[0]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[416]) );
  DFEC1 regs_reg_12__31_ ( .D(i_data_Rd[31]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(i_data_Rd[30]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(i_data_Rd[29]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(i_data_Rd[28]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(i_data_Rd[27]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(i_data_Rd[26]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(i_data_Rd[25]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(i_data_Rd[24]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(i_data_Rd[23]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(i_data_Rd[22]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(i_data_Rd[21]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(i_data_Rd[20]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(i_data_Rd[19]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(i_data_Rd[18]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(i_data_Rd[17]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(i_data_Rd[16]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(i_data_Rd[15]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(i_data_Rd[13]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(i_data_Rd[12]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(i_data_Rd[11]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(i_data_Rd[9]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(i_data_Rd[8]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(i_data_Rd[7]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(i_data_Rd[6]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(i_data_Rd[5]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(i_data_Rd[4]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(i_data_Rd[3]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(i_data_Rd[2]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(i_data_Rd[1]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(i_data_Rd[0]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[384]) );
  DFEC1 regs_reg_11__31_ ( .D(i_data_Rd[31]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(i_data_Rd[30]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(i_data_Rd[29]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(i_data_Rd[28]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(i_data_Rd[27]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(i_data_Rd[26]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(i_data_Rd[25]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(i_data_Rd[24]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(i_data_Rd[23]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(i_data_Rd[22]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(i_data_Rd[21]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(i_data_Rd[20]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(i_data_Rd[19]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(i_data_Rd[18]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(i_data_Rd[17]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(i_data_Rd[16]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(i_data_Rd[15]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(i_data_Rd[13]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(i_data_Rd[12]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(i_data_Rd[11]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(i_data_Rd[10]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(i_data_Rd[9]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(i_data_Rd[8]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(i_data_Rd[7]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(i_data_Rd[6]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(i_data_Rd[5]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(i_data_Rd[4]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(i_data_Rd[3]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(i_data_Rd[2]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(i_data_Rd[1]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(i_data_Rd[0]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[352]) );
  DFEC1 regs_reg_10__31_ ( .D(i_data_Rd[31]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(i_data_Rd[30]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(i_data_Rd[29]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(i_data_Rd[28]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(i_data_Rd[27]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(i_data_Rd[26]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(i_data_Rd[25]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(i_data_Rd[24]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(i_data_Rd[23]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(i_data_Rd[22]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(i_data_Rd[21]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(i_data_Rd[20]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(i_data_Rd[19]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(i_data_Rd[18]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(i_data_Rd[17]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(i_data_Rd[16]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(i_data_Rd[15]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(i_data_Rd[13]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(i_data_Rd[12]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(i_data_Rd[11]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(i_data_Rd[9]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(i_data_Rd[8]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(i_data_Rd[7]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(i_data_Rd[6]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(i_data_Rd[5]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(i_data_Rd[4]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(i_data_Rd[3]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(i_data_Rd[2]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(i_data_Rd[1]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(i_data_Rd[0]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[320]) );
  DFEC1 regs_reg_9__31_ ( .D(i_data_Rd[31]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(i_data_Rd[30]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(i_data_Rd[29]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(i_data_Rd[28]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(i_data_Rd[27]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(i_data_Rd[26]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(i_data_Rd[25]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(i_data_Rd[24]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(i_data_Rd[23]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(i_data_Rd[22]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(i_data_Rd[21]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(i_data_Rd[20]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(i_data_Rd[19]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(i_data_Rd[18]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(i_data_Rd[17]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(i_data_Rd[16]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(i_data_Rd[15]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(i_data_Rd[14]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(i_data_Rd[13]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(i_data_Rd[12]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(i_data_Rd[11]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(i_data_Rd[10]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(i_data_Rd[9]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(i_data_Rd[8]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(i_data_Rd[7]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(i_data_Rd[6]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(i_data_Rd[5]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(i_data_Rd[4]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(i_data_Rd[3]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(i_data_Rd[2]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(i_data_Rd[1]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(i_data_Rd[0]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[288]) );
  DFEC1 regs_reg_8__31_ ( .D(i_data_Rd[31]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(i_data_Rd[30]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(i_data_Rd[29]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(i_data_Rd[28]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(i_data_Rd[27]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(i_data_Rd[26]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(i_data_Rd[25]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(i_data_Rd[24]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(i_data_Rd[23]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(i_data_Rd[22]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(i_data_Rd[21]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(i_data_Rd[20]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(i_data_Rd[19]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(i_data_Rd[18]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(i_data_Rd[17]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(i_data_Rd[16]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(i_data_Rd[15]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(i_data_Rd[14]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(i_data_Rd[13]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(i_data_Rd[12]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(i_data_Rd[11]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(i_data_Rd[10]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(i_data_Rd[9]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(i_data_Rd[8]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(i_data_Rd[7]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(i_data_Rd[6]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(i_data_Rd[5]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(i_data_Rd[4]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(i_data_Rd[3]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(i_data_Rd[2]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(i_data_Rd[1]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(i_data_Rd[0]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[256]) );
  DFEC1 regs_reg_7__31_ ( .D(i_data_Rd[31]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(i_data_Rd[30]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(i_data_Rd[29]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(i_data_Rd[28]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(i_data_Rd[27]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(i_data_Rd[26]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(i_data_Rd[25]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(i_data_Rd[24]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(i_data_Rd[23]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(i_data_Rd[22]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(i_data_Rd[21]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(i_data_Rd[20]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(i_data_Rd[19]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(i_data_Rd[18]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(i_data_Rd[17]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(i_data_Rd[16]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(i_data_Rd[15]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(i_data_Rd[14]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(i_data_Rd[13]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(i_data_Rd[12]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(i_data_Rd[11]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(i_data_Rd[10]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(i_data_Rd[9]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(i_data_Rd[8]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(i_data_Rd[7]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(i_data_Rd[6]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(i_data_Rd[5]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(i_data_Rd[4]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(i_data_Rd[3]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(i_data_Rd[2]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(i_data_Rd[1]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(i_data_Rd[0]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[224]) );
  DFEC1 regs_reg_6__31_ ( .D(i_data_Rd[31]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(i_data_Rd[30]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(i_data_Rd[29]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(i_data_Rd[28]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(i_data_Rd[27]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(i_data_Rd[26]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(i_data_Rd[25]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(i_data_Rd[24]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(i_data_Rd[23]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(i_data_Rd[22]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(i_data_Rd[21]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(i_data_Rd[20]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(i_data_Rd[19]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(i_data_Rd[18]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(i_data_Rd[17]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(i_data_Rd[16]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(i_data_Rd[15]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(i_data_Rd[14]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(i_data_Rd[13]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(i_data_Rd[12]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(i_data_Rd[11]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(i_data_Rd[10]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(i_data_Rd[9]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(i_data_Rd[8]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(i_data_Rd[7]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(i_data_Rd[6]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(i_data_Rd[5]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(i_data_Rd[4]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(i_data_Rd[3]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(i_data_Rd[2]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(i_data_Rd[1]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(i_data_Rd[0]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[192]) );
  DFEC1 regs_reg_5__31_ ( .D(i_data_Rd[31]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(i_data_Rd[30]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(i_data_Rd[29]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(i_data_Rd[28]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[188]) );
  DFEC1 regs_reg_5__27_ ( .D(i_data_Rd[27]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(i_data_Rd[26]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(i_data_Rd[25]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(i_data_Rd[24]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(i_data_Rd[23]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(i_data_Rd[22]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(i_data_Rd[21]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(i_data_Rd[20]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(i_data_Rd[19]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(i_data_Rd[18]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(i_data_Rd[17]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(i_data_Rd[16]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(i_data_Rd[15]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(i_data_Rd[14]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(i_data_Rd[13]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(i_data_Rd[12]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(i_data_Rd[11]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(i_data_Rd[10]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(i_data_Rd[9]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(i_data_Rd[8]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(i_data_Rd[7]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(i_data_Rd[6]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(i_data_Rd[5]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(i_data_Rd[4]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(i_data_Rd[3]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(i_data_Rd[2]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(i_data_Rd[1]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(i_data_Rd[0]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[160]) );
  DFEC1 regs_reg_4__31_ ( .D(i_data_Rd[31]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(i_data_Rd[30]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(i_data_Rd[29]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(i_data_Rd[28]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(i_data_Rd[27]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(i_data_Rd[26]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(i_data_Rd[25]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(i_data_Rd[24]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(i_data_Rd[23]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(i_data_Rd[22]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(i_data_Rd[21]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(i_data_Rd[20]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(i_data_Rd[19]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(i_data_Rd[18]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(i_data_Rd[17]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(i_data_Rd[16]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(i_data_Rd[15]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(i_data_Rd[14]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(i_data_Rd[13]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(i_data_Rd[12]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(i_data_Rd[11]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(i_data_Rd[10]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(i_data_Rd[9]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(i_data_Rd[8]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(i_data_Rd[7]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(i_data_Rd[6]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(i_data_Rd[5]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(i_data_Rd[4]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(i_data_Rd[3]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(i_data_Rd[2]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(i_data_Rd[1]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(i_data_Rd[0]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[128]) );
  DFEC1 regs_reg_3__31_ ( .D(i_data_Rd[31]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(i_data_Rd[30]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(i_data_Rd[29]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(i_data_Rd[28]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(i_data_Rd[27]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(i_data_Rd[26]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(i_data_Rd[25]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(i_data_Rd[24]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(i_data_Rd[23]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(i_data_Rd[22]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(i_data_Rd[21]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(i_data_Rd[20]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(i_data_Rd[19]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(i_data_Rd[18]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(i_data_Rd[17]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(i_data_Rd[16]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(i_data_Rd[15]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(i_data_Rd[14]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(i_data_Rd[13]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(i_data_Rd[12]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(i_data_Rd[11]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(i_data_Rd[10]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(i_data_Rd[9]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(i_data_Rd[8]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(i_data_Rd[7]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(i_data_Rd[6]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(i_data_Rd[5]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(i_data_Rd[4]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(i_data_Rd[3]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(i_data_Rd[2]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(i_data_Rd[1]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(i_data_Rd[0]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[96]) );
  DFEC1 regs_reg_2__31_ ( .D(i_data_Rd[31]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(i_data_Rd[30]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(i_data_Rd[29]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(i_data_Rd[28]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(i_data_Rd[27]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(i_data_Rd[26]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(i_data_Rd[25]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(i_data_Rd[24]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(i_data_Rd[23]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(i_data_Rd[22]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(i_data_Rd[21]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(i_data_Rd[20]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(i_data_Rd[19]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(i_data_Rd[18]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(i_data_Rd[17]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(i_data_Rd[16]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(i_data_Rd[15]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(i_data_Rd[14]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(i_data_Rd[13]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(i_data_Rd[12]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(i_data_Rd[11]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(i_data_Rd[10]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(i_data_Rd[9]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(i_data_Rd[8]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(i_data_Rd[7]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(i_data_Rd[6]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(i_data_Rd[5]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(i_data_Rd[4]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(i_data_Rd[3]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(i_data_Rd[2]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(i_data_Rd[1]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(i_data_Rd[0]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[64]) );
  DFEC1 regs_reg_1__31_ ( .D(n1), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(n64), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(n63), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(n62), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(n61), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(n60), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(n59), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(n58), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(n57), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(n56), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(n55), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(n54), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(n53), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(n52), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(n51), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(n50), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(n49), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(n48), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(n47), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(n46), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(n45), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(n33), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(n24), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(n19), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(n14), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(n12), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(n10), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(n8), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(n7), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(n4), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(n3), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(n2), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[32]) );
  DFEC1 regs_reg_0__31_ ( .D(n1), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(n64), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(n63), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(n62), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(n61), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(n60), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(n59), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(n58), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(n57), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(n56), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(n55), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(n54), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(n53), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(n52), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(n51), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(n50), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(n49), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(n48), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(n47), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(n46), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(n45), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(n33), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(n24), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(n19), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(n14), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(n12), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(n10), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(n8), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(n7), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(n4), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(n3), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(n2), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[0]) );
  MUX21 regs_reg_31__31__U4 ( .A(regs[1023]), .B(i_data_Rd[31]), .S(n31), .Q(
        n65) );
  DFC1 regs_reg_31__31_ ( .D(n65), .C(i_clk), .RN(i_rst_n), .Q(regs[1023]) );
  BUF6 U2 ( .A(n1563), .Q(n73) );
  BUF6 U3 ( .A(n1561), .Q(n74) );
  BUF8 U4 ( .A(n1568), .Q(n68) );
  BUF8 U5 ( .A(n1567), .Q(n114) );
  BUF6 U6 ( .A(n1564), .Q(n113) );
  BUF6 U7 ( .A(n1562), .Q(n112) );
  BUF6 U8 ( .A(n839), .Q(n67) );
  BUF6 U9 ( .A(n845), .Q(n110) );
  BUF6 U10 ( .A(n842), .Q(n109) );
  BUF2 U11 ( .A(i_data_Rd[31]), .Q(n1) );
  BUF2 U12 ( .A(i_data_Rd[0]), .Q(n2) );
  BUF2 U13 ( .A(i_data_Rd[1]), .Q(n3) );
  BUF2 U14 ( .A(i_data_Rd[2]), .Q(n4) );
  BUF2 U15 ( .A(i_data_Rd[3]), .Q(n7) );
  BUF2 U16 ( .A(i_data_Rd[4]), .Q(n8) );
  BUF2 U17 ( .A(i_data_Rd[5]), .Q(n10) );
  BUF2 U18 ( .A(i_data_Rd[6]), .Q(n12) );
  BUF2 U19 ( .A(i_data_Rd[7]), .Q(n14) );
  BUF2 U20 ( .A(i_data_Rd[8]), .Q(n19) );
  BUF2 U21 ( .A(i_data_Rd[9]), .Q(n24) );
  BUF2 U22 ( .A(i_data_Rd[10]), .Q(n33) );
  BUF2 U23 ( .A(i_data_Rd[11]), .Q(n45) );
  BUF2 U24 ( .A(i_data_Rd[12]), .Q(n46) );
  BUF2 U25 ( .A(i_data_Rd[13]), .Q(n47) );
  BUF2 U26 ( .A(i_data_Rd[14]), .Q(n48) );
  BUF2 U27 ( .A(i_data_Rd[15]), .Q(n49) );
  BUF2 U28 ( .A(i_data_Rd[16]), .Q(n50) );
  BUF2 U29 ( .A(i_data_Rd[17]), .Q(n51) );
  BUF2 U30 ( .A(i_data_Rd[18]), .Q(n52) );
  BUF2 U31 ( .A(i_data_Rd[19]), .Q(n53) );
  BUF2 U32 ( .A(i_data_Rd[20]), .Q(n54) );
  BUF2 U33 ( .A(i_data_Rd[21]), .Q(n55) );
  BUF2 U34 ( .A(i_data_Rd[22]), .Q(n56) );
  BUF2 U35 ( .A(i_data_Rd[23]), .Q(n57) );
  BUF2 U36 ( .A(i_data_Rd[24]), .Q(n58) );
  BUF2 U37 ( .A(i_data_Rd[25]), .Q(n59) );
  BUF2 U38 ( .A(i_data_Rd[26]), .Q(n60) );
  BUF2 U39 ( .A(i_data_Rd[27]), .Q(n61) );
  BUF2 U40 ( .A(i_data_Rd[28]), .Q(n62) );
  BUF2 U41 ( .A(i_data_Rd[29]), .Q(n63) );
  BUF2 U42 ( .A(i_data_Rd[30]), .Q(n64) );
  NAND21 U43 ( .A(n800), .B(n799), .Q(o_data_Rt[29]) );
  AOI221 U44 ( .A(n834), .B(n590), .C(n832), .D(n589), .Q(n602) );
  AOI220 U45 ( .A(n834), .B(n282), .C(n832), .D(n281), .Q(n294) );
  AOI220 U46 ( .A(n834), .B(n722), .C(n832), .D(n721), .Q(n734) );
  AOI220 U47 ( .A(n854), .B(n798), .C(n852), .D(n797), .Q(n799) );
  AOI220 U48 ( .A(n834), .B(n678), .C(n832), .D(n677), .Q(n690) );
  AOI220 U49 ( .A(n834), .B(n348), .C(n832), .D(n347), .Q(n360) );
  AOI220 U50 ( .A(n834), .B(n216), .C(n832), .D(n215), .Q(n228) );
  AOI220 U51 ( .A(n834), .B(n194), .C(n832), .D(n193), .Q(n206) );
  AOI221 U52 ( .A(n834), .B(n568), .C(n832), .D(n567), .Q(n580) );
  AOI221 U53 ( .A(n1556), .B(n1004), .C(n1554), .D(n1003), .Q(n1016) );
  AOI221 U54 ( .A(n1556), .B(n938), .C(n1554), .D(n937), .Q(n950) );
  AOI221 U55 ( .A(n1556), .B(n1334), .C(n1554), .D(n1333), .Q(n1346) );
  AOI220 U56 ( .A(n834), .B(n172), .C(n832), .D(n171), .Q(n184) );
  AOI221 U57 ( .A(n1556), .B(n1488), .C(n1554), .D(n1487), .Q(n1500) );
  AOI220 U58 ( .A(n1556), .B(n1268), .C(n1554), .D(n1267), .Q(n1280) );
  AOI221 U59 ( .A(n1556), .B(n1290), .C(n1554), .D(n1289), .Q(n1302) );
  AOI220 U60 ( .A(n109), .B(regs[221]), .C(n71), .D(regs[157]), .Q(n795) );
  AOI220 U61 ( .A(n109), .B(regs[479]), .C(n71), .D(regs[415]), .Q(n829) );
  AOI220 U62 ( .A(n70), .B(regs[1022]), .C(n67), .D(regs[958]), .Q(n804) );
  AOI220 U63 ( .A(n70), .B(regs[765]), .C(n67), .D(regs[701]), .Q(n792) );
  AOI220 U64 ( .A(n70), .B(regs[253]), .C(n67), .D(regs[189]), .Q(n796) );
  AOI220 U65 ( .A(n109), .B(regs[733]), .C(n71), .D(regs[669]), .Q(n791) );
  AOI220 U66 ( .A(regs[704]), .B(n109), .C(regs[640]), .D(n71), .Q(n153) );
  AOI220 U67 ( .A(n70), .B(regs[761]), .C(n67), .D(regs[697]), .Q(n704) );
  AOI220 U68 ( .A(n70), .B(regs[238]), .C(n67), .D(regs[174]), .Q(n466) );
  AOI220 U69 ( .A(n109), .B(regs[478]), .C(n71), .D(regs[414]), .Q(n807) );
  AOI220 U70 ( .A(n1556), .B(n916), .C(n1554), .D(n915), .Q(n928) );
  AOI220 U71 ( .A(n109), .B(regs[222]), .C(n71), .D(regs[158]), .Q(n817) );
  AOI220 U72 ( .A(n842), .B(regs[215]), .C(n71), .D(regs[151]), .Q(n663) );
  AOI220 U73 ( .A(n70), .B(regs[249]), .C(n67), .D(regs[185]), .Q(n708) );
  AOI220 U74 ( .A(n842), .B(regs[984]), .C(n71), .D(regs[920]), .Q(n671) );
  AOI221 U75 ( .A(n70), .B(regs[743]), .C(n67), .D(regs[679]), .Q(n308) );
  AOI221 U76 ( .A(n70), .B(regs[231]), .C(n67), .D(regs[167]), .Q(n312) );
  AOI220 U77 ( .A(n109), .B(regs[735]), .C(n71), .D(regs[671]), .Q(n837) );
  AOI220 U78 ( .A(n109), .B(regs[991]), .C(n71), .D(regs[927]), .Q(n825) );
  AOI220 U79 ( .A(n109), .B(regs[734]), .C(n71), .D(regs[670]), .Q(n813) );
  AOI220 U80 ( .A(regs[736]), .B(n70), .C(regs[672]), .D(n67), .Q(n154) );
  AOI220 U81 ( .A(n70), .B(regs[504]), .C(n839), .D(regs[440]), .Q(n676) );
  AOI221 U82 ( .A(n109), .B(regs[965]), .C(n71), .D(regs[901]), .Q(n253) );
  AOI220 U83 ( .A(n109), .B(regs[960]), .C(n71), .D(regs[896]), .Q(n141) );
  AOI221 U84 ( .A(n109), .B(regs[453]), .C(n71), .D(regs[389]), .Q(n257) );
  AOI220 U85 ( .A(n70), .B(regs[248]), .C(n67), .D(regs[184]), .Q(n686) );
  AOI220 U86 ( .A(n70), .B(regs[752]), .C(n67), .D(regs[688]), .Q(n506) );
  AOI220 U87 ( .A(n70), .B(regs[508]), .C(n67), .D(regs[444]), .Q(n764) );
  AOI221 U88 ( .A(n109), .B(regs[706]), .C(n71), .D(regs[642]), .Q(n197) );
  AOI220 U89 ( .A(n109), .B(regs[989]), .C(n71), .D(regs[925]), .Q(n781) );
  AOI220 U90 ( .A(n109), .B(regs[214]), .C(n71), .D(regs[150]), .Q(n641) );
  AOI221 U91 ( .A(n70), .B(regs[1000]), .C(n67), .D(regs[936]), .Q(n320) );
  AOI220 U92 ( .A(n70), .B(regs[1021]), .C(n67), .D(regs[957]), .Q(n782) );
  AOI221 U93 ( .A(n109), .B(regs[196]), .C(n71), .D(regs[132]), .Q(n245) );
  AOI220 U94 ( .A(n109), .B(regs[726]), .C(n71), .D(regs[662]), .Q(n637) );
  AOI220 U95 ( .A(n842), .B(regs[732]), .C(n71), .D(regs[668]), .Q(n769) );
  AOI220 U96 ( .A(n109), .B(regs[708]), .C(n71), .D(regs[644]), .Q(n241) );
  AOI220 U97 ( .A(n842), .B(regs[451]), .C(n71), .D(regs[387]), .Q(n213) );
  AOI220 U98 ( .A(n109), .B(regs[470]), .C(n71), .D(regs[406]), .Q(n631) );
  AOI221 U99 ( .A(n109), .B(regs[194]), .C(n71), .D(regs[130]), .Q(n201) );
  AOI221 U100 ( .A(n70), .B(regs[484]), .C(n67), .D(regs[420]), .Q(n236) );
  AOI220 U101 ( .A(n70), .B(regs[483]), .C(n67), .D(regs[419]), .Q(n214) );
  AOI221 U102 ( .A(n70), .B(regs[996]), .C(n67), .D(regs[932]), .Q(n232) );
  AOI220 U103 ( .A(n1556), .B(n982), .C(n1554), .D(n981), .Q(n994) );
  AOI221 U104 ( .A(n70), .B(regs[742]), .C(n839), .D(regs[678]), .Q(n286) );
  AOI220 U105 ( .A(n70), .B(regs[252]), .C(n67), .D(regs[188]), .Q(n774) );
  AOI221 U106 ( .A(n70), .B(regs[227]), .C(n67), .D(regs[163]), .Q(n224) );
  AOI220 U107 ( .A(n109), .B(regs[727]), .C(n71), .D(regs[663]), .Q(n659) );
  AOI221 U108 ( .A(n70), .B(regs[738]), .C(n839), .D(regs[674]), .Q(n198) );
  AOI220 U109 ( .A(n842), .B(regs[983]), .C(n71), .D(regs[919]), .Q(n649) );
  AOI220 U110 ( .A(n109), .B(regs[477]), .C(n71), .D(regs[413]), .Q(n785) );
  AOI220 U111 ( .A(n70), .B(regs[1009]), .C(n67), .D(regs[945]), .Q(n518) );
  AOI220 U112 ( .A(n70), .B(regs[509]), .C(n67), .D(regs[445]), .Q(n786) );
  AOI221 U113 ( .A(n70), .B(regs[739]), .C(n839), .D(regs[675]), .Q(n220) );
  AOI220 U114 ( .A(n70), .B(regs[764]), .C(n67), .D(regs[700]), .Q(n770) );
  AOI220 U115 ( .A(n109), .B(regs[476]), .C(n71), .D(regs[412]), .Q(n763) );
  AOI221 U116 ( .A(n1556), .B(n960), .C(n1554), .D(n959), .Q(n972) );
  AOI220 U117 ( .A(n109), .B(regs[962]), .C(n71), .D(regs[898]), .Q(n187) );
  AOI220 U118 ( .A(regs[1000]), .B(n1562), .C(regs[936]), .D(n74), .Q(n1042)
         );
  AOI220 U119 ( .A(regs[971]), .B(n113), .C(regs[907]), .D(n73), .Q(n1107) );
  AOI220 U120 ( .A(regs[976]), .B(n113), .C(regs[912]), .D(n73), .Q(n1217) );
  AOI220 U121 ( .A(regs[508]), .B(n112), .C(regs[444]), .D(n74), .Q(n1486) );
  AOI220 U122 ( .A(regs[201]), .B(n113), .C(regs[137]), .D(n73), .Q(n1077) );
  AOI220 U123 ( .A(regs[755]), .B(n112), .C(regs[691]), .D(n74), .Q(n1294) );
  AOI220 U124 ( .A(regs[1011]), .B(n112), .C(regs[947]), .D(n74), .Q(n1284) );
  AOI220 U125 ( .A(regs[754]), .B(n112), .C(regs[690]), .D(n74), .Q(n1272) );
  AOI220 U126 ( .A(regs[202]), .B(n1564), .C(regs[138]), .D(n73), .Q(n1099) );
  AOI220 U127 ( .A(regs[459]), .B(n1564), .C(regs[395]), .D(n73), .Q(n1111) );
  AOI220 U128 ( .A(regs[200]), .B(n113), .C(regs[136]), .D(n73), .Q(n1055) );
  AOI220 U129 ( .A(n109), .B(regs[217]), .C(n71), .D(regs[153]), .Q(n707) );
  AOI221 U130 ( .A(n111), .B(regs[72]), .C(n110), .D(regs[8]), .Q(n331) );
  AOI220 U131 ( .A(n111), .B(regs[71]), .C(n110), .D(regs[7]), .Q(n309) );
  AOI220 U132 ( .A(regs[966]), .B(n113), .C(regs[902]), .D(n73), .Q(n997) );
  AOI220 U133 ( .A(regs[503]), .B(n112), .C(regs[439]), .D(n74), .Q(n1376) );
  AOI220 U134 ( .A(regs[743]), .B(n112), .C(regs[679]), .D(n74), .Q(n1030) );
  AOI220 U135 ( .A(regs[480]), .B(n1562), .C(regs[416]), .D(n74), .Q(n869) );
  AOI221 U136 ( .A(n111), .B(regs[584]), .C(n110), .D(regs[520]), .Q(n327) );
  AOI220 U137 ( .A(n109), .B(regs[986]), .C(n71), .D(regs[922]), .Q(n715) );
  AOI220 U138 ( .A(n111), .B(regs[344]), .C(n110), .D(regs[280]), .Q(n673) );
  AOI220 U139 ( .A(n109), .B(regs[471]), .C(n71), .D(regs[407]), .Q(n653) );
  AOI220 U140 ( .A(regs[981]), .B(n113), .C(regs[917]), .D(n73), .Q(n1327) );
  AOI220 U141 ( .A(n111), .B(regs[858]), .C(n110), .D(regs[794]), .Q(n713) );
  AOI220 U142 ( .A(regs[985]), .B(n1564), .C(regs[921]), .D(n73), .Q(n1415) );
  AOI220 U143 ( .A(n109), .B(regs[474]), .C(n71), .D(regs[410]), .Q(n719) );
  AOI220 U144 ( .A(regs[1015]), .B(n112), .C(regs[951]), .D(n74), .Q(n1372) );
  AOI220 U145 ( .A(n111), .B(regs[74]), .C(n110), .D(regs[10]), .Q(n375) );
  AOI220 U146 ( .A(n70), .B(regs[245]), .C(n839), .D(regs[181]), .Q(n620) );
  AOI220 U147 ( .A(n109), .B(regs[730]), .C(n71), .D(regs[666]), .Q(n725) );
  AOI220 U148 ( .A(n109), .B(regs[472]), .C(n71), .D(regs[408]), .Q(n675) );
  AOI220 U149 ( .A(n109), .B(regs[985]), .C(n71), .D(regs[921]), .Q(n693) );
  AOI221 U150 ( .A(n111), .B(regs[73]), .C(n110), .D(regs[9]), .Q(n353) );
  AOI220 U151 ( .A(n111), .B(regs[88]), .C(n110), .D(regs[24]), .Q(n683) );
  AOI220 U152 ( .A(n111), .B(regs[857]), .C(n110), .D(regs[793]), .Q(n691) );
  AOI220 U153 ( .A(regs[469]), .B(n113), .C(regs[405]), .D(n73), .Q(n1331) );
  AOI220 U154 ( .A(n111), .B(regs[327]), .C(n110), .D(regs[263]), .Q(n299) );
  AOI221 U155 ( .A(n111), .B(regs[585]), .C(n110), .D(regs[521]), .Q(n349) );
  AOI220 U156 ( .A(n109), .B(regs[216]), .C(n71), .D(regs[152]), .Q(n685) );
  AOI221 U157 ( .A(n111), .B(regs[842]), .C(n110), .D(regs[778]), .Q(n361) );
  AOI220 U158 ( .A(regs[449]), .B(n113), .C(regs[385]), .D(n73), .Q(n891) );
  AOI221 U159 ( .A(n111), .B(regs[345]), .C(n110), .D(regs[281]), .Q(n695) );
  AOI221 U160 ( .A(n111), .B(regs[329]), .C(n110), .D(regs[265]), .Q(n343) );
  AOI220 U161 ( .A(n111), .B(regs[600]), .C(n110), .D(regs[536]), .Q(n679) );
  AOI221 U162 ( .A(n111), .B(regs[330]), .C(n110), .D(regs[266]), .Q(n365) );
  AOI221 U163 ( .A(n111), .B(regs[841]), .C(n110), .D(regs[777]), .Q(n339) );
  AOI220 U164 ( .A(n111), .B(regs[601]), .C(n110), .D(regs[537]), .Q(n701) );
  AOI220 U165 ( .A(regs[742]), .B(n112), .C(regs[678]), .D(n74), .Q(n1008) );
  AOI220 U166 ( .A(n109), .B(regs[475]), .C(n71), .D(regs[411]), .Q(n741) );
  AOI220 U167 ( .A(n111), .B(regs[844]), .C(n110), .D(regs[780]), .Q(n405) );
  AOI220 U168 ( .A(n109), .B(regs[731]), .C(n71), .D(regs[667]), .Q(n747) );
  AOI220 U169 ( .A(n109), .B(regs[988]), .C(n71), .D(regs[924]), .Q(n759) );
  AOI220 U170 ( .A(n111), .B(regs[583]), .C(n110), .D(regs[519]), .Q(n305) );
  AOI220 U171 ( .A(n111), .B(regs[331]), .C(n110), .D(regs[267]), .Q(n387) );
  AOI220 U172 ( .A(n109), .B(regs[219]), .C(n71), .D(regs[155]), .Q(n751) );
  AOI220 U173 ( .A(regs[246]), .B(n112), .C(regs[182]), .D(n74), .Q(n1364) );
  AOI220 U174 ( .A(regs[504]), .B(n112), .C(regs[440]), .D(n74), .Q(n1398) );
  AOI220 U175 ( .A(regs[729]), .B(n113), .C(regs[665]), .D(n73), .Q(n1425) );
  AOI220 U176 ( .A(regs[724]), .B(n113), .C(regs[660]), .D(n73), .Q(n1315) );
  AOI220 U177 ( .A(n111), .B(regs[587]), .C(n110), .D(regs[523]), .Q(n393) );
  AOI220 U178 ( .A(n109), .B(regs[987]), .C(n71), .D(regs[923]), .Q(n737) );
  AOI220 U179 ( .A(regs[244]), .B(n112), .C(regs[180]), .D(n74), .Q(n1320) );
  AOI220 U180 ( .A(n109), .B(regs[218]), .C(n71), .D(regs[154]), .Q(n729) );
  AOI220 U181 ( .A(regs[470]), .B(n113), .C(regs[406]), .D(n73), .Q(n1353) );
  AOI220 U182 ( .A(regs[632]), .B(n69), .C(regs[568]), .D(n72), .Q(n1402) );
  AOI220 U183 ( .A(regs[893]), .B(n1566), .C(regs[829]), .D(n72), .Q(n1502) );
  AOI220 U184 ( .A(regs[116]), .B(n69), .C(regs[52]), .D(n72), .Q(n1318) );
  AOI220 U185 ( .A(regs[727]), .B(n113), .C(regs[663]), .D(n73), .Q(n1381) );
  AOI220 U186 ( .A(regs[738]), .B(n112), .C(regs[674]), .D(n74), .Q(n920) );
  AOI220 U187 ( .A(regs[766]), .B(n112), .C(regs[702]), .D(n74), .Q(n1536) );
  AOI220 U188 ( .A(regs[706]), .B(n113), .C(regs[642]), .D(n73), .Q(n919) );
  AOI220 U189 ( .A(regs[99]), .B(n69), .C(regs[35]), .D(n72), .Q(n944) );
  AOI220 U190 ( .A(regs[984]), .B(n113), .C(regs[920]), .D(n73), .Q(n1393) );
  AOI220 U191 ( .A(regs[883]), .B(n1566), .C(regs[819]), .D(n72), .Q(n1282) );
  AOI220 U192 ( .A(regs[611]), .B(n1566), .C(regs[547]), .D(n72), .Q(n940) );
  AOI220 U193 ( .A(regs[979]), .B(n113), .C(regs[915]), .D(n73), .Q(n1283) );
  AOI220 U194 ( .A(regs[226]), .B(n112), .C(regs[162]), .D(n74), .Q(n924) );
  AOI220 U195 ( .A(regs[472]), .B(n113), .C(regs[408]), .D(n73), .Q(n1397) );
  AOI220 U196 ( .A(regs[983]), .B(n113), .C(regs[919]), .D(n73), .Q(n1371) );
  AOI220 U197 ( .A(regs[735]), .B(n113), .C(regs[671]), .D(n73), .Q(n1559) );
  AOI220 U198 ( .A(regs[1009]), .B(n112), .C(regs[945]), .D(n74), .Q(n1240) );
  BUF12 U199 ( .A(n840), .Q(n70) );
  AOI220 U200 ( .A(regs[380]), .B(n69), .C(regs[316]), .D(n72), .Q(n1484) );
  AOI220 U201 ( .A(regs[467]), .B(n113), .C(regs[403]), .D(n73), .Q(n1287) );
  AOI220 U202 ( .A(regs[369]), .B(n69), .C(regs[305]), .D(n72), .Q(n1242) );
  AOI220 U203 ( .A(regs[1008]), .B(n112), .C(regs[944]), .D(n74), .Q(n1218) );
  AOI220 U204 ( .A(regs[890]), .B(n69), .C(regs[826]), .D(n72), .Q(n1436) );
  AOI220 U205 ( .A(regs[888]), .B(n69), .C(regs[824]), .D(n72), .Q(n1392) );
  AOI220 U206 ( .A(regs[723]), .B(n113), .C(regs[659]), .D(n73), .Q(n1293) );
  AOI220 U207 ( .A(regs[240]), .B(n112), .C(regs[176]), .D(n74), .Q(n1232) );
  AOI220 U208 ( .A(regs[636]), .B(n69), .C(regs[572]), .D(n72), .Q(n1490) );
  AOI220 U209 ( .A(regs[476]), .B(n113), .C(regs[412]), .D(n73), .Q(n1485) );
  BUF6 U210 ( .A(n843), .Q(n75) );
  AOI220 U211 ( .A(regs[765]), .B(n112), .C(regs[701]), .D(n74), .Q(n1514) );
  AOI220 U212 ( .A(regs[119]), .B(n69), .C(regs[55]), .D(n72), .Q(n1384) );
  AOI220 U213 ( .A(regs[502]), .B(n112), .C(regs[438]), .D(n74), .Q(n1354) );
  AOI220 U214 ( .A(regs[353]), .B(n1566), .C(regs[289]), .D(n72), .Q(n890) );
  AOI220 U215 ( .A(regs[871]), .B(n69), .C(regs[807]), .D(n72), .Q(n1018) );
  AOI220 U216 ( .A(regs[1001]), .B(n112), .C(regs[937]), .D(n74), .Q(n1064) );
  AOI220 U217 ( .A(regs[493]), .B(n112), .C(regs[429]), .D(n74), .Q(n1156) );
  AOI220 U218 ( .A(regs[712]), .B(n113), .C(regs[648]), .D(n73), .Q(n1051) );
  AOI220 U219 ( .A(regs[361]), .B(n69), .C(regs[297]), .D(n72), .Q(n1066) );
  AOI220 U220 ( .A(regs[617]), .B(n1566), .C(regs[553]), .D(n72), .Q(n1072) );
  AOI220 U221 ( .A(regs[363]), .B(n1566), .C(regs[299]), .D(n72), .Q(n1110) );
  AOI220 U222 ( .A(regs[749]), .B(n112), .C(regs[685]), .D(n74), .Q(n1162) );
  AOI220 U223 ( .A(regs[621]), .B(n1566), .C(regs[557]), .D(n72), .Q(n1160) );
  AOI220 U224 ( .A(regs[237]), .B(n112), .C(regs[173]), .D(n74), .Q(n1166) );
  AOI220 U225 ( .A(regs[358]), .B(n1566), .C(regs[294]), .D(n72), .Q(n1000) );
  AOI220 U226 ( .A(regs[96]), .B(n1566), .C(regs[32]), .D(n72), .Q(n878) );
  AOI220 U227 ( .A(regs[492]), .B(n112), .C(regs[428]), .D(n74), .Q(n1134) );
  AOI220 U228 ( .A(regs[711]), .B(n113), .C(regs[647]), .D(n73), .Q(n1029) );
  AOI220 U229 ( .A(regs[615]), .B(n69), .C(regs[551]), .D(n72), .Q(n1028) );
  AOI220 U230 ( .A(regs[870]), .B(n1566), .C(regs[806]), .D(n72), .Q(n996) );
  AOI220 U231 ( .A(regs[1003]), .B(n112), .C(regs[939]), .D(n74), .Q(n1108) );
  AOI220 U232 ( .A(regs[708]), .B(n113), .C(regs[644]), .D(n73), .Q(n963) );
  AOI220 U233 ( .A(regs[356]), .B(n69), .C(regs[292]), .D(n72), .Q(n956) );
  AOI220 U234 ( .A(regs[236]), .B(n112), .C(regs[172]), .D(n74), .Q(n1144) );
  AOI220 U235 ( .A(regs[110]), .B(n69), .C(regs[46]), .D(n72), .Q(n1186) );
  NOR22 U236 ( .A(n1588), .B(n1581), .Q(n40) );
  AOI220 U237 ( .A(regs[490]), .B(n112), .C(regs[426]), .D(n74), .Q(n1090) );
  AOI220 U238 ( .A(regs[960]), .B(n113), .C(regs[896]), .D(n73), .Q(n863) );
  AOI220 U239 ( .A(regs[618]), .B(n1566), .C(regs[554]), .D(n72), .Q(n1094) );
  AOI220 U240 ( .A(regs[874]), .B(n1566), .C(regs[810]), .D(n72), .Q(n1084) );
  AOI220 U241 ( .A(regs[232]), .B(n112), .C(regs[168]), .D(n74), .Q(n1056) );
  AOI220 U242 ( .A(regs[108]), .B(n69), .C(regs[44]), .D(n72), .Q(n1142) );
  NOR22 U243 ( .A(n1584), .B(n1581), .Q(n37) );
  BUF6 U244 ( .A(n841), .Q(n71) );
  BUF15 U245 ( .A(n844), .Q(n66) );
  NOR22 U246 ( .A(n1590), .B(n1582), .Q(n29) );
  NOR22 U247 ( .A(n1588), .B(n1582), .Q(n31) );
  NOR22 U248 ( .A(n1589), .B(n1582), .Q(n30) );
  NOR22 U249 ( .A(n1584), .B(n1582), .Q(n28) );
  BUF8 U250 ( .A(n1565), .Q(n72) );
  BUF6 U251 ( .A(n1566), .Q(n69) );
  NAND22 U252 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[1]), .Q(n858) );
  AOI220 U253 ( .A(n834), .B(n524), .C(n832), .D(n523), .Q(n536) );
  AOI220 U254 ( .A(n834), .B(n833), .C(n832), .D(n831), .Q(n856) );
  AOI220 U255 ( .A(n834), .B(n480), .C(n832), .D(n479), .Q(n492) );
  AOI220 U256 ( .A(n834), .B(n502), .C(n832), .D(n501), .Q(n514) );
  AOI220 U257 ( .A(n834), .B(n656), .C(n832), .D(n655), .Q(n668) );
  AOI220 U258 ( .A(n834), .B(n546), .C(n832), .D(n545), .Q(n558) );
  AOI220 U259 ( .A(n834), .B(n304), .C(n832), .D(n303), .Q(n316) );
  AOI220 U260 ( .A(n834), .B(n458), .C(n832), .D(n457), .Q(n470) );
  AOI220 U261 ( .A(n834), .B(n436), .C(n832), .D(n435), .Q(n448) );
  AOI220 U262 ( .A(n834), .B(n766), .C(n832), .D(n765), .Q(n778) );
  AOI220 U263 ( .A(n834), .B(n700), .C(n832), .D(n699), .Q(n712) );
  AOI220 U264 ( .A(n834), .B(n149), .C(n832), .D(n148), .Q(n162) );
  AOI220 U265 ( .A(n834), .B(n810), .C(n832), .D(n809), .Q(n822) );
  AOI220 U266 ( .A(n834), .B(n788), .C(n832), .D(n787), .Q(n800) );
  AOI220 U267 ( .A(n834), .B(n392), .C(n832), .D(n391), .Q(n404) );
  AOI220 U268 ( .A(n834), .B(n744), .C(n832), .D(n743), .Q(n756) );
  AOI220 U269 ( .A(n109), .B(regs[967]), .C(n841), .D(regs[903]), .Q(n297) );
  AOI220 U270 ( .A(n66), .B(regs[894]), .C(n75), .D(regs[830]), .Q(n802) );
  AOI220 U271 ( .A(n66), .B(regs[620]), .C(n75), .D(regs[556]), .Q(n416) );
  AOI220 U272 ( .A(n66), .B(regs[380]), .C(n75), .D(regs[316]), .Q(n762) );
  AOI220 U273 ( .A(n66), .B(regs[375]), .C(n75), .D(regs[311]), .Q(n652) );
  AOI220 U274 ( .A(n66), .B(regs[627]), .C(n75), .D(regs[563]), .Q(n570) );
  AOI220 U275 ( .A(n66), .B(regs[125]), .C(n75), .D(regs[61]), .Q(n794) );
  AOI220 U276 ( .A(n66), .B(regs[371]), .C(n75), .D(regs[307]), .Q(n564) );
  AOI220 U277 ( .A(n66), .B(regs[636]), .C(n75), .D(regs[572]), .Q(n768) );
  AOI220 U278 ( .A(n66), .B(regs[883]), .C(n75), .D(regs[819]), .Q(n560) );
  AOI221 U279 ( .A(n111), .B(regs[332]), .C(n845), .D(regs[268]), .Q(n409) );
  AOI220 U280 ( .A(n66), .B(regs[381]), .C(n75), .D(regs[317]), .Q(n784) );
  AOI220 U281 ( .A(n66), .B(regs[124]), .C(n75), .D(regs[60]), .Q(n772) );
  AOI220 U282 ( .A(n66), .B(regs[373]), .C(n75), .D(regs[309]), .Q(n608) );
  AOI220 U283 ( .A(n66), .B(regs[126]), .C(n75), .D(regs[62]), .Q(n816) );
  AOI220 U284 ( .A(n66), .B(regs[895]), .C(n75), .D(regs[831]), .Q(n824) );
  AOI220 U285 ( .A(n66), .B(regs[629]), .C(n75), .D(regs[565]), .Q(n614) );
  AOI220 U286 ( .A(n66), .B(regs[383]), .C(n75), .D(regs[319]), .Q(n828) );
  AOI220 U287 ( .A(n66), .B(regs[639]), .C(n75), .D(regs[575]), .Q(n836) );
  AOI220 U288 ( .A(n66), .B(regs[630]), .C(n75), .D(regs[566]), .Q(n636) );
  AOI220 U289 ( .A(n66), .B(regs[626]), .C(n75), .D(regs[562]), .Q(n548) );
  AOI220 U290 ( .A(regs[608]), .B(n66), .C(regs[544]), .D(n75), .Q(n152) );
  AOI220 U291 ( .A(n66), .B(regs[621]), .C(n75), .D(regs[557]), .Q(n438) );
  AOI220 U292 ( .A(n66), .B(regs[109]), .C(n75), .D(regs[45]), .Q(n442) );
  AOI220 U293 ( .A(n66), .B(regs[370]), .C(n75), .D(regs[306]), .Q(n542) );
  AOI220 U294 ( .A(n66), .B(regs[878]), .C(n75), .D(regs[814]), .Q(n450) );
  AOI220 U295 ( .A(n66), .B(regs[631]), .C(n75), .D(regs[567]), .Q(n658) );
  AOI220 U296 ( .A(n66), .B(regs[376]), .C(n75), .D(regs[312]), .Q(n674) );
  AOI220 U297 ( .A(n66), .B(regs[633]), .C(n75), .D(regs[569]), .Q(n702) );
  AOI220 U298 ( .A(n66), .B(regs[366]), .C(n75), .D(regs[302]), .Q(n454) );
  AOI220 U299 ( .A(n111), .B(regs[89]), .C(n110), .D(regs[25]), .Q(n705) );
  AOI220 U300 ( .A(n66), .B(regs[108]), .C(n75), .D(regs[44]), .Q(n420) );
  AOI220 U301 ( .A(n66), .B(regs[119]), .C(n75), .D(regs[55]), .Q(n662) );
  AOI220 U302 ( .A(n111), .B(regs[834]), .C(n110), .D(regs[770]), .Q(n185) );
  AOI220 U303 ( .A(n66), .B(regs[114]), .C(n75), .D(regs[50]), .Q(n552) );
  AOI220 U304 ( .A(n66), .B(regs[877]), .C(n75), .D(regs[813]), .Q(n428) );
  AOI220 U305 ( .A(n111), .B(regs[322]), .C(n110), .D(regs[258]), .Q(n189) );
  AOI220 U306 ( .A(regs[593]), .B(n68), .C(regs[529]), .D(n114), .Q(n1247) );
  AOI220 U307 ( .A(regs[848]), .B(n68), .C(regs[784]), .D(n114), .Q(n1215) );
  AOI220 U308 ( .A(regs[852]), .B(n68), .C(regs[788]), .D(n114), .Q(n1303) );
  AOI220 U309 ( .A(regs[81]), .B(n68), .C(regs[17]), .D(n114), .Q(n1251) );
  AOI220 U310 ( .A(regs[596]), .B(n68), .C(regs[532]), .D(n114), .Q(n1313) );
  AOI220 U311 ( .A(regs[597]), .B(n68), .C(regs[533]), .D(n114), .Q(n1335) );
  AOI220 U312 ( .A(regs[84]), .B(n68), .C(regs[20]), .D(n114), .Q(n1317) );
  AOI220 U313 ( .A(regs[853]), .B(n68), .C(regs[789]), .D(n114), .Q(n1325) );
  AOI220 U314 ( .A(regs[851]), .B(n68), .C(regs[787]), .D(n114), .Q(n1281) );
  AOI220 U315 ( .A(regs[339]), .B(n68), .C(regs[275]), .D(n114), .Q(n1285) );
  AOI220 U316 ( .A(regs[595]), .B(n68), .C(regs[531]), .D(n114), .Q(n1291) );
  AOI220 U317 ( .A(regs[598]), .B(n68), .C(regs[534]), .D(n114), .Q(n1357) );
  AOI220 U318 ( .A(regs[83]), .B(n68), .C(regs[19]), .D(n114), .Q(n1295) );
  AOI220 U319 ( .A(regs[850]), .B(n68), .C(regs[786]), .D(n114), .Q(n1259) );
  AOI220 U320 ( .A(regs[338]), .B(n68), .C(regs[274]), .D(n114), .Q(n1263) );
  AOI220 U321 ( .A(regs[594]), .B(n68), .C(regs[530]), .D(n114), .Q(n1269) );
  AOI220 U322 ( .A(regs[82]), .B(n68), .C(regs[18]), .D(n114), .Q(n1273) );
  NOR22 U323 ( .A(n1591), .B(n1584), .Q(n5) );
  AOI220 U324 ( .A(regs[849]), .B(n68), .C(regs[785]), .D(n114), .Q(n1237) );
  AOI220 U325 ( .A(regs[863]), .B(n68), .C(regs[799]), .D(n114), .Q(n1545) );
  AOI220 U326 ( .A(regs[604]), .B(n68), .C(regs[540]), .D(n114), .Q(n1489) );
  AOI220 U327 ( .A(regs[92]), .B(n68), .C(regs[28]), .D(n114), .Q(n1493) );
  NOR22 U328 ( .A(n1591), .B(n1588), .Q(n11) );
  AOI220 U329 ( .A(regs[76]), .B(n68), .C(regs[12]), .D(n114), .Q(n1141) );
  AOI220 U330 ( .A(regs[93]), .B(n68), .C(regs[29]), .D(n114), .Q(n1515) );
  AOI220 U331 ( .A(regs[605]), .B(n68), .C(regs[541]), .D(n114), .Q(n1511) );
  AOI220 U332 ( .A(regs[861]), .B(n68), .C(regs[797]), .D(n114), .Q(n1501) );
  AOI220 U333 ( .A(regs[94]), .B(n68), .C(regs[30]), .D(n114), .Q(n1537) );
  AOI220 U334 ( .A(regs[606]), .B(n68), .C(regs[542]), .D(n114), .Q(n1533) );
  NOR22 U335 ( .A(n1581), .B(n1590), .Q(n38) );
  NOR22 U336 ( .A(n1581), .B(n1589), .Q(n39) );
  AOI220 U337 ( .A(regs[862]), .B(n68), .C(regs[798]), .D(n114), .Q(n1523) );
  AOI220 U338 ( .A(regs[860]), .B(n68), .C(regs[796]), .D(n114), .Q(n1479) );
  AOI220 U339 ( .A(regs[607]), .B(n68), .C(regs[543]), .D(n114), .Q(n1557) );
  AOI220 U340 ( .A(regs[588]), .B(n68), .C(regs[524]), .D(n114), .Q(n1137) );
  AOI220 U341 ( .A(regs[845]), .B(n68), .C(regs[781]), .D(n114), .Q(n1149) );
  BUF6 U342 ( .A(n846), .Q(n111) );
  AOI220 U343 ( .A(regs[78]), .B(n68), .C(regs[14]), .D(n114), .Q(n1185) );
  AOI220 U344 ( .A(regs[333]), .B(n68), .C(regs[269]), .D(n114), .Q(n1153) );
  AOI220 U345 ( .A(regs[79]), .B(n68), .C(regs[15]), .D(n114), .Q(n1207) );
  AOI220 U346 ( .A(regs[589]), .B(n68), .C(regs[525]), .D(n114), .Q(n1159) );
  NOR22 U347 ( .A(n1591), .B(n1590), .Q(n6) );
  AOI220 U348 ( .A(regs[77]), .B(n68), .C(regs[13]), .D(n114), .Q(n1163) );
  AOI220 U349 ( .A(regs[80]), .B(n68), .C(regs[16]), .D(n114), .Q(n1229) );
  NOR22 U350 ( .A(n1591), .B(n1589), .Q(n9) );
  NOR22 U351 ( .A(n143), .B(n150), .Q(n834) );
  NOR22 U352 ( .A(i_addr_Rt_4_), .B(n143), .Q(n832) );
  NOR22 U353 ( .A(i_addr_Rs[4]), .B(n865), .Q(n1554) );
  NOR22 U354 ( .A(i_addr_Rs[3]), .B(i_addr_Rs[4]), .Q(n1574) );
  NOR22 U355 ( .A(i_addr_Rt_3_), .B(i_addr_Rt_4_), .Q(n852) );
  AOI221 U356 ( .A(n1576), .B(n1498), .C(n1574), .D(n1497), .Q(n1499) );
  AOI221 U357 ( .A(n1576), .B(n1146), .C(n1574), .D(n1145), .Q(n1147) );
  AOI221 U358 ( .A(n1576), .B(n1322), .C(n1574), .D(n1321), .Q(n1323) );
  AOI221 U359 ( .A(n1576), .B(n948), .C(n1574), .D(n947), .Q(n949) );
  AOI221 U360 ( .A(n1576), .B(n882), .C(n1574), .D(n881), .Q(n883) );
  AOI221 U361 ( .A(n1576), .B(n970), .C(n1574), .D(n969), .Q(n971) );
  AOI221 U362 ( .A(n1576), .B(n1124), .C(n1574), .D(n1123), .Q(n1125) );
  AOI221 U363 ( .A(n1576), .B(n1366), .C(n1574), .D(n1365), .Q(n1367) );
  AOI220 U364 ( .A(n70), .B(regs[490]), .C(n67), .D(regs[426]), .Q(n368) );
  AOI220 U365 ( .A(n109), .B(regs[460]), .C(n71), .D(regs[396]), .Q(n411) );
  AOI220 U366 ( .A(n109), .B(regs[458]), .C(n71), .D(regs[394]), .Q(n367) );
  AOI220 U367 ( .A(n109), .B(regs[201]), .C(n71), .D(regs[137]), .Q(n355) );
  AOI220 U368 ( .A(n70), .B(regs[1003]), .C(n67), .D(regs[939]), .Q(n386) );
  AOI220 U369 ( .A(n70), .B(regs[748]), .C(n67), .D(regs[684]), .Q(n418) );
  AOI220 U370 ( .A(n109), .B(regs[452]), .C(n71), .D(regs[388]), .Q(n235) );
  AOI220 U371 ( .A(n70), .B(regs[1001]), .C(n67), .D(regs[937]), .Q(n342) );
  AOI220 U372 ( .A(n111), .B(regs[607]), .C(n110), .D(regs[543]), .Q(n835) );
  AOI220 U373 ( .A(n109), .B(regs[982]), .C(n71), .D(regs[918]), .Q(n627) );
  AOI220 U374 ( .A(n109), .B(regs[966]), .C(n71), .D(regs[902]), .Q(n275) );
  AOI220 U375 ( .A(n109), .B(regs[970]), .C(n71), .D(regs[906]), .Q(n363) );
  AOI220 U376 ( .A(n109), .B(regs[961]), .C(n71), .D(regs[897]), .Q(n165) );
  AOI220 U377 ( .A(n70), .B(regs[236]), .C(n67), .D(regs[172]), .Q(n422) );
  AOI220 U378 ( .A(n70), .B(regs[745]), .C(n67), .D(regs[681]), .Q(n352) );
  AOI220 U379 ( .A(n111), .B(regs[94]), .C(n110), .D(regs[30]), .Q(n815) );
  AOI220 U380 ( .A(n109), .B(regs[971]), .C(n71), .D(regs[907]), .Q(n385) );
  AOI220 U381 ( .A(n70), .B(regs[1002]), .C(n67), .D(regs[938]), .Q(n364) );
  AOI220 U382 ( .A(n109), .B(regs[200]), .C(n71), .D(regs[136]), .Q(n333) );
  AOI220 U383 ( .A(n109), .B(regs[705]), .C(n71), .D(regs[641]), .Q(n175) );
  AOI220 U384 ( .A(n109), .B(regs[969]), .C(n71), .D(regs[905]), .Q(n341) );
  AOI220 U385 ( .A(n109), .B(regs[448]), .C(n71), .D(regs[384]), .Q(n146) );
  AOI220 U386 ( .A(n109), .B(regs[972]), .C(n71), .D(regs[908]), .Q(n407) );
  AOI220 U387 ( .A(n70), .B(regs[1004]), .C(n67), .D(regs[940]), .Q(n408) );
  AOI220 U388 ( .A(n70), .B(regs[491]), .C(n67), .D(regs[427]), .Q(n390) );
  AOI220 U389 ( .A(n70), .B(regs[255]), .C(n67), .D(regs[191]), .Q(n850) );
  AOI220 U390 ( .A(n111), .B(regs[351]), .C(n110), .D(regs[287]), .Q(n827) );
  AOI220 U391 ( .A(n70), .B(regs[746]), .C(n67), .D(regs[682]), .Q(n374) );
  AOI220 U392 ( .A(n109), .B(regs[203]), .C(n71), .D(regs[139]), .Q(n399) );
  AOI220 U393 ( .A(n109), .B(regs[459]), .C(n71), .D(regs[395]), .Q(n389) );
  AOI221 U394 ( .A(n1576), .B(n904), .C(n1574), .D(n903), .Q(n905) );
  AOI220 U395 ( .A(n109), .B(regs[202]), .C(n71), .D(regs[138]), .Q(n377) );
  AOI220 U396 ( .A(n70), .B(regs[233]), .C(n67), .D(regs[169]), .Q(n356) );
  AOI220 U397 ( .A(n109), .B(regs[714]), .C(n841), .D(regs[650]), .Q(n373) );
  AOI220 U398 ( .A(n109), .B(regs[715]), .C(n841), .D(regs[651]), .Q(n395) );
  AOI220 U399 ( .A(n109), .B(regs[709]), .C(n71), .D(regs[645]), .Q(n263) );
  AOI220 U400 ( .A(n109), .B(regs[713]), .C(n71), .D(regs[649]), .Q(n351) );
  AOI220 U401 ( .A(n70), .B(regs[747]), .C(n67), .D(regs[683]), .Q(n396) );
  AOI220 U402 ( .A(n70), .B(regs[489]), .C(n67), .D(regs[425]), .Q(n346) );
  AOI220 U403 ( .A(n70), .B(regs[234]), .C(n67), .D(regs[170]), .Q(n378) );
  AOI220 U404 ( .A(n109), .B(regs[197]), .C(n71), .D(regs[133]), .Q(n267) );
  AOI220 U405 ( .A(n109), .B(regs[449]), .C(n71), .D(regs[385]), .Q(n169) );
  AOI220 U406 ( .A(n109), .B(regs[457]), .C(n71), .D(regs[393]), .Q(n345) );
  AOI220 U407 ( .A(n842), .B(regs[199]), .C(n71), .D(regs[135]), .Q(n311) );
  AOI220 U408 ( .A(n109), .B(regs[712]), .C(n71), .D(regs[648]), .Q(n329) );
  AOI220 U409 ( .A(n109), .B(regs[724]), .C(n71), .D(regs[660]), .Q(n593) );
  AOI220 U410 ( .A(n70), .B(regs[744]), .C(n67), .D(regs[680]), .Q(n330) );
  AOI220 U411 ( .A(n70), .B(regs[750]), .C(n67), .D(regs[686]), .Q(n462) );
  AOI220 U412 ( .A(n842), .B(regs[466]), .C(n71), .D(regs[402]), .Q(n543) );
  AOI220 U413 ( .A(n842), .B(regs[456]), .C(n71), .D(regs[392]), .Q(n323) );
  AOI220 U414 ( .A(n109), .B(regs[980]), .C(n71), .D(regs[916]), .Q(n583) );
  AOI220 U415 ( .A(n109), .B(regs[464]), .C(n71), .D(regs[400]), .Q(n499) );
  AOI220 U416 ( .A(n70), .B(regs[1007]), .C(n67), .D(regs[943]), .Q(n474) );
  AOI220 U417 ( .A(n109), .B(regs[722]), .C(n841), .D(regs[658]), .Q(n549) );
  AOI220 U418 ( .A(n109), .B(regs[211]), .C(n71), .D(regs[147]), .Q(n575) );
  AOI220 U419 ( .A(n842), .B(regs[198]), .C(n71), .D(regs[134]), .Q(n289) );
  AOI220 U420 ( .A(n70), .B(regs[496]), .C(n67), .D(regs[432]), .Q(n500) );
  AOI220 U421 ( .A(n109), .B(regs[220]), .C(n841), .D(regs[156]), .Q(n773) );
  AOI220 U422 ( .A(n109), .B(regs[723]), .C(n841), .D(regs[659]), .Q(n571) );
  AOI220 U423 ( .A(n70), .B(regs[495]), .C(n67), .D(regs[431]), .Q(n478) );
  AOI220 U424 ( .A(n842), .B(regs[968]), .C(n71), .D(regs[904]), .Q(n319) );
  AOI220 U425 ( .A(n109), .B(regs[467]), .C(n71), .D(regs[403]), .Q(n565) );
  AOI220 U426 ( .A(n842), .B(regs[990]), .C(n841), .D(regs[926]), .Q(n803) );
  AOI220 U427 ( .A(n109), .B(regs[450]), .C(n71), .D(regs[386]), .Q(n191) );
  AOI220 U428 ( .A(n842), .B(regs[210]), .C(n71), .D(regs[146]), .Q(n553) );
  AOI220 U429 ( .A(n109), .B(regs[979]), .C(n71), .D(regs[915]), .Q(n561) );
  AOI220 U430 ( .A(n70), .B(regs[1008]), .C(n67), .D(regs[944]), .Q(n496) );
  AOI220 U431 ( .A(n109), .B(regs[192]), .C(n71), .D(regs[128]), .Q(n157) );
  AOI220 U432 ( .A(n70), .B(regs[749]), .C(n67), .D(regs[685]), .Q(n440) );
  AOI220 U433 ( .A(n109), .B(regs[454]), .C(n71), .D(regs[390]), .Q(n279) );
  AOI220 U434 ( .A(n70), .B(regs[995]), .C(n67), .D(regs[931]), .Q(n210) );
  AOI220 U435 ( .A(n842), .B(regs[455]), .C(n71), .D(regs[391]), .Q(n301) );
  AOI220 U436 ( .A(n70), .B(regs[232]), .C(n67), .D(regs[168]), .Q(n334) );
  AOI220 U437 ( .A(n109), .B(regs[711]), .C(n71), .D(regs[647]), .Q(n307) );
  AOI220 U438 ( .A(n70), .B(regs[241]), .C(n67), .D(regs[177]), .Q(n532) );
  AOI220 U439 ( .A(n109), .B(regs[193]), .C(n71), .D(regs[129]), .Q(n179) );
  AOI220 U440 ( .A(n842), .B(regs[195]), .C(n71), .D(regs[131]), .Q(n223) );
  AOI220 U441 ( .A(n109), .B(regs[707]), .C(n71), .D(regs[643]), .Q(n219) );
  AOI220 U442 ( .A(n842), .B(regs[963]), .C(n71), .D(regs[899]), .Q(n209) );
  AOI220 U443 ( .A(n109), .B(regs[725]), .C(n841), .D(regs[661]), .Q(n615) );
  AOI220 U444 ( .A(n109), .B(regs[981]), .C(n71), .D(regs[917]), .Q(n605) );
  AOI220 U445 ( .A(n842), .B(regs[212]), .C(n71), .D(regs[148]), .Q(n597) );
  AOI220 U446 ( .A(n109), .B(regs[465]), .C(n71), .D(regs[401]), .Q(n521) );
  AOI220 U447 ( .A(n70), .B(regs[1006]), .C(n67), .D(regs[942]), .Q(n452) );
  AOI220 U448 ( .A(n109), .B(regs[710]), .C(n841), .D(regs[646]), .Q(n285) );
  AOI220 U449 ( .A(n70), .B(regs[1010]), .C(n67), .D(regs[946]), .Q(n540) );
  AOI220 U450 ( .A(n70), .B(regs[493]), .C(n67), .D(regs[429]), .Q(n434) );
  AOI220 U451 ( .A(n111), .B(regs[321]), .C(n110), .D(regs[257]), .Q(n167) );
  AOI220 U452 ( .A(regs[987]), .B(n113), .C(regs[923]), .D(n73), .Q(n1459) );
  AOI220 U453 ( .A(regs[887]), .B(n69), .C(regs[823]), .D(n72), .Q(n1370) );
  AOI220 U454 ( .A(regs[233]), .B(n112), .C(regs[169]), .D(n74), .Q(n1078) );
  AOI220 U455 ( .A(regs[216]), .B(n113), .C(regs[152]), .D(n73), .Q(n1407) );
  AOI220 U456 ( .A(regs[375]), .B(n69), .C(regs[311]), .D(n72), .Q(n1374) );
  AOI220 U457 ( .A(regs[103]), .B(n69), .C(regs[39]), .D(n72), .Q(n1032) );
  AOI220 U458 ( .A(regs[471]), .B(n113), .C(regs[407]), .D(n73), .Q(n1375) );
  AOI220 U459 ( .A(regs[231]), .B(n112), .C(regs[167]), .D(n74), .Q(n1034) );
  AOI220 U460 ( .A(regs[199]), .B(n113), .C(regs[135]), .D(n73), .Q(n1033) );
  AOI220 U461 ( .A(regs[744]), .B(n112), .C(regs[680]), .D(n74), .Q(n1052) );
  AOI220 U462 ( .A(regs[121]), .B(n69), .C(regs[57]), .D(n72), .Q(n1428) );
  AOI220 U463 ( .A(regs[576]), .B(n111), .C(regs[512]), .D(n110), .Q(n151) );
  AOI220 U464 ( .A(regs[634]), .B(n69), .C(regs[570]), .D(n72), .Q(n1446) );
  AOI220 U465 ( .A(regs[1014]), .B(n112), .C(regs[950]), .D(n74), .Q(n1350) );
  AOI220 U466 ( .A(regs[120]), .B(n69), .C(regs[56]), .D(n72), .Q(n1406) );
  AOI220 U467 ( .A(regs[217]), .B(n1564), .C(regs[153]), .D(n73), .Q(n1429) );
  AOI220 U468 ( .A(regs[125]), .B(n69), .C(regs[61]), .D(n72), .Q(n1516) );
  AOI220 U469 ( .A(regs[381]), .B(n69), .C(regs[317]), .D(n72), .Q(n1506) );
  AOI220 U470 ( .A(regs[248]), .B(n112), .C(regs[184]), .D(n74), .Q(n1408) );
  AOI220 U471 ( .A(regs[122]), .B(n69), .C(regs[58]), .D(n72), .Q(n1450) );
  AOI220 U472 ( .A(regs[759]), .B(n112), .C(regs[695]), .D(n74), .Q(n1382) );
  AOI220 U473 ( .A(regs[379]), .B(n69), .C(regs[315]), .D(n72), .Q(n1462) );
  AOI220 U474 ( .A(regs[986]), .B(n1564), .C(regs[922]), .D(n73), .Q(n1437) );
  AOI220 U475 ( .A(regs[455]), .B(n113), .C(regs[391]), .D(n73), .Q(n1023) );
  AOI220 U476 ( .A(n111), .B(regs[64]), .C(n110), .D(regs[0]), .Q(n155) );
  AOI220 U477 ( .A(regs[968]), .B(n113), .C(regs[904]), .D(n73), .Q(n1041) );
  AOI220 U478 ( .A(regs[456]), .B(n113), .C(regs[392]), .D(n73), .Q(n1045) );
  AOI220 U479 ( .A(regs[633]), .B(n69), .C(regs[569]), .D(n72), .Q(n1424) );
  AOI220 U480 ( .A(regs[1018]), .B(n112), .C(regs[954]), .D(n74), .Q(n1438) );
  AOI220 U481 ( .A(regs[487]), .B(n1562), .C(regs[423]), .D(n74), .Q(n1024) );
  AOI220 U482 ( .A(regs[764]), .B(n112), .C(regs[700]), .D(n74), .Q(n1492) );
  AOI220 U483 ( .A(regs[631]), .B(n69), .C(regs[567]), .D(n72), .Q(n1380) );
  AOI220 U484 ( .A(n111), .B(regs[832]), .C(n110), .D(regs[768]), .Q(n139) );
  AOI220 U485 ( .A(regs[967]), .B(n113), .C(regs[903]), .D(n73), .Q(n1019) );
  AOI220 U486 ( .A(regs[731]), .B(n113), .C(regs[667]), .D(n73), .Q(n1469) );
  AOI220 U487 ( .A(regs[733]), .B(n113), .C(regs[669]), .D(n73), .Q(n1513) );
  AOI220 U488 ( .A(regs[728]), .B(n113), .C(regs[664]), .D(n73), .Q(n1403) );
  AOI220 U489 ( .A(regs[761]), .B(n112), .C(regs[697]), .D(n74), .Q(n1426) );
  AOI220 U490 ( .A(regs[760]), .B(n112), .C(regs[696]), .D(n74), .Q(n1404) );
  AOI220 U491 ( .A(regs[1017]), .B(n112), .C(regs[953]), .D(n74), .Q(n1416) );
  AOI220 U492 ( .A(regs[635]), .B(n69), .C(regs[571]), .D(n72), .Q(n1468) );
  AOI220 U493 ( .A(n111), .B(regs[320]), .C(n110), .D(regs[256]), .Q(n144) );
  AOI220 U494 ( .A(regs[999]), .B(n1562), .C(regs[935]), .D(n74), .Q(n1020) );
  AOI220 U495 ( .A(regs[377]), .B(n69), .C(regs[313]), .D(n72), .Q(n1418) );
  AOI220 U496 ( .A(regs[889]), .B(n69), .C(regs[825]), .D(n72), .Q(n1414) );
  AOI220 U497 ( .A(regs[124]), .B(n69), .C(regs[60]), .D(n72), .Q(n1494) );
  AOI220 U498 ( .A(n111), .B(regs[65]), .C(n110), .D(regs[1]), .Q(n177) );
  AOI220 U499 ( .A(n111), .B(regs[833]), .C(n110), .D(regs[769]), .Q(n163) );
  AOI220 U500 ( .A(regs[344]), .B(n68), .C(regs[280]), .D(n114), .Q(n1395) );
  AOI220 U501 ( .A(n111), .B(regs[577]), .C(n110), .D(regs[513]), .Q(n173) );
  AOI220 U502 ( .A(regs[215]), .B(n113), .C(regs[151]), .D(n73), .Q(n1385) );
  AOI220 U503 ( .A(regs[488]), .B(n1562), .C(regs[424]), .D(n74), .Q(n1046) );
  AOI220 U504 ( .A(regs[473]), .B(n1564), .C(regs[409]), .D(n73), .Q(n1419) );
  AOI220 U505 ( .A(regs[1020]), .B(n1562), .C(regs[956]), .D(n74), .Q(n1482)
         );
  AOI220 U506 ( .A(n111), .B(regs[66]), .C(n110), .D(regs[2]), .Q(n199) );
  AOI220 U507 ( .A(n846), .B(regs[578]), .C(n110), .D(regs[514]), .Q(n195) );
  AOI220 U508 ( .A(regs[247]), .B(n112), .C(regs[183]), .D(n74), .Q(n1386) );
  AOI220 U509 ( .A(n109), .B(regs[204]), .C(n71), .D(regs[140]), .Q(n421) );
  AOI220 U510 ( .A(regs[238]), .B(n112), .C(regs[174]), .D(n74), .Q(n1188) );
  AOI220 U511 ( .A(n111), .B(regs[342]), .C(n110), .D(regs[278]), .Q(n629) );
  AOI220 U512 ( .A(n109), .B(regs[716]), .C(n841), .D(regs[652]), .Q(n417) );
  AOI220 U513 ( .A(n846), .B(regs[598]), .C(n110), .D(regs[534]), .Q(n635) );
  AOI220 U514 ( .A(regs[718]), .B(n1564), .C(regs[654]), .D(n73), .Q(n1183) );
  AOI220 U515 ( .A(regs[750]), .B(n112), .C(regs[686]), .D(n74), .Q(n1184) );
  AOI220 U516 ( .A(n111), .B(regs[86]), .C(n110), .D(regs[22]), .Q(n639) );
  AOI220 U517 ( .A(n846), .B(regs[855]), .C(n110), .D(regs[791]), .Q(n647) );
  AOI220 U518 ( .A(n111), .B(regs[343]), .C(n110), .D(regs[279]), .Q(n651) );
  AOI220 U519 ( .A(n846), .B(regs[599]), .C(n110), .D(regs[535]), .Q(n657) );
  AOI220 U520 ( .A(n111), .B(regs[87]), .C(n110), .D(regs[23]), .Q(n661) );
  AOI220 U521 ( .A(regs[747]), .B(n112), .C(regs[683]), .D(n74), .Q(n1118) );
  AOI220 U522 ( .A(n846), .B(regs[856]), .C(n110), .D(regs[792]), .Q(n669) );
  AOI220 U523 ( .A(regs[715]), .B(n113), .C(regs[651]), .D(n73), .Q(n1117) );
  AOI220 U524 ( .A(regs[1006]), .B(n112), .C(regs[942]), .D(n74), .Q(n1174) );
  AOI220 U525 ( .A(regs[235]), .B(n112), .C(regs[171]), .D(n74), .Q(n1122) );
  AOI220 U526 ( .A(regs[203]), .B(n113), .C(regs[139]), .D(n73), .Q(n1121) );
  AOI220 U527 ( .A(regs[207]), .B(n113), .C(regs[143]), .D(n73), .Q(n1209) );
  AOI220 U528 ( .A(regs[239]), .B(n112), .C(regs[175]), .D(n74), .Q(n1210) );
  AOI220 U529 ( .A(regs[751]), .B(n1562), .C(regs[687]), .D(n74), .Q(n1206) );
  AOI220 U530 ( .A(regs[1002]), .B(n112), .C(regs[938]), .D(n74), .Q(n1086) );
  AOI220 U531 ( .A(n109), .B(regs[973]), .C(n71), .D(regs[909]), .Q(n429) );
  AOI220 U532 ( .A(n109), .B(regs[721]), .C(n841), .D(regs[657]), .Q(n527) );
  AOI220 U533 ( .A(n109), .B(regs[208]), .C(n71), .D(regs[144]), .Q(n509) );
  AOI220 U534 ( .A(n109), .B(regs[209]), .C(n71), .D(regs[145]), .Q(n531) );
  AOI220 U535 ( .A(n109), .B(regs[720]), .C(n841), .D(regs[656]), .Q(n505) );
  AOI220 U536 ( .A(n111), .B(regs[338]), .C(n110), .D(regs[274]), .Q(n541) );
  AOI220 U537 ( .A(n846), .B(regs[594]), .C(n110), .D(regs[530]), .Q(n547) );
  AOI220 U538 ( .A(n109), .B(regs[976]), .C(n71), .D(regs[912]), .Q(n495) );
  AOI220 U539 ( .A(n111), .B(regs[82]), .C(n110), .D(regs[18]), .Q(n551) );
  AOI220 U540 ( .A(n109), .B(regs[207]), .C(n71), .D(regs[143]), .Q(n487) );
  AOI220 U541 ( .A(regs[364]), .B(n69), .C(regs[300]), .D(n72), .Q(n1132) );
  AOI220 U542 ( .A(n111), .B(regs[851]), .C(n110), .D(regs[787]), .Q(n559) );
  AOI220 U543 ( .A(n109), .B(regs[719]), .C(n841), .D(regs[655]), .Q(n483) );
  AOI220 U544 ( .A(n111), .B(regs[339]), .C(n110), .D(regs[275]), .Q(n563) );
  AOI220 U545 ( .A(n109), .B(regs[463]), .C(n71), .D(regs[399]), .Q(n477) );
  AOI220 U546 ( .A(n111), .B(regs[595]), .C(n110), .D(regs[531]), .Q(n569) );
  AOI220 U547 ( .A(regs[748]), .B(n112), .C(regs[684]), .D(n74), .Q(n1140) );
  AOI220 U548 ( .A(n109), .B(regs[975]), .C(n71), .D(regs[911]), .Q(n473) );
  AOI220 U549 ( .A(n111), .B(regs[83]), .C(n110), .D(regs[19]), .Q(n573) );
  AOI220 U550 ( .A(n109), .B(regs[206]), .C(n71), .D(regs[142]), .Q(n465) );
  AOI220 U551 ( .A(n111), .B(regs[852]), .C(n110), .D(regs[788]), .Q(n581) );
  AOI220 U552 ( .A(n109), .B(regs[718]), .C(n841), .D(regs[654]), .Q(n461) );
  AOI220 U553 ( .A(n109), .B(regs[462]), .C(n71), .D(regs[398]), .Q(n455) );
  AOI220 U554 ( .A(regs[1005]), .B(n112), .C(regs[941]), .D(n74), .Q(n1152) );
  AOI220 U555 ( .A(n111), .B(regs[596]), .C(n110), .D(regs[532]), .Q(n591) );
  AOI220 U556 ( .A(n109), .B(regs[974]), .C(n71), .D(regs[910]), .Q(n451) );
  AOI220 U557 ( .A(n109), .B(regs[205]), .C(n71), .D(regs[141]), .Q(n443) );
  AOI220 U558 ( .A(n109), .B(regs[717]), .C(n841), .D(regs[653]), .Q(n439) );
  AOI220 U559 ( .A(n109), .B(regs[461]), .C(n71), .D(regs[397]), .Q(n433) );
  AOI220 U560 ( .A(n111), .B(regs[597]), .C(n110), .D(regs[533]), .Q(n613) );
  AOI220 U561 ( .A(regs[722]), .B(n113), .C(regs[658]), .D(n73), .Q(n1271) );
  AOI220 U562 ( .A(regs[969]), .B(n113), .C(regs[905]), .D(n73), .Q(n1063) );
  AOI220 U563 ( .A(n111), .B(regs[580]), .C(n110), .D(regs[516]), .Q(n239) );
  AOI220 U564 ( .A(n111), .B(regs[324]), .C(n110), .D(regs[260]), .Q(n233) );
  AOI220 U565 ( .A(regs[115]), .B(n69), .C(regs[51]), .D(n72), .Q(n1296) );
  AOI220 U566 ( .A(regs[211]), .B(n113), .C(regs[147]), .D(n73), .Q(n1297) );
  AOI220 U567 ( .A(regs[243]), .B(n112), .C(regs[179]), .D(n74), .Q(n1298) );
  AOI220 U568 ( .A(n111), .B(regs[836]), .C(n110), .D(regs[772]), .Q(n229) );
  AOI220 U569 ( .A(regs[499]), .B(n112), .C(regs[435]), .D(n74), .Q(n1288) );
  AOI220 U570 ( .A(regs[489]), .B(n112), .C(regs[425]), .D(n74), .Q(n1068) );
  AOI220 U571 ( .A(regs[963]), .B(n113), .C(regs[899]), .D(n73), .Q(n931) );
  AOI220 U572 ( .A(regs[457]), .B(n113), .C(regs[393]), .D(n73), .Q(n1067) );
  AOI220 U573 ( .A(n111), .B(regs[67]), .C(n110), .D(regs[3]), .Q(n221) );
  AOI220 U574 ( .A(n111), .B(regs[579]), .C(n110), .D(regs[515]), .Q(n217) );
  AOI220 U575 ( .A(regs[212]), .B(n113), .C(regs[148]), .D(n73), .Q(n1319) );
  AOI220 U576 ( .A(regs[707]), .B(n113), .C(regs[643]), .D(n73), .Q(n941) );
  AOI220 U577 ( .A(regs[756]), .B(n112), .C(regs[692]), .D(n74), .Q(n1316) );
  AOI220 U578 ( .A(regs[884]), .B(n69), .C(regs[820]), .D(n72), .Q(n1304) );
  AOI220 U579 ( .A(regs[980]), .B(n113), .C(regs[916]), .D(n73), .Q(n1305) );
  AOI220 U580 ( .A(regs[1012]), .B(n112), .C(regs[948]), .D(n74), .Q(n1306) );
  AOI220 U581 ( .A(regs[213]), .B(n113), .C(regs[149]), .D(n73), .Q(n1341) );
  AOI220 U582 ( .A(regs[245]), .B(n112), .C(regs[181]), .D(n74), .Q(n1342) );
  AOI220 U583 ( .A(regs[639]), .B(n69), .C(regs[575]), .D(n72), .Q(n1558) );
  AOI220 U584 ( .A(n111), .B(regs[323]), .C(n110), .D(regs[259]), .Q(n211) );
  AOI220 U585 ( .A(regs[757]), .B(n112), .C(regs[693]), .D(n74), .Q(n1338) );
  AOI220 U586 ( .A(regs[745]), .B(n112), .C(regs[681]), .D(n74), .Q(n1074) );
  AOI220 U587 ( .A(regs[127]), .B(n69), .C(regs[63]), .D(n72), .Q(n1570) );
  AOI220 U588 ( .A(regs[501]), .B(n112), .C(regs[437]), .D(n74), .Q(n1332) );
  AOI220 U589 ( .A(regs[197]), .B(n113), .C(regs[133]), .D(n73), .Q(n989) );
  AOI220 U590 ( .A(regs[1013]), .B(n112), .C(regs[949]), .D(n74), .Q(n1328) );
  AOI220 U591 ( .A(regs[709]), .B(n113), .C(regs[645]), .D(n73), .Q(n985) );
  AOI220 U592 ( .A(regs[198]), .B(n113), .C(regs[134]), .D(n73), .Q(n1011) );
  AOI220 U593 ( .A(regs[710]), .B(n113), .C(regs[646]), .D(n73), .Q(n1007) );
  AOI220 U594 ( .A(regs[118]), .B(n69), .C(regs[54]), .D(n72), .Q(n1362) );
  AOI220 U595 ( .A(regs[214]), .B(n113), .C(regs[150]), .D(n73), .Q(n1363) );
  AOI220 U596 ( .A(n846), .B(regs[835]), .C(n110), .D(regs[771]), .Q(n207) );
  AOI220 U597 ( .A(regs[713]), .B(n113), .C(regs[649]), .D(n73), .Q(n1073) );
  AOI220 U598 ( .A(regs[758]), .B(n112), .C(regs[694]), .D(n74), .Q(n1360) );
  AOI220 U599 ( .A(regs[254]), .B(n112), .C(regs[190]), .D(n74), .Q(n1540) );
  AOI220 U600 ( .A(regs[126]), .B(n69), .C(regs[62]), .D(n72), .Q(n1538) );
  AOI220 U601 ( .A(regs[970]), .B(n113), .C(regs[906]), .D(n73), .Q(n1085) );
  AOI220 U602 ( .A(regs[448]), .B(n113), .C(regs[384]), .D(n73), .Q(n868) );
  AOI220 U603 ( .A(regs[879]), .B(n69), .C(regs[815]), .D(n72), .Q(n1194) );
  AOI220 U604 ( .A(regs[458]), .B(n113), .C(regs[394]), .D(n73), .Q(n1089) );
  AOI220 U605 ( .A(regs[208]), .B(n113), .C(regs[144]), .D(n73), .Q(n1231) );
  AOI220 U606 ( .A(regs[746]), .B(n112), .C(regs[682]), .D(n74), .Q(n1096) );
  AOI220 U607 ( .A(regs[714]), .B(n1564), .C(regs[650]), .D(n73), .Q(n1095) );
  AOI220 U608 ( .A(regs[720]), .B(n113), .C(regs[656]), .D(n73), .Q(n1227) );
  AOI220 U609 ( .A(n111), .B(regs[350]), .C(n110), .D(regs[286]), .Q(n805) );
  AOI220 U610 ( .A(n111), .B(regs[326]), .C(n110), .D(regs[262]), .Q(n277) );
  AOI220 U611 ( .A(n111), .B(regs[606]), .C(n110), .D(regs[542]), .Q(n811) );
  AOI220 U612 ( .A(n111), .B(regs[863]), .C(n110), .D(regs[799]), .Q(n823) );
  AOI220 U613 ( .A(n109), .B(regs[223]), .C(n71), .D(regs[159]), .Q(n849) );
  AOI220 U614 ( .A(n111), .B(regs[325]), .C(n110), .D(regs[261]), .Q(n255) );
  AOI220 U615 ( .A(regs[992]), .B(n112), .C(regs[928]), .D(n74), .Q(n864) );
  AOI220 U616 ( .A(regs[209]), .B(n113), .C(regs[145]), .D(n73), .Q(n1253) );
  AOI220 U617 ( .A(regs[241]), .B(n112), .C(regs[177]), .D(n74), .Q(n1254) );
  AOI220 U618 ( .A(regs[625]), .B(n69), .C(regs[561]), .D(n72), .Q(n1248) );
  AOI220 U619 ( .A(regs[721]), .B(n113), .C(regs[657]), .D(n73), .Q(n1249) );
  AOI220 U620 ( .A(regs[753]), .B(n112), .C(regs[689]), .D(n74), .Q(n1250) );
  AOI220 U621 ( .A(regs[481]), .B(n1562), .C(regs[417]), .D(n74), .Q(n892) );
  AOI220 U622 ( .A(regs[881]), .B(n69), .C(regs[817]), .D(n72), .Q(n1238) );
  AOI220 U623 ( .A(regs[977]), .B(n113), .C(regs[913]), .D(n73), .Q(n1239) );
  AOI220 U624 ( .A(regs[704]), .B(n113), .C(regs[640]), .D(n73), .Q(n875) );
  AOI220 U625 ( .A(regs[736]), .B(n112), .C(regs[672]), .D(n74), .Q(n876) );
  AOI220 U626 ( .A(regs[343]), .B(n68), .C(regs[279]), .D(n114), .Q(n1373) );
  AOI220 U627 ( .A(regs[855]), .B(n68), .C(regs[791]), .D(n114), .Q(n1369) );
  AOI220 U628 ( .A(regs[841]), .B(n68), .C(regs[777]), .D(n114), .Q(n1061) );
  AOI220 U629 ( .A(regs[599]), .B(n68), .C(regs[535]), .D(n114), .Q(n1379) );
  AOI220 U630 ( .A(regs[858]), .B(n68), .C(regs[794]), .D(n114), .Q(n1435) );
  AOI220 U631 ( .A(regs[840]), .B(n68), .C(regs[776]), .D(n114), .Q(n1039) );
  AOI220 U632 ( .A(regs[329]), .B(n68), .C(regs[265]), .D(n114), .Q(n1065) );
  AOI220 U633 ( .A(regs[873]), .B(n69), .C(regs[809]), .D(n72), .Q(n1062) );
  AOI220 U634 ( .A(regs[88]), .B(n68), .C(regs[24]), .D(n114), .Q(n1405) );
  AOI220 U635 ( .A(regs[877]), .B(n1566), .C(regs[813]), .D(n72), .Q(n1150) );
  AOI220 U636 ( .A(regs[600]), .B(n68), .C(regs[536]), .D(n114), .Q(n1401) );
  AOI220 U637 ( .A(regs[624]), .B(n69), .C(regs[560]), .D(n72), .Q(n1226) );
  AOI220 U638 ( .A(regs[872]), .B(n1566), .C(regs[808]), .D(n72), .Q(n1040) );
  AOI220 U639 ( .A(regs[843]), .B(n68), .C(regs[779]), .D(n114), .Q(n1105) );
  AOI220 U640 ( .A(regs[585]), .B(n68), .C(regs[521]), .D(n114), .Q(n1071) );
  AOI220 U641 ( .A(regs[856]), .B(n68), .C(regs[792]), .D(n114), .Q(n1391) );
  AOI220 U642 ( .A(regs[875]), .B(n1566), .C(regs[811]), .D(n72), .Q(n1106) );
  AOI220 U643 ( .A(regs[857]), .B(n68), .C(regs[793]), .D(n114), .Q(n1413) );
  AOI220 U644 ( .A(regs[365]), .B(n69), .C(regs[301]), .D(n72), .Q(n1154) );
  AOI220 U645 ( .A(regs[105]), .B(n69), .C(regs[41]), .D(n72), .Q(n1076) );
  AOI220 U646 ( .A(regs[345]), .B(n68), .C(regs[281]), .D(n114), .Q(n1417) );
  AOI220 U647 ( .A(regs[73]), .B(n68), .C(regs[9]), .D(n114), .Q(n1075) );
  AOI220 U648 ( .A(regs[89]), .B(n68), .C(regs[25]), .D(n114), .Q(n1427) );
  AOI220 U649 ( .A(regs[601]), .B(n68), .C(regs[537]), .D(n114), .Q(n1423) );
  AOI220 U650 ( .A(regs[627]), .B(n69), .C(regs[563]), .D(n72), .Q(n1292) );
  AOI220 U651 ( .A(regs[867]), .B(n69), .C(regs[803]), .D(n72), .Q(n930) );
  AOI220 U652 ( .A(regs[610]), .B(n69), .C(regs[546]), .D(n72), .Q(n918) );
  AOI220 U653 ( .A(regs[844]), .B(n68), .C(regs[780]), .D(n114), .Q(n1127) );
  AOI220 U654 ( .A(regs[111]), .B(n69), .C(regs[47]), .D(n72), .Q(n1208) );
  AOI220 U655 ( .A(regs[623]), .B(n69), .C(regs[559]), .D(n72), .Q(n1204) );
  AOI220 U656 ( .A(regs[842]), .B(n68), .C(regs[778]), .D(n114), .Q(n1083) );
  AOI220 U657 ( .A(regs[876]), .B(n1566), .C(regs[812]), .D(n72), .Q(n1128) );
  AOI220 U658 ( .A(regs[354]), .B(n69), .C(regs[290]), .D(n72), .Q(n912) );
  AOI220 U659 ( .A(regs[372]), .B(n69), .C(regs[308]), .D(n72), .Q(n1308) );
  AOI220 U660 ( .A(regs[75]), .B(n68), .C(regs[11]), .D(n114), .Q(n1119) );
  AOI220 U661 ( .A(regs[834]), .B(n68), .C(regs[770]), .D(n114), .Q(n907) );
  AOI220 U662 ( .A(regs[107]), .B(n1566), .C(regs[43]), .D(n72), .Q(n1120) );
  AOI220 U663 ( .A(regs[330]), .B(n68), .C(regs[266]), .D(n114), .Q(n1087) );
  AOI220 U664 ( .A(regs[629]), .B(n69), .C(regs[565]), .D(n72), .Q(n1336) );
  AOI220 U665 ( .A(regs[98]), .B(n69), .C(regs[34]), .D(n72), .Q(n922) );
  AOI220 U666 ( .A(regs[586]), .B(n68), .C(regs[522]), .D(n114), .Q(n1093) );
  AOI220 U667 ( .A(regs[626]), .B(n69), .C(regs[562]), .D(n72), .Q(n1270) );
  AOI220 U668 ( .A(regs[587]), .B(n68), .C(regs[523]), .D(n114), .Q(n1115) );
  AOI220 U669 ( .A(regs[885]), .B(n69), .C(regs[821]), .D(n72), .Q(n1326) );
  AOI220 U670 ( .A(regs[86]), .B(n68), .C(regs[22]), .D(n114), .Q(n1361) );
  AOI220 U671 ( .A(regs[619]), .B(n1566), .C(regs[555]), .D(n72), .Q(n1116) );
  AOI220 U672 ( .A(regs[106]), .B(n1566), .C(regs[42]), .D(n72), .Q(n1098) );
  AOI220 U673 ( .A(regs[74]), .B(n68), .C(regs[10]), .D(n114), .Q(n1097) );
  AOI220 U674 ( .A(regs[630]), .B(n1566), .C(regs[566]), .D(n72), .Q(n1358) );
  AOI220 U675 ( .A(regs[886]), .B(n1566), .C(regs[822]), .D(n72), .Q(n1348) );
  AOI220 U676 ( .A(regs[366]), .B(n69), .C(regs[302]), .D(n72), .Q(n1176) );
  AOI220 U677 ( .A(regs[331]), .B(n68), .C(regs[267]), .D(n114), .Q(n1109) );
  AOI220 U678 ( .A(regs[87]), .B(n68), .C(regs[23]), .D(n114), .Q(n1383) );
  AOI220 U679 ( .A(regs[321]), .B(n68), .C(regs[257]), .D(n114), .Q(n889) );
  AOI220 U680 ( .A(regs[869]), .B(n69), .C(regs[805]), .D(n72), .Q(n974) );
  AOI220 U681 ( .A(regs[616]), .B(n69), .C(regs[552]), .D(n72), .Q(n1050) );
  AOI220 U682 ( .A(regs[100]), .B(n69), .C(regs[36]), .D(n72), .Q(n966) );
  AOI220 U683 ( .A(regs[584]), .B(n68), .C(regs[520]), .D(n114), .Q(n1049) );
  AOI220 U684 ( .A(regs[837]), .B(n68), .C(regs[773]), .D(n114), .Q(n973) );
  AOI220 U685 ( .A(regs[609]), .B(n69), .C(regs[545]), .D(n72), .Q(n896) );
  AOI220 U686 ( .A(regs[104]), .B(n69), .C(regs[40]), .D(n72), .Q(n1054) );
  AOI220 U687 ( .A(regs[72]), .B(n68), .C(regs[8]), .D(n114), .Q(n1053) );
  AOI220 U688 ( .A(regs[357]), .B(n1566), .C(regs[293]), .D(n72), .Q(n978) );
  AOI220 U689 ( .A(regs[97]), .B(n69), .C(regs[33]), .D(n72), .Q(n900) );
  AOI220 U690 ( .A(regs[64]), .B(n68), .C(regs[0]), .D(n114), .Q(n877) );
  AOI220 U691 ( .A(regs[612]), .B(n69), .C(regs[548]), .D(n72), .Q(n962) );
  AOI220 U692 ( .A(regs[320]), .B(n68), .C(regs[256]), .D(n114), .Q(n866) );
  AOI220 U693 ( .A(regs[839]), .B(n68), .C(regs[775]), .D(n114), .Q(n1017) );
  AOI220 U694 ( .A(regs[832]), .B(n68), .C(regs[768]), .D(n114), .Q(n861) );
  AOI220 U695 ( .A(regs[613]), .B(n69), .C(regs[549]), .D(n72), .Q(n984) );
  AOI220 U696 ( .A(regs[359]), .B(n69), .C(regs[295]), .D(n72), .Q(n1022) );
  AOI220 U697 ( .A(regs[327]), .B(n68), .C(regs[263]), .D(n114), .Q(n1021) );
  AOI220 U698 ( .A(regs[71]), .B(n68), .C(regs[7]), .D(n114), .Q(n1031) );
  AOI220 U699 ( .A(regs[101]), .B(n1566), .C(regs[37]), .D(n72), .Q(n988) );
  AOI220 U700 ( .A(regs[608]), .B(n69), .C(regs[544]), .D(n72), .Q(n874) );
  AOI220 U701 ( .A(regs[836]), .B(n68), .C(regs[772]), .D(n114), .Q(n951) );
  AOI220 U702 ( .A(regs[868]), .B(n69), .C(regs[804]), .D(n72), .Q(n952) );
  AOI220 U703 ( .A(regs[583]), .B(n68), .C(regs[519]), .D(n114), .Q(n1027) );
  AOI220 U704 ( .A(regs[102]), .B(n1566), .C(regs[38]), .D(n72), .Q(n1010) );
  AOI220 U705 ( .A(regs[328]), .B(n68), .C(regs[264]), .D(n114), .Q(n1043) );
  AOI220 U706 ( .A(regs[614]), .B(n1566), .C(regs[550]), .D(n72), .Q(n1006) );
  NAND22 U707 ( .A(n1580), .B(i_addr_Rd[3]), .Q(n1591) );
  NOR22 U708 ( .A(i_addr_Rt_3_), .B(n150), .Q(n854) );
  NOR22 U709 ( .A(i_addr_Rs[2]), .B(n858), .Q(n1566) );
  NOR31 U710 ( .A(i_addr_Rs[0]), .B(n860), .C(n857), .Q(n1564) );
  NOR22 U711 ( .A(n865), .B(n872), .Q(n1556) );
  NAND31 U712 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n108), .Q(n1588) );
  NOR31 U713 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .C(i_addr_Rt_2_), .Q(n845)
         );
  NAND31 U714 ( .A(n108), .B(n1586), .C(n1585), .Q(n1584) );
  NOR22 U715 ( .A(i_addr_Rs[3]), .B(n872), .Q(n1576) );
  NAND31 U716 ( .A(i_addr_Rd[1]), .B(n108), .C(n1586), .Q(n1589) );
  NOR21 U717 ( .A(i_addr_Rd[4]), .B(n1579), .Q(n1580) );
  NAND31 U718 ( .A(i_addr_Rd[0]), .B(n108), .C(n1585), .Q(n1590) );
  INV3 U719 ( .A(i_addr_Rs[4]), .Q(n872) );
  INV2 U720 ( .A(i_addr_Rs[0]), .Q(n859) );
  INV3 U721 ( .A(i_addr_Rs[2]), .Q(n857) );
  NOR31 U722 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[1]), .C(i_addr_Rs[2]), .Q(n1567)
         );
  INV3 U723 ( .A(i_addr_Rt_2_), .Q(n135) );
  INV2 U724 ( .A(i_addr_Rs[1]), .Q(n860) );
  INV3 U725 ( .A(i_addr_Rs[3]), .Q(n865) );
  INV3 U726 ( .A(i_addr_Rt_3_), .Q(n143) );
  INV2 U727 ( .A(i_con_RegWr), .Q(n1579) );
  INV3 U728 ( .A(i_addr_Rt_4_), .Q(n150) );
  NOR32 U729 ( .A(i_addr_Rt_1_), .B(i_addr_Rt_2_), .C(n137), .Q(n843) );
  NAND31 U730 ( .A(i_con_RegWr), .B(i_addr_Rd[4]), .C(n1583), .Q(n1587) );
  INV3 U731 ( .A(i_addr_Rd[3]), .Q(n1583) );
  NAND31 U732 ( .A(i_addr_Rd[4]), .B(i_con_RegWr), .C(i_addr_Rd[3]), .Q(n1582)
         );
  INV3 U733 ( .A(i_addr_Rd[0]), .Q(n1586) );
  INV3 U734 ( .A(i_addr_Rd[1]), .Q(n1585) );
  NOR21 U735 ( .A(i_addr_Rt_2_), .B(n136), .Q(n844) );
  NOR31 U736 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_2_), .C(n138), .Q(n846) );
  AOI220 U737 ( .A(n111), .B(regs[91]), .C(n110), .D(regs[27]), .Q(n749) );
  AOI220 U738 ( .A(n111), .B(regs[603]), .C(n110), .D(regs[539]), .Q(n745) );
  AOI220 U739 ( .A(n111), .B(regs[347]), .C(n110), .D(regs[283]), .Q(n739) );
  AOI220 U740 ( .A(n111), .B(regs[859]), .C(n110), .D(regs[795]), .Q(n735) );
  AOI220 U741 ( .A(n109), .B(regs[729]), .C(n841), .D(regs[665]), .Q(n703) );
  AOI220 U742 ( .A(n109), .B(regs[473]), .C(n841), .D(regs[409]), .Q(n697) );
  AOI220 U743 ( .A(n842), .B(regs[213]), .C(n71), .D(regs[149]), .Q(n619) );
  AOI220 U744 ( .A(n842), .B(regs[469]), .C(n71), .D(regs[405]), .Q(n609) );
  AOI220 U745 ( .A(n70), .B(regs[501]), .C(n839), .D(regs[437]), .Q(n610) );
  AOI220 U746 ( .A(n70), .B(regs[244]), .C(n839), .D(regs[180]), .Q(n598) );
  AOI220 U747 ( .A(n842), .B(regs[468]), .C(n71), .D(regs[404]), .Q(n587) );
  AOI220 U748 ( .A(n70), .B(regs[500]), .C(n839), .D(regs[436]), .Q(n588) );
  AOI220 U749 ( .A(n109), .B(regs[728]), .C(n841), .D(regs[664]), .Q(n681) );
  AOI220 U750 ( .A(n111), .B(regs[862]), .C(n110), .D(regs[798]), .Q(n801) );
  AOI220 U751 ( .A(n111), .B(regs[95]), .C(n110), .D(regs[31]), .Q(n847) );
  AOI220 U752 ( .A(n111), .B(regs[93]), .C(n110), .D(regs[29]), .Q(n793) );
  AOI220 U753 ( .A(n111), .B(regs[605]), .C(n110), .D(regs[541]), .Q(n789) );
  AOI220 U754 ( .A(n111), .B(regs[349]), .C(n110), .D(regs[285]), .Q(n783) );
  AOI220 U755 ( .A(n111), .B(regs[861]), .C(n110), .D(regs[797]), .Q(n779) );
  AOI220 U756 ( .A(n111), .B(regs[92]), .C(n110), .D(regs[28]), .Q(n771) );
  AOI220 U757 ( .A(n111), .B(regs[604]), .C(n110), .D(regs[540]), .Q(n767) );
  AOI220 U758 ( .A(n111), .B(regs[348]), .C(n110), .D(regs[284]), .Q(n761) );
  AOI220 U759 ( .A(n111), .B(regs[860]), .C(n110), .D(regs[796]), .Q(n757) );
  AOI220 U760 ( .A(n111), .B(regs[90]), .C(n110), .D(regs[26]), .Q(n727) );
  AOI220 U761 ( .A(n111), .B(regs[602]), .C(n110), .D(regs[538]), .Q(n723) );
  AOI220 U762 ( .A(n111), .B(regs[346]), .C(n110), .D(regs[282]), .Q(n717) );
  AOI220 U763 ( .A(n70), .B(regs[506]), .C(n839), .D(regs[442]), .Q(n720) );
  AOI220 U764 ( .A(n842), .B(regs[978]), .C(n841), .D(regs[914]), .Q(n539) );
  AOI220 U765 ( .A(n111), .B(regs[333]), .C(n110), .D(regs[269]), .Q(n431) );
  AOI220 U766 ( .A(n111), .B(regs[76]), .C(n110), .D(regs[12]), .Q(n419) );
  AOI220 U767 ( .A(n846), .B(regs[588]), .C(n110), .D(regs[524]), .Q(n415) );
  AOI220 U768 ( .A(n111), .B(regs[335]), .C(n110), .D(regs[271]), .Q(n475) );
  AOI220 U769 ( .A(n111), .B(regs[847]), .C(n110), .D(regs[783]), .Q(n471) );
  AOI220 U770 ( .A(n111), .B(regs[78]), .C(n110), .D(regs[14]), .Q(n463) );
  AOI220 U771 ( .A(n111), .B(regs[334]), .C(n110), .D(regs[270]), .Q(n453) );
  AOI220 U772 ( .A(n111), .B(regs[846]), .C(n110), .D(regs[782]), .Q(n449) );
  AOI220 U773 ( .A(n111), .B(regs[81]), .C(n110), .D(regs[17]), .Q(n529) );
  AOI220 U774 ( .A(n846), .B(regs[593]), .C(n110), .D(regs[529]), .Q(n525) );
  AOI220 U775 ( .A(n111), .B(regs[337]), .C(n110), .D(regs[273]), .Q(n519) );
  AOI220 U776 ( .A(n842), .B(regs[977]), .C(n841), .D(regs[913]), .Q(n517) );
  AOI220 U777 ( .A(n111), .B(regs[80]), .C(n110), .D(regs[16]), .Q(n507) );
  AOI220 U778 ( .A(n846), .B(regs[592]), .C(n110), .D(regs[528]), .Q(n503) );
  AOI220 U779 ( .A(n111), .B(regs[336]), .C(n110), .D(regs[272]), .Q(n497) );
  AOI220 U780 ( .A(n111), .B(regs[848]), .C(n110), .D(regs[784]), .Q(n493) );
  AOI220 U781 ( .A(n109), .B(regs[964]), .C(n841), .D(regs[900]), .Q(n231) );
  AOI220 U782 ( .A(regs[225]), .B(n112), .C(regs[161]), .D(n74), .Q(n902) );
  AOI220 U783 ( .A(regs[737]), .B(n112), .C(regs[673]), .D(n74), .Q(n898) );
  AOI220 U784 ( .A(regs[739]), .B(n112), .C(regs[675]), .D(n74), .Q(n942) );
  AOI220 U785 ( .A(regs[230]), .B(n112), .C(regs[166]), .D(n74), .Q(n1012) );
  AOI220 U786 ( .A(regs[486]), .B(n112), .C(regs[422]), .D(n74), .Q(n1002) );
  AOI220 U787 ( .A(regs[998]), .B(n112), .C(regs[934]), .D(n74), .Q(n998) );
  AOI220 U788 ( .A(regs[482]), .B(n112), .C(regs[418]), .D(n74), .Q(n914) );
  AOI220 U789 ( .A(regs[994]), .B(n112), .C(regs[930]), .D(n74), .Q(n910) );
  AOI220 U790 ( .A(regs[228]), .B(n112), .C(regs[164]), .D(n74), .Q(n968) );
  AOI220 U791 ( .A(regs[740]), .B(n112), .C(regs[676]), .D(n74), .Q(n964) );
  AOI220 U792 ( .A(regs[484]), .B(n112), .C(regs[420]), .D(n74), .Q(n958) );
  AOI220 U793 ( .A(regs[996]), .B(n112), .C(regs[932]), .D(n74), .Q(n954) );
  AOI220 U794 ( .A(regs[229]), .B(n112), .C(regs[165]), .D(n74), .Q(n990) );
  AOI220 U795 ( .A(regs[741]), .B(n112), .C(regs[677]), .D(n74), .Q(n986) );
  AOI220 U796 ( .A(regs[485]), .B(n112), .C(regs[421]), .D(n74), .Q(n980) );
  AOI220 U797 ( .A(regs[997]), .B(n112), .C(regs[933]), .D(n74), .Q(n976) );
  AOI220 U798 ( .A(regs[252]), .B(n112), .C(regs[188]), .D(n74), .Q(n1496) );
  AOI220 U799 ( .A(regs[255]), .B(n112), .C(regs[191]), .D(n74), .Q(n1572) );
  AOI220 U800 ( .A(regs[767]), .B(n112), .C(regs[703]), .D(n74), .Q(n1560) );
  AOI220 U801 ( .A(regs[511]), .B(n112), .C(regs[447]), .D(n74), .Q(n1552) );
  AOI220 U802 ( .A(regs[495]), .B(n112), .C(regs[431]), .D(n74), .Q(n1200) );
  AOI220 U803 ( .A(regs[1007]), .B(n112), .C(regs[943]), .D(n74), .Q(n1196) );
  AOI220 U804 ( .A(regs[752]), .B(n112), .C(regs[688]), .D(n74), .Q(n1228) );
  AOI220 U805 ( .A(regs[1022]), .B(n112), .C(regs[958]), .D(n74), .Q(n1526) );
  AOI220 U806 ( .A(regs[250]), .B(n112), .C(regs[186]), .D(n74), .Q(n1452) );
  AOI220 U807 ( .A(regs[762]), .B(n112), .C(regs[698]), .D(n74), .Q(n1448) );
  AOI220 U808 ( .A(regs[506]), .B(n112), .C(regs[442]), .D(n74), .Q(n1442) );
  AOI220 U809 ( .A(regs[251]), .B(n112), .C(regs[187]), .D(n74), .Q(n1474) );
  AOI220 U810 ( .A(regs[763]), .B(n112), .C(regs[699]), .D(n74), .Q(n1470) );
  AOI220 U811 ( .A(regs[507]), .B(n112), .C(regs[443]), .D(n74), .Q(n1464) );
  AOI220 U812 ( .A(regs[1019]), .B(n112), .C(regs[955]), .D(n74), .Q(n1460) );
  AOI220 U813 ( .A(regs[500]), .B(n112), .C(regs[436]), .D(n74), .Q(n1310) );
  AOI221 U814 ( .A(n66), .B(regs[887]), .C(n843), .D(regs[823]), .Q(n648) );
  AOI221 U815 ( .A(n66), .B(regs[118]), .C(n75), .D(regs[54]), .Q(n640) );
  AOI221 U816 ( .A(n66), .B(regs[628]), .C(n843), .D(regs[564]), .Q(n592) );
  AOI221 U817 ( .A(n70), .B(regs[251]), .C(n67), .D(regs[187]), .Q(n752) );
  AOI221 U818 ( .A(n70), .B(regs[763]), .C(n67), .D(regs[699]), .Q(n748) );
  AOI221 U819 ( .A(n70), .B(regs[507]), .C(n67), .D(regs[443]), .Q(n742) );
  AOI221 U820 ( .A(n70), .B(regs[1019]), .C(n67), .D(regs[955]), .Q(n738) );
  AOI221 U821 ( .A(n66), .B(regs[115]), .C(n843), .D(regs[51]), .Q(n574) );
  AOI221 U822 ( .A(n66), .B(regs[121]), .C(n843), .D(regs[57]), .Q(n706) );
  AOI221 U823 ( .A(n66), .B(regs[377]), .C(n75), .D(regs[313]), .Q(n696) );
  AOI221 U824 ( .A(n66), .B(regs[374]), .C(n75), .D(regs[310]), .Q(n630) );
  AOI221 U825 ( .A(n66), .B(regs[884]), .C(n75), .D(regs[820]), .Q(n582) );
  AOI221 U826 ( .A(n66), .B(regs[632]), .C(n843), .D(regs[568]), .Q(n680) );
  AOI221 U827 ( .A(n66), .B(regs[888]), .C(n75), .D(regs[824]), .Q(n670) );
  AOI221 U828 ( .A(n66), .B(regs[638]), .C(n843), .D(regs[574]), .Q(n812) );
  AOI221 U829 ( .A(n66), .B(regs[382]), .C(n75), .D(regs[318]), .Q(n806) );
  AOI221 U830 ( .A(n66), .B(regs[637]), .C(n75), .D(regs[573]), .Q(n790) );
  AOI221 U831 ( .A(n66), .B(regs[893]), .C(n75), .D(regs[829]), .Q(n780) );
  AOI221 U832 ( .A(n70), .B(regs[1020]), .C(n67), .D(regs[956]), .Q(n760) );
  AOI221 U833 ( .A(n70), .B(regs[250]), .C(n67), .D(regs[186]), .Q(n730) );
  AOI221 U834 ( .A(n70), .B(regs[762]), .C(n67), .D(regs[698]), .Q(n726) );
  AOI221 U835 ( .A(n66), .B(regs[101]), .C(n75), .D(regs[37]), .Q(n266) );
  AOI221 U836 ( .A(n66), .B(regs[613]), .C(n75), .D(regs[549]), .Q(n262) );
  AOI221 U837 ( .A(n66), .B(regs[357]), .C(n75), .D(regs[293]), .Q(n256) );
  AOI221 U838 ( .A(n66), .B(regs[869]), .C(n75), .D(regs[805]), .Q(n252) );
  AOI221 U839 ( .A(n66), .B(regs[103]), .C(n75), .D(regs[39]), .Q(n310) );
  AOI221 U840 ( .A(n66), .B(regs[615]), .C(n75), .D(regs[551]), .Q(n306) );
  AOI221 U841 ( .A(n66), .B(regs[359]), .C(n75), .D(regs[295]), .Q(n300) );
  AOI221 U842 ( .A(n66), .B(regs[871]), .C(n843), .D(regs[807]), .Q(n296) );
  AOI221 U843 ( .A(n66), .B(regs[875]), .C(n75), .D(regs[811]), .Q(n384) );
  AOI221 U844 ( .A(n66), .B(regs[99]), .C(n75), .D(regs[35]), .Q(n222) );
  AOI221 U845 ( .A(n66), .B(regs[867]), .C(n75), .D(regs[803]), .Q(n208) );
  AOI221 U846 ( .A(n66), .B(regs[97]), .C(n75), .D(regs[33]), .Q(n178) );
  AOI221 U847 ( .A(n66), .B(regs[609]), .C(n75), .D(regs[545]), .Q(n174) );
  AOI221 U848 ( .A(n66), .B(regs[353]), .C(n75), .D(regs[289]), .Q(n168) );
  AOI221 U849 ( .A(n66), .B(regs[865]), .C(n75), .D(regs[801]), .Q(n164) );
  AOI221 U850 ( .A(n66), .B(regs[102]), .C(n843), .D(regs[38]), .Q(n288) );
  AOI221 U851 ( .A(n66), .B(regs[614]), .C(n843), .D(regs[550]), .Q(n284) );
  AOI221 U852 ( .A(n66), .B(regs[358]), .C(n75), .D(regs[294]), .Q(n278) );
  AOI221 U853 ( .A(n66), .B(regs[870]), .C(n75), .D(regs[806]), .Q(n274) );
  AOI221 U854 ( .A(n66), .B(regs[96]), .C(n75), .D(regs[32]), .Q(n156) );
  AOI221 U855 ( .A(n66), .B(regs[352]), .C(n75), .D(regs[288]), .Q(n145) );
  AOI221 U856 ( .A(n66), .B(regs[864]), .C(n843), .D(regs[800]), .Q(n140) );
  AOI221 U857 ( .A(n66), .B(regs[106]), .C(n843), .D(regs[42]), .Q(n376) );
  AOI221 U858 ( .A(n66), .B(regs[618]), .C(n843), .D(regs[554]), .Q(n372) );
  AOI221 U859 ( .A(n66), .B(regs[362]), .C(n75), .D(regs[298]), .Q(n366) );
  AOI221 U860 ( .A(n66), .B(regs[876]), .C(n75), .D(regs[812]), .Q(n406) );
  AOI221 U861 ( .A(n66), .B(regs[105]), .C(n75), .D(regs[41]), .Q(n354) );
  AOI221 U862 ( .A(n66), .B(regs[617]), .C(n75), .D(regs[553]), .Q(n350) );
  AOI221 U863 ( .A(n66), .B(regs[361]), .C(n75), .D(regs[297]), .Q(n344) );
  AOI221 U864 ( .A(n66), .B(regs[873]), .C(n843), .D(regs[809]), .Q(n340) );
  AOI221 U865 ( .A(n66), .B(regs[879]), .C(n75), .D(regs[815]), .Q(n472) );
  AOI221 U866 ( .A(n66), .B(regs[610]), .C(n75), .D(regs[546]), .Q(n196) );
  AOI221 U867 ( .A(n66), .B(regs[354]), .C(n75), .D(regs[290]), .Q(n190) );
  AOI221 U868 ( .A(n66), .B(regs[866]), .C(n75), .D(regs[802]), .Q(n186) );
  AOI221 U869 ( .A(n66), .B(regs[369]), .C(n75), .D(regs[305]), .Q(n520) );
  AOI221 U870 ( .A(n66), .B(regs[881]), .C(n75), .D(regs[817]), .Q(n516) );
  AOI221 U871 ( .A(n66), .B(regs[100]), .C(n75), .D(regs[36]), .Q(n244) );
  AOI221 U872 ( .A(n66), .B(regs[612]), .C(n75), .D(regs[548]), .Q(n240) );
  AOI221 U873 ( .A(n66), .B(regs[104]), .C(n843), .D(regs[40]), .Q(n332) );
  AOI221 U874 ( .A(n66), .B(regs[616]), .C(n843), .D(regs[552]), .Q(n328) );
  AOI221 U875 ( .A(n66), .B(regs[360]), .C(n75), .D(regs[296]), .Q(n322) );
  AOI220 U876 ( .A(regs[70]), .B(n68), .C(regs[6]), .D(n114), .Q(n1009) );
  AOI220 U877 ( .A(regs[582]), .B(n68), .C(regs[518]), .D(n114), .Q(n1005) );
  AOI220 U878 ( .A(regs[581]), .B(n68), .C(regs[517]), .D(n114), .Q(n983) );
  AOI220 U879 ( .A(regs[348]), .B(n68), .C(regs[284]), .D(n114), .Q(n1483) );
  AOI220 U880 ( .A(regs[351]), .B(n68), .C(regs[287]), .D(n114), .Q(n1549) );
  AOI220 U881 ( .A(regs[349]), .B(n68), .C(regs[285]), .D(n114), .Q(n1505) );
  AOI220 U882 ( .A(regs[350]), .B(n68), .C(regs[286]), .D(n114), .Q(n1527) );
  AOI221 U883 ( .A(n66), .B(regs[889]), .C(n75), .D(regs[825]), .Q(n692) );
  AOI221 U884 ( .A(n66), .B(regs[120]), .C(n75), .D(regs[56]), .Q(n684) );
  AOI221 U885 ( .A(n66), .B(regs[127]), .C(n75), .D(regs[63]), .Q(n848) );
  AOI221 U886 ( .A(n66), .B(regs[882]), .C(n843), .D(regs[818]), .Q(n538) );
  AOI221 U887 ( .A(n66), .B(regs[111]), .C(n75), .D(regs[47]), .Q(n486) );
  AOI221 U888 ( .A(n66), .B(regs[623]), .C(n843), .D(regs[559]), .Q(n482) );
  AOI221 U889 ( .A(n66), .B(regs[367]), .C(n75), .D(regs[303]), .Q(n476) );
  AOI221 U890 ( .A(n66), .B(regs[110]), .C(n843), .D(regs[46]), .Q(n464) );
  AOI221 U891 ( .A(n66), .B(regs[622]), .C(n75), .D(regs[558]), .Q(n460) );
  AOI221 U892 ( .A(n66), .B(regs[113]), .C(n75), .D(regs[49]), .Q(n530) );
  AOI221 U893 ( .A(n66), .B(regs[625]), .C(n75), .D(regs[561]), .Q(n526) );
  AOI221 U894 ( .A(n66), .B(regs[112]), .C(n75), .D(regs[48]), .Q(n508) );
  AOI221 U895 ( .A(n66), .B(regs[624]), .C(n843), .D(regs[560]), .Q(n504) );
  AOI221 U896 ( .A(n66), .B(regs[368]), .C(n75), .D(regs[304]), .Q(n498) );
  AOI221 U897 ( .A(n66), .B(regs[880]), .C(n75), .D(regs[816]), .Q(n494) );
  AOI221 U898 ( .A(regs[355]), .B(n69), .C(regs[291]), .D(n72), .Q(n934) );
  AOI221 U899 ( .A(regs[866]), .B(n69), .C(regs[802]), .D(n72), .Q(n908) );
  AOI221 U900 ( .A(regs[360]), .B(n69), .C(regs[296]), .D(n72), .Q(n1044) );
  AOI221 U901 ( .A(regs[622]), .B(n69), .C(regs[558]), .D(n72), .Q(n1182) );
  AOI221 U902 ( .A(regs[112]), .B(n69), .C(regs[48]), .D(n72), .Q(n1230) );
  AOI221 U903 ( .A(regs[880]), .B(n69), .C(regs[816]), .D(n72), .Q(n1216) );
  AOI221 U904 ( .A(regs[109]), .B(n69), .C(regs[45]), .D(n72), .Q(n1164) );
  AOI221 U905 ( .A(regs[637]), .B(n69), .C(regs[573]), .D(n72), .Q(n1512) );
  AOI221 U906 ( .A(regs[638]), .B(n69), .C(regs[574]), .D(n72), .Q(n1534) );
  NOR30 U907 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[2]), .C(n860), .Q(n1568) );
  AOI221 U908 ( .A(n70), .B(regs[247]), .C(n67), .D(regs[183]), .Q(n664) );
  AOI221 U909 ( .A(n70), .B(regs[759]), .C(n67), .D(regs[695]), .Q(n660) );
  AOI221 U910 ( .A(n70), .B(regs[503]), .C(n67), .D(regs[439]), .Q(n654) );
  AOI221 U911 ( .A(n70), .B(regs[1015]), .C(n67), .D(regs[951]), .Q(n650) );
  AOI221 U912 ( .A(n70), .B(regs[243]), .C(n67), .D(regs[179]), .Q(n576) );
  AOI221 U913 ( .A(n70), .B(regs[755]), .C(n67), .D(regs[691]), .Q(n572) );
  AOI221 U914 ( .A(n70), .B(regs[499]), .C(n67), .D(regs[435]), .Q(n566) );
  AOI221 U915 ( .A(n70), .B(regs[1011]), .C(n67), .D(regs[947]), .Q(n562) );
  AOI221 U916 ( .A(n70), .B(regs[246]), .C(n67), .D(regs[182]), .Q(n642) );
  AOI221 U917 ( .A(n70), .B(regs[758]), .C(n67), .D(regs[694]), .Q(n638) );
  AOI221 U918 ( .A(n70), .B(regs[502]), .C(n67), .D(regs[438]), .Q(n632) );
  AOI221 U919 ( .A(n70), .B(regs[1014]), .C(n67), .D(regs[950]), .Q(n628) );
  AOI221 U920 ( .A(n70), .B(regs[756]), .C(n67), .D(regs[692]), .Q(n594) );
  AOI221 U921 ( .A(n70), .B(regs[1012]), .C(n67), .D(regs[948]), .Q(n584) );
  AOI221 U922 ( .A(n70), .B(regs[1016]), .C(n67), .D(regs[952]), .Q(n672) );
  AOI221 U923 ( .A(n70), .B(regs[242]), .C(n67), .D(regs[178]), .Q(n554) );
  AOI221 U924 ( .A(n70), .B(regs[754]), .C(n67), .D(regs[690]), .Q(n550) );
  AOI221 U925 ( .A(n70), .B(regs[498]), .C(n67), .D(regs[434]), .Q(n544) );
  AOI221 U926 ( .A(n111), .B(regs[69]), .C(n110), .D(regs[5]), .Q(n265) );
  AOI221 U927 ( .A(n111), .B(regs[581]), .C(n110), .D(regs[517]), .Q(n261) );
  AOI221 U928 ( .A(n70), .B(regs[237]), .C(n67), .D(regs[173]), .Q(n444) );
  AOI221 U929 ( .A(n70), .B(regs[751]), .C(n67), .D(regs[687]), .Q(n484) );
  AOI221 U930 ( .A(regs[892]), .B(n69), .C(regs[828]), .D(n72), .Q(n1480) );
  AOI221 U931 ( .A(regs[620]), .B(n69), .C(regs[556]), .D(n72), .Q(n1138) );
  AOI221 U932 ( .A(regs[378]), .B(n69), .C(regs[314]), .D(n72), .Q(n1440) );
  AOI221 U933 ( .A(regs[123]), .B(n69), .C(regs[59]), .D(n72), .Q(n1472) );
  AOI221 U934 ( .A(regs[891]), .B(n69), .C(regs[827]), .D(n72), .Q(n1458) );
  AOI221 U935 ( .A(regs[628]), .B(n69), .C(regs[564]), .D(n72), .Q(n1314) );
  BUF2 U936 ( .A(n25), .Q(n125) );
  BUF2 U937 ( .A(n26), .Q(n124) );
  BUF2 U938 ( .A(n23), .Q(n126) );
  BUF2 U939 ( .A(n15), .Q(n133) );
  BUF2 U940 ( .A(n16), .Q(n132) );
  BUF2 U941 ( .A(n13), .Q(n134) );
  BUF2 U942 ( .A(n42), .Q(n117) );
  BUF2 U943 ( .A(n41), .Q(n118) );
  BUF2 U944 ( .A(n43), .Q(n116) );
  BUF2 U945 ( .A(n35), .Q(n120) );
  BUF2 U946 ( .A(n32), .Q(n122) );
  BUF2 U947 ( .A(n34), .Q(n121) );
  BUF2 U948 ( .A(i_addr_Rd[2]), .Q(n108) );
  AOI221 U949 ( .A(n70), .B(regs[757]), .C(n67), .D(regs[693]), .Q(n616) );
  AOI221 U950 ( .A(n70), .B(regs[1013]), .C(n67), .D(regs[949]), .Q(n606) );
  AOI221 U951 ( .A(n70), .B(regs[760]), .C(n67), .D(regs[696]), .Q(n682) );
  AOI221 U952 ( .A(n70), .B(regs[511]), .C(n67), .D(regs[447]), .Q(n830) );
  AOI221 U953 ( .A(n70), .B(regs[1018]), .C(n839), .D(regs[954]), .Q(n716) );
  AOI221 U954 ( .A(n70), .B(regs[229]), .C(n67), .D(regs[165]), .Q(n268) );
  AOI221 U955 ( .A(n70), .B(regs[741]), .C(n67), .D(regs[677]), .Q(n264) );
  AOI221 U956 ( .A(n70), .B(regs[485]), .C(n67), .D(regs[421]), .Q(n258) );
  AOI221 U957 ( .A(n111), .B(regs[837]), .C(n110), .D(regs[773]), .Q(n251) );
  AOI221 U958 ( .A(n70), .B(regs[997]), .C(n67), .D(regs[933]), .Q(n254) );
  AOI221 U959 ( .A(n70), .B(regs[487]), .C(n839), .D(regs[423]), .Q(n302) );
  AOI221 U960 ( .A(n111), .B(regs[839]), .C(n845), .D(regs[775]), .Q(n295) );
  AOI221 U961 ( .A(n70), .B(regs[999]), .C(n839), .D(regs[935]), .Q(n298) );
  AOI221 U962 ( .A(n111), .B(regs[75]), .C(n845), .D(regs[11]), .Q(n397) );
  AOI221 U963 ( .A(n111), .B(regs[843]), .C(n110), .D(regs[779]), .Q(n383) );
  AOI221 U964 ( .A(n70), .B(regs[225]), .C(n67), .D(regs[161]), .Q(n180) );
  AOI221 U965 ( .A(n70), .B(regs[737]), .C(n67), .D(regs[673]), .Q(n176) );
  AOI221 U966 ( .A(n70), .B(regs[481]), .C(n67), .D(regs[417]), .Q(n170) );
  AOI221 U967 ( .A(n70), .B(regs[993]), .C(n67), .D(regs[929]), .Q(n166) );
  AOI221 U968 ( .A(n70), .B(regs[230]), .C(n67), .D(regs[166]), .Q(n290) );
  AOI221 U969 ( .A(n70), .B(regs[486]), .C(n67), .D(regs[422]), .Q(n280) );
  AOI221 U970 ( .A(n111), .B(regs[838]), .C(n110), .D(regs[774]), .Q(n273) );
  AOI221 U971 ( .A(n70), .B(regs[998]), .C(n67), .D(regs[934]), .Q(n276) );
  AOI221 U972 ( .A(n70), .B(regs[480]), .C(n67), .D(regs[416]), .Q(n147) );
  AOI221 U973 ( .A(n111), .B(regs[586]), .C(n110), .D(regs[522]), .Q(n371) );
  AOI221 U974 ( .A(n70), .B(regs[482]), .C(n67), .D(regs[418]), .Q(n192) );
  AOI221 U975 ( .A(n834), .B(n238), .C(n832), .D(n237), .Q(n250) );
  AOI221 U976 ( .A(n70), .B(regs[488]), .C(n67), .D(regs[424]), .Q(n324) );
  NOR31 U977 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .C(n135), .Q(n841) );
  NOR31 U978 ( .A(i_addr_Rt_1_), .B(n137), .C(n135), .Q(n839) );
  NOR21 U979 ( .A(n136), .B(n135), .Q(n840) );
  NOR31 U980 ( .A(i_addr_Rs[1]), .B(n859), .C(n857), .Q(n1561) );
  NOR21 U981 ( .A(n858), .B(n857), .Q(n1562) );
  BUF2 U982 ( .A(n21), .Q(n128) );
  BUF2 U983 ( .A(n20), .Q(n129) );
  BUF2 U984 ( .A(n18), .Q(n130) );
  BUF2 U985 ( .A(n22), .Q(n127) );
  BUF2 U986 ( .A(n27), .Q(n123) );
  BUF2 U987 ( .A(n17), .Q(n131) );
  BUF2 U988 ( .A(n44), .Q(n115) );
  NOR40 U989 ( .A(n108), .B(n1586), .C(n1591), .D(n1585), .Q(n44) );
  AOI221 U990 ( .A(n854), .B(n182), .C(n852), .D(n181), .Q(n183) );
  AOI221 U991 ( .A(n854), .B(n292), .C(n852), .D(n291), .Q(n293) );
  AOI221 U992 ( .A(n854), .B(n446), .C(n852), .D(n445), .Q(n447) );
  AOI221 U993 ( .A(n854), .B(n490), .C(n852), .D(n489), .Q(n491) );
  AOI221 U994 ( .A(n854), .B(n468), .C(n852), .D(n467), .Q(n469) );
  AOI221 U995 ( .A(n854), .B(n204), .C(n852), .D(n203), .Q(n205) );
  AOI221 U996 ( .A(n854), .B(n534), .C(n852), .D(n533), .Q(n535) );
  AOI221 U997 ( .A(n854), .B(n512), .C(n852), .D(n511), .Q(n513) );
  AOI221 U998 ( .A(n854), .B(n248), .C(n852), .D(n247), .Q(n249) );
  AOI221 U999 ( .A(n854), .B(n336), .C(n852), .D(n335), .Q(n337) );
  AOI221 U1000 ( .A(n834), .B(n326), .C(n832), .D(n325), .Q(n338) );
  NOR31 U1001 ( .A(i_addr_Rt_0_), .B(n138), .C(n135), .Q(n842) );
  AOI221 U1002 ( .A(n1576), .B(n992), .C(n1574), .D(n991), .Q(n993) );
  AOI221 U1003 ( .A(n1576), .B(n1036), .C(n1574), .D(n1035), .Q(n1037) );
  AOI221 U1004 ( .A(n1556), .B(n1092), .C(n1554), .D(n1091), .Q(n1104) );
  AOI221 U1005 ( .A(n1576), .B(n1300), .C(n1574), .D(n1299), .Q(n1301) );
  AOI221 U1006 ( .A(n1576), .B(n1190), .C(n1574), .D(n1189), .Q(n1191) );
  AOI221 U1007 ( .A(n1576), .B(n1168), .C(n1574), .D(n1167), .Q(n1169) );
  AOI221 U1008 ( .A(n1576), .B(n1278), .C(n1574), .D(n1277), .Q(n1279) );
  AOI221 U1009 ( .A(n1556), .B(n1114), .C(n1554), .D(n1113), .Q(n1126) );
  AOI221 U1010 ( .A(n1556), .B(n1510), .C(n1554), .D(n1509), .Q(n1522) );
  AOI221 U1011 ( .A(n1556), .B(n1444), .C(n1554), .D(n1443), .Q(n1456) );
  AOI221 U1012 ( .A(n1556), .B(n1466), .C(n1554), .D(n1465), .Q(n1478) );
  AOI221 U1013 ( .A(n1556), .B(n1422), .C(n1554), .D(n1421), .Q(n1434) );
  NOR31 U1014 ( .A(i_addr_Rs[1]), .B(i_addr_Rs[2]), .C(n859), .Q(n1565) );
  NOR31 U1015 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[1]), .C(n857), .Q(n1563) );
  NOR40 U1016 ( .A(n108), .B(n1585), .C(n1586), .D(n1582), .Q(n27) );
  NOR40 U1017 ( .A(n108), .B(i_addr_Rd[1]), .C(n1586), .D(n1582), .Q(n25) );
  NOR40 U1018 ( .A(n108), .B(n1585), .C(n1586), .D(n1587), .Q(n17) );
  NOR40 U1019 ( .A(n108), .B(i_addr_Rd[1]), .C(n1586), .D(n1587), .Q(n15) );
  NOR40 U1020 ( .A(i_addr_Rd[1]), .B(n108), .C(n1586), .D(n1591), .Q(n42) );
  NOR40 U1021 ( .A(i_addr_Rd[0]), .B(n108), .C(n1591), .D(n1585), .Q(n43) );
  NOR40 U1022 ( .A(i_addr_Rd[0]), .B(n108), .C(n1585), .D(n1581), .Q(n35) );
  NOR40 U1023 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n108), .D(n1581), .Q(
        n32) );
  NOR40 U1024 ( .A(n108), .B(i_addr_Rd[1]), .C(n1586), .D(n1581), .Q(n34) );
  BUF2 U1025 ( .A(n36), .Q(n119) );
  NOR40 U1026 ( .A(n108), .B(n1585), .C(n1586), .D(n1581), .Q(n36) );
  NAND22 U1027 ( .A(n1580), .B(n1583), .Q(n1581) );
  AOI221 U1028 ( .A(n1576), .B(n926), .C(n1574), .D(n925), .Q(n927) );
  NOR40 U1029 ( .A(i_addr_Rd[0]), .B(n108), .C(n1585), .D(n1582), .Q(n26) );
  NOR40 U1030 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n108), .D(n1582), .Q(
        n23) );
  NOR40 U1031 ( .A(i_addr_Rd[0]), .B(n108), .C(n1585), .D(n1587), .Q(n16) );
  NOR40 U1032 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n108), .D(n1587), .Q(
        n13) );
  NOR40 U1033 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[0]), .C(n108), .D(n1591), .Q(
        n41) );
  NAND22 U1034 ( .A(n756), .B(n755), .Q(o_data_Rt[27]) );
  AOI221 U1035 ( .A(n854), .B(n754), .C(n852), .D(n753), .Q(n755) );
  NAND41 U1036 ( .A(n752), .B(n751), .C(n750), .D(n749), .Q(n753) );
  NAND41 U1037 ( .A(n748), .B(n747), .C(n746), .D(n745), .Q(n754) );
  NAND41 U1038 ( .A(n742), .B(n741), .C(n740), .D(n739), .Q(n743) );
  NAND41 U1039 ( .A(n738), .B(n737), .C(n736), .D(n735), .Q(n744) );
  NAND22 U1040 ( .A(n668), .B(n667), .Q(o_data_Rt[23]) );
  AOI221 U1041 ( .A(n854), .B(n666), .C(n852), .D(n665), .Q(n667) );
  NAND41 U1042 ( .A(n664), .B(n663), .C(n662), .D(n661), .Q(n665) );
  NAND41 U1043 ( .A(n660), .B(n659), .C(n658), .D(n657), .Q(n666) );
  NAND41 U1044 ( .A(n654), .B(n653), .C(n652), .D(n651), .Q(n655) );
  NAND41 U1045 ( .A(n650), .B(n649), .C(n648), .D(n647), .Q(n656) );
  NAND22 U1046 ( .A(n580), .B(n579), .Q(o_data_Rt[19]) );
  AOI221 U1047 ( .A(n854), .B(n578), .C(n852), .D(n577), .Q(n579) );
  NAND41 U1048 ( .A(n576), .B(n575), .C(n574), .D(n573), .Q(n577) );
  NAND41 U1049 ( .A(n572), .B(n571), .C(n570), .D(n569), .Q(n578) );
  NAND41 U1050 ( .A(n566), .B(n565), .C(n564), .D(n563), .Q(n567) );
  NAND41 U1051 ( .A(n562), .B(n561), .C(n560), .D(n559), .Q(n568) );
  NAND22 U1052 ( .A(n712), .B(n711), .Q(o_data_Rt[25]) );
  AOI221 U1053 ( .A(n854), .B(n710), .C(n852), .D(n709), .Q(n711) );
  NAND41 U1054 ( .A(n708), .B(n707), .C(n706), .D(n705), .Q(n709) );
  NAND41 U1055 ( .A(n704), .B(n703), .C(n702), .D(n701), .Q(n710) );
  NAND41 U1056 ( .A(n698), .B(n697), .C(n696), .D(n695), .Q(n699) );
  AOI221 U1057 ( .A(n70), .B(regs[505]), .C(n839), .D(regs[441]), .Q(n698) );
  NAND41 U1058 ( .A(n694), .B(n693), .C(n692), .D(n691), .Q(n700) );
  AOI221 U1059 ( .A(n70), .B(regs[1017]), .C(n839), .D(regs[953]), .Q(n694) );
  NAND22 U1060 ( .A(n624), .B(n623), .Q(o_data_Rt[21]) );
  AOI221 U1061 ( .A(n854), .B(n622), .C(n852), .D(n621), .Q(n623) );
  NAND41 U1062 ( .A(n620), .B(n619), .C(n618), .D(n617), .Q(n621) );
  NAND41 U1063 ( .A(n616), .B(n615), .C(n614), .D(n613), .Q(n622) );
  AOI221 U1064 ( .A(n834), .B(n612), .C(n832), .D(n611), .Q(n624) );
  NAND41 U1065 ( .A(n610), .B(n609), .C(n608), .D(n607), .Q(n611) );
  NAND41 U1066 ( .A(n606), .B(n605), .C(n604), .D(n603), .Q(n612) );
  NAND22 U1067 ( .A(n646), .B(n645), .Q(o_data_Rt[22]) );
  AOI221 U1068 ( .A(n854), .B(n644), .C(n852), .D(n643), .Q(n645) );
  NAND41 U1069 ( .A(n642), .B(n641), .C(n640), .D(n639), .Q(n643) );
  NAND41 U1070 ( .A(n638), .B(n637), .C(n636), .D(n635), .Q(n644) );
  AOI221 U1071 ( .A(n834), .B(n634), .C(n832), .D(n633), .Q(n646) );
  NAND41 U1072 ( .A(n632), .B(n631), .C(n630), .D(n629), .Q(n633) );
  NAND41 U1073 ( .A(n628), .B(n627), .C(n626), .D(n625), .Q(n634) );
  NAND22 U1074 ( .A(n602), .B(n601), .Q(o_data_Rt[20]) );
  AOI221 U1075 ( .A(n854), .B(n600), .C(n852), .D(n599), .Q(n601) );
  NAND41 U1076 ( .A(n598), .B(n597), .C(n596), .D(n595), .Q(n599) );
  NAND41 U1077 ( .A(n594), .B(n593), .C(n592), .D(n591), .Q(n600) );
  NAND41 U1078 ( .A(n588), .B(n587), .C(n586), .D(n585), .Q(n589) );
  NAND41 U1079 ( .A(n584), .B(n583), .C(n582), .D(n581), .Q(n590) );
  NAND22 U1080 ( .A(n690), .B(n689), .Q(o_data_Rt[24]) );
  AOI221 U1081 ( .A(n854), .B(n688), .C(n852), .D(n687), .Q(n689) );
  NAND41 U1082 ( .A(n686), .B(n685), .C(n684), .D(n683), .Q(n687) );
  NAND41 U1083 ( .A(n682), .B(n681), .C(n680), .D(n679), .Q(n688) );
  NAND41 U1084 ( .A(n676), .B(n675), .C(n674), .D(n673), .Q(n677) );
  NAND41 U1085 ( .A(n672), .B(n671), .C(n670), .D(n669), .Q(n678) );
  NAND22 U1086 ( .A(n822), .B(n821), .Q(o_data_Rt[30]) );
  AOI221 U1087 ( .A(n854), .B(n820), .C(n852), .D(n819), .Q(n821) );
  NAND41 U1088 ( .A(n818), .B(n817), .C(n816), .D(n815), .Q(n819) );
  AOI221 U1089 ( .A(n70), .B(regs[254]), .C(n839), .D(regs[190]), .Q(n818) );
  NAND41 U1090 ( .A(n814), .B(n813), .C(n812), .D(n811), .Q(n820) );
  AOI221 U1091 ( .A(n70), .B(regs[766]), .C(n67), .D(regs[702]), .Q(n814) );
  NAND41 U1092 ( .A(n808), .B(n807), .C(n806), .D(n805), .Q(n809) );
  AOI221 U1093 ( .A(n70), .B(regs[510]), .C(n67), .D(regs[446]), .Q(n808) );
  NAND41 U1094 ( .A(n804), .B(n803), .C(n802), .D(n801), .Q(n810) );
  NAND22 U1095 ( .A(n856), .B(n855), .Q(o_data_Rt[31]) );
  AOI221 U1096 ( .A(n854), .B(n853), .C(n852), .D(n851), .Q(n855) );
  NAND41 U1097 ( .A(n850), .B(n849), .C(n848), .D(n847), .Q(n851) );
  NAND41 U1098 ( .A(n838), .B(n837), .C(n836), .D(n835), .Q(n853) );
  AOI221 U1099 ( .A(n70), .B(regs[767]), .C(n67), .D(regs[703]), .Q(n838) );
  NAND41 U1100 ( .A(n830), .B(n829), .C(n828), .D(n827), .Q(n831) );
  NAND41 U1101 ( .A(n826), .B(n825), .C(n824), .D(n823), .Q(n833) );
  AOI221 U1102 ( .A(n70), .B(regs[1023]), .C(n839), .D(regs[959]), .Q(n826) );
  NAND41 U1103 ( .A(n796), .B(n795), .C(n794), .D(n793), .Q(n797) );
  NAND41 U1104 ( .A(n792), .B(n791), .C(n790), .D(n789), .Q(n798) );
  NAND41 U1105 ( .A(n786), .B(n785), .C(n784), .D(n783), .Q(n787) );
  NAND41 U1106 ( .A(n782), .B(n781), .C(n780), .D(n779), .Q(n788) );
  NAND22 U1107 ( .A(n778), .B(n777), .Q(o_data_Rt[28]) );
  AOI221 U1108 ( .A(n854), .B(n776), .C(n852), .D(n775), .Q(n777) );
  NAND41 U1109 ( .A(n774), .B(n773), .C(n772), .D(n771), .Q(n775) );
  NAND41 U1110 ( .A(n770), .B(n769), .C(n768), .D(n767), .Q(n776) );
  NAND41 U1111 ( .A(n764), .B(n763), .C(n762), .D(n761), .Q(n765) );
  NAND41 U1112 ( .A(n760), .B(n759), .C(n758), .D(n757), .Q(n766) );
  NAND22 U1113 ( .A(n734), .B(n733), .Q(o_data_Rt[26]) );
  AOI221 U1114 ( .A(n854), .B(n732), .C(n852), .D(n731), .Q(n733) );
  NAND41 U1115 ( .A(n730), .B(n729), .C(n728), .D(n727), .Q(n731) );
  NAND41 U1116 ( .A(n726), .B(n725), .C(n724), .D(n723), .Q(n732) );
  NAND41 U1117 ( .A(n720), .B(n719), .C(n718), .D(n717), .Q(n721) );
  NAND41 U1118 ( .A(n716), .B(n715), .C(n714), .D(n713), .Q(n722) );
  NAND22 U1119 ( .A(n558), .B(n557), .Q(o_data_Rt[18]) );
  AOI221 U1120 ( .A(n854), .B(n556), .C(n852), .D(n555), .Q(n557) );
  NAND41 U1121 ( .A(n554), .B(n553), .C(n552), .D(n551), .Q(n555) );
  NAND41 U1122 ( .A(n550), .B(n549), .C(n548), .D(n547), .Q(n556) );
  NAND41 U1123 ( .A(n544), .B(n543), .C(n542), .D(n541), .Q(n545) );
  NAND41 U1124 ( .A(n540), .B(n539), .C(n538), .D(n537), .Q(n546) );
  NAND22 U1125 ( .A(n272), .B(n271), .Q(o_data_Rt[5]) );
  AOI221 U1126 ( .A(n854), .B(n270), .C(n852), .D(n269), .Q(n271) );
  NAND41 U1127 ( .A(n268), .B(n267), .C(n266), .D(n265), .Q(n269) );
  NAND41 U1128 ( .A(n264), .B(n263), .C(n262), .D(n261), .Q(n270) );
  AOI221 U1129 ( .A(n834), .B(n260), .C(n832), .D(n259), .Q(n272) );
  NAND41 U1130 ( .A(n258), .B(n257), .C(n256), .D(n255), .Q(n259) );
  NAND41 U1131 ( .A(n254), .B(n253), .C(n252), .D(n251), .Q(n260) );
  NAND22 U1132 ( .A(n316), .B(n315), .Q(o_data_Rt[7]) );
  AOI221 U1133 ( .A(n854), .B(n314), .C(n852), .D(n313), .Q(n315) );
  NAND41 U1134 ( .A(n312), .B(n311), .C(n310), .D(n309), .Q(n313) );
  NAND41 U1135 ( .A(n308), .B(n307), .C(n306), .D(n305), .Q(n314) );
  NAND41 U1136 ( .A(n302), .B(n301), .C(n300), .D(n299), .Q(n303) );
  NAND41 U1137 ( .A(n298), .B(n297), .C(n296), .D(n295), .Q(n304) );
  NAND22 U1138 ( .A(n404), .B(n403), .Q(o_data_Rt[11]) );
  AOI221 U1139 ( .A(n854), .B(n402), .C(n852), .D(n401), .Q(n403) );
  NAND41 U1140 ( .A(n400), .B(n399), .C(n398), .D(n397), .Q(n401) );
  NAND41 U1141 ( .A(n396), .B(n395), .C(n394), .D(n393), .Q(n402) );
  NAND41 U1142 ( .A(n390), .B(n389), .C(n388), .D(n387), .Q(n391) );
  NAND41 U1143 ( .A(n386), .B(n385), .C(n384), .D(n383), .Q(n392) );
  NAND22 U1144 ( .A(n228), .B(n227), .Q(o_data_Rt[3]) );
  AOI221 U1145 ( .A(n854), .B(n226), .C(n852), .D(n225), .Q(n227) );
  NAND41 U1146 ( .A(n224), .B(n223), .C(n222), .D(n221), .Q(n225) );
  NAND41 U1147 ( .A(n220), .B(n219), .C(n218), .D(n217), .Q(n226) );
  NAND41 U1148 ( .A(n214), .B(n213), .C(n212), .D(n211), .Q(n215) );
  NAND41 U1149 ( .A(n210), .B(n209), .C(n208), .D(n207), .Q(n216) );
  NAND22 U1150 ( .A(n184), .B(n183), .Q(o_data_Rt[1]) );
  NAND41 U1151 ( .A(n180), .B(n179), .C(n178), .D(n177), .Q(n181) );
  NAND41 U1152 ( .A(n176), .B(n175), .C(n174), .D(n173), .Q(n182) );
  NAND41 U1153 ( .A(n170), .B(n169), .C(n168), .D(n167), .Q(n171) );
  NAND41 U1154 ( .A(n166), .B(n165), .C(n164), .D(n163), .Q(n172) );
  NAND22 U1155 ( .A(n294), .B(n293), .Q(o_data_Rt[6]) );
  NAND41 U1156 ( .A(n290), .B(n289), .C(n288), .D(n287), .Q(n291) );
  AOI221 U1157 ( .A(n111), .B(regs[70]), .C(n845), .D(regs[6]), .Q(n287) );
  NAND41 U1158 ( .A(n286), .B(n285), .C(n284), .D(n283), .Q(n292) );
  AOI221 U1159 ( .A(n111), .B(regs[582]), .C(n110), .D(regs[518]), .Q(n283) );
  NAND41 U1160 ( .A(n280), .B(n279), .C(n278), .D(n277), .Q(n281) );
  NAND41 U1161 ( .A(n276), .B(n275), .C(n274), .D(n273), .Q(n282) );
  NAND22 U1162 ( .A(n162), .B(n161), .Q(o_data_Rt[0]) );
  AOI221 U1163 ( .A(n854), .B(n160), .C(n852), .D(n159), .Q(n161) );
  NAND41 U1164 ( .A(n158), .B(n157), .C(n156), .D(n155), .Q(n159) );
  AOI221 U1165 ( .A(n70), .B(regs[224]), .C(n67), .D(regs[160]), .Q(n158) );
  NAND41 U1166 ( .A(n154), .B(n153), .C(n152), .D(n151), .Q(n160) );
  NAND41 U1167 ( .A(n147), .B(n146), .C(n145), .D(n144), .Q(n148) );
  NAND41 U1168 ( .A(n142), .B(n141), .C(n140), .D(n139), .Q(n149) );
  AOI221 U1169 ( .A(n70), .B(regs[992]), .C(n839), .D(regs[928]), .Q(n142) );
  NAND22 U1170 ( .A(n448), .B(n447), .Q(o_data_Rt[13]) );
  NAND41 U1171 ( .A(n444), .B(n443), .C(n442), .D(n441), .Q(n445) );
  AOI221 U1172 ( .A(n111), .B(regs[77]), .C(n845), .D(regs[13]), .Q(n441) );
  NAND41 U1173 ( .A(n440), .B(n439), .C(n438), .D(n437), .Q(n446) );
  NAND41 U1174 ( .A(n434), .B(n433), .C(n432), .D(n431), .Q(n435) );
  NAND41 U1175 ( .A(n430), .B(n429), .C(n428), .D(n427), .Q(n436) );
  AOI221 U1176 ( .A(n111), .B(regs[845]), .C(n845), .D(regs[781]), .Q(n427) );
  NAND22 U1177 ( .A(n382), .B(n381), .Q(o_data_Rt[10]) );
  AOI221 U1178 ( .A(n854), .B(n380), .C(n852), .D(n379), .Q(n381) );
  NAND41 U1179 ( .A(n378), .B(n377), .C(n376), .D(n375), .Q(n379) );
  NAND41 U1180 ( .A(n374), .B(n373), .C(n372), .D(n371), .Q(n380) );
  AOI221 U1181 ( .A(n834), .B(n370), .C(n832), .D(n369), .Q(n382) );
  NAND41 U1182 ( .A(n368), .B(n367), .C(n366), .D(n365), .Q(n369) );
  NAND41 U1183 ( .A(n364), .B(n363), .C(n362), .D(n361), .Q(n370) );
  NAND22 U1184 ( .A(n426), .B(n425), .Q(o_data_Rt[12]) );
  AOI221 U1185 ( .A(n854), .B(n424), .C(n852), .D(n423), .Q(n425) );
  NAND41 U1186 ( .A(n422), .B(n421), .C(n420), .D(n419), .Q(n423) );
  NAND41 U1187 ( .A(n418), .B(n417), .C(n416), .D(n415), .Q(n424) );
  AOI221 U1188 ( .A(n834), .B(n414), .C(n832), .D(n413), .Q(n426) );
  NAND41 U1189 ( .A(n412), .B(n411), .C(n410), .D(n409), .Q(n413) );
  NAND41 U1190 ( .A(n408), .B(n407), .C(n406), .D(n405), .Q(n414) );
  NAND22 U1191 ( .A(n360), .B(n359), .Q(o_data_Rt[9]) );
  AOI221 U1192 ( .A(n854), .B(n358), .C(n852), .D(n357), .Q(n359) );
  NAND41 U1193 ( .A(n356), .B(n355), .C(n354), .D(n353), .Q(n357) );
  NAND41 U1194 ( .A(n352), .B(n351), .C(n350), .D(n349), .Q(n358) );
  NAND41 U1195 ( .A(n346), .B(n345), .C(n344), .D(n343), .Q(n347) );
  NAND41 U1196 ( .A(n342), .B(n341), .C(n340), .D(n339), .Q(n348) );
  NAND22 U1197 ( .A(n492), .B(n491), .Q(o_data_Rt[15]) );
  NAND41 U1198 ( .A(n488), .B(n487), .C(n486), .D(n485), .Q(n489) );
  AOI221 U1199 ( .A(n111), .B(regs[79]), .C(n845), .D(regs[15]), .Q(n485) );
  NAND41 U1200 ( .A(n484), .B(n483), .C(n482), .D(n481), .Q(n490) );
  NAND41 U1201 ( .A(n478), .B(n477), .C(n476), .D(n475), .Q(n479) );
  NAND41 U1202 ( .A(n474), .B(n473), .C(n472), .D(n471), .Q(n480) );
  NAND22 U1203 ( .A(n470), .B(n469), .Q(o_data_Rt[14]) );
  NAND41 U1204 ( .A(n466), .B(n465), .C(n464), .D(n463), .Q(n467) );
  NAND41 U1205 ( .A(n462), .B(n461), .C(n460), .D(n459), .Q(n468) );
  NAND41 U1206 ( .A(n456), .B(n455), .C(n454), .D(n453), .Q(n457) );
  AOI221 U1207 ( .A(n70), .B(regs[494]), .C(n67), .D(regs[430]), .Q(n456) );
  NAND41 U1208 ( .A(n452), .B(n451), .C(n450), .D(n449), .Q(n458) );
  NAND22 U1209 ( .A(n206), .B(n205), .Q(o_data_Rt[2]) );
  NAND41 U1210 ( .A(n202), .B(n201), .C(n200), .D(n199), .Q(n203) );
  NAND41 U1211 ( .A(n198), .B(n197), .C(n196), .D(n195), .Q(n204) );
  NAND41 U1212 ( .A(n192), .B(n191), .C(n190), .D(n189), .Q(n193) );
  NAND41 U1213 ( .A(n188), .B(n187), .C(n186), .D(n185), .Q(n194) );
  NAND22 U1214 ( .A(n536), .B(n535), .Q(o_data_Rt[17]) );
  NAND41 U1215 ( .A(n532), .B(n531), .C(n530), .D(n529), .Q(n533) );
  NAND41 U1216 ( .A(n528), .B(n527), .C(n526), .D(n525), .Q(n534) );
  AOI221 U1217 ( .A(n70), .B(regs[753]), .C(n839), .D(regs[689]), .Q(n528) );
  NAND41 U1218 ( .A(n522), .B(n521), .C(n520), .D(n519), .Q(n523) );
  NAND41 U1219 ( .A(n518), .B(n517), .C(n516), .D(n515), .Q(n524) );
  NAND22 U1220 ( .A(n514), .B(n513), .Q(o_data_Rt[16]) );
  NAND41 U1221 ( .A(n510), .B(n509), .C(n508), .D(n507), .Q(n511) );
  NAND41 U1222 ( .A(n506), .B(n505), .C(n504), .D(n503), .Q(n512) );
  NAND41 U1223 ( .A(n500), .B(n499), .C(n498), .D(n497), .Q(n501) );
  NAND41 U1224 ( .A(n496), .B(n495), .C(n494), .D(n493), .Q(n502) );
  NAND22 U1225 ( .A(n250), .B(n249), .Q(o_data_Rt[4]) );
  NAND41 U1226 ( .A(n246), .B(n245), .C(n244), .D(n243), .Q(n247) );
  AOI221 U1227 ( .A(n111), .B(regs[68]), .C(n110), .D(regs[4]), .Q(n243) );
  AOI221 U1228 ( .A(n70), .B(regs[228]), .C(n67), .D(regs[164]), .Q(n246) );
  NAND41 U1229 ( .A(n242), .B(n241), .C(n240), .D(n239), .Q(n248) );
  AOI221 U1230 ( .A(n70), .B(regs[740]), .C(n67), .D(regs[676]), .Q(n242) );
  NAND41 U1231 ( .A(n236), .B(n235), .C(n234), .D(n233), .Q(n237) );
  NAND41 U1232 ( .A(n232), .B(n231), .C(n230), .D(n229), .Q(n238) );
  NAND22 U1233 ( .A(n338), .B(n337), .Q(o_data_Rt[8]) );
  NAND41 U1234 ( .A(n334), .B(n333), .C(n332), .D(n331), .Q(n335) );
  NAND41 U1235 ( .A(n330), .B(n329), .C(n328), .D(n327), .Q(n336) );
  NAND41 U1236 ( .A(n324), .B(n323), .C(n322), .D(n321), .Q(n325) );
  AOI221 U1237 ( .A(n111), .B(regs[328]), .C(n845), .D(regs[264]), .Q(n321) );
  NAND41 U1238 ( .A(n320), .B(n319), .C(n318), .D(n317), .Q(n326) );
  AOI221 U1239 ( .A(n111), .B(regs[840]), .C(n845), .D(regs[776]), .Q(n317) );
  NAND22 U1240 ( .A(n884), .B(n883), .Q(o_data_Rs[0]) );
  NAND41 U1241 ( .A(n880), .B(n879), .C(n878), .D(n877), .Q(n881) );
  NAND41 U1242 ( .A(n876), .B(n875), .C(n874), .D(n873), .Q(n882) );
  AOI221 U1243 ( .A(n1556), .B(n871), .C(n1554), .D(n870), .Q(n884) );
  NAND41 U1244 ( .A(n869), .B(n868), .C(n867), .D(n866), .Q(n870) );
  NAND41 U1245 ( .A(n864), .B(n863), .C(n862), .D(n861), .Q(n871) );
  NAND22 U1246 ( .A(n906), .B(n905), .Q(o_data_Rs[1]) );
  NAND41 U1247 ( .A(n902), .B(n901), .C(n900), .D(n899), .Q(n903) );
  NAND41 U1248 ( .A(n898), .B(n897), .C(n896), .D(n895), .Q(n904) );
  AOI221 U1249 ( .A(n1556), .B(n894), .C(n1554), .D(n893), .Q(n906) );
  NAND41 U1250 ( .A(n892), .B(n891), .C(n890), .D(n889), .Q(n893) );
  NAND41 U1251 ( .A(n888), .B(n887), .C(n886), .D(n885), .Q(n894) );
  NAND22 U1252 ( .A(n950), .B(n949), .Q(o_data_Rs[3]) );
  NAND41 U1253 ( .A(n946), .B(n945), .C(n944), .D(n943), .Q(n947) );
  NAND41 U1254 ( .A(n942), .B(n941), .C(n940), .D(n939), .Q(n948) );
  NAND41 U1255 ( .A(n936), .B(n935), .C(n934), .D(n933), .Q(n937) );
  NAND41 U1256 ( .A(n932), .B(n931), .C(n930), .D(n929), .Q(n938) );
  NAND22 U1257 ( .A(n1016), .B(n1015), .Q(o_data_Rs[6]) );
  AOI221 U1258 ( .A(n1576), .B(n1014), .C(n1574), .D(n1013), .Q(n1015) );
  NAND41 U1259 ( .A(n1012), .B(n1011), .C(n1010), .D(n1009), .Q(n1013) );
  NAND41 U1260 ( .A(n1008), .B(n1007), .C(n1006), .D(n1005), .Q(n1014) );
  NAND41 U1261 ( .A(n1002), .B(n1001), .C(n1000), .D(n999), .Q(n1003) );
  NAND41 U1262 ( .A(n998), .B(n997), .C(n996), .D(n995), .Q(n1004) );
  NAND22 U1263 ( .A(n928), .B(n927), .Q(o_data_Rs[2]) );
  NAND41 U1264 ( .A(n924), .B(n923), .C(n922), .D(n921), .Q(n925) );
  NAND41 U1265 ( .A(n920), .B(n919), .C(n918), .D(n917), .Q(n926) );
  NAND41 U1266 ( .A(n914), .B(n913), .C(n912), .D(n911), .Q(n915) );
  NAND41 U1267 ( .A(n910), .B(n909), .C(n908), .D(n907), .Q(n916) );
  NAND22 U1268 ( .A(n972), .B(n971), .Q(o_data_Rs[4]) );
  NAND41 U1269 ( .A(n968), .B(n967), .C(n966), .D(n965), .Q(n969) );
  NAND41 U1270 ( .A(n964), .B(n963), .C(n962), .D(n961), .Q(n970) );
  NAND41 U1271 ( .A(n958), .B(n957), .C(n956), .D(n955), .Q(n959) );
  NAND41 U1272 ( .A(n954), .B(n953), .C(n952), .D(n951), .Q(n960) );
  NAND22 U1273 ( .A(n994), .B(n993), .Q(o_data_Rs[5]) );
  NAND41 U1274 ( .A(n990), .B(n989), .C(n988), .D(n987), .Q(n991) );
  NAND41 U1275 ( .A(n986), .B(n985), .C(n984), .D(n983), .Q(n992) );
  NAND41 U1276 ( .A(n980), .B(n979), .C(n978), .D(n977), .Q(n981) );
  NAND41 U1277 ( .A(n976), .B(n975), .C(n974), .D(n973), .Q(n982) );
  NAND22 U1278 ( .A(n1500), .B(n1499), .Q(o_data_Rs[28]) );
  NAND41 U1279 ( .A(n1496), .B(n1495), .C(n1494), .D(n1493), .Q(n1497) );
  NAND41 U1280 ( .A(n1492), .B(n1491), .C(n1490), .D(n1489), .Q(n1498) );
  NAND41 U1281 ( .A(n1486), .B(n1485), .C(n1484), .D(n1483), .Q(n1487) );
  NAND41 U1282 ( .A(n1482), .B(n1481), .C(n1480), .D(n1479), .Q(n1488) );
  NAND22 U1283 ( .A(n1060), .B(n1059), .Q(o_data_Rs[8]) );
  AOI221 U1284 ( .A(n1576), .B(n1058), .C(n1574), .D(n1057), .Q(n1059) );
  NAND41 U1285 ( .A(n1056), .B(n1055), .C(n1054), .D(n1053), .Q(n1057) );
  NAND41 U1286 ( .A(n1052), .B(n1051), .C(n1050), .D(n1049), .Q(n1058) );
  AOI221 U1287 ( .A(n1556), .B(n1048), .C(n1554), .D(n1047), .Q(n1060) );
  NAND41 U1288 ( .A(n1046), .B(n1045), .C(n1044), .D(n1043), .Q(n1047) );
  NAND41 U1289 ( .A(n1042), .B(n1041), .C(n1040), .D(n1039), .Q(n1048) );
  NAND22 U1290 ( .A(n1038), .B(n1037), .Q(o_data_Rs[7]) );
  NAND41 U1291 ( .A(n1034), .B(n1033), .C(n1032), .D(n1031), .Q(n1035) );
  NAND41 U1292 ( .A(n1030), .B(n1029), .C(n1028), .D(n1027), .Q(n1036) );
  AOI221 U1293 ( .A(n1556), .B(n1026), .C(n1554), .D(n1025), .Q(n1038) );
  NAND41 U1294 ( .A(n1024), .B(n1023), .C(n1022), .D(n1021), .Q(n1025) );
  NAND41 U1295 ( .A(n1020), .B(n1019), .C(n1018), .D(n1017), .Q(n1026) );
  NAND22 U1296 ( .A(n1104), .B(n1103), .Q(o_data_Rs[10]) );
  AOI221 U1297 ( .A(n1576), .B(n1102), .C(n1574), .D(n1101), .Q(n1103) );
  NAND41 U1298 ( .A(n1100), .B(n1099), .C(n1098), .D(n1097), .Q(n1101) );
  NAND41 U1299 ( .A(n1096), .B(n1095), .C(n1094), .D(n1093), .Q(n1102) );
  NAND41 U1300 ( .A(n1090), .B(n1089), .C(n1088), .D(n1087), .Q(n1091) );
  NAND41 U1301 ( .A(n1086), .B(n1085), .C(n1084), .D(n1083), .Q(n1092) );
  NAND22 U1302 ( .A(n1302), .B(n1301), .Q(o_data_Rs[19]) );
  NAND41 U1303 ( .A(n1298), .B(n1297), .C(n1296), .D(n1295), .Q(n1299) );
  NAND41 U1304 ( .A(n1294), .B(n1293), .C(n1292), .D(n1291), .Q(n1300) );
  NAND41 U1305 ( .A(n1288), .B(n1287), .C(n1286), .D(n1285), .Q(n1289) );
  NAND41 U1306 ( .A(n1284), .B(n1283), .C(n1282), .D(n1281), .Q(n1290) );
  NAND22 U1307 ( .A(n1192), .B(n1191), .Q(o_data_Rs[14]) );
  NAND41 U1308 ( .A(n1188), .B(n1187), .C(n1186), .D(n1185), .Q(n1189) );
  NAND41 U1309 ( .A(n1184), .B(n1183), .C(n1182), .D(n1181), .Q(n1190) );
  AOI221 U1310 ( .A(n1556), .B(n1180), .C(n1554), .D(n1179), .Q(n1192) );
  NAND41 U1311 ( .A(n1178), .B(n1177), .C(n1176), .D(n1175), .Q(n1179) );
  NAND41 U1312 ( .A(n1174), .B(n1173), .C(n1172), .D(n1171), .Q(n1180) );
  NAND22 U1313 ( .A(n1258), .B(n1257), .Q(o_data_Rs[17]) );
  AOI221 U1314 ( .A(n1576), .B(n1256), .C(n1574), .D(n1255), .Q(n1257) );
  NAND41 U1315 ( .A(n1254), .B(n1253), .C(n1252), .D(n1251), .Q(n1255) );
  NAND41 U1316 ( .A(n1250), .B(n1249), .C(n1248), .D(n1247), .Q(n1256) );
  AOI221 U1317 ( .A(n1556), .B(n1246), .C(n1554), .D(n1245), .Q(n1258) );
  NAND41 U1318 ( .A(n1244), .B(n1243), .C(n1242), .D(n1241), .Q(n1245) );
  NAND41 U1319 ( .A(n1240), .B(n1239), .C(n1238), .D(n1237), .Q(n1246) );
  NAND22 U1320 ( .A(n1578), .B(n1577), .Q(o_data_Rs[31]) );
  AOI221 U1321 ( .A(n1576), .B(n1575), .C(n1574), .D(n1573), .Q(n1577) );
  NAND41 U1322 ( .A(n1572), .B(n1571), .C(n1570), .D(n1569), .Q(n1573) );
  NAND41 U1323 ( .A(n1560), .B(n1559), .C(n1558), .D(n1557), .Q(n1575) );
  AOI221 U1324 ( .A(n1556), .B(n1555), .C(n1554), .D(n1553), .Q(n1578) );
  NAND41 U1325 ( .A(n1552), .B(n1551), .C(n1550), .D(n1549), .Q(n1553) );
  NAND41 U1326 ( .A(n1548), .B(n1547), .C(n1546), .D(n1545), .Q(n1555) );
  NAND22 U1327 ( .A(n1214), .B(n1213), .Q(o_data_Rs[15]) );
  AOI221 U1328 ( .A(n1576), .B(n1212), .C(n1574), .D(n1211), .Q(n1213) );
  NAND41 U1329 ( .A(n1210), .B(n1209), .C(n1208), .D(n1207), .Q(n1211) );
  NAND41 U1330 ( .A(n1206), .B(n1205), .C(n1204), .D(n1203), .Q(n1212) );
  AOI221 U1331 ( .A(n1556), .B(n1202), .C(n1554), .D(n1201), .Q(n1214) );
  NAND41 U1332 ( .A(n1200), .B(n1199), .C(n1198), .D(n1197), .Q(n1201) );
  NAND41 U1333 ( .A(n1196), .B(n1195), .C(n1194), .D(n1193), .Q(n1202) );
  NAND22 U1334 ( .A(n1236), .B(n1235), .Q(o_data_Rs[16]) );
  AOI221 U1335 ( .A(n1576), .B(n1234), .C(n1574), .D(n1233), .Q(n1235) );
  NAND41 U1336 ( .A(n1232), .B(n1231), .C(n1230), .D(n1229), .Q(n1233) );
  NAND41 U1337 ( .A(n1228), .B(n1227), .C(n1226), .D(n1225), .Q(n1234) );
  AOI221 U1338 ( .A(n1556), .B(n1224), .C(n1554), .D(n1223), .Q(n1236) );
  NAND41 U1339 ( .A(n1222), .B(n1221), .C(n1220), .D(n1219), .Q(n1223) );
  NAND41 U1340 ( .A(n1218), .B(n1217), .C(n1216), .D(n1215), .Q(n1224) );
  NAND22 U1341 ( .A(n1170), .B(n1169), .Q(o_data_Rs[13]) );
  NAND41 U1342 ( .A(n1166), .B(n1165), .C(n1164), .D(n1163), .Q(n1167) );
  NAND41 U1343 ( .A(n1162), .B(n1161), .C(n1160), .D(n1159), .Q(n1168) );
  AOI221 U1344 ( .A(n1556), .B(n1158), .C(n1554), .D(n1157), .Q(n1170) );
  NAND41 U1345 ( .A(n1156), .B(n1155), .C(n1154), .D(n1153), .Q(n1157) );
  NAND41 U1346 ( .A(n1152), .B(n1151), .C(n1150), .D(n1149), .Q(n1158) );
  NAND22 U1347 ( .A(n1280), .B(n1279), .Q(o_data_Rs[18]) );
  NAND41 U1348 ( .A(n1276), .B(n1275), .C(n1274), .D(n1273), .Q(n1277) );
  NAND41 U1349 ( .A(n1272), .B(n1271), .C(n1270), .D(n1269), .Q(n1278) );
  NAND41 U1350 ( .A(n1266), .B(n1265), .C(n1264), .D(n1263), .Q(n1267) );
  NAND41 U1351 ( .A(n1262), .B(n1261), .C(n1260), .D(n1259), .Q(n1268) );
  NAND22 U1352 ( .A(n1148), .B(n1147), .Q(o_data_Rs[12]) );
  NAND41 U1353 ( .A(n1144), .B(n1143), .C(n1142), .D(n1141), .Q(n1145) );
  NAND41 U1354 ( .A(n1140), .B(n1139), .C(n1138), .D(n1137), .Q(n1146) );
  AOI221 U1355 ( .A(n1556), .B(n1136), .C(n1554), .D(n1135), .Q(n1148) );
  NAND41 U1356 ( .A(n1134), .B(n1133), .C(n1132), .D(n1131), .Q(n1135) );
  NAND41 U1357 ( .A(n1130), .B(n1129), .C(n1128), .D(n1127), .Q(n1136) );
  NAND22 U1358 ( .A(n1126), .B(n1125), .Q(o_data_Rs[11]) );
  NAND41 U1359 ( .A(n1122), .B(n1121), .C(n1120), .D(n1119), .Q(n1123) );
  NAND41 U1360 ( .A(n1118), .B(n1117), .C(n1116), .D(n1115), .Q(n1124) );
  NAND41 U1361 ( .A(n1112), .B(n1111), .C(n1110), .D(n1109), .Q(n1113) );
  NAND41 U1362 ( .A(n1108), .B(n1107), .C(n1106), .D(n1105), .Q(n1114) );
  NAND22 U1363 ( .A(n1522), .B(n1521), .Q(o_data_Rs[29]) );
  AOI221 U1364 ( .A(n1576), .B(n1520), .C(n1574), .D(n1519), .Q(n1521) );
  NAND41 U1365 ( .A(n1518), .B(n1517), .C(n1516), .D(n1515), .Q(n1519) );
  NAND41 U1366 ( .A(n1514), .B(n1513), .C(n1512), .D(n1511), .Q(n1520) );
  NAND41 U1367 ( .A(n1508), .B(n1507), .C(n1506), .D(n1505), .Q(n1509) );
  NAND41 U1368 ( .A(n1504), .B(n1503), .C(n1502), .D(n1501), .Q(n1510) );
  NAND22 U1369 ( .A(n1544), .B(n1543), .Q(o_data_Rs[30]) );
  AOI221 U1370 ( .A(n1576), .B(n1542), .C(n1574), .D(n1541), .Q(n1543) );
  NAND41 U1371 ( .A(n1540), .B(n1539), .C(n1538), .D(n1537), .Q(n1541) );
  NAND41 U1372 ( .A(n1536), .B(n1535), .C(n1534), .D(n1533), .Q(n1542) );
  AOI221 U1373 ( .A(n1556), .B(n1532), .C(n1554), .D(n1531), .Q(n1544) );
  NAND41 U1374 ( .A(n1530), .B(n1529), .C(n1528), .D(n1527), .Q(n1531) );
  NAND41 U1375 ( .A(n1526), .B(n1525), .C(n1524), .D(n1523), .Q(n1532) );
  NAND22 U1376 ( .A(n1082), .B(n1081), .Q(o_data_Rs[9]) );
  AOI221 U1377 ( .A(n1576), .B(n1080), .C(n1574), .D(n1079), .Q(n1081) );
  NAND41 U1378 ( .A(n1078), .B(n1077), .C(n1076), .D(n1075), .Q(n1079) );
  NAND41 U1379 ( .A(n1074), .B(n1073), .C(n1072), .D(n1071), .Q(n1080) );
  AOI221 U1380 ( .A(n1556), .B(n1070), .C(n1554), .D(n1069), .Q(n1082) );
  NAND41 U1381 ( .A(n1068), .B(n1067), .C(n1066), .D(n1065), .Q(n1069) );
  NAND41 U1382 ( .A(n1064), .B(n1063), .C(n1062), .D(n1061), .Q(n1070) );
  NAND22 U1383 ( .A(n1368), .B(n1367), .Q(o_data_Rs[22]) );
  NAND41 U1384 ( .A(n1364), .B(n1363), .C(n1362), .D(n1361), .Q(n1365) );
  NAND41 U1385 ( .A(n1360), .B(n1359), .C(n1358), .D(n1357), .Q(n1366) );
  AOI221 U1386 ( .A(n1556), .B(n1356), .C(n1554), .D(n1355), .Q(n1368) );
  NAND41 U1387 ( .A(n1354), .B(n1353), .C(n1352), .D(n1351), .Q(n1355) );
  NAND41 U1388 ( .A(n1350), .B(n1349), .C(n1348), .D(n1347), .Q(n1356) );
  NAND22 U1389 ( .A(n1456), .B(n1455), .Q(o_data_Rs[26]) );
  AOI221 U1390 ( .A(n1576), .B(n1454), .C(n1574), .D(n1453), .Q(n1455) );
  NAND41 U1391 ( .A(n1452), .B(n1451), .C(n1450), .D(n1449), .Q(n1453) );
  NAND41 U1392 ( .A(n1448), .B(n1447), .C(n1446), .D(n1445), .Q(n1454) );
  NAND41 U1393 ( .A(n1442), .B(n1441), .C(n1440), .D(n1439), .Q(n1443) );
  NAND41 U1394 ( .A(n1438), .B(n1437), .C(n1436), .D(n1435), .Q(n1444) );
  NAND22 U1395 ( .A(n1478), .B(n1477), .Q(o_data_Rs[27]) );
  AOI221 U1396 ( .A(n1576), .B(n1476), .C(n1574), .D(n1475), .Q(n1477) );
  NAND41 U1397 ( .A(n1474), .B(n1473), .C(n1472), .D(n1471), .Q(n1475) );
  NAND41 U1398 ( .A(n1470), .B(n1469), .C(n1468), .D(n1467), .Q(n1476) );
  NAND41 U1399 ( .A(n1464), .B(n1463), .C(n1462), .D(n1461), .Q(n1465) );
  NAND41 U1400 ( .A(n1460), .B(n1459), .C(n1458), .D(n1457), .Q(n1466) );
  NAND22 U1401 ( .A(n1346), .B(n1345), .Q(o_data_Rs[21]) );
  AOI221 U1402 ( .A(n1576), .B(n1344), .C(n1574), .D(n1343), .Q(n1345) );
  NAND41 U1403 ( .A(n1342), .B(n1341), .C(n1340), .D(n1339), .Q(n1343) );
  NAND41 U1404 ( .A(n1338), .B(n1337), .C(n1336), .D(n1335), .Q(n1344) );
  NAND41 U1405 ( .A(n1332), .B(n1331), .C(n1330), .D(n1329), .Q(n1333) );
  NAND41 U1406 ( .A(n1328), .B(n1327), .C(n1326), .D(n1325), .Q(n1334) );
  NAND22 U1407 ( .A(n1434), .B(n1433), .Q(o_data_Rs[25]) );
  AOI221 U1408 ( .A(n1576), .B(n1432), .C(n1574), .D(n1431), .Q(n1433) );
  NAND41 U1409 ( .A(n1430), .B(n1429), .C(n1428), .D(n1427), .Q(n1431) );
  NAND41 U1410 ( .A(n1426), .B(n1425), .C(n1424), .D(n1423), .Q(n1432) );
  NAND41 U1411 ( .A(n1420), .B(n1419), .C(n1418), .D(n1417), .Q(n1421) );
  NAND41 U1412 ( .A(n1416), .B(n1415), .C(n1414), .D(n1413), .Q(n1422) );
  NAND22 U1413 ( .A(n1390), .B(n1389), .Q(o_data_Rs[23]) );
  AOI221 U1414 ( .A(n1576), .B(n1388), .C(n1574), .D(n1387), .Q(n1389) );
  NAND41 U1415 ( .A(n1386), .B(n1385), .C(n1384), .D(n1383), .Q(n1387) );
  NAND41 U1416 ( .A(n1382), .B(n1381), .C(n1380), .D(n1379), .Q(n1388) );
  AOI221 U1417 ( .A(n1556), .B(n1378), .C(n1554), .D(n1377), .Q(n1390) );
  NAND41 U1418 ( .A(n1376), .B(n1375), .C(n1374), .D(n1373), .Q(n1377) );
  NAND41 U1419 ( .A(n1372), .B(n1371), .C(n1370), .D(n1369), .Q(n1378) );
  NAND22 U1420 ( .A(n1324), .B(n1323), .Q(o_data_Rs[20]) );
  NAND41 U1421 ( .A(n1320), .B(n1319), .C(n1318), .D(n1317), .Q(n1321) );
  NAND41 U1422 ( .A(n1316), .B(n1315), .C(n1314), .D(n1313), .Q(n1322) );
  AOI221 U1423 ( .A(n1556), .B(n1312), .C(n1554), .D(n1311), .Q(n1324) );
  NAND41 U1424 ( .A(n1310), .B(n1309), .C(n1308), .D(n1307), .Q(n1311) );
  NAND41 U1425 ( .A(n1306), .B(n1305), .C(n1304), .D(n1303), .Q(n1312) );
  NAND22 U1426 ( .A(n1412), .B(n1411), .Q(o_data_Rs[24]) );
  AOI221 U1427 ( .A(n1576), .B(n1410), .C(n1574), .D(n1409), .Q(n1411) );
  NAND41 U1428 ( .A(n1408), .B(n1407), .C(n1406), .D(n1405), .Q(n1409) );
  NAND41 U1429 ( .A(n1404), .B(n1403), .C(n1402), .D(n1401), .Q(n1410) );
  AOI221 U1430 ( .A(n1556), .B(n1400), .C(n1554), .D(n1399), .Q(n1412) );
  NAND41 U1431 ( .A(n1398), .B(n1397), .C(n1396), .D(n1395), .Q(n1399) );
  NAND41 U1432 ( .A(n1394), .B(n1393), .C(n1392), .D(n1391), .Q(n1400) );
  NAND22 U1433 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .Q(n136) );
  NOR21 U1434 ( .A(n1589), .B(n1587), .Q(n21) );
  NOR21 U1435 ( .A(n1590), .B(n1587), .Q(n20) );
  NOR21 U1436 ( .A(n1584), .B(n1587), .Q(n18) );
  NOR21 U1437 ( .A(n1588), .B(n1587), .Q(n22) );
  INV3 U1438 ( .A(i_addr_Rt_1_), .Q(n138) );
  INV3 U1439 ( .A(i_addr_Rt_0_), .Q(n137) );
  AOI220 U1440 ( .A(n840), .B(regs[994]), .C(n67), .D(regs[930]), .Q(n188) );
  AOI220 U1441 ( .A(n840), .B(regs[226]), .C(n67), .D(regs[162]), .Q(n202) );
  AOI220 U1442 ( .A(n844), .B(regs[98]), .C(n843), .D(regs[34]), .Q(n200) );
  AOI220 U1443 ( .A(n844), .B(regs[355]), .C(n75), .D(regs[291]), .Q(n212) );
  AOI220 U1444 ( .A(n844), .B(regs[611]), .C(n75), .D(regs[547]), .Q(n218) );
  AOI220 U1445 ( .A(n66), .B(regs[868]), .C(n843), .D(regs[804]), .Q(n230) );
  AOI220 U1446 ( .A(n844), .B(regs[356]), .C(n75), .D(regs[292]), .Q(n234) );
  AOI220 U1447 ( .A(n66), .B(regs[872]), .C(n843), .D(regs[808]), .Q(n318) );
  AOI220 U1448 ( .A(n844), .B(regs[874]), .C(n75), .D(regs[810]), .Q(n362) );
  AOI220 U1449 ( .A(n844), .B(regs[363]), .C(n75), .D(regs[299]), .Q(n388) );
  AOI220 U1450 ( .A(n844), .B(regs[619]), .C(n75), .D(regs[555]), .Q(n394) );
  AOI220 U1451 ( .A(n840), .B(regs[235]), .C(n67), .D(regs[171]), .Q(n400) );
  AOI220 U1452 ( .A(n66), .B(regs[107]), .C(n843), .D(regs[43]), .Q(n398) );
  AOI220 U1453 ( .A(n840), .B(regs[492]), .C(n67), .D(regs[428]), .Q(n412) );
  AOI220 U1454 ( .A(n66), .B(regs[364]), .C(n843), .D(regs[300]), .Q(n410) );
  AOI220 U1455 ( .A(n840), .B(regs[1005]), .C(n67), .D(regs[941]), .Q(n430) );
  AOI220 U1456 ( .A(n66), .B(regs[365]), .C(n843), .D(regs[301]), .Q(n432) );
  AOI220 U1457 ( .A(n846), .B(regs[589]), .C(n845), .D(regs[525]), .Q(n437) );
  AOI220 U1458 ( .A(n846), .B(regs[590]), .C(n845), .D(regs[526]), .Q(n459) );
  AOI220 U1459 ( .A(n846), .B(regs[591]), .C(n845), .D(regs[527]), .Q(n481) );
  AOI220 U1460 ( .A(n840), .B(regs[239]), .C(n67), .D(regs[175]), .Q(n488) );
  AOI220 U1461 ( .A(n840), .B(regs[240]), .C(n67), .D(regs[176]), .Q(n510) );
  AOI220 U1462 ( .A(n846), .B(regs[849]), .C(n845), .D(regs[785]), .Q(n515) );
  AOI220 U1463 ( .A(n840), .B(regs[497]), .C(n67), .D(regs[433]), .Q(n522) );
  AOI220 U1464 ( .A(n846), .B(regs[850]), .C(n845), .D(regs[786]), .Q(n537) );
  AOI220 U1465 ( .A(n66), .B(regs[372]), .C(n843), .D(regs[308]), .Q(n586) );
  AOI220 U1466 ( .A(n846), .B(regs[340]), .C(n110), .D(regs[276]), .Q(n585) );
  AOI220 U1467 ( .A(n66), .B(regs[116]), .C(n843), .D(regs[52]), .Q(n596) );
  AOI220 U1468 ( .A(n846), .B(regs[84]), .C(n110), .D(regs[20]), .Q(n595) );
  AOI220 U1469 ( .A(n66), .B(regs[885]), .C(n843), .D(regs[821]), .Q(n604) );
  AOI220 U1470 ( .A(n846), .B(regs[853]), .C(n110), .D(regs[789]), .Q(n603) );
  AOI220 U1471 ( .A(n846), .B(regs[341]), .C(n110), .D(regs[277]), .Q(n607) );
  AOI220 U1472 ( .A(n66), .B(regs[117]), .C(n843), .D(regs[53]), .Q(n618) );
  AOI220 U1473 ( .A(n846), .B(regs[85]), .C(n110), .D(regs[21]), .Q(n617) );
  AOI220 U1474 ( .A(n66), .B(regs[886]), .C(n843), .D(regs[822]), .Q(n626) );
  AOI220 U1475 ( .A(n846), .B(regs[854]), .C(n110), .D(regs[790]), .Q(n625) );
  AOI220 U1476 ( .A(n66), .B(regs[890]), .C(n843), .D(regs[826]), .Q(n714) );
  AOI220 U1477 ( .A(n66), .B(regs[378]), .C(n843), .D(regs[314]), .Q(n718) );
  AOI220 U1478 ( .A(n66), .B(regs[634]), .C(n843), .D(regs[570]), .Q(n724) );
  AOI220 U1479 ( .A(n66), .B(regs[122]), .C(n843), .D(regs[58]), .Q(n728) );
  AOI220 U1480 ( .A(n66), .B(regs[891]), .C(n843), .D(regs[827]), .Q(n736) );
  AOI220 U1481 ( .A(n66), .B(regs[379]), .C(n843), .D(regs[315]), .Q(n740) );
  AOI220 U1482 ( .A(n66), .B(regs[635]), .C(n843), .D(regs[571]), .Q(n746) );
  AOI220 U1483 ( .A(n66), .B(regs[123]), .C(n843), .D(regs[59]), .Q(n750) );
  AOI220 U1484 ( .A(n66), .B(regs[892]), .C(n843), .D(regs[828]), .Q(n758) );
  AOI220 U1485 ( .A(regs[864]), .B(n1566), .C(regs[800]), .D(n1565), .Q(n862)
         );
  AOI220 U1486 ( .A(regs[352]), .B(n1566), .C(regs[288]), .D(n1565), .Q(n867)
         );
  AOI220 U1487 ( .A(regs[576]), .B(n68), .C(regs[512]), .D(n114), .Q(n873) );
  AOI220 U1488 ( .A(regs[224]), .B(n1562), .C(regs[160]), .D(n74), .Q(n880) );
  AOI220 U1489 ( .A(regs[192]), .B(n1564), .C(regs[128]), .D(n73), .Q(n879) );
  AOI220 U1490 ( .A(regs[993]), .B(n1562), .C(regs[929]), .D(n74), .Q(n888) );
  AOI220 U1491 ( .A(regs[961]), .B(n1564), .C(regs[897]), .D(n73), .Q(n887) );
  AOI220 U1492 ( .A(regs[865]), .B(n1566), .C(regs[801]), .D(n1565), .Q(n886)
         );
  AOI220 U1493 ( .A(regs[833]), .B(n68), .C(regs[769]), .D(n114), .Q(n885) );
  AOI220 U1494 ( .A(regs[705]), .B(n113), .C(regs[641]), .D(n73), .Q(n897) );
  AOI220 U1495 ( .A(regs[577]), .B(n68), .C(regs[513]), .D(n114), .Q(n895) );
  AOI220 U1496 ( .A(regs[193]), .B(n113), .C(regs[129]), .D(n73), .Q(n901) );
  AOI220 U1497 ( .A(regs[65]), .B(n68), .C(regs[1]), .D(n114), .Q(n899) );
  AOI220 U1498 ( .A(regs[962]), .B(n113), .C(regs[898]), .D(n73), .Q(n909) );
  AOI220 U1499 ( .A(regs[450]), .B(n113), .C(regs[386]), .D(n73), .Q(n913) );
  AOI220 U1500 ( .A(regs[322]), .B(n68), .C(regs[258]), .D(n1567), .Q(n911) );
  AOI220 U1501 ( .A(regs[578]), .B(n68), .C(regs[514]), .D(n114), .Q(n917) );
  AOI220 U1502 ( .A(regs[194]), .B(n113), .C(regs[130]), .D(n73), .Q(n923) );
  AOI220 U1503 ( .A(regs[66]), .B(n68), .C(regs[2]), .D(n114), .Q(n921) );
  AOI220 U1504 ( .A(regs[995]), .B(n112), .C(regs[931]), .D(n1561), .Q(n932)
         );
  AOI220 U1505 ( .A(regs[835]), .B(n68), .C(regs[771]), .D(n114), .Q(n929) );
  AOI220 U1506 ( .A(regs[483]), .B(n112), .C(regs[419]), .D(n1561), .Q(n936)
         );
  AOI220 U1507 ( .A(regs[451]), .B(n113), .C(regs[387]), .D(n1563), .Q(n935)
         );
  AOI220 U1508 ( .A(regs[323]), .B(n68), .C(regs[259]), .D(n1567), .Q(n933) );
  AOI220 U1509 ( .A(regs[579]), .B(n68), .C(regs[515]), .D(n114), .Q(n939) );
  AOI220 U1510 ( .A(regs[227]), .B(n1562), .C(regs[163]), .D(n74), .Q(n946) );
  AOI220 U1511 ( .A(regs[195]), .B(n113), .C(regs[131]), .D(n73), .Q(n945) );
  AOI220 U1512 ( .A(regs[67]), .B(n68), .C(regs[3]), .D(n114), .Q(n943) );
  AOI220 U1513 ( .A(regs[964]), .B(n113), .C(regs[900]), .D(n73), .Q(n953) );
  AOI220 U1514 ( .A(regs[452]), .B(n113), .C(regs[388]), .D(n73), .Q(n957) );
  AOI220 U1515 ( .A(regs[324]), .B(n68), .C(regs[260]), .D(n114), .Q(n955) );
  AOI220 U1516 ( .A(regs[580]), .B(n68), .C(regs[516]), .D(n114), .Q(n961) );
  AOI220 U1517 ( .A(regs[196]), .B(n113), .C(regs[132]), .D(n73), .Q(n967) );
  AOI220 U1518 ( .A(regs[68]), .B(n68), .C(regs[4]), .D(n1567), .Q(n965) );
  AOI220 U1519 ( .A(regs[965]), .B(n113), .C(regs[901]), .D(n1563), .Q(n975)
         );
  AOI220 U1520 ( .A(regs[453]), .B(n113), .C(regs[389]), .D(n73), .Q(n979) );
  AOI220 U1521 ( .A(regs[325]), .B(n68), .C(regs[261]), .D(n1567), .Q(n977) );
  AOI220 U1522 ( .A(regs[69]), .B(n68), .C(regs[5]), .D(n1567), .Q(n987) );
  AOI220 U1523 ( .A(regs[838]), .B(n68), .C(regs[774]), .D(n1567), .Q(n995) );
  AOI220 U1524 ( .A(regs[454]), .B(n113), .C(regs[390]), .D(n73), .Q(n1001) );
  AOI220 U1525 ( .A(regs[326]), .B(n68), .C(regs[262]), .D(n1567), .Q(n999) );
  AOI220 U1526 ( .A(regs[362]), .B(n1566), .C(regs[298]), .D(n1565), .Q(n1088)
         );
  AOI220 U1527 ( .A(regs[234]), .B(n112), .C(regs[170]), .D(n1561), .Q(n1100)
         );
  AOI220 U1528 ( .A(regs[491]), .B(n112), .C(regs[427]), .D(n1561), .Q(n1112)
         );
  AOI220 U1529 ( .A(regs[1004]), .B(n112), .C(regs[940]), .D(n1561), .Q(n1130)
         );
  AOI220 U1530 ( .A(regs[972]), .B(n113), .C(regs[908]), .D(n1563), .Q(n1129)
         );
  AOI220 U1531 ( .A(regs[460]), .B(n113), .C(regs[396]), .D(n73), .Q(n1133) );
  AOI220 U1532 ( .A(regs[332]), .B(n1568), .C(regs[268]), .D(n114), .Q(n1131)
         );
  AOI220 U1533 ( .A(regs[716]), .B(n113), .C(regs[652]), .D(n73), .Q(n1139) );
  AOI220 U1534 ( .A(regs[204]), .B(n113), .C(regs[140]), .D(n73), .Q(n1143) );
  AOI220 U1535 ( .A(regs[973]), .B(n113), .C(regs[909]), .D(n73), .Q(n1151) );
  AOI220 U1536 ( .A(regs[461]), .B(n113), .C(regs[397]), .D(n73), .Q(n1155) );
  AOI220 U1537 ( .A(regs[717]), .B(n113), .C(regs[653]), .D(n73), .Q(n1161) );
  AOI220 U1538 ( .A(regs[205]), .B(n113), .C(regs[141]), .D(n73), .Q(n1165) );
  AOI220 U1539 ( .A(regs[974]), .B(n1564), .C(regs[910]), .D(n73), .Q(n1173)
         );
  AOI220 U1540 ( .A(regs[878]), .B(n1566), .C(regs[814]), .D(n72), .Q(n1172)
         );
  AOI220 U1541 ( .A(regs[846]), .B(n68), .C(regs[782]), .D(n114), .Q(n1171) );
  AOI220 U1542 ( .A(regs[494]), .B(n1562), .C(regs[430]), .D(n74), .Q(n1178)
         );
  AOI220 U1543 ( .A(regs[462]), .B(n113), .C(regs[398]), .D(n73), .Q(n1177) );
  AOI220 U1544 ( .A(regs[334]), .B(n68), .C(regs[270]), .D(n114), .Q(n1175) );
  AOI220 U1545 ( .A(regs[590]), .B(n68), .C(regs[526]), .D(n114), .Q(n1181) );
  AOI220 U1546 ( .A(regs[206]), .B(n113), .C(regs[142]), .D(n73), .Q(n1187) );
  AOI220 U1547 ( .A(regs[975]), .B(n1564), .C(regs[911]), .D(n73), .Q(n1195)
         );
  AOI220 U1548 ( .A(regs[847]), .B(n68), .C(regs[783]), .D(n1567), .Q(n1193)
         );
  AOI220 U1549 ( .A(regs[463]), .B(n1564), .C(regs[399]), .D(n73), .Q(n1199)
         );
  AOI220 U1550 ( .A(regs[367]), .B(n1566), .C(regs[303]), .D(n72), .Q(n1198)
         );
  AOI220 U1551 ( .A(regs[335]), .B(n68), .C(regs[271]), .D(n114), .Q(n1197) );
  AOI220 U1552 ( .A(regs[719]), .B(n113), .C(regs[655]), .D(n73), .Q(n1205) );
  AOI220 U1553 ( .A(regs[591]), .B(n68), .C(regs[527]), .D(n114), .Q(n1203) );
  AOI220 U1554 ( .A(regs[496]), .B(n112), .C(regs[432]), .D(n1561), .Q(n1222)
         );
  AOI220 U1555 ( .A(regs[464]), .B(n1564), .C(regs[400]), .D(n1563), .Q(n1221)
         );
  AOI220 U1556 ( .A(regs[368]), .B(n1566), .C(regs[304]), .D(n1565), .Q(n1220)
         );
  AOI220 U1557 ( .A(regs[336]), .B(n1568), .C(regs[272]), .D(n114), .Q(n1219)
         );
  AOI220 U1558 ( .A(regs[592]), .B(n68), .C(regs[528]), .D(n114), .Q(n1225) );
  AOI220 U1559 ( .A(regs[497]), .B(n112), .C(regs[433]), .D(n1561), .Q(n1244)
         );
  AOI220 U1560 ( .A(regs[465]), .B(n1564), .C(regs[401]), .D(n1563), .Q(n1243)
         );
  AOI220 U1561 ( .A(regs[337]), .B(n1568), .C(regs[273]), .D(n114), .Q(n1241)
         );
  AOI220 U1562 ( .A(regs[113]), .B(n1566), .C(regs[49]), .D(n1565), .Q(n1252)
         );
  AOI220 U1563 ( .A(regs[1010]), .B(n112), .C(regs[946]), .D(n1561), .Q(n1262)
         );
  AOI220 U1564 ( .A(regs[978]), .B(n113), .C(regs[914]), .D(n1563), .Q(n1261)
         );
  AOI220 U1565 ( .A(regs[882]), .B(n69), .C(regs[818]), .D(n1565), .Q(n1260)
         );
  AOI220 U1566 ( .A(regs[498]), .B(n112), .C(regs[434]), .D(n1561), .Q(n1266)
         );
  AOI220 U1567 ( .A(regs[466]), .B(n113), .C(regs[402]), .D(n1563), .Q(n1265)
         );
  AOI220 U1568 ( .A(regs[370]), .B(n69), .C(regs[306]), .D(n1565), .Q(n1264)
         );
  AOI220 U1569 ( .A(regs[242]), .B(n112), .C(regs[178]), .D(n1561), .Q(n1276)
         );
  AOI220 U1570 ( .A(regs[210]), .B(n113), .C(regs[146]), .D(n1563), .Q(n1275)
         );
  AOI220 U1571 ( .A(regs[114]), .B(n1566), .C(regs[50]), .D(n1565), .Q(n1274)
         );
  AOI220 U1572 ( .A(regs[371]), .B(n1566), .C(regs[307]), .D(n72), .Q(n1286)
         );
  AOI220 U1573 ( .A(regs[468]), .B(n113), .C(regs[404]), .D(n73), .Q(n1309) );
  AOI220 U1574 ( .A(regs[340]), .B(n68), .C(regs[276]), .D(n114), .Q(n1307) );
  AOI220 U1575 ( .A(regs[373]), .B(n1566), .C(regs[309]), .D(n72), .Q(n1330)
         );
  AOI220 U1576 ( .A(regs[341]), .B(n68), .C(regs[277]), .D(n114), .Q(n1329) );
  AOI220 U1577 ( .A(regs[725]), .B(n113), .C(regs[661]), .D(n73), .Q(n1337) );
  AOI220 U1578 ( .A(regs[117]), .B(n1566), .C(regs[53]), .D(n72), .Q(n1340) );
  AOI220 U1579 ( .A(regs[85]), .B(n1568), .C(regs[21]), .D(n114), .Q(n1339) );
  AOI220 U1580 ( .A(regs[982]), .B(n113), .C(regs[918]), .D(n73), .Q(n1349) );
  AOI220 U1581 ( .A(regs[854]), .B(n1568), .C(regs[790]), .D(n114), .Q(n1347)
         );
  AOI220 U1582 ( .A(regs[374]), .B(n1566), .C(regs[310]), .D(n72), .Q(n1352)
         );
  AOI220 U1583 ( .A(regs[342]), .B(n68), .C(regs[278]), .D(n114), .Q(n1351) );
  AOI220 U1584 ( .A(regs[726]), .B(n113), .C(regs[662]), .D(n73), .Q(n1359) );
  AOI220 U1585 ( .A(regs[1016]), .B(n112), .C(regs[952]), .D(n1561), .Q(n1394)
         );
  AOI220 U1586 ( .A(regs[376]), .B(n69), .C(regs[312]), .D(n1565), .Q(n1396)
         );
  AOI220 U1587 ( .A(regs[505]), .B(n112), .C(regs[441]), .D(n1561), .Q(n1420)
         );
  AOI220 U1588 ( .A(regs[249]), .B(n112), .C(regs[185]), .D(n1561), .Q(n1430)
         );
  AOI220 U1589 ( .A(regs[474]), .B(n113), .C(regs[410]), .D(n1563), .Q(n1441)
         );
  AOI220 U1590 ( .A(regs[346]), .B(n68), .C(regs[282]), .D(n114), .Q(n1439) );
  AOI220 U1591 ( .A(regs[730]), .B(n113), .C(regs[666]), .D(n1563), .Q(n1447)
         );
  AOI220 U1592 ( .A(regs[602]), .B(n68), .C(regs[538]), .D(n114), .Q(n1445) );
  AOI220 U1593 ( .A(regs[218]), .B(n113), .C(regs[154]), .D(n1563), .Q(n1451)
         );
  AOI220 U1594 ( .A(regs[90]), .B(n68), .C(regs[26]), .D(n114), .Q(n1449) );
  AOI220 U1595 ( .A(regs[859]), .B(n68), .C(regs[795]), .D(n114), .Q(n1457) );
  AOI220 U1596 ( .A(regs[475]), .B(n113), .C(regs[411]), .D(n1563), .Q(n1463)
         );
  AOI220 U1597 ( .A(regs[347]), .B(n68), .C(regs[283]), .D(n114), .Q(n1461) );
  AOI220 U1598 ( .A(regs[603]), .B(n68), .C(regs[539]), .D(n114), .Q(n1467) );
  AOI220 U1599 ( .A(regs[219]), .B(n113), .C(regs[155]), .D(n1563), .Q(n1473)
         );
  AOI220 U1600 ( .A(regs[91]), .B(n68), .C(regs[27]), .D(n114), .Q(n1471) );
  AOI220 U1601 ( .A(regs[988]), .B(n1564), .C(regs[924]), .D(n73), .Q(n1481)
         );
  AOI220 U1602 ( .A(regs[732]), .B(n113), .C(regs[668]), .D(n73), .Q(n1491) );
  AOI220 U1603 ( .A(regs[220]), .B(n1564), .C(regs[156]), .D(n73), .Q(n1495)
         );
  AOI220 U1604 ( .A(regs[1021]), .B(n1562), .C(regs[957]), .D(n74), .Q(n1504)
         );
  AOI220 U1605 ( .A(regs[989]), .B(n113), .C(regs[925]), .D(n73), .Q(n1503) );
  AOI220 U1606 ( .A(regs[509]), .B(n1562), .C(regs[445]), .D(n74), .Q(n1508)
         );
  AOI220 U1607 ( .A(regs[477]), .B(n113), .C(regs[413]), .D(n73), .Q(n1507) );
  AOI220 U1608 ( .A(regs[253]), .B(n1562), .C(regs[189]), .D(n74), .Q(n1518)
         );
  AOI220 U1609 ( .A(regs[221]), .B(n113), .C(regs[157]), .D(n73), .Q(n1517) );
  AOI220 U1610 ( .A(regs[990]), .B(n1564), .C(regs[926]), .D(n73), .Q(n1525)
         );
  AOI220 U1611 ( .A(regs[894]), .B(n69), .C(regs[830]), .D(n1565), .Q(n1524)
         );
  AOI220 U1612 ( .A(regs[510]), .B(n112), .C(regs[446]), .D(n1561), .Q(n1530)
         );
  AOI220 U1613 ( .A(regs[478]), .B(n113), .C(regs[414]), .D(n1563), .Q(n1529)
         );
  AOI220 U1614 ( .A(regs[382]), .B(n69), .C(regs[318]), .D(n1565), .Q(n1528)
         );
  AOI220 U1615 ( .A(regs[734]), .B(n113), .C(regs[670]), .D(n73), .Q(n1535) );
  AOI220 U1616 ( .A(regs[222]), .B(n113), .C(regs[158]), .D(n73), .Q(n1539) );
  AOI220 U1617 ( .A(regs[1023]), .B(n1562), .C(regs[959]), .D(n74), .Q(n1548)
         );
  AOI220 U1618 ( .A(regs[991]), .B(n113), .C(regs[927]), .D(n73), .Q(n1547) );
  AOI220 U1619 ( .A(regs[895]), .B(n69), .C(regs[831]), .D(n1565), .Q(n1546)
         );
  AOI220 U1620 ( .A(regs[479]), .B(n113), .C(regs[415]), .D(n73), .Q(n1551) );
  AOI220 U1621 ( .A(regs[383]), .B(n1566), .C(regs[319]), .D(n1565), .Q(n1550)
         );
  AOI220 U1622 ( .A(regs[223]), .B(n113), .C(regs[159]), .D(n73), .Q(n1571) );
  AOI220 U1623 ( .A(regs[95]), .B(n1568), .C(regs[31]), .D(n114), .Q(n1569) );
endmodule


module decode ( i_clk, i_nrst, i_addr_pc4, i_con_Wregwrite, i_data_Wregwrite, 
        i_addr_Wregwrite, i_addr_Erd, i_addr_Mrd, i_con_Eregwrite, 
        i_con_Mregwrite, i_addr_rtM, i_addr_rtW, i_con_memreadM, 
        i_con_memreadW, i_data_Wmemout, o_data_rs, o_data_rt, o_addr_rd, 
        o_addr_rt, o_data_jr, o_con_jump, o_addr_pc4, o_addr_branch, 
        o_con_Ealuop, o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite, 
        o_con_Malupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall, 
        o_con_Ebop, o_data_signext, o_con_Efamux, o_con_Efbmux, o_data_Fmemout, 
        o_addr_jump_31_, o_addr_jump_30_, o_addr_jump_29_, o_addr_jump_28_, 
        o_addr_jump_27_, o_addr_jump_26_, o_addr_jump_25_, o_addr_jump_24_, 
        o_addr_jump_23_, o_addr_jump_22_, o_addr_jump_21_, o_addr_jump_20_, 
        o_addr_jump_19_, o_addr_jump_17_, o_addr_jump_16_, o_addr_jump_15_, 
        o_addr_jump_14_, o_addr_jump_13_, o_addr_jump_12_, o_addr_jump_11_, 
        o_addr_jump_10_, o_addr_jump_9_, o_addr_jump_8_, o_addr_jump_7_, 
        o_addr_jump_6_, o_addr_jump_5_, o_addr_jump_4_, o_addr_jump_3_, 
        o_addr_jump_2_, o_addr_jump_1_, o_addr_jump_0_, i_data_instr_31_, 
        i_data_instr_30_, i_data_instr_29_, i_data_instr_28_, i_data_instr_27_, 
        i_data_instr_26_, i_data_instr_25_, i_data_instr_24_, i_data_instr_23_, 
        i_data_instr_22_, i_data_instr_21_, i_data_instr_20_, i_data_instr_19_, 
        i_data_instr_18_, i_data_instr_17_, i_data_instr_14_, i_data_instr_13_, 
        i_data_instr_12_, i_data_instr_11_, i_data_instr_10_, i_data_instr_9_, 
        i_data_instr_8_, i_data_instr_7_, i_data_instr_6_, i_data_instr_5_, 
        i_data_instr_4_, i_data_instr_3_, i_data_instr_2_, i_data_instr_1_, 
        i_data_instr_0_, o_addr_jump_18_, i_data_instr_16_, 
        i_data_instr_15__BAR, o_con_Ealusrc_BAR );
  input [31:0] i_addr_pc4;
  input [31:0] i_data_Wregwrite;
  input [4:0] i_addr_Wregwrite;
  input [4:0] i_addr_Erd;
  input [4:0] i_addr_Mrd;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  input [31:0] i_data_Wmemout;
  output [31:0] o_data_rs;
  output [31:0] o_data_rt;
  output [4:0] o_addr_rd;
  output [4:0] o_addr_rt;
  output [31:0] o_data_jr;
  output [1:0] o_con_jump;
  output [31:0] o_addr_pc4;
  output [31:0] o_addr_branch;
  output [5:0] o_con_Ealuop;
  output [2:0] o_con_Ebop;
  output [31:0] o_data_signext;
  output [2:0] o_con_Efamux;
  output [2:0] o_con_Efbmux;
  output [31:0] o_data_Fmemout;
  input i_clk, i_nrst, i_con_Wregwrite, i_con_Eregwrite, i_con_Mregwrite,
         i_con_memreadM, i_con_memreadW, i_data_instr_31_, i_data_instr_30_,
         i_data_instr_29_, i_data_instr_28_, i_data_instr_27_,
         i_data_instr_26_, i_data_instr_25_, i_data_instr_24_,
         i_data_instr_23_, i_data_instr_22_, i_data_instr_21_,
         i_data_instr_20_, i_data_instr_19_, i_data_instr_18_,
         i_data_instr_17_, i_data_instr_14_, i_data_instr_13_,
         i_data_instr_12_, i_data_instr_11_, i_data_instr_10_, i_data_instr_9_,
         i_data_instr_8_, i_data_instr_7_, i_data_instr_6_, i_data_instr_5_,
         i_data_instr_4_, i_data_instr_3_, i_data_instr_2_, i_data_instr_1_,
         i_data_instr_0_, i_data_instr_16_, i_data_instr_15__BAR;
  output o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8,
         o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall, o_addr_jump_31_,
         o_addr_jump_30_, o_addr_jump_29_, o_addr_jump_28_, o_addr_jump_27_,
         o_addr_jump_26_, o_addr_jump_25_, o_addr_jump_24_, o_addr_jump_23_,
         o_addr_jump_22_, o_addr_jump_21_, o_addr_jump_20_, o_addr_jump_19_,
         o_addr_jump_17_, o_addr_jump_16_, o_addr_jump_15_, o_addr_jump_14_,
         o_addr_jump_13_, o_addr_jump_12_, o_addr_jump_11_, o_addr_jump_10_,
         o_addr_jump_9_, o_addr_jump_8_, o_addr_jump_7_, o_addr_jump_6_,
         o_addr_jump_5_, o_addr_jump_4_, o_addr_jump_3_, o_addr_jump_2_,
         o_addr_jump_1_, o_addr_jump_0_, o_addr_jump_18_, o_con_Ealusrc_BAR;
  wire   i_data_instr_25_, i_data_instr_24_, i_data_instr_23_,
         i_data_instr_22_, i_data_instr_21_, i_data_instr_20_,
         i_data_instr_19_, i_data_instr_18_, i_data_instr_17_,
         i_data_instr_16_, i_data_instr_14_, i_data_instr_13_,
         i_data_instr_12_, i_data_instr_11_, i_data_instr_10_, i_data_instr_9_,
         i_data_instr_8_, i_data_instr_7_, i_data_instr_6_, i_data_instr_5_,
         i_data_instr_4_, i_data_instr_3_, i_data_instr_2_, i_data_instr_1_,
         i_data_instr_0_, n177, control_o_con_alusrc, control_o_con_regdst,
         jbcon_o_con_aluPC4, control_o_con_memread, control_o_con_memwrite,
         control_o_con_memtoreg, control_o_con_regwrite,
         pcadd_o_addr_pcbranchE_31_, pcadd_o_addr_pcbranchE_30_,
         pcadd_o_addr_pcbranchE_29_, pcadd_o_addr_pcbranchE_28_,
         pcadd_o_addr_pcbranchE_27_, pcadd_o_addr_pcbranchE_26_,
         pcadd_o_addr_pcbranchE_25_, pcadd_o_addr_pcbranchE_24_,
         pcadd_o_addr_pcbranchE_23_, pcadd_o_addr_pcbranchE_22_,
         pcadd_o_addr_pcbranchE_21_, pcadd_o_addr_pcbranchE_20_,
         pcadd_o_addr_pcbranchE_19_, pcadd_o_addr_pcbranchE_18_,
         pcadd_o_addr_pcbranchE_17_, pcadd_o_addr_pcbranchE_16_,
         pcadd_o_addr_pcbranchE_15_, pcadd_o_addr_pcbranchE_14_,
         pcadd_o_addr_pcbranchE_13_, pcadd_o_addr_pcbranchE_12_,
         pcadd_o_addr_pcbranchE_11_, pcadd_o_addr_pcbranchE_10_,
         pcadd_o_addr_pcbranchE_9_, pcadd_o_addr_pcbranchE_8_,
         pcadd_o_addr_pcbranchE_7_, pcadd_o_addr_pcbranchE_6_,
         pcadd_o_addr_pcbranchE_5_, pcadd_o_addr_pcbranchE_4_,
         pcadd_o_addr_pcbranchE_3_, pcadd_o_addr_pcbranchE_2_, n1, n6,
         add_x_16_n30, add_x_16_n29, add_x_16_n28, add_x_16_n27, add_x_16_n26,
         add_x_16_n25, add_x_16_n24, add_x_16_n23, add_x_16_n22, add_x_16_n21,
         add_x_16_n20, add_x_16_n19, add_x_16_n18, add_x_16_n17, add_x_16_n16,
         add_x_16_n15, add_x_16_n14, add_x_16_n13, add_x_16_n12, add_x_16_n11,
         add_x_16_n10, add_x_16_n9, add_x_16_n8, add_x_16_n7, add_x_16_n6,
         add_x_16_n5, add_x_16_n4, add_x_16_n3, add_x_16_n2, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176;
  wire   [31:0] regbank_o_data_Rt;
  wire   [5:0] control_o_con_aluop;
  wire   [2:0] for_o_con_fa;
  wire   [2:0] for_o_con_fb;
  wire   [1:0] jbcon_o_con_bop;
  assign o_addr_jump_31_ = i_addr_pc4[31];
  assign o_addr_jump_30_ = i_addr_pc4[30];
  assign o_addr_jump_29_ = i_addr_pc4[29];
  assign o_addr_jump_28_ = i_addr_pc4[28];
  assign o_addr_branch[1] = o_addr_pc4[1];
  assign o_addr_branch[0] = o_addr_pc4[0];
  assign o_addr_jump_27_ = i_data_instr_25_;
  assign o_addr_jump_26_ = i_data_instr_24_;
  assign o_addr_jump_25_ = i_data_instr_23_;
  assign o_addr_jump_24_ = i_data_instr_22_;
  assign o_addr_jump_23_ = i_data_instr_21_;
  assign o_addr_jump_22_ = i_data_instr_20_;
  assign o_addr_jump_21_ = i_data_instr_19_;
  assign o_addr_jump_20_ = i_data_instr_18_;
  assign o_addr_jump_19_ = i_data_instr_17_;
  assign o_addr_jump_18_ = i_data_instr_16_;
  assign o_addr_jump_16_ = i_data_instr_14_;
  assign o_addr_jump_15_ = i_data_instr_13_;
  assign o_addr_jump_14_ = i_data_instr_12_;
  assign o_addr_jump_13_ = i_data_instr_11_;
  assign o_addr_jump_12_ = i_data_instr_10_;
  assign o_addr_jump_11_ = i_data_instr_9_;
  assign o_addr_jump_10_ = i_data_instr_8_;
  assign o_addr_jump_9_ = i_data_instr_7_;
  assign o_addr_jump_8_ = i_data_instr_6_;
  assign o_addr_jump_7_ = i_data_instr_5_;
  assign o_addr_jump_6_ = i_data_instr_4_;
  assign o_addr_jump_5_ = i_data_instr_3_;
  assign o_addr_jump_4_ = i_data_instr_2_;
  assign o_addr_jump_3_ = i_data_instr_1_;
  assign o_addr_jump_2_ = i_data_instr_0_;

  D_register_bank u_regbank ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_addr_Rs({
        i_data_instr_25_, i_data_instr_24_, i_data_instr_23_, i_data_instr_22_, 
        i_data_instr_21_}), .i_con_RegWr(i_con_Wregwrite), .i_addr_Rd(
        i_addr_Wregwrite), .i_data_Rd(i_data_Wregwrite), .o_data_Rs(o_data_jr), 
        .o_data_Rt(regbank_o_data_Rt), .i_addr_Rt_4_(i_data_instr_20_), 
        .i_addr_Rt_3_(i_data_instr_19_), .i_addr_Rt_2_(i_data_instr_18_), 
        .i_addr_Rt_1_(i_data_instr_17_), .i_addr_Rt_0_(i_data_instr_16_) );
  DFC1 pipe_bop_reg_2_ ( .D(n6), .C(i_clk), .RN(i_nrst), .Q(o_con_Ebop[2]) );
  DFC1 pipe_bop_reg_1_ ( .D(jbcon_o_con_bop[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[1]) );
  DFC1 pipe_bop_reg_0_ ( .D(jbcon_o_con_bop[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[0]) );
  DFC1 pipe_data_rs_reg_31_ ( .D(o_data_jr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[31]) );
  DFC1 pipe_data_rs_reg_30_ ( .D(o_data_jr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[30]) );
  DFC1 pipe_data_rs_reg_29_ ( .D(o_data_jr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[29]) );
  DFC1 pipe_data_rs_reg_28_ ( .D(o_data_jr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[28]) );
  DFC1 pipe_data_rs_reg_27_ ( .D(o_data_jr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[27]) );
  DFC1 pipe_data_rs_reg_26_ ( .D(o_data_jr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[26]) );
  DFC1 pipe_data_rs_reg_25_ ( .D(o_data_jr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[25]) );
  DFC1 pipe_data_rs_reg_24_ ( .D(o_data_jr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[24]) );
  DFC1 pipe_data_rs_reg_23_ ( .D(o_data_jr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[23]) );
  DFC1 pipe_data_rs_reg_22_ ( .D(o_data_jr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[22]) );
  DFC1 pipe_data_rs_reg_21_ ( .D(o_data_jr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[21]) );
  DFC1 pipe_data_rs_reg_20_ ( .D(o_data_jr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[20]) );
  DFC1 pipe_data_rs_reg_19_ ( .D(o_data_jr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[19]) );
  DFC1 pipe_data_rs_reg_18_ ( .D(o_data_jr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[18]) );
  DFC1 pipe_data_rs_reg_17_ ( .D(o_data_jr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[17]) );
  DFC1 pipe_data_rs_reg_16_ ( .D(o_data_jr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[16]) );
  DFC1 pipe_data_rs_reg_15_ ( .D(o_data_jr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[15]) );
  DFC1 pipe_data_rs_reg_14_ ( .D(o_data_jr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[14]) );
  DFC1 pipe_data_rs_reg_13_ ( .D(o_data_jr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[13]) );
  DFC1 pipe_data_rs_reg_12_ ( .D(o_data_jr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[12]) );
  DFC1 pipe_data_rs_reg_11_ ( .D(o_data_jr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[11]) );
  DFC1 pipe_data_rs_reg_10_ ( .D(o_data_jr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[10]) );
  DFC1 pipe_data_rs_reg_9_ ( .D(o_data_jr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[9]) );
  DFC1 pipe_data_rs_reg_8_ ( .D(o_data_jr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[8]) );
  DFC1 pipe_data_rs_reg_7_ ( .D(o_data_jr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[7]) );
  DFC1 pipe_data_rs_reg_6_ ( .D(o_data_jr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[6]) );
  DFC1 pipe_data_rs_reg_5_ ( .D(o_data_jr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[5]) );
  DFC1 pipe_data_rs_reg_4_ ( .D(o_data_jr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[4]) );
  DFC1 pipe_data_rs_reg_3_ ( .D(o_data_jr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[3]) );
  DFC1 pipe_data_rs_reg_2_ ( .D(o_data_jr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[2]) );
  DFC1 pipe_data_rs_reg_1_ ( .D(o_data_jr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[1]) );
  DFC1 pipe_data_rs_reg_0_ ( .D(o_data_jr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[0]) );
  DFC1 pipe_data_rt_reg_31_ ( .D(regbank_o_data_Rt[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[31]) );
  DFC1 pipe_data_rt_reg_30_ ( .D(regbank_o_data_Rt[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC1 pipe_data_rt_reg_29_ ( .D(regbank_o_data_Rt[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[29]) );
  DFC1 pipe_data_rt_reg_28_ ( .D(regbank_o_data_Rt[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28]) );
  DFC1 pipe_data_rt_reg_27_ ( .D(regbank_o_data_Rt[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27]) );
  DFC1 pipe_data_rt_reg_26_ ( .D(regbank_o_data_Rt[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26]) );
  DFC1 pipe_data_rt_reg_25_ ( .D(regbank_o_data_Rt[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25]) );
  DFC1 pipe_data_rt_reg_24_ ( .D(regbank_o_data_Rt[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24]) );
  DFC1 pipe_data_rt_reg_23_ ( .D(regbank_o_data_Rt[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23]) );
  DFC1 pipe_data_rt_reg_22_ ( .D(regbank_o_data_Rt[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC1 pipe_data_rt_reg_21_ ( .D(regbank_o_data_Rt[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21]) );
  DFC1 pipe_data_rt_reg_20_ ( .D(regbank_o_data_Rt[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20]) );
  DFC1 pipe_data_rt_reg_19_ ( .D(regbank_o_data_Rt[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19]) );
  DFC1 pipe_data_rt_reg_18_ ( .D(regbank_o_data_Rt[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18]) );
  DFC1 pipe_data_rt_reg_17_ ( .D(regbank_o_data_Rt[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17]) );
  DFC1 pipe_data_rt_reg_16_ ( .D(regbank_o_data_Rt[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC1 pipe_data_rt_reg_15_ ( .D(regbank_o_data_Rt[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15]) );
  DFC1 pipe_data_rt_reg_14_ ( .D(regbank_o_data_Rt[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14]) );
  DFC1 pipe_data_rt_reg_13_ ( .D(regbank_o_data_Rt[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC1 pipe_data_rt_reg_12_ ( .D(regbank_o_data_Rt[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12]) );
  DFC1 pipe_data_rt_reg_11_ ( .D(regbank_o_data_Rt[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11]) );
  DFC1 pipe_data_rt_reg_10_ ( .D(regbank_o_data_Rt[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC1 pipe_data_rt_reg_9_ ( .D(regbank_o_data_Rt[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[9]) );
  DFC1 pipe_data_rt_reg_8_ ( .D(regbank_o_data_Rt[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[8]) );
  DFC1 pipe_data_rt_reg_7_ ( .D(regbank_o_data_Rt[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[7]) );
  DFC1 pipe_data_rt_reg_6_ ( .D(regbank_o_data_Rt[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[6]) );
  DFC1 pipe_data_rt_reg_5_ ( .D(regbank_o_data_Rt[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[5]) );
  DFC1 pipe_data_rt_reg_4_ ( .D(regbank_o_data_Rt[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[4]) );
  DFC1 pipe_data_rt_reg_3_ ( .D(regbank_o_data_Rt[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[3]) );
  DFC1 pipe_data_rt_reg_2_ ( .D(regbank_o_data_Rt[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[2]) );
  DFC1 pipe_data_rt_reg_1_ ( .D(regbank_o_data_Rt[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[1]) );
  DFC1 pipe_data_rt_reg_0_ ( .D(regbank_o_data_Rt[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[0]) );
  DFC1 pipe_addr_rt_reg_4_ ( .D(i_data_instr_20_), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[4]) );
  DFC1 pipe_addr_rt_reg_3_ ( .D(i_data_instr_19_), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[3]) );
  DFC1 pipe_addr_rt_reg_2_ ( .D(i_data_instr_18_), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[2]) );
  DFC1 pipe_addr_rt_reg_1_ ( .D(i_data_instr_17_), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[1]) );
  DFC1 pipe_addr_rt_reg_0_ ( .D(i_data_instr_16_), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[0]) );
  DFC1 pipe_addr_pc4_reg_31_ ( .D(i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC1 pipe_addr_pc4_reg_30_ ( .D(i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC1 pipe_addr_pc4_reg_29_ ( .D(i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC1 pipe_addr_pc4_reg_28_ ( .D(i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC1 pipe_addr_pc4_reg_27_ ( .D(i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC1 pipe_addr_pc4_reg_26_ ( .D(i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC1 pipe_addr_pc4_reg_25_ ( .D(i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC1 pipe_addr_pc4_reg_24_ ( .D(i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC1 pipe_addr_pc4_reg_23_ ( .D(i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC1 pipe_addr_pc4_reg_22_ ( .D(i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC1 pipe_addr_pc4_reg_21_ ( .D(i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC1 pipe_addr_pc4_reg_20_ ( .D(i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC1 pipe_addr_pc4_reg_19_ ( .D(i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC1 pipe_addr_pc4_reg_18_ ( .D(i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC1 pipe_addr_pc4_reg_17_ ( .D(i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC1 pipe_addr_pc4_reg_16_ ( .D(i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC1 pipe_addr_pc4_reg_15_ ( .D(i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC1 pipe_addr_pc4_reg_14_ ( .D(i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC1 pipe_addr_pc4_reg_13_ ( .D(i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC1 pipe_addr_pc4_reg_12_ ( .D(i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC1 pipe_addr_pc4_reg_11_ ( .D(i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC1 pipe_addr_pc4_reg_10_ ( .D(i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC1 pipe_addr_pc4_reg_9_ ( .D(i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC1 pipe_addr_pc4_reg_8_ ( .D(i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC1 pipe_addr_pc4_reg_7_ ( .D(i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC1 pipe_addr_pc4_reg_6_ ( .D(i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC1 pipe_addr_pc4_reg_5_ ( .D(i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC1 pipe_addr_pc4_reg_4_ ( .D(i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC1 pipe_addr_pc4_reg_3_ ( .D(i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC1 pipe_addr_pc4_reg_2_ ( .D(i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC1 pipe_con_Ealuop_reg_5_ ( .D(control_o_con_aluop[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[5]) );
  DFC1 pipe_con_Ealuop_reg_4_ ( .D(control_o_con_aluop[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[4]) );
  DFC1 pipe_con_Ealuop_reg_3_ ( .D(control_o_con_aluop[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[3]) );
  DFC1 pipe_con_Ealuop_reg_2_ ( .D(control_o_con_aluop[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[2]) );
  DFC1 pipe_con_Ealuop_reg_1_ ( .D(control_o_con_aluop[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[1]) );
  DFC1 pipe_con_Ealuop_reg_0_ ( .D(control_o_con_aluop[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[0]) );
  DFC1 pipe_con_Ealusrc_reg ( .D(control_o_con_alusrc), .C(i_clk), .RN(i_nrst), 
        .QN(o_con_Ealusrc_BAR) );
  DFC1 pipe_con_Eregdst_reg ( .D(control_o_con_regdst), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Eregdst) );
  DFC1 pipe_con_MaluPC4_reg ( .D(jbcon_o_con_aluPC4), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Malupc8) );
  DFC1 pipe_con_Mmemread_reg ( .D(control_o_con_memread), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemread) );
  DFC1 pipe_con_Mmemwrite_reg ( .D(control_o_con_memwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemwrite) );
  DFC1 pipe_con_Wmemtoreg_reg ( .D(control_o_con_memtoreg), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wmemtoreg) );
  DFC1 pipe_con_Wregwrite_reg ( .D(control_o_con_regwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wregwrite) );
  DFC1 pipe_signext_o_data_immD_reg_15_ ( .D(o_addr_jump_17_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[15]) );
  DFC1 pipe_signext_o_data_immD_reg_14_ ( .D(i_data_instr_14_), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[14]) );
  DFC1 pipe_signext_o_data_immD_reg_13_ ( .D(i_data_instr_13_), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[13]) );
  DFC1 pipe_signext_o_data_immD_reg_12_ ( .D(i_data_instr_12_), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[12]) );
  DFC1 pipe_signext_o_data_immD_reg_11_ ( .D(i_data_instr_11_), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[11]) );
  DFC1 pipe_signext_o_data_immD_reg_9_ ( .D(i_data_instr_9_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[9]) );
  DFC1 pipe_signext_o_data_immD_reg_7_ ( .D(i_data_instr_7_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[7]) );
  DFC1 pipe_signext_o_data_immD_reg_6_ ( .D(i_data_instr_6_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[6]) );
  DFC1 pipe_signext_o_data_immD_reg_5_ ( .D(i_data_instr_5_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[5]) );
  DFC1 pipe_signext_o_data_immD_reg_4_ ( .D(i_data_instr_4_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[4]) );
  DFC1 pipe_signext_o_data_immD_reg_3_ ( .D(i_data_instr_3_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[3]) );
  DFC1 pipe_signext_o_data_immD_reg_2_ ( .D(i_data_instr_2_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[2]) );
  DFC1 pipe_signext_o_data_immD_reg_1_ ( .D(i_data_instr_1_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[1]) );
  DFC1 pipe_signext_o_data_immD_reg_0_ ( .D(i_data_instr_0_), .C(i_clk), .RN(
        i_nrst), .Q(o_data_signext[0]) );
  DFC1 pipe_con_Efamux_reg_2_ ( .D(for_o_con_fa[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[2]) );
  DFC1 pipe_con_Efamux_reg_1_ ( .D(for_o_con_fa[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[1]) );
  DFC1 pipe_FWmemout_reg_31_ ( .D(i_data_Wmemout[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[31]) );
  DFC1 pipe_FWmemout_reg_30_ ( .D(i_data_Wmemout[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[30]) );
  DFC1 pipe_FWmemout_reg_29_ ( .D(i_data_Wmemout[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[29]) );
  DFC1 pipe_FWmemout_reg_28_ ( .D(i_data_Wmemout[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[28]) );
  DFC1 pipe_FWmemout_reg_27_ ( .D(i_data_Wmemout[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[27]) );
  DFC1 pipe_FWmemout_reg_26_ ( .D(i_data_Wmemout[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[26]) );
  DFC1 pipe_FWmemout_reg_25_ ( .D(i_data_Wmemout[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[25]) );
  DFC1 pipe_FWmemout_reg_24_ ( .D(i_data_Wmemout[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[24]) );
  DFC1 pipe_FWmemout_reg_23_ ( .D(i_data_Wmemout[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[23]) );
  DFC1 pipe_FWmemout_reg_22_ ( .D(i_data_Wmemout[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[22]) );
  DFC1 pipe_FWmemout_reg_21_ ( .D(i_data_Wmemout[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[21]) );
  DFC1 pipe_FWmemout_reg_20_ ( .D(i_data_Wmemout[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[20]) );
  DFC1 pipe_FWmemout_reg_19_ ( .D(i_data_Wmemout[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[19]) );
  DFC1 pipe_FWmemout_reg_18_ ( .D(i_data_Wmemout[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[18]) );
  DFC1 pipe_FWmemout_reg_17_ ( .D(i_data_Wmemout[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[17]) );
  DFC1 pipe_FWmemout_reg_16_ ( .D(i_data_Wmemout[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[16]) );
  DFC1 pipe_FWmemout_reg_15_ ( .D(i_data_Wmemout[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[15]) );
  DFC1 pipe_FWmemout_reg_14_ ( .D(i_data_Wmemout[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[14]) );
  DFC1 pipe_FWmemout_reg_13_ ( .D(i_data_Wmemout[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[13]) );
  DFC1 pipe_FWmemout_reg_12_ ( .D(i_data_Wmemout[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[12]) );
  DFC1 pipe_FWmemout_reg_11_ ( .D(i_data_Wmemout[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[11]) );
  DFC1 pipe_FWmemout_reg_10_ ( .D(i_data_Wmemout[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[10]) );
  DFC1 pipe_FWmemout_reg_9_ ( .D(i_data_Wmemout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[9]) );
  DFC1 pipe_FWmemout_reg_8_ ( .D(i_data_Wmemout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[8]) );
  DFC1 pipe_FWmemout_reg_7_ ( .D(i_data_Wmemout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[7]) );
  DFC1 pipe_FWmemout_reg_6_ ( .D(i_data_Wmemout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[6]) );
  DFC1 pipe_FWmemout_reg_5_ ( .D(i_data_Wmemout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[5]) );
  DFC1 pipe_FWmemout_reg_4_ ( .D(i_data_Wmemout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[4]) );
  DFC1 pipe_FWmemout_reg_3_ ( .D(i_data_Wmemout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[3]) );
  DFC1 pipe_FWmemout_reg_2_ ( .D(i_data_Wmemout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[2]) );
  DFC1 pipe_FWmemout_reg_1_ ( .D(i_data_Wmemout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[1]) );
  DFC1 pipe_FWmemout_reg_0_ ( .D(i_data_Wmemout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[0]) );
  DFC1 pipe_addr_branch_reg_31_ ( .D(pcadd_o_addr_pcbranchE_31_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[31]) );
  DFC1 pipe_addr_branch_reg_30_ ( .D(pcadd_o_addr_pcbranchE_30_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[30]) );
  DFC1 pipe_addr_branch_reg_29_ ( .D(pcadd_o_addr_pcbranchE_29_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[29]) );
  DFC1 pipe_addr_branch_reg_28_ ( .D(pcadd_o_addr_pcbranchE_28_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[28]) );
  DFC1 pipe_addr_branch_reg_27_ ( .D(pcadd_o_addr_pcbranchE_27_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[27]) );
  DFC1 pipe_addr_branch_reg_26_ ( .D(pcadd_o_addr_pcbranchE_26_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[26]) );
  DFC1 pipe_addr_branch_reg_25_ ( .D(pcadd_o_addr_pcbranchE_25_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[25]) );
  DFC1 pipe_addr_branch_reg_24_ ( .D(pcadd_o_addr_pcbranchE_24_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[24]) );
  DFC1 pipe_addr_branch_reg_23_ ( .D(pcadd_o_addr_pcbranchE_23_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[23]) );
  DFC1 pipe_addr_branch_reg_22_ ( .D(pcadd_o_addr_pcbranchE_22_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[22]) );
  DFC1 pipe_addr_branch_reg_21_ ( .D(pcadd_o_addr_pcbranchE_21_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[21]) );
  DFC1 pipe_addr_branch_reg_20_ ( .D(pcadd_o_addr_pcbranchE_20_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[20]) );
  DFC1 pipe_addr_branch_reg_19_ ( .D(pcadd_o_addr_pcbranchE_19_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[19]) );
  DFC1 pipe_addr_branch_reg_18_ ( .D(pcadd_o_addr_pcbranchE_18_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[18]) );
  DFC1 pipe_addr_branch_reg_17_ ( .D(pcadd_o_addr_pcbranchE_17_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[17]) );
  DFC1 pipe_addr_branch_reg_16_ ( .D(pcadd_o_addr_pcbranchE_16_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[16]) );
  DFC1 pipe_addr_branch_reg_15_ ( .D(pcadd_o_addr_pcbranchE_15_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[15]) );
  DFC1 pipe_addr_branch_reg_14_ ( .D(pcadd_o_addr_pcbranchE_14_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[14]) );
  DFC1 pipe_addr_branch_reg_13_ ( .D(pcadd_o_addr_pcbranchE_13_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[13]) );
  DFC1 pipe_addr_branch_reg_12_ ( .D(pcadd_o_addr_pcbranchE_12_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[12]) );
  DFC1 pipe_addr_branch_reg_11_ ( .D(pcadd_o_addr_pcbranchE_11_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[11]) );
  DFC1 pipe_addr_branch_reg_10_ ( .D(pcadd_o_addr_pcbranchE_10_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[10]) );
  DFC1 pipe_addr_branch_reg_9_ ( .D(pcadd_o_addr_pcbranchE_9_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[9]) );
  DFC1 pipe_addr_branch_reg_8_ ( .D(pcadd_o_addr_pcbranchE_8_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[8]) );
  DFC1 pipe_addr_branch_reg_7_ ( .D(pcadd_o_addr_pcbranchE_7_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[7]) );
  DFC1 pipe_addr_branch_reg_6_ ( .D(pcadd_o_addr_pcbranchE_6_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[6]) );
  DFC1 pipe_addr_branch_reg_5_ ( .D(pcadd_o_addr_pcbranchE_5_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[5]) );
  DFC1 pipe_addr_branch_reg_4_ ( .D(pcadd_o_addr_pcbranchE_4_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[4]) );
  DFC1 pipe_addr_branch_reg_3_ ( .D(pcadd_o_addr_pcbranchE_3_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[3]) );
  DFC1 pipe_addr_branch_reg_2_ ( .D(pcadd_o_addr_pcbranchE_2_), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[2]) );
  DFC1 pipe_addr_branch_reg_1_ ( .D(i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_pc4[1]) );
  DFC1 pipe_addr_branch_reg_0_ ( .D(i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_pc4[0]) );
  DFC3 pipe_signext_o_data_immD_reg_16_ ( .D(n1), .C(i_clk), .RN(i_nrst), .Q(
        o_data_signext[16]) );
  DFC3 pipe_con_Efbmux_reg_1_ ( .D(for_o_con_fb[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[1]) );
  DFC3 pipe_signext_o_data_immD_reg_10_ ( .D(i_data_instr_10_), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[10]) );
  DFC3 pipe_con_Efbmux_reg_2_ ( .D(for_o_con_fb[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[2]) );
  DFC3 pipe_con_Efbmux_reg_0_ ( .D(for_o_con_fb[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[0]) );
  DFC3 pipe_con_Efamux_reg_0_ ( .D(for_o_con_fa[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[0]) );
  DFC3 pipe_signext_o_data_immD_reg_8_ ( .D(i_data_instr_8_), .C(i_clk), .RN(
        i_nrst), .Q(n177) );
  ADD22 add_x_16_U31 ( .A(i_addr_pc4[2]), .B(i_data_instr_0_), .CO(
        add_x_16_n30), .S(pcadd_o_addr_pcbranchE_2_) );
  INV3 U3 ( .A(i_data_instr_15__BAR), .Q(o_addr_jump_17_) );
  XOR30 U4 ( .A(add_x_16_n17), .B(i_data_instr_14_), .C(i_addr_pc4[16]), .Q(
        pcadd_o_addr_pcbranchE_16_) );
  XOR30 U5 ( .A(add_x_16_n18), .B(i_data_instr_13_), .C(i_addr_pc4[15]), .Q(
        pcadd_o_addr_pcbranchE_15_) );
  XOR30 U6 ( .A(add_x_16_n26), .B(i_data_instr_5_), .C(i_addr_pc4[7]), .Q(
        pcadd_o_addr_pcbranchE_7_) );
  NAND20 U7 ( .A(o_addr_jump_17_), .B(i_addr_pc4[30]), .Q(n58) );
  NAND21 U8 ( .A(o_addr_jump_17_), .B(i_addr_pc4[27]), .Q(n55) );
  INV2 U9 ( .A(i_data_instr_28_), .Q(n172) );
  NAND31 U10 ( .A(n60), .B(n59), .C(n58), .Q(add_x_16_n2) );
  NAND22 U11 ( .A(add_x_16_n3), .B(i_addr_pc4[30]), .Q(n59) );
  NAND22 U12 ( .A(add_x_16_n6), .B(i_addr_pc4[27]), .Q(n56) );
  NAND22 U13 ( .A(add_x_16_n16), .B(o_addr_jump_17_), .Q(n54) );
  NAND22 U14 ( .A(add_x_16_n16), .B(i_addr_pc4[17]), .Q(n53) );
  INV2 U15 ( .A(control_o_con_aluop[4]), .Q(n175) );
  AOI210 U16 ( .A(n76), .B(n75), .C(control_o_con_aluop[1]), .Q(n77) );
  OAI210 U17 ( .A(i_addr_Erd[2]), .B(n90), .C(n106), .Q(n91) );
  INV2 U18 ( .A(n75), .Q(n74) );
  AOI311 U19 ( .A(i_data_instr_3_), .B(n165), .C(n164), .D(i_data_instr_26_), 
        .Q(n166) );
  INV0 U20 ( .A(o_addr_jump_17_), .Q(n174) );
  INV1 U21 ( .A(i_data_instr_19_), .Q(n143) );
  INV1 U22 ( .A(i_data_instr_18_), .Q(n148) );
  NAND21 U23 ( .A(i_data_instr_3_), .B(i_addr_pc4[5]), .Q(n46) );
  XOR21 U24 ( .A(add_x_16_n3), .B(n61), .Q(pcadd_o_addr_pcbranchE_30_) );
  NAND22 U25 ( .A(add_x_16_n3), .B(o_addr_jump_17_), .Q(n60) );
  NAND33 U26 ( .A(n57), .B(n56), .C(n55), .Q(add_x_16_n5) );
  NAND22 U27 ( .A(add_x_16_n6), .B(o_addr_jump_17_), .Q(n57) );
  NAND33 U28 ( .A(n54), .B(n53), .C(n52), .Q(add_x_16_n15) );
  NAND33 U29 ( .A(n45), .B(n44), .C(n43), .Q(add_x_16_n16) );
  NAND22 U30 ( .A(add_x_16_n18), .B(i_data_instr_13_), .Q(n51) );
  NAND22 U31 ( .A(add_x_16_n18), .B(i_addr_pc4[15]), .Q(n50) );
  NAND31 U32 ( .A(n42), .B(n41), .C(n40), .Q(add_x_16_n25) );
  OAI210 U33 ( .A(n67), .B(n66), .C(n175), .Q(control_o_con_aluop[3]) );
  OAI2111 U34 ( .A(i_addr_Mrd[1]), .B(n100), .C(n99), .D(n98), .Q(n114) );
  NAND33 U35 ( .A(n39), .B(n38), .C(n37), .Q(add_x_16_n26) );
  OAI211 U36 ( .A(n157), .B(n156), .C(n155), .Q(for_o_con_fb[2]) );
  INV2 U37 ( .A(n118), .Q(n119) );
  INV2 U38 ( .A(n156), .Q(n154) );
  NAND22 U39 ( .A(add_x_16_n27), .B(i_addr_pc4[6]), .Q(n38) );
  NAND31 U40 ( .A(n48), .B(n47), .C(n46), .Q(add_x_16_n27) );
  INV2 U41 ( .A(n115), .Q(n117) );
  INV2 U42 ( .A(n77), .Q(control_o_con_regwrite) );
  INV1 U43 ( .A(control_o_con_aluop[5]), .Q(n65) );
  NAND30 U44 ( .A(control_o_con_aluop[0]), .B(n172), .C(n158), .Q(n63) );
  NAND31 U45 ( .A(i_con_memreadW), .B(n125), .C(n124), .Q(n156) );
  NAND41 U46 ( .A(i_con_memreadM), .B(n150), .C(n151), .D(n149), .Q(n155) );
  NAND31 U47 ( .A(i_con_Eregwrite), .B(n135), .C(n134), .Q(n153) );
  AOI310 U48 ( .A(n173), .B(n172), .C(n171), .D(control_o_con_memtoreg), .Q(
        n176) );
  OAI220 U49 ( .A(n162), .B(n161), .C(n160), .D(n159), .Q(jbcon_o_con_bop[1])
         );
  NAND41 U50 ( .A(i_con_memreadW), .B(n84), .C(n83), .D(n101), .Q(n116) );
  OAI212 U51 ( .A(i_data_instr_28_), .B(n167), .C(n169), .Q(o_con_jump[0]) );
  NAND21 U52 ( .A(i_con_Eregwrite), .B(n89), .Q(n94) );
  OAI211 U53 ( .A(n160), .B(n69), .C(n68), .Q(control_o_con_memread) );
  NOR21 U54 ( .A(i_data_instr_27_), .B(n166), .Q(n167) );
  NAND21 U55 ( .A(i_data_instr_26_), .B(n64), .Q(n69) );
  IMUX20 U56 ( .A(n142), .B(i_data_instr_17_), .S(i_addr_Erd[1]), .Q(n132) );
  NOR20 U57 ( .A(n73), .B(n168), .Q(control_o_con_regdst) );
  IMUX20 U58 ( .A(n140), .B(i_data_instr_16_), .S(i_addr_Erd[0]), .Q(n130) );
  INV2 U59 ( .A(n64), .Q(n66) );
  OAI212 U60 ( .A(i_data_instr_28_), .B(n163), .C(n169), .Q(o_con_ifstall) );
  NAND41 U61 ( .A(i_con_memreadM), .B(n109), .C(n108), .D(n107), .Q(n110) );
  INV2 U62 ( .A(n101), .Q(n113) );
  NOR21 U63 ( .A(i_data_instr_27_), .B(n158), .Q(n163) );
  INV1 U64 ( .A(n169), .Q(n73) );
  NAND22 U65 ( .A(o_addr_jump_17_), .B(i_addr_pc4[17]), .Q(n52) );
  INV2 U66 ( .A(i_data_instr_16_), .Q(n140) );
  NOR21 U67 ( .A(n72), .B(i_data_instr_30_), .Q(n173) );
  INV2 U68 ( .A(i_data_instr_17_), .Q(n142) );
  INV1 U69 ( .A(i_data_instr_25_), .Q(n104) );
  INV2 U70 ( .A(i_data_instr_29_), .Q(n72) );
  INV1 U71 ( .A(i_con_Mregwrite), .Q(n126) );
  NOR21 U72 ( .A(i_data_instr_26_), .B(i_data_instr_27_), .Q(n67) );
  INV2 U73 ( .A(i_data_instr_5_), .Q(n164) );
  NAND22 U74 ( .A(i_data_instr_14_), .B(i_addr_pc4[16]), .Q(n43) );
  NAND22 U75 ( .A(i_data_instr_13_), .B(i_addr_pc4[15]), .Q(n49) );
  INV1 U76 ( .A(i_data_instr_31_), .Q(n71) );
  NAND21 U77 ( .A(i_data_instr_5_), .B(i_addr_pc4[7]), .Q(n40) );
  INV1 U78 ( .A(i_data_instr_20_), .Q(n141) );
  INV3 U79 ( .A(i_data_instr_26_), .Q(n158) );
  NOR31 U80 ( .A(i_data_instr_30_), .B(i_data_instr_29_), .C(i_data_instr_31_), 
        .Q(n169) );
  INV2 U81 ( .A(i_data_instr_27_), .Q(n160) );
  BUF6 U82 ( .A(n177), .Q(o_data_signext[8]) );
  XOR31 U83 ( .A(i_addr_pc4[31]), .B(o_addr_jump_17_), .C(add_x_16_n2), .Q(
        pcadd_o_addr_pcbranchE_31_) );
  XOR31 U84 ( .A(add_x_16_n27), .B(i_data_instr_4_), .C(i_addr_pc4[6]), .Q(
        pcadd_o_addr_pcbranchE_6_) );
  XOR31 U85 ( .A(add_x_16_n28), .B(i_data_instr_3_), .C(i_addr_pc4[5]), .Q(
        pcadd_o_addr_pcbranchE_5_) );
  NAND22 U86 ( .A(add_x_16_n28), .B(i_addr_pc4[5]), .Q(n47) );
  NAND22 U87 ( .A(add_x_16_n26), .B(i_data_instr_5_), .Q(n42) );
  NAND22 U88 ( .A(add_x_16_n26), .B(i_addr_pc4[7]), .Q(n41) );
  NAND33 U89 ( .A(n51), .B(n50), .C(n49), .Q(add_x_16_n17) );
  NAND22 U90 ( .A(add_x_16_n17), .B(i_data_instr_14_), .Q(n45) );
  NAND22 U91 ( .A(add_x_16_n17), .B(i_addr_pc4[16]), .Q(n44) );
  NAND22 U92 ( .A(add_x_16_n28), .B(i_data_instr_3_), .Q(n48) );
  NAND22 U93 ( .A(add_x_16_n27), .B(i_data_instr_4_), .Q(n39) );
  NAND22 U94 ( .A(i_data_instr_4_), .B(i_addr_pc4[6]), .Q(n37) );
  ADD32 U95 ( .A(i_addr_pc4[13]), .B(i_data_instr_11_), .CI(add_x_16_n20), 
        .CO(add_x_16_n19), .S(pcadd_o_addr_pcbranchE_13_) );
  ADD32 U96 ( .A(i_addr_pc4[14]), .B(i_data_instr_12_), .CI(add_x_16_n19), 
        .CO(add_x_16_n18), .S(pcadd_o_addr_pcbranchE_14_) );
  ADD32 U97 ( .A(o_addr_jump_17_), .B(i_addr_pc4[28]), .CI(add_x_16_n5), .CO(
        add_x_16_n4), .S(pcadd_o_addr_pcbranchE_28_) );
  ADD32 U98 ( .A(o_addr_jump_17_), .B(i_addr_pc4[29]), .CI(add_x_16_n4), .CO(
        add_x_16_n3), .S(pcadd_o_addr_pcbranchE_29_) );
  ADD32 U99 ( .A(o_addr_jump_17_), .B(i_addr_pc4[21]), .CI(add_x_16_n12), .CO(
        add_x_16_n11), .S(pcadd_o_addr_pcbranchE_21_) );
  ADD32 U100 ( .A(o_addr_jump_17_), .B(i_addr_pc4[22]), .CI(add_x_16_n11), 
        .CO(add_x_16_n10), .S(pcadd_o_addr_pcbranchE_22_) );
  ADD32 U101 ( .A(i_addr_pc4[3]), .B(i_data_instr_1_), .CI(add_x_16_n30), .CO(
        add_x_16_n29), .S(pcadd_o_addr_pcbranchE_3_) );
  ADD32 U102 ( .A(i_addr_pc4[4]), .B(i_data_instr_2_), .CI(add_x_16_n29), .CO(
        add_x_16_n28), .S(pcadd_o_addr_pcbranchE_4_) );
  ADD32 U103 ( .A(o_addr_jump_17_), .B(i_addr_pc4[19]), .CI(add_x_16_n14), 
        .CO(add_x_16_n13), .S(pcadd_o_addr_pcbranchE_19_) );
  ADD32 U104 ( .A(o_addr_jump_17_), .B(i_addr_pc4[20]), .CI(add_x_16_n13), 
        .CO(add_x_16_n12), .S(pcadd_o_addr_pcbranchE_20_) );
  ADD32 U105 ( .A(o_addr_jump_17_), .B(i_addr_pc4[26]), .CI(add_x_16_n7), .CO(
        add_x_16_n6), .S(pcadd_o_addr_pcbranchE_26_) );
  ADD32 U106 ( .A(i_addr_pc4[11]), .B(i_data_instr_9_), .CI(add_x_16_n22), 
        .CO(add_x_16_n21), .S(pcadd_o_addr_pcbranchE_11_) );
  ADD32 U107 ( .A(i_addr_pc4[12]), .B(i_data_instr_10_), .CI(add_x_16_n21), 
        .CO(add_x_16_n20), .S(pcadd_o_addr_pcbranchE_12_) );
  ADD32 U108 ( .A(o_addr_jump_17_), .B(i_addr_pc4[23]), .CI(add_x_16_n10), 
        .CO(add_x_16_n9), .S(pcadd_o_addr_pcbranchE_23_) );
  ADD32 U109 ( .A(o_addr_jump_17_), .B(i_addr_pc4[18]), .CI(add_x_16_n15), 
        .CO(add_x_16_n14), .S(pcadd_o_addr_pcbranchE_18_) );
  ADD32 U110 ( .A(o_addr_jump_17_), .B(i_addr_pc4[24]), .CI(add_x_16_n9), .CO(
        add_x_16_n8), .S(pcadd_o_addr_pcbranchE_24_) );
  ADD32 U111 ( .A(o_addr_jump_17_), .B(i_addr_pc4[25]), .CI(add_x_16_n8), .CO(
        add_x_16_n7), .S(pcadd_o_addr_pcbranchE_25_) );
  ADD32 U112 ( .A(i_addr_pc4[9]), .B(i_data_instr_7_), .CI(add_x_16_n24), .CO(
        add_x_16_n23), .S(pcadd_o_addr_pcbranchE_9_) );
  ADD32 U113 ( .A(i_addr_pc4[10]), .B(i_data_instr_8_), .CI(add_x_16_n23), 
        .CO(add_x_16_n22), .S(pcadd_o_addr_pcbranchE_10_) );
  ADD32 U114 ( .A(i_addr_pc4[8]), .B(i_data_instr_6_), .CI(add_x_16_n25), .CO(
        add_x_16_n24), .S(pcadd_o_addr_pcbranchE_8_) );
  XOR31 U115 ( .A(add_x_16_n16), .B(o_addr_jump_17_), .C(i_addr_pc4[17]), .Q(
        pcadd_o_addr_pcbranchE_17_) );
  XOR31 U116 ( .A(add_x_16_n6), .B(o_addr_jump_17_), .C(i_addr_pc4[27]), .Q(
        pcadd_o_addr_pcbranchE_27_) );
  XOR20 U117 ( .A(o_addr_jump_17_), .B(i_addr_pc4[30]), .Q(n61) );
  NAND20 U118 ( .A(n169), .B(n163), .Q(n161) );
  OAI210 U119 ( .A(n163), .B(n66), .C(n65), .Q(control_o_con_aluop[2]) );
  NOR40 U120 ( .A(n113), .B(n112), .C(n111), .D(n110), .Q(n115) );
  NOR30 U121 ( .A(n158), .B(n160), .C(i_data_instr_28_), .Q(n75) );
  NOR40 U122 ( .A(n96), .B(n95), .C(n94), .D(n93), .Q(n118) );
  INV0 U123 ( .A(i_data_instr_21_), .Q(n103) );
  INV0 U124 ( .A(i_data_instr_22_), .Q(n102) );
  NOR21 U125 ( .A(n71), .B(n70), .Q(control_o_con_memwrite) );
  NOR21 U126 ( .A(n74), .B(n73), .Q(jbcon_o_con_aluPC4) );
  AOI211 U127 ( .A(n156), .B(n152), .C(n157), .Q(for_o_con_fb[0]) );
  NAND41 U128 ( .A(n138), .B(n153), .C(n137), .D(n136), .Q(n152) );
  NOR31 U129 ( .A(n154), .B(n157), .C(n153), .Q(for_o_con_fb[1]) );
  NAND22 U130 ( .A(n139), .B(n141), .Q(n151) );
  NOR21 U131 ( .A(n119), .B(for_o_con_fa[2]), .Q(for_o_con_fa[1]) );
  NAND22 U132 ( .A(n117), .B(n116), .Q(for_o_con_fa[2]) );
  AOI211 U133 ( .A(n176), .B(n175), .C(n174), .Q(n1) );
  AOI211 U134 ( .A(n63), .B(n69), .C(n160), .Q(control_o_con_aluop[4]) );
  AOI211 U135 ( .A(n116), .B(n114), .C(n115), .Q(for_o_con_fa[0]) );
  OAI2111 U136 ( .A(i_addr_Erd[2]), .B(n106), .C(n92), .D(n91), .Q(n93) );
  IMUX20 U137 ( .A(i_data_instr_21_), .B(n103), .S(i_addr_Erd[0]), .Q(n92) );
  NAND22 U138 ( .A(n82), .B(n104), .Q(n101) );
  INV0 U139 ( .A(i_data_instr_24_), .Q(n105) );
  NAND22 U140 ( .A(n67), .B(n172), .Q(n168) );
  NAND22 U141 ( .A(n151), .B(n155), .Q(n157) );
  INV3 U142 ( .A(n173), .Q(n70) );
  INV0 U143 ( .A(i_data_instr_23_), .Q(n106) );
  NAND22 U144 ( .A(n169), .B(n168), .Q(o_con_jump[1]) );
  NOR20 U145 ( .A(i_data_instr_31_), .B(n70), .Q(control_o_con_aluop[0]) );
  NOR40 U146 ( .A(i_data_instr_30_), .B(i_data_instr_31_), .C(n72), .D(n172), 
        .Q(n64) );
  NAND20 U147 ( .A(i_data_instr_26_), .B(i_data_instr_27_), .Q(n171) );
  NOR40 U148 ( .A(i_data_instr_28_), .B(i_data_instr_31_), .C(n171), .D(n70), 
        .Q(control_o_con_aluop[5]) );
  AOI2110 U149 ( .A(n72), .B(n168), .C(i_data_instr_30_), .D(i_data_instr_31_), 
        .Q(control_o_con_aluop[1]) );
  OAI310 U150 ( .A(i_data_instr_30_), .B(n74), .C(n71), .D(n70), .Q(
        control_o_con_alusrc) );
  NOR20 U151 ( .A(i_data_instr_30_), .B(i_data_instr_29_), .Q(n76) );
  NAND30 U152 ( .A(n76), .B(n75), .C(i_data_instr_31_), .Q(n68) );
  AOI2110 U153 ( .A(n72), .B(n74), .C(i_data_instr_30_), .D(n71), .Q(
        control_o_con_memtoreg) );
  IMUX20 U154 ( .A(n102), .B(i_data_instr_22_), .S(i_addr_rtW[1]), .Q(n81) );
  IMUX20 U155 ( .A(n103), .B(i_data_instr_21_), .S(i_addr_rtW[0]), .Q(n80) );
  IMUX20 U156 ( .A(n104), .B(i_data_instr_25_), .S(i_addr_rtW[4]), .Q(n79) );
  IMUX20 U157 ( .A(n106), .B(i_data_instr_23_), .S(i_addr_rtW[2]), .Q(n78) );
  NOR40 U158 ( .A(n81), .B(n80), .C(n79), .D(n78), .Q(n84) );
  IMUX20 U159 ( .A(i_data_instr_24_), .B(n105), .S(i_addr_rtW[3]), .Q(n83) );
  NOR40 U160 ( .A(i_data_instr_21_), .B(i_data_instr_23_), .C(i_data_instr_24_), .D(i_data_instr_22_), .Q(n82) );
  NOR40 U161 ( .A(i_addr_Mrd[0]), .B(i_addr_Mrd[4]), .C(i_addr_Mrd[2]), .D(
        i_addr_Mrd[3]), .Q(n85) );
  NOR20 U162 ( .A(i_data_instr_22_), .B(n85), .Q(n100) );
  IMUX20 U163 ( .A(n103), .B(i_data_instr_21_), .S(i_addr_Mrd[0]), .Q(n88) );
  IMUX20 U164 ( .A(n105), .B(i_data_instr_24_), .S(i_addr_Mrd[3]), .Q(n87) );
  IMUX20 U165 ( .A(n104), .B(i_data_instr_25_), .S(i_addr_Mrd[4]), .Q(n86) );
  NOR40 U166 ( .A(n88), .B(n87), .C(n86), .D(n126), .Q(n99) );
  IMUX20 U167 ( .A(n102), .B(i_data_instr_22_), .S(i_addr_Erd[1]), .Q(n96) );
  IMUX20 U168 ( .A(n105), .B(i_data_instr_24_), .S(i_addr_Erd[3]), .Q(n95) );
  IMUX20 U169 ( .A(i_data_instr_25_), .B(n104), .S(i_addr_Erd[4]), .Q(n89) );
  NOR40 U170 ( .A(i_addr_Erd[1]), .B(i_addr_Erd[3]), .C(i_addr_Erd[0]), .D(
        i_data_instr_25_), .Q(n90) );
  IMUX20 U171 ( .A(n106), .B(i_data_instr_23_), .S(i_addr_Mrd[2]), .Q(n97) );
  AOI2110 U172 ( .A(i_addr_Mrd[1]), .B(n102), .C(n118), .D(n97), .Q(n98) );
  IMUX20 U173 ( .A(n102), .B(i_data_instr_22_), .S(i_addr_rtM[1]), .Q(n112) );
  IMUX20 U174 ( .A(n103), .B(i_data_instr_21_), .S(i_addr_rtM[0]), .Q(n111) );
  IMUX20 U175 ( .A(i_data_instr_25_), .B(n104), .S(i_addr_rtM[4]), .Q(n109) );
  IMUX20 U176 ( .A(i_data_instr_24_), .B(n105), .S(i_addr_rtM[3]), .Q(n108) );
  IMUX20 U177 ( .A(i_data_instr_23_), .B(n106), .S(i_addr_rtM[2]), .Q(n107) );
  IMUX20 U178 ( .A(n143), .B(i_data_instr_19_), .S(i_addr_rtW[3]), .Q(n123) );
  IMUX20 U179 ( .A(n148), .B(i_data_instr_18_), .S(i_addr_rtW[2]), .Q(n122) );
  IMUX20 U180 ( .A(n142), .B(i_data_instr_17_), .S(i_addr_rtW[1]), .Q(n121) );
  IMUX20 U181 ( .A(n140), .B(i_data_instr_16_), .S(i_addr_rtW[0]), .Q(n120) );
  NOR40 U182 ( .A(n123), .B(n122), .C(n121), .D(n120), .Q(n125) );
  IMUX20 U183 ( .A(i_data_instr_20_), .B(n141), .S(i_addr_rtW[4]), .Q(n124) );
  IMUX20 U184 ( .A(n141), .B(i_data_instr_20_), .S(i_addr_Mrd[4]), .Q(n129) );
  IMUX20 U185 ( .A(n148), .B(i_data_instr_18_), .S(i_addr_Mrd[2]), .Q(n128) );
  IMUX20 U186 ( .A(n143), .B(i_data_instr_19_), .S(i_addr_Mrd[3]), .Q(n127) );
  NOR40 U187 ( .A(n129), .B(n128), .C(n127), .D(n126), .Q(n138) );
  IMUX20 U188 ( .A(n141), .B(i_data_instr_20_), .S(i_addr_Erd[4]), .Q(n133) );
  IMUX20 U189 ( .A(n143), .B(i_data_instr_19_), .S(i_addr_Erd[3]), .Q(n131) );
  NOR40 U190 ( .A(n133), .B(n132), .C(n131), .D(n130), .Q(n135) );
  IMUX20 U191 ( .A(i_data_instr_18_), .B(n148), .S(i_addr_Erd[2]), .Q(n134) );
  IMUX20 U192 ( .A(i_data_instr_17_), .B(n142), .S(i_addr_Mrd[1]), .Q(n137) );
  IMUX20 U193 ( .A(i_data_instr_16_), .B(n140), .S(i_addr_Mrd[0]), .Q(n136) );
  NOR40 U194 ( .A(i_data_instr_17_), .B(i_data_instr_19_), .C(i_data_instr_16_), .D(i_data_instr_18_), .Q(n139) );
  IMUX20 U195 ( .A(n140), .B(i_data_instr_16_), .S(i_addr_rtM[0]), .Q(n147) );
  IMUX20 U196 ( .A(n141), .B(i_data_instr_20_), .S(i_addr_rtM[4]), .Q(n146) );
  IMUX20 U197 ( .A(n142), .B(i_data_instr_17_), .S(i_addr_rtM[1]), .Q(n145) );
  IMUX20 U198 ( .A(n143), .B(i_data_instr_19_), .S(i_addr_rtM[3]), .Q(n144) );
  NOR40 U199 ( .A(n147), .B(n146), .C(n145), .D(n144), .Q(n150) );
  IMUX20 U200 ( .A(i_data_instr_18_), .B(n148), .S(i_addr_rtM[2]), .Q(n149) );
  NAND30 U201 ( .A(i_data_instr_28_), .B(n169), .C(n158), .Q(n159) );
  OAI310 U202 ( .A(i_data_instr_16_), .B(i_data_instr_28_), .C(n161), .D(n159), 
        .Q(jbcon_o_con_bop[0]) );
  NOR20 U203 ( .A(i_data_instr_16_), .B(i_data_instr_28_), .Q(n162) );
  NOR40 U204 ( .A(i_data_instr_0_), .B(i_data_instr_1_), .C(i_data_instr_2_), 
        .D(i_data_instr_4_), .Q(n165) );
  OAI2110 U205 ( .A(n172), .B(i_data_instr_27_), .C(n169), .D(i_data_instr_26_), .Q(n170) );
  AOI210 U206 ( .A(n172), .B(i_data_instr_27_), .C(n170), .Q(n6) );
endmodule


module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Efamux, i_con_Efbmux, 
        i_con_Ealuop, i_con_Eregdst, i_con_Mmemread, i_con_Mmemwrite, 
        i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, i_con_bop, 
        o_data_alures, o_data_rt, o_addr_regdst, o_con_Mmemread, 
        o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, o_con_Wregwrite, 
        o_addr_Erd, o_addr_Mrt, o_con_ifbranch, i_con_Ealusrc_BAR, 
        o_data_pc4_31_, o_data_pc4_30_, o_data_pc4_29__BAR, o_data_pc4_28_, 
        o_data_pc4_26_, o_data_pc4_24_, o_data_pc4_22_, o_data_pc4_20_, 
        o_data_pc4_18_, o_data_pc4_16_, o_data_pc4_14_, o_data_pc4_12_, 
        o_data_pc4_10_, o_data_pc4_8_, o_data_pc4_6_, o_data_pc4_4_, 
        o_data_pc4_3_, o_data_pc4_2_, o_data_pc4_1_, o_data_pc4_0_, 
        o_data_pc4_27__BAR, o_data_pc4_25__BAR, o_data_pc4_23__BAR, 
        o_data_pc4_21__BAR, o_data_pc4_19__BAR, o_data_pc4_17__BAR, 
        o_data_pc4_15__BAR, o_data_pc4_13__BAR, o_data_pc4_11__BAR, 
        o_data_pc4_9__BAR, o_data_pc4_7__BAR, o_data_pc4_5__BAR );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [5:0] i_con_Ealuop;
  input [2:0] i_con_bop;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Eregdst, i_con_Mmemread, i_con_Mmemwrite,
         i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, i_con_Ealusrc_BAR;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch, o_data_pc4_31_, o_data_pc4_30_,
         o_data_pc4_29__BAR, o_data_pc4_28_, o_data_pc4_26_, o_data_pc4_24_,
         o_data_pc4_22_, o_data_pc4_20_, o_data_pc4_18_, o_data_pc4_16_,
         o_data_pc4_14_, o_data_pc4_12_, o_data_pc4_10_, o_data_pc4_8_,
         o_data_pc4_6_, o_data_pc4_4_, o_data_pc4_3_, o_data_pc4_2_,
         o_data_pc4_1_, o_data_pc4_0_, o_data_pc4_27__BAR, o_data_pc4_25__BAR,
         o_data_pc4_23__BAR, o_data_pc4_21__BAR, o_data_pc4_19__BAR,
         o_data_pc4_17__BAR, o_data_pc4_15__BAR, o_data_pc4_13__BAR,
         o_data_pc4_11__BAR, o_data_pc4_9__BAR, o_data_pc4_7__BAR,
         o_data_pc4_5__BAR;
  wire   u_alu_N306, u_alu_N256, u_alu_N255, u_alu_N254, u_alu_N253,
         u_alu_N252, u_alu_N250, u_alu_N249, u_alu_N248, u_alu_N247,
         u_alu_N246, u_alu_N245, u_alu_N244, u_alu_N243, u_alu_N242,
         u_alu_N241, u_alu_N236, u_alu_N235, u_alu_N234, u_alu_N233,
         u_alu_N232, u_alu_N231, u_alu_N230, u_alu_N229, u_alu_N228,
         u_alu_N227, u_alu_N226, u_alu_N225, u_alu_N224, u_alu_N223,
         u_alu_N222, u_alu_N221, u_alu_N220, u_alu_N219, u_alu_N218,
         u_alu_N217, u_alu_N216, u_alu_N215, u_alu_N214, u_alu_N213,
         u_alu_N212, u_alu_N211, u_alu_N210, u_alu_N209, u_alu_N204,
         u_alu_N203, u_alu_N202, u_alu_N201, u_alu_N200, u_alu_N199,
         u_alu_N198, u_alu_N197, u_alu_N196, u_alu_N195, u_alu_N194,
         u_alu_N193, u_alu_N173, u_alu_N172, u_alu_N171, u_alu_N170,
         u_alu_N169, u_alu_N168, u_alu_N167, u_alu_N166, u_alu_N165,
         u_alu_half_sub_0_, u_alu_half_sub_1_, u_alu_half_sub_2_,
         u_alu_half_sub_3_, u_alu_half_sub_4_, u_alu_half_sub_5_,
         u_alu_half_sub_6_, u_alu_half_sub_7_, u_alu_half_sub_8_,
         u_alu_half_sub_9_, u_alu_half_sub_10_, u_alu_half_sub_11_,
         u_alu_half_sub_12_, u_alu_half_sub_13_, u_alu_half_sub_14_,
         u_alu_half_sub_15_, u_alu_half_sub_16_, u_alu_sum_1_0_,
         u_alu_sum_1_1_, u_alu_sum_1_2_, u_alu_sum_1_3_, u_alu_sum_1_4_,
         u_alu_sum_1_5_, u_alu_sum_1_6_, u_alu_sum_1_7_, u_alu_sum_1_8_,
         u_alu_ashr_4_SH_3_, u_alu_ashr_4_SH_1_, u_alu_DP_OP_85J3_126_1427_n46,
         u_alu_DP_OP_85J3_126_1427_n45, u_alu_DP_OP_85J3_126_1427_n44,
         u_alu_DP_OP_85J3_126_1427_n43, u_alu_DP_OP_85J3_126_1427_n42,
         u_alu_DP_OP_85J3_126_1427_n41, u_alu_DP_OP_85J3_126_1427_n40,
         u_alu_DP_OP_85J3_126_1427_n39, u_alu_DP_OP_85J3_126_1427_n38,
         u_alu_DP_OP_85J3_126_1427_n37, u_alu_DP_OP_85J3_126_1427_n36,
         u_alu_DP_OP_85J3_126_1427_n35, u_alu_DP_OP_85J3_126_1427_n34,
         u_alu_DP_OP_85J3_126_1427_n33, u_alu_DP_OP_85J3_126_1427_n32,
         u_alu_DP_OP_84J3_125_2615_n15, u_alu_DP_OP_84J3_125_2615_n14,
         u_alu_DP_OP_84J3_125_2615_n13, u_alu_DP_OP_84J3_125_2615_n12,
         u_alu_DP_OP_84J3_125_2615_n11, u_alu_DP_OP_84J3_125_2615_n10,
         u_alu_DP_OP_84J3_125_2615_n9, u_alu_DP_OP_84J3_125_2615_n6,
         u_alu_DP_OP_84J3_125_2615_n5, u_alu_DP_OP_84J3_125_2615_n4,
         u_alu_DP_OP_84J3_125_2615_n3, u_alu_DP_OP_84J3_125_2615_n2,
         u_alu_DP_OP_84J3_125_2615_n1, u_alu_DP_OP_83J3_124_3384_n15,
         u_alu_DP_OP_83J3_124_3384_n14, u_alu_DP_OP_83J3_124_3384_n13,
         u_alu_DP_OP_83J3_124_3384_n12, u_alu_DP_OP_83J3_124_3384_n11,
         u_alu_DP_OP_83J3_124_3384_n10, u_alu_DP_OP_83J3_124_3384_n9,
         u_alu_DP_OP_83J3_124_3384_n7, u_alu_DP_OP_83J3_124_3384_n6,
         u_alu_DP_OP_83J3_124_3384_n5, u_alu_DP_OP_83J3_124_3384_n4,
         u_alu_DP_OP_83J3_124_3384_n3, u_alu_DP_OP_83J3_124_3384_n2,
         u_alu_DP_OP_83J3_124_3384_n1, u_alu_lt_x_11_B_2_, u_alu_sub_x_2_n17,
         u_alu_sub_x_2_n16, u_alu_sub_x_2_n15, u_alu_sub_x_2_n14,
         u_alu_sub_x_2_n13, u_alu_sub_x_2_n12, u_alu_sub_x_2_n11,
         u_alu_sub_x_2_n10, u_alu_sub_x_2_n9, u_alu_sub_x_2_n8,
         u_alu_sub_x_2_n7, u_alu_sub_x_2_n6, u_alu_sub_x_2_n5,
         u_alu_sub_x_2_n4, u_alu_sub_x_2_n3, u_alu_sub_x_2_n2,
         u_alu_add_x_1_n8, u_alu_add_x_1_n7, u_alu_add_x_1_n6,
         u_alu_add_x_1_n5, u_alu_add_x_1_n4, u_alu_add_x_1_n3,
         u_alu_add_x_1_n2, DP_OP_77J3_127_5954_I3, DP_OP_77J3_127_5954_n46,
         DP_OP_77J3_127_5954_n45, DP_OP_77J3_127_5954_n44,
         DP_OP_77J3_127_5954_n43, DP_OP_77J3_127_5954_n42,
         DP_OP_77J3_127_5954_n41, DP_OP_77J3_127_5954_n40,
         DP_OP_77J3_127_5954_n39, DP_OP_77J3_127_5954_n23,
         DP_OP_77J3_127_5954_n22, DP_OP_77J3_127_5954_n21,
         DP_OP_77J3_127_5954_n20, DP_OP_77J3_127_5954_n19,
         DP_OP_77J3_127_5954_n18, DP_OP_77J3_127_5954_n17,
         DP_OP_77J3_127_5954_n16, DP_OP_77J3_127_5954_n15,
         DP_OP_77J3_127_5954_n14, DP_OP_77J3_127_5954_n13,
         DP_OP_77J3_127_5954_n12, DP_OP_77J3_127_5954_n11,
         DP_OP_77J3_127_5954_n10, DP_OP_77J3_127_5954_n8,
         DP_OP_77J3_127_5954_n7, DP_OP_77J3_127_5954_n6,
         DP_OP_77J3_127_5954_n5, DP_OP_77J3_127_5954_n4,
         DP_OP_77J3_127_5954_n3, DP_OP_77J3_127_5954_n2,
         DP_OP_77J3_127_5954_n1, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275;
  wire   [31:0] alu_o_data_AluRes;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;
  wire   [15:0] u_alu_pre_subb;
  wire   [15:1] u_alu_pre_suba;
  wire   [6:1] u_alu_pre_sum_4b;
  wire   [7:0] u_alu_pre_sum_4a;
  wire   [8:1] u_alu_pre_sum_3b;
  wire   [8:0] u_alu_pre_sum_3a;

  DFC1 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC1 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC1 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC1 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC1 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC1 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_31_) );
  DFC1 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_30_) );
  DFC1 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_29__BAR) );
  DFC1 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_28_) );
  DFC1 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_27__BAR) );
  DFC1 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_26_) );
  DFC1 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_25__BAR) );
  DFC1 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_24_) );
  DFC1 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_23__BAR) );
  DFC1 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_22_) );
  DFC1 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_21__BAR) );
  DFC1 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_20_) );
  DFC1 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_19__BAR) );
  DFC1 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_18_) );
  DFC1 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_17__BAR) );
  DFC1 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_16_) );
  DFC1 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_15__BAR) );
  DFC1 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_14_) );
  DFC1 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_13__BAR) );
  DFC1 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_12_) );
  DFC1 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_11__BAR) );
  DFC1 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_10_) );
  DFC1 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_9__BAR) );
  DFC1 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_8_) );
  DFC1 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_7__BAR) );
  DFC1 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_6_) );
  DFC1 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_5__BAR) );
  DFC1 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_4_) );
  DFC1 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_3_) );
  DFC1 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_2_) );
  DFC1 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_1_) );
  DFC1 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_0_) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  DFC1 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC1 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC1 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC1 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC1 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC1 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC1 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC1 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC1 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC1 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC1 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC1 pipe_alures_reg_15_ ( .D(alu_o_data_AluRes[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[15]) );
  DFC1 pipe_alures_reg_14_ ( .D(alu_o_data_AluRes[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[14]) );
  DFC1 pipe_alures_reg_13_ ( .D(alu_o_data_AluRes[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[13]) );
  DFC1 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC1 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC1 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC1 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC1 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC1 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC1 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC1 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC1 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC1 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC1 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC1 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC1 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC1 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC1 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC1 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC1 pipe_rt_reg_28_ ( .D(compare_i_data_rt[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[28]) );
  DFC1 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  DFC1 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC1 pipe_rt_reg_25_ ( .D(compare_i_data_rt[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[25]) );
  DFC1 pipe_rt_reg_24_ ( .D(compare_i_data_rt[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[24]) );
  DFC1 pipe_rt_reg_23_ ( .D(compare_i_data_rt[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[23]) );
  DFC1 pipe_rt_reg_22_ ( .D(compare_i_data_rt[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[22]) );
  DFC1 pipe_rt_reg_21_ ( .D(compare_i_data_rt[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[21]) );
  DFC1 pipe_rt_reg_20_ ( .D(compare_i_data_rt[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[20]) );
  DFC1 pipe_rt_reg_19_ ( .D(compare_i_data_rt[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[19]) );
  DFC1 pipe_rt_reg_18_ ( .D(compare_i_data_rt[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[18]) );
  DFC1 pipe_rt_reg_17_ ( .D(compare_i_data_rt[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[17]) );
  DFC1 pipe_rt_reg_16_ ( .D(compare_i_data_rt[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[16]) );
  DFC1 pipe_rt_reg_15_ ( .D(compare_i_data_rt[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[15]) );
  DFC1 pipe_rt_reg_14_ ( .D(compare_i_data_rt[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[14]) );
  DFC1 pipe_rt_reg_13_ ( .D(compare_i_data_rt[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[13]) );
  DFC1 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC1 pipe_rt_reg_11_ ( .D(compare_i_data_rt[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[11]) );
  DFC1 pipe_rt_reg_10_ ( .D(compare_i_data_rt[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[10]) );
  DFC1 pipe_rt_reg_9_ ( .D(compare_i_data_rt[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[9]) );
  DFC1 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC1 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC1 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC1 pipe_rt_reg_5_ ( .D(compare_i_data_rt[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[5]) );
  DFC1 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC1 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC1 pipe_rt_reg_2_ ( .D(compare_i_data_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[2]) );
  DFC1 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC1 pipe_rt_reg_0_ ( .D(compare_i_data_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[0]) );
  DFC1 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC1 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC1 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC1 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC1 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC1 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC1 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC1 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC1 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_con_Malupc8_reg ( .D(i_con_Malupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Malupc8) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U47 ( .A(n77), .B(compare_i_data_rs[30]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n33), .CO(u_alu_DP_OP_85J3_126_1427_n32), 
        .S(u_alu_pre_suba[14]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U48 ( .A(n79), .B(compare_i_data_rs[29]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n34), .CO(u_alu_DP_OP_85J3_126_1427_n33), 
        .S(u_alu_pre_suba[13]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U49 ( .A(n90), .B(compare_i_data_rs[28]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n35), .CO(u_alu_DP_OP_85J3_126_1427_n34), 
        .S(u_alu_pre_suba[12]) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U11 ( .A(compare_i_data_rs[30]), .B(
        alu_i_data_B[30]), .CI(u_alu_DP_OP_84J3_125_2615_n10), .CO(
        u_alu_DP_OP_84J3_125_2615_n9), .S(u_alu_pre_sum_4a[6]) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U12 ( .A(compare_i_data_rs[29]), .B(
        alu_i_data_B[29]), .CI(u_alu_DP_OP_84J3_125_2615_n11), .CO(
        u_alu_DP_OP_84J3_125_2615_n10), .S(u_alu_pre_sum_4a[5]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U2 ( .A(u_alu_pre_sum_4a[6]), .B(
        u_alu_DP_OP_84J3_125_2615_n2), .CO(u_alu_DP_OP_84J3_125_2615_n1), .S(
        u_alu_pre_sum_4b[6]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U3 ( .A(u_alu_pre_sum_4a[5]), .B(
        u_alu_DP_OP_84J3_125_2615_n3), .CO(u_alu_DP_OP_84J3_125_2615_n2), .S(
        u_alu_pre_sum_4b[5]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U7 ( .A(u_alu_pre_sum_4a[1]), .B(
        u_alu_pre_sum_4a[0]), .CO(u_alu_DP_OP_84J3_125_2615_n6), .S(
        u_alu_pre_sum_4b[1]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U4 ( .A(u_alu_pre_sum_4a[4]), .B(
        u_alu_DP_OP_84J3_125_2615_n4), .CO(u_alu_DP_OP_84J3_125_2615_n3), .S(
        u_alu_pre_sum_4b[4]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U5 ( .A(u_alu_pre_sum_4a[3]), .B(
        u_alu_DP_OP_84J3_125_2615_n5), .CO(u_alu_DP_OP_84J3_125_2615_n4), .S(
        u_alu_pre_sum_4b[3]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U6 ( .A(u_alu_pre_sum_4a[2]), .B(
        u_alu_DP_OP_84J3_125_2615_n6), .CO(u_alu_DP_OP_84J3_125_2615_n5), .S(
        u_alu_pre_sum_4b[2]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U17 ( .A(compare_i_data_rs[24]), .B(
        alu_i_data_B[24]), .CO(u_alu_DP_OP_84J3_125_2615_n15), .S(
        u_alu_pre_sum_4a[0]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U5 ( .A(u_alu_pre_sum_3a[4]), .B(
        u_alu_DP_OP_83J3_124_3384_n5), .CO(u_alu_DP_OP_83J3_124_3384_n4), .S(
        u_alu_pre_sum_3b[4]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U6 ( .A(u_alu_pre_sum_3a[3]), .B(
        u_alu_DP_OP_83J3_124_3384_n6), .CO(u_alu_DP_OP_83J3_124_3384_n5), .S(
        u_alu_pre_sum_3b[3]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U7 ( .A(u_alu_pre_sum_3a[2]), .B(
        u_alu_DP_OP_83J3_124_3384_n7), .CO(u_alu_DP_OP_83J3_124_3384_n6), .S(
        u_alu_pre_sum_3b[2]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U8 ( .A(u_alu_pre_sum_3a[1]), .B(
        u_alu_pre_sum_3a[0]), .CO(u_alu_DP_OP_83J3_124_3384_n7), .S(
        u_alu_pre_sum_3b[1]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U10 ( .A(compare_i_data_rs[23]), .B(
        alu_i_data_B[23]), .CI(u_alu_DP_OP_83J3_124_3384_n9), .CO(
        u_alu_pre_sum_3a[8]), .S(u_alu_pre_sum_3a[7]) );
  ADD31 u_alu_sub_x_2_U14 ( .A(n121), .B(compare_i_data_rs[3]), .CI(
        u_alu_sub_x_2_n15), .CO(u_alu_sub_x_2_n14), .S(u_alu_half_sub_3_) );
  ADD31 u_alu_sub_x_2_U13 ( .A(n93), .B(compare_i_data_rs[4]), .CI(
        u_alu_sub_x_2_n14), .CO(u_alu_sub_x_2_n13), .S(u_alu_half_sub_4_) );
  ADD31 u_alu_sub_x_2_U12 ( .A(n122), .B(compare_i_data_rs[5]), .CI(
        u_alu_sub_x_2_n13), .CO(u_alu_sub_x_2_n12), .S(u_alu_half_sub_5_) );
  AOI221 DP_OP_77J3_127_5954_U25 ( .A(DP_OP_77J3_127_5954_I3), .B(
        compare_i_data_rs[9]), .C(DP_OP_77J3_127_5954_n39), .D(n120), .Q(
        DP_OP_77J3_127_5954_n16) );
  AOI221 DP_OP_77J3_127_5954_U23 ( .A(DP_OP_77J3_127_5954_I3), .B(
        compare_i_data_rs[10]), .C(DP_OP_77J3_127_5954_n40), .D(n120), .Q(
        DP_OP_77J3_127_5954_n15) );
  ADD22 DP_OP_77J3_127_5954_U30 ( .A(DP_OP_77J3_127_5954_n20), .B(
        compare_i_data_rs[13]), .CO(DP_OP_77J3_127_5954_n19), .S(
        DP_OP_77J3_127_5954_n43) );
  AOI221 DP_OP_77J3_127_5954_U13 ( .A(DP_OP_77J3_127_5954_I3), .B(
        compare_i_data_rs[15]), .C(DP_OP_77J3_127_5954_n45), .D(n120), .Q(
        DP_OP_77J3_127_5954_n10) );
  ADD22 DP_OP_77J3_127_5954_U29 ( .A(DP_OP_77J3_127_5954_n19), .B(
        compare_i_data_rs[14]), .CO(DP_OP_77J3_127_5954_n18), .S(
        DP_OP_77J3_127_5954_n44) );
  AOI221 DP_OP_77J3_127_5954_U21 ( .A(DP_OP_77J3_127_5954_I3), .B(
        compare_i_data_rs[11]), .C(DP_OP_77J3_127_5954_n41), .D(n120), .Q(
        DP_OP_77J3_127_5954_n14) );
  ADD22 DP_OP_77J3_127_5954_U28 ( .A(DP_OP_77J3_127_5954_n18), .B(
        compare_i_data_rs[15]), .CO(DP_OP_77J3_127_5954_n46), .S(
        DP_OP_77J3_127_5954_n45) );
  AOI221 DP_OP_77J3_127_5954_U19 ( .A(DP_OP_77J3_127_5954_I3), .B(
        compare_i_data_rs[12]), .C(DP_OP_77J3_127_5954_n42), .D(n120), .Q(
        DP_OP_77J3_127_5954_n13) );
  AOI221 DP_OP_77J3_127_5954_U17 ( .A(DP_OP_77J3_127_5954_I3), .B(
        compare_i_data_rs[13]), .C(DP_OP_77J3_127_5954_n43), .D(n120), .Q(
        DP_OP_77J3_127_5954_n12) );
  AOI221 DP_OP_77J3_127_5954_U15 ( .A(DP_OP_77J3_127_5954_I3), .B(
        compare_i_data_rs[14]), .C(DP_OP_77J3_127_5954_n44), .D(n120), .Q(
        DP_OP_77J3_127_5954_n11) );
  ADD22 DP_OP_77J3_127_5954_U34 ( .A(compare_i_data_rs[8]), .B(
        compare_i_data_rs[9]), .CO(DP_OP_77J3_127_5954_n23), .S(
        DP_OP_77J3_127_5954_n39) );
  ADD22 DP_OP_77J3_127_5954_U33 ( .A(DP_OP_77J3_127_5954_n23), .B(
        compare_i_data_rs[10]), .CO(DP_OP_77J3_127_5954_n22), .S(
        DP_OP_77J3_127_5954_n40) );
  ADD22 DP_OP_77J3_127_5954_U32 ( .A(DP_OP_77J3_127_5954_n22), .B(
        compare_i_data_rs[11]), .CO(DP_OP_77J3_127_5954_n21), .S(
        DP_OP_77J3_127_5954_n41) );
  ADD22 DP_OP_77J3_127_5954_U31 ( .A(DP_OP_77J3_127_5954_n21), .B(
        compare_i_data_rs[12]), .CO(DP_OP_77J3_127_5954_n20), .S(
        DP_OP_77J3_127_5954_n42) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U16 ( .A(compare_i_data_rs[25]), .B(
        alu_i_data_B[25]), .CI(u_alu_DP_OP_84J3_125_2615_n15), .CO(
        u_alu_DP_OP_84J3_125_2615_n14), .S(u_alu_pre_sum_4a[1]) );
  ADD32 u_alu_add_x_1_U8 ( .A(compare_i_data_rs[1]), .B(n71), .CI(
        u_alu_add_x_1_n8), .CO(u_alu_add_x_1_n7), .S(u_alu_sum_1_1_) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U15 ( .A(compare_i_data_rs[26]), .B(
        alu_i_data_B[26]), .CI(u_alu_DP_OP_84J3_125_2615_n14), .CO(
        u_alu_DP_OP_84J3_125_2615_n13), .S(u_alu_pre_sum_4a[2]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U59 ( .A(n73), .B(compare_i_data_rs[18]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n45), .CO(u_alu_DP_OP_85J3_126_1427_n44), 
        .S(u_alu_pre_suba[2]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U15 ( .A(compare_i_data_rs[18]), .B(
        alu_i_data_B[18]), .CI(u_alu_DP_OP_83J3_124_3384_n14), .CO(
        u_alu_DP_OP_83J3_124_3384_n13), .S(u_alu_pre_sum_3a[2]) );
  ADD32 u_alu_add_x_1_U7 ( .A(compare_i_data_rs[2]), .B(u_alu_lt_x_11_B_2_), 
        .CI(u_alu_add_x_1_n7), .CO(u_alu_add_x_1_n6), .S(u_alu_sum_1_2_) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U14 ( .A(compare_i_data_rs[27]), .B(
        alu_i_data_B[27]), .CI(u_alu_DP_OP_84J3_125_2615_n13), .CO(
        u_alu_DP_OP_84J3_125_2615_n12), .S(u_alu_pre_sum_4a[3]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U14 ( .A(compare_i_data_rs[19]), .B(
        alu_i_data_B[19]), .CI(u_alu_DP_OP_83J3_124_3384_n13), .CO(
        u_alu_DP_OP_83J3_124_3384_n12), .S(u_alu_pre_sum_3a[3]) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U13 ( .A(compare_i_data_rs[28]), .B(
        alu_i_data_B[28]), .CI(u_alu_DP_OP_84J3_125_2615_n12), .CO(
        u_alu_DP_OP_84J3_125_2615_n11), .S(u_alu_pre_sum_4a[4]) );
  ADD32 u_alu_add_x_1_U6 ( .A(compare_i_data_rs[3]), .B(n229), .CI(
        u_alu_add_x_1_n6), .CO(u_alu_add_x_1_n5), .S(u_alu_sum_1_3_) );
  ADD32 u_alu_add_x_1_U5 ( .A(compare_i_data_rs[4]), .B(alu_i_data_B[4]), .CI(
        u_alu_add_x_1_n5), .CO(u_alu_add_x_1_n4), .S(u_alu_sum_1_4_) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U13 ( .A(compare_i_data_rs[20]), .B(
        alu_i_data_B[20]), .CI(u_alu_DP_OP_83J3_124_3384_n12), .CO(
        u_alu_DP_OP_83J3_124_3384_n11), .S(u_alu_pre_sum_3a[4]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U56 ( .A(n72), .B(compare_i_data_rs[21]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n42), .CO(u_alu_DP_OP_85J3_126_1427_n41), 
        .S(u_alu_pre_suba[5]) );
  ADD32 u_alu_add_x_1_U4 ( .A(compare_i_data_rs[5]), .B(alu_i_data_B[5]), .CI(
        u_alu_add_x_1_n4), .CO(u_alu_add_x_1_n3), .S(u_alu_sum_1_5_) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U12 ( .A(compare_i_data_rs[21]), .B(
        alu_i_data_B[21]), .CI(u_alu_DP_OP_83J3_124_3384_n11), .CO(
        u_alu_DP_OP_83J3_124_3384_n10), .S(u_alu_pre_sum_3a[5]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U4 ( .A(u_alu_pre_sum_3a[5]), .B(
        u_alu_DP_OP_83J3_124_3384_n4), .CO(u_alu_DP_OP_83J3_124_3384_n3), .S(
        u_alu_pre_sum_3b[5]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U11 ( .A(compare_i_data_rs[22]), .B(
        alu_i_data_B[22]), .CI(u_alu_DP_OP_83J3_124_3384_n10), .CO(
        u_alu_DP_OP_83J3_124_3384_n9), .S(u_alu_pre_sum_3a[6]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U3 ( .A(u_alu_pre_sum_3a[6]), .B(
        u_alu_DP_OP_83J3_124_3384_n3), .CO(u_alu_DP_OP_83J3_124_3384_n2), .S(
        u_alu_pre_sum_3b[6]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U2 ( .A(u_alu_pre_sum_3a[7]), .B(
        u_alu_DP_OP_83J3_124_3384_n2), .CO(u_alu_DP_OP_83J3_124_3384_n1), .S(
        u_alu_pre_sum_3b[7]) );
  ADD32 u_alu_sub_x_2_U8 ( .A(n124), .B(compare_i_data_rs[9]), .CI(
        u_alu_sub_x_2_n9), .CO(u_alu_sub_x_2_n8), .S(u_alu_half_sub_9_) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U51 ( .A(n78), .B(compare_i_data_rs[26]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n37), .CO(u_alu_DP_OP_85J3_126_1427_n36), 
        .S(u_alu_pre_suba[10]) );
  ADD22 DP_OP_77J3_127_5954_U9 ( .A(n112), .B(alu_i_data_B[8]), .CO(
        DP_OP_77J3_127_5954_n8), .S(u_alu_N165) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U50 ( .A(n76), .B(compare_i_data_rs[27]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n36), .CO(u_alu_DP_OP_85J3_126_1427_n35), 
        .S(u_alu_pre_suba[11]) );
  ADD32 DP_OP_77J3_127_5954_U8 ( .A(n113), .B(alu_i_data_B[9]), .CI(
        DP_OP_77J3_127_5954_n8), .CO(DP_OP_77J3_127_5954_n7), .S(u_alu_N166)
         );
  ADD32 DP_OP_77J3_127_5954_U7 ( .A(n114), .B(alu_i_data_B[10]), .CI(
        DP_OP_77J3_127_5954_n7), .CO(DP_OP_77J3_127_5954_n6), .S(u_alu_N167)
         );
  ADD32 u_alu_sub_x_2_U4 ( .A(n126), .B(compare_i_data_rs[13]), .CI(
        u_alu_sub_x_2_n5), .CO(u_alu_sub_x_2_n4), .S(u_alu_half_sub_13_) );
  ADD32 DP_OP_77J3_127_5954_U6 ( .A(n115), .B(alu_i_data_B[11]), .CI(
        DP_OP_77J3_127_5954_n6), .CO(DP_OP_77J3_127_5954_n5), .S(u_alu_N168)
         );
  ADD32 u_alu_sub_x_2_U3 ( .A(n127), .B(compare_i_data_rs[14]), .CI(
        u_alu_sub_x_2_n4), .CO(u_alu_sub_x_2_n3), .S(u_alu_half_sub_14_) );
  ADD32 u_alu_sub_x_2_U2 ( .A(n80), .B(compare_i_data_rs[15]), .CI(
        u_alu_sub_x_2_n3), .CO(u_alu_sub_x_2_n2), .S(u_alu_half_sub_15_) );
  ADD32 u_alu_sub_x_2_U16 ( .A(n83), .B(compare_i_data_rs[1]), .CI(
        u_alu_sub_x_2_n17), .CO(u_alu_sub_x_2_n16), .S(u_alu_half_sub_1_) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U58 ( .A(n86), .B(compare_i_data_rs[19]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n44), .CO(u_alu_DP_OP_85J3_126_1427_n43), 
        .S(u_alu_pre_suba[3]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U57 ( .A(n87), .B(compare_i_data_rs[20]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n43), .CO(u_alu_DP_OP_85J3_126_1427_n42), 
        .S(u_alu_pre_suba[4]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U55 ( .A(n85), .B(compare_i_data_rs[22]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n41), .CO(u_alu_DP_OP_85J3_126_1427_n40), 
        .S(u_alu_pre_suba[6]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U54 ( .A(n84), .B(compare_i_data_rs[23]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n40), .CO(u_alu_DP_OP_85J3_126_1427_n39), 
        .S(u_alu_pre_suba[7]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U53 ( .A(n89), .B(compare_i_data_rs[24]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n39), .CO(u_alu_DP_OP_85J3_126_1427_n38), 
        .S(u_alu_pre_suba[8]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U52 ( .A(n88), .B(compare_i_data_rs[25]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n38), .CO(u_alu_DP_OP_85J3_126_1427_n37), 
        .S(u_alu_pre_suba[9]) );
  ADD32 u_alu_sub_x_2_U5 ( .A(n94), .B(compare_i_data_rs[12]), .CI(
        u_alu_sub_x_2_n6), .CO(u_alu_sub_x_2_n5), .S(u_alu_half_sub_12_) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U16 ( .A(compare_i_data_rs[17]), .B(
        alu_i_data_B[17]), .CI(u_alu_DP_OP_83J3_124_3384_n15), .CO(
        u_alu_DP_OP_83J3_124_3384_n14), .S(u_alu_pre_sum_3a[1]) );
  ADD32 u_alu_sub_x_2_U15 ( .A(n95), .B(compare_i_data_rs[2]), .CI(
        u_alu_sub_x_2_n16), .CO(u_alu_sub_x_2_n15), .S(u_alu_half_sub_2_) );
  ADD32 u_alu_sub_x_2_U11 ( .A(n123), .B(compare_i_data_rs[6]), .CI(
        u_alu_sub_x_2_n12), .CO(u_alu_sub_x_2_n11), .S(u_alu_half_sub_6_) );
  NOR23 U3 ( .A(n526), .B(n513), .Q(n624) );
  INV3 U4 ( .A(n513), .Q(n512) );
  INV3 U5 ( .A(n515), .Q(n514) );
  INV3 U6 ( .A(i_con_Ealusrc_BAR), .Q(n70) );
  NOR21 U7 ( .A(n1143), .B(n231), .Q(n1056) );
  INV3 U8 ( .A(compare_i_data_rt[0]), .Q(n852) );
  INV3 U9 ( .A(n763), .Q(n111) );
  INV3 U10 ( .A(n111), .Q(n516) );
  INV3 U11 ( .A(n518), .Q(n517) );
  NAND31 U12 ( .A(n620), .B(n619), .C(n618), .Q(compare_i_data_rs[2]) );
  IMUX21 U13 ( .A(n842), .B(n1210), .S(n70), .Q(alu_i_data_B[5]) );
  BUF2 U14 ( .A(n1078), .Q(n519) );
  INV3 U15 ( .A(n959), .Q(n956) );
  NAND41 U16 ( .A(n1028), .B(n1027), .C(n1026), .D(n1025), .Q(
        alu_o_data_AluRes[28]) );
  IMUX20 U17 ( .A(n1076), .B(n1079), .S(compare_i_data_rs[12]), .Q(n1) );
  CLKIN0 U18 ( .A(u_alu_half_sub_12_), .Q(n2) );
  IMUX20 U19 ( .A(n467), .B(n432), .S(u_alu_ashr_4_SH_3_), .Q(n3) );
  IMUX20 U20 ( .A(n3), .B(n445), .S(i_data_immext[10]), .Q(n4) );
  AOI220 U21 ( .A(n4), .B(n1077), .C(n859), .D(u_alu_N169), .Q(n5) );
  CLKIN0 U22 ( .A(n372), .Q(n6) );
  NAND30 U23 ( .A(n519), .B(n327), .C(n6), .Q(n7) );
  OAI2110 U24 ( .A(n861), .B(n2), .C(n5), .D(n7), .Q(n8) );
  AOI210 U25 ( .A(compare_i_data_rs[12]), .B(n82), .C(n8), .Q(n9) );
  IMUX20 U26 ( .A(n1086), .B(n1087), .S(compare_i_data_rs[12]), .Q(n10) );
  OAI210 U27 ( .A(n82), .B(n10), .C(alu_i_data_B[12]), .Q(n11) );
  OAI2110 U28 ( .A(alu_i_data_B[12]), .B(n1), .C(n9), .D(n11), .Q(
        alu_o_data_AluRes[12]) );
  NAND20 U29 ( .A(DP_OP_77J3_127_5954_n46), .B(n120), .Q(n12) );
  XNR21 U30 ( .A(DP_OP_77J3_127_5954_n1), .B(n12), .Q(u_alu_N173) );
  IMUX20 U31 ( .A(n1076), .B(n1079), .S(compare_i_data_rs[13]), .Q(n13) );
  CLKIN0 U32 ( .A(n1077), .Q(n14) );
  IMUX20 U33 ( .A(n474), .B(n434), .S(u_alu_ashr_4_SH_3_), .Q(n15) );
  IMUX20 U34 ( .A(n15), .B(n446), .S(i_data_immext[10]), .Q(n16) );
  CLKIN0 U35 ( .A(n861), .Q(n17) );
  AOI220 U36 ( .A(n859), .B(u_alu_N170), .C(u_alu_half_sub_13_), .D(n17), .Q(
        n18) );
  CLKIN0 U37 ( .A(n372), .Q(n19) );
  NAND30 U38 ( .A(n519), .B(n334), .C(n19), .Q(n20) );
  OAI2110 U39 ( .A(n14), .B(n16), .C(n18), .D(n20), .Q(n21) );
  AOI210 U40 ( .A(compare_i_data_rs[13]), .B(n82), .C(n21), .Q(n22) );
  IMUX20 U41 ( .A(n1086), .B(n1087), .S(compare_i_data_rs[13]), .Q(n23) );
  OAI210 U42 ( .A(n82), .B(n23), .C(alu_i_data_B[13]), .Q(n24) );
  OAI2110 U43 ( .A(alu_i_data_B[13]), .B(n13), .C(n22), .D(n24), .Q(
        alu_o_data_AluRes[13]) );
  IMUX20 U44 ( .A(n1076), .B(n1079), .S(compare_i_data_rs[14]), .Q(n25) );
  CLKIN0 U45 ( .A(u_alu_half_sub_14_), .Q(n26) );
  IMUX20 U46 ( .A(n478), .B(n437), .S(u_alu_ashr_4_SH_3_), .Q(n27) );
  IMUX20 U47 ( .A(n27), .B(n456), .S(i_data_immext[10]), .Q(n28) );
  AOI220 U48 ( .A(n28), .B(n1077), .C(n859), .D(u_alu_N171), .Q(n29) );
  CLKIN0 U49 ( .A(n372), .Q(n30) );
  NAND30 U50 ( .A(n519), .B(n343), .C(n30), .Q(n31) );
  OAI2110 U51 ( .A(n861), .B(n26), .C(n29), .D(n31), .Q(n32) );
  AOI210 U52 ( .A(compare_i_data_rs[14]), .B(n82), .C(n32), .Q(n33) );
  IMUX20 U53 ( .A(n1086), .B(n1087), .S(compare_i_data_rs[14]), .Q(n34) );
  OAI210 U54 ( .A(n82), .B(n34), .C(alu_i_data_B[14]), .Q(n35) );
  OAI2110 U55 ( .A(alu_i_data_B[14]), .B(n25), .C(n33), .D(n35), .Q(
        alu_o_data_AluRes[14]) );
  NOR20 U56 ( .A(compare_i_data_rs[18]), .B(n73), .Q(n36) );
  IMAJ30 U57 ( .A(n103), .B(alu_i_data_B[19]), .C(n36), .Q(n37) );
  IMAJ30 U58 ( .A(n74), .B(u_alu_DP_OP_85J3_126_1427_n46), .C(
        compare_i_data_rs[17]), .Q(n38) );
  NAND20 U59 ( .A(n184), .B(n38), .Q(n39) );
  AOI210 U60 ( .A(n37), .B(n39), .C(n185), .Q(n40) );
  CLKIN0 U61 ( .A(n40), .Q(n186) );
  NAND20 U62 ( .A(u_alu_pre_sum_4a[7]), .B(u_alu_DP_OP_84J3_125_2615_n1), .Q(
        n41) );
  OAI2110 U63 ( .A(u_alu_pre_sum_4a[7]), .B(u_alu_DP_OP_84J3_125_2615_n1), .C(
        n1070), .D(n41), .Q(n1073) );
  CLKIN0 U64 ( .A(n861), .Q(n42) );
  AOI220 U65 ( .A(n859), .B(u_alu_N172), .C(u_alu_half_sub_15_), .D(n42), .Q(
        n43) );
  CLKIN0 U66 ( .A(n372), .Q(n44) );
  AOI210 U67 ( .A(n80), .B(n1079), .C(n82), .Q(n45) );
  AOI210 U68 ( .A(compare_i_data_rs[15]), .B(n521), .C(n82), .Q(n46) );
  OAI210 U69 ( .A(n1086), .B(compare_i_data_rs[15]), .C(n46), .Q(n47) );
  IMUX20 U70 ( .A(n483), .B(n440), .S(u_alu_ashr_4_SH_3_), .Q(n48) );
  IMUX20 U71 ( .A(n48), .B(n457), .S(i_data_immext[10]), .Q(n49) );
  AOI220 U72 ( .A(alu_i_data_B[15]), .B(n47), .C(n49), .D(n1077), .Q(n50) );
  NAND30 U73 ( .A(n80), .B(n1076), .C(n858), .Q(n51) );
  OAI2110 U74 ( .A(n858), .B(n45), .C(n50), .D(n51), .Q(n52) );
  AOI310 U75 ( .A(n1078), .B(n351), .C(n44), .D(n52), .Q(n53) );
  NAND20 U76 ( .A(n43), .B(n53), .Q(alu_o_data_AluRes[15]) );
  CLKIN0 U77 ( .A(n372), .Q(n54) );
  NAND30 U78 ( .A(n1077), .B(n443), .C(n54), .Q(n998) );
  IMUX20 U79 ( .A(n959), .B(n962), .S(u_alu_pre_sum_3a[0]), .Q(n55) );
  AOI2110 U80 ( .A(n1069), .B(u_alu_pre_subb[0]), .C(n872), .D(n55), .Q(n56)
         );
  CLKIN0 U81 ( .A(n56), .Q(alu_o_data_AluRes[16]) );
  AOI222 U82 ( .A(DP_OP_77J3_127_5954_I3), .B(compare_i_data_rs[8]), .C(n107), 
        .D(n120), .Q(DP_OP_77J3_127_5954_n17) );
  NAND26 U83 ( .A(n860), .B(n859), .Q(n962) );
  NOR24 U84 ( .A(n634), .B(n111), .Q(n776) );
  NOR32 U85 ( .A(n528), .B(i_con_Efamux[1]), .C(i_con_Efamux[2]), .Q(n625) );
  NOR32 U86 ( .A(n527), .B(i_con_Efamux[1]), .C(i_con_Efamux[0]), .Q(n626) );
  NOR32 U87 ( .A(n635), .B(i_con_Efbmux[1]), .C(i_con_Efbmux[0]), .Q(n778) );
  NOR32 U88 ( .A(n636), .B(i_con_Efbmux[1]), .C(i_con_Efbmux[2]), .Q(n777) );
  IMUX23 U89 ( .A(n831), .B(n1206), .S(n70), .Q(n71) );
  BUF8 U90 ( .A(u_alu_sum_1_8_), .Q(n120) );
  AOI2111 U91 ( .A(n1077), .B(u_alu_N250), .C(n982), .D(n981), .Q(n986) );
  AOI2111 U92 ( .A(n1077), .B(u_alu_N246), .C(n926), .D(n925), .Q(n930) );
  OAI211 U93 ( .A(n162), .B(n161), .C(n160), .Q(n176) );
  AOI2111 U94 ( .A(n1077), .B(u_alu_N247), .C(n938), .D(n937), .Q(n942) );
  AOI2111 U95 ( .A(n1077), .B(u_alu_N254), .C(n1034), .D(n1033), .Q(n1038) );
  AOI2111 U96 ( .A(n1077), .B(u_alu_N248), .C(n950), .D(n949), .Q(n954) );
  AOI2111 U97 ( .A(n1077), .B(u_alu_N245), .C(n913), .D(n912), .Q(n917) );
  AOI2111 U98 ( .A(n1077), .B(u_alu_N252), .C(n1008), .D(n1007), .Q(n1012) );
  NOR21 U99 ( .A(i_data_immext[10]), .B(n506), .Q(u_alu_N244) );
  IMUX20 U100 ( .A(n221), .B(u_alu_pre_subb[0]), .S(u_alu_pre_suba[1]), .Q(
        u_alu_pre_subb[1]) );
  NAND30 U101 ( .A(n1076), .B(n865), .C(n81), .Q(n867) );
  INV1 U102 ( .A(n1087), .Q(n521) );
  NOR21 U103 ( .A(n372), .B(n445), .Q(u_alu_N253) );
  IMAJ30 U104 ( .A(n76), .B(compare_i_data_rs[27]), .C(n205), .Q(n134) );
  NAND21 U105 ( .A(compare_i_data_rs[21]), .B(n72), .Q(n142) );
  CLKIN0 U106 ( .A(alu_i_data_B[16]), .Q(n865) );
  NOR20 U107 ( .A(compare_i_data_rs[30]), .B(n77), .Q(n137) );
  NOR20 U108 ( .A(compare_i_data_rs[26]), .B(n78), .Q(n133) );
  NAND21 U109 ( .A(compare_i_data_rs[29]), .B(n79), .Q(n131) );
  INV3 U110 ( .A(alu_i_data_B[17]), .Q(n74) );
  INV2 U111 ( .A(alu_i_data_B[5]), .Q(n122) );
  INV3 U112 ( .A(alu_i_data_B[29]), .Q(n79) );
  INV3 U113 ( .A(alu_i_data_B[26]), .Q(n78) );
  INV3 U114 ( .A(alu_i_data_B[27]), .Q(n76) );
  INV3 U115 ( .A(alu_i_data_B[30]), .Q(n77) );
  XNR20 U116 ( .A(compare_i_data_rs[26]), .B(alu_i_data_B[26]), .Q(n992) );
  INV3 U117 ( .A(alu_i_data_B[8]), .Q(n75) );
  NAND20 U118 ( .A(alu_i_data_B[14]), .B(n106), .Q(n164) );
  MUX22 U119 ( .A(compare_i_data_rt[4]), .B(i_data_immext[4]), .S(n70), .Q(
        alu_i_data_B[4]) );
  NAND21 U120 ( .A(compare_i_data_rt[17]), .B(n711), .Q(n712) );
  INV3 U121 ( .A(compare_i_data_rs[15]), .Q(n858) );
  INV3 U122 ( .A(compare_i_data_rs[18]), .Q(n887) );
  CLKIN3 U123 ( .A(compare_i_data_rs[16]), .Q(n81) );
  INV3 U124 ( .A(compare_i_data_rs[19]), .Q(n103) );
  INV3 U125 ( .A(compare_i_data_rs[29]), .Q(n1032) );
  INV2 U126 ( .A(compare_i_data_rs[14]), .Q(n106) );
  OAI212 U127 ( .A(n517), .B(n1237), .C(n748), .Q(compare_i_data_rt[8]) );
  AOI210 U128 ( .A(n624), .B(i_data_rs[4]), .C(n612), .Q(n613) );
  NAND22 U129 ( .A(n624), .B(i_data_rs[0]), .Q(n629) );
  OAI210 U130 ( .A(n516), .B(n658), .C(n657), .Q(n659) );
  OAI211 U131 ( .A(n512), .B(n750), .C(n601), .Q(n602) );
  OAI211 U132 ( .A(n512), .B(n688), .C(n559), .Q(n560) );
  OAI210 U133 ( .A(n516), .B(n698), .C(n697), .Q(n699) );
  OAI211 U134 ( .A(n512), .B(n718), .C(n577), .Q(n578) );
  OAI211 U135 ( .A(n512), .B(n722), .C(n580), .Q(n581) );
  OAI210 U136 ( .A(n516), .B(n668), .C(n667), .Q(n669) );
  OAI210 U137 ( .A(n516), .B(n648), .C(n647), .Q(n649) );
  OAI211 U138 ( .A(n512), .B(n726), .C(n583), .Q(n584) );
  OAI210 U139 ( .A(n516), .B(n663), .C(n662), .Q(n664) );
  AOI220 U140 ( .A(n777), .B(i_data_FMalures[3]), .C(n111), .D(
        i_data_FEalures[3]), .Q(n768) );
  AOI221 U141 ( .A(n626), .B(i_data_FMmemout[31]), .C(n625), .D(
        i_data_FMalures[31]), .Q(n529) );
  INV2 U142 ( .A(n1200), .Q(n1171) );
  NAND22 U143 ( .A(n633), .B(i_con_Efbmux[1]), .Q(n763) );
  INV2 U144 ( .A(u_alu_ashr_4_SH_1_), .Q(n373) );
  AOI220 U145 ( .A(i_con_Ealuop[4]), .B(n1179), .C(i_con_Ealuop[5]), .D(n1176), 
        .Q(n1177) );
  INV3 U146 ( .A(i_data_FEalures[22]), .Q(n683) );
  INV3 U147 ( .A(i_data_FEalures[23]), .Q(n678) );
  INV1 U148 ( .A(i_con_Efamux[0]), .Q(n528) );
  NAND41 U149 ( .A(n973), .B(n972), .C(n971), .D(n970), .Q(n974) );
  NOR22 U150 ( .A(n964), .B(n963), .Q(n1071) );
  NAND21 U151 ( .A(u_alu_pre_subb[14]), .B(n1069), .Q(n1054) );
  NOR22 U152 ( .A(n861), .B(u_alu_half_sub_16_), .Q(n1068) );
  AOI210 U153 ( .A(compare_i_data_rs[11]), .B(n82), .C(n1148), .Q(n1145) );
  INV3 U154 ( .A(u_alu_sub_x_2_n2), .Q(u_alu_half_sub_16_) );
  AOI210 U155 ( .A(compare_i_data_rs[10]), .B(n82), .C(n1153), .Q(n1150) );
  OAI211 U156 ( .A(n1089), .B(compare_i_data_rs[8]), .C(n1090), .Q(
        alu_o_data_AluRes[8]) );
  AOI210 U157 ( .A(alu_i_data_B[9]), .B(n82), .C(n1088), .Q(n1083) );
  NAND20 U158 ( .A(u_alu_N165), .B(n859), .Q(n796) );
  AOI210 U159 ( .A(alu_i_data_B[7]), .B(n82), .C(n1098), .Q(n1095) );
  INV3 U160 ( .A(u_alu_pre_suba[9]), .Q(n226) );
  NAND21 U161 ( .A(u_alu_half_sub_8_), .B(n826), .Q(n798) );
  INV3 U162 ( .A(u_alu_sum_1_8_), .Q(DP_OP_77J3_127_5954_I3) );
  INV3 U163 ( .A(u_alu_pre_suba[7]), .Q(n225) );
  NAND20 U164 ( .A(u_alu_sum_1_7_), .B(n859), .Q(n802) );
  NAND20 U165 ( .A(u_alu_sum_1_6_), .B(n859), .Q(n805) );
  NAND20 U166 ( .A(u_alu_N209), .B(n519), .Q(n866) );
  AOI220 U167 ( .A(n1077), .B(u_alu_N229), .C(u_alu_half_sub_4_), .D(n826), 
        .Q(n809) );
  NAND20 U168 ( .A(u_alu_sum_1_5_), .B(n859), .Q(n808) );
  INV2 U169 ( .A(u_alu_pre_sum_3a[5]), .Q(n933) );
  INV2 U170 ( .A(u_alu_pre_sum_3a[4]), .Q(n920) );
  AOI2111 U171 ( .A(n1077), .B(u_alu_N244), .C(n901), .D(n900), .Q(n905) );
  INV2 U172 ( .A(u_alu_pre_sum_3a[3]), .Q(n908) );
  INV3 U173 ( .A(u_alu_pre_suba[3]), .Q(n223) );
  INV3 U174 ( .A(n520), .Q(n82) );
  INV2 U175 ( .A(u_alu_pre_sum_3a[2]), .Q(n896) );
  NAND31 U176 ( .A(n1267), .B(n1266), .C(n1265), .Q(n1270) );
  INV2 U177 ( .A(n861), .Q(n826) );
  INV1 U178 ( .A(n1056), .Q(n868) );
  MUX22 U179 ( .A(n409), .B(n408), .S(i_data_immext[8]), .Q(n437) );
  MUX22 U180 ( .A(n413), .B(n412), .S(i_data_immext[8]), .Q(n440) );
  IMAJ30 U181 ( .A(n96), .B(alu_i_data_B[23]), .C(n203), .Q(n187) );
  NOR20 U182 ( .A(compare_i_data_rs[24]), .B(n89), .Q(n132) );
  IMAJ30 U183 ( .A(n100), .B(alu_i_data_B[13]), .C(n163), .Q(n174) );
  OAI211 U184 ( .A(alu_i_data_B[14]), .B(n106), .C(n144), .Q(n173) );
  INV3 U185 ( .A(alu_i_data_B[23]), .Q(n84) );
  INV3 U186 ( .A(alu_i_data_B[22]), .Q(n85) );
  NOR20 U187 ( .A(alu_i_data_B[24]), .B(n110), .Q(n193) );
  NOR20 U188 ( .A(alu_i_data_B[25]), .B(n102), .Q(n192) );
  INV3 U189 ( .A(alu_i_data_B[20]), .Q(n87) );
  INV3 U190 ( .A(alu_i_data_B[19]), .Q(n86) );
  NOR20 U191 ( .A(alu_i_data_B[13]), .B(n100), .Q(n145) );
  NOR20 U192 ( .A(alu_i_data_B[31]), .B(n99), .Q(n129) );
  INV3 U193 ( .A(alu_i_data_B[21]), .Q(n72) );
  INV3 U194 ( .A(alu_i_data_B[18]), .Q(n73) );
  INV1 U195 ( .A(alu_i_data_B[6]), .Q(n123) );
  NAND20 U196 ( .A(n101), .B(alu_i_data_B[28]), .Q(n130) );
  INV3 U197 ( .A(compare_i_data_rs[30]), .Q(n1042) );
  INV3 U198 ( .A(alu_i_data_B[0]), .Q(n1154) );
  INV3 U199 ( .A(compare_i_data_rt[1]), .Q(n831) );
  INV3 U200 ( .A(compare_i_data_rs[17]), .Q(n98) );
  INV3 U201 ( .A(alu_i_data_B[15]), .Q(n80) );
  INV3 U202 ( .A(compare_i_data_rs[28]), .Q(n101) );
  NAND22 U203 ( .A(compare_i_data_rt[20]), .B(n711), .Q(n696) );
  INV3 U204 ( .A(compare_i_data_rs[13]), .Q(n100) );
  INV3 U205 ( .A(compare_i_data_rs[11]), .Q(n97) );
  INV3 U206 ( .A(compare_i_data_rs[25]), .Q(n102) );
  CLKIN3 U207 ( .A(compare_i_data_rs[0]), .Q(n128) );
  INV2 U208 ( .A(u_alu_lt_x_11_B_2_), .Q(n95) );
  OAI211 U209 ( .A(n517), .B(n1226), .C(n670), .Q(compare_i_data_rt[25]) );
  IMUX23 U210 ( .A(n843), .B(n1209), .S(n70), .Q(n229) );
  NAND31 U211 ( .A(n617), .B(n616), .C(n615), .Q(compare_i_data_rs[3]) );
  OAI211 U212 ( .A(n517), .B(n1225), .C(n675), .Q(compare_i_data_rt[24]) );
  IMUX23 U213 ( .A(n836), .B(n1207), .S(n70), .Q(u_alu_lt_x_11_B_2_) );
  NAND20 U214 ( .A(compare_i_data_rt[31]), .B(n711), .Q(n641) );
  NAND33 U215 ( .A(n629), .B(n628), .C(n627), .Q(compare_i_data_rs[0]) );
  AOI211 U216 ( .A(n624), .B(i_data_rs[21]), .C(n560), .Q(n561) );
  AOI211 U217 ( .A(n624), .B(i_data_rs[15]), .C(n578), .Q(n579) );
  AOI211 U218 ( .A(n624), .B(i_data_rs[30]), .C(n533), .Q(n534) );
  AOI211 U219 ( .A(n624), .B(i_data_rs[23]), .C(n554), .Q(n555) );
  AOI211 U220 ( .A(n624), .B(i_data_rs[28]), .C(n539), .Q(n540) );
  AOI211 U221 ( .A(n624), .B(i_data_rs[29]), .C(n536), .Q(n537) );
  AOI211 U222 ( .A(n624), .B(i_data_rs[26]), .C(n545), .Q(n546) );
  AOI211 U223 ( .A(n624), .B(i_data_rs[27]), .C(n542), .Q(n543) );
  AOI211 U224 ( .A(n624), .B(i_data_rs[25]), .C(n548), .Q(n549) );
  AOI211 U225 ( .A(n624), .B(i_data_rs[14]), .C(n581), .Q(n582) );
  AOI210 U226 ( .A(n624), .B(i_data_rs[8]), .C(n599), .Q(n600) );
  AOI211 U227 ( .A(n624), .B(i_data_rs[10]), .C(n593), .Q(n594) );
  AOI211 U228 ( .A(n624), .B(i_data_rs[12]), .C(n587), .Q(n588) );
  OAI210 U229 ( .A(n512), .B(n693), .C(n562), .Q(n563) );
  NAND21 U230 ( .A(n776), .B(i_data_rt[2]), .Q(n772) );
  AOI220 U231 ( .A(n778), .B(i_data_FMmemout[4]), .C(n777), .D(
        i_data_FMalures[4]), .Q(n761) );
  AOI220 U232 ( .A(n778), .B(i_data_FMmemout[5]), .C(n777), .D(
        i_data_FMalures[5]), .Q(n757) );
  INV3 U233 ( .A(n611), .Q(n513) );
  INV2 U234 ( .A(i_data_immext[8]), .Q(n509) );
  NOR21 U235 ( .A(i_con_Efbmux[1]), .B(n633), .Q(n634) );
  INV3 U236 ( .A(i_data_FEalures[31]), .Q(n638) );
  INV2 U237 ( .A(i_data_FEalures[17]), .Q(n708) );
  INV3 U238 ( .A(i_data_FEalures[8]), .Q(n746) );
  INV2 U239 ( .A(i_con_Efbmux[0]), .Q(n636) );
  INV2 U240 ( .A(i_con_Efamux[1]), .Q(n524) );
  INV2 U241 ( .A(i_data_immext[0]), .Q(n1205) );
  INV1 U242 ( .A(i_con_Efamux[2]), .Q(n527) );
  INV2 U243 ( .A(i_con_Efbmux[2]), .Q(n635) );
  INV3 U244 ( .A(i_data_FEalures[9]), .Q(n742) );
  INV3 U245 ( .A(i_con_Efbmux[1]), .Q(n632) );
  NOR21 U246 ( .A(i_con_Efbmux[2]), .B(i_con_Efbmux[0]), .Q(n633) );
  INV3 U247 ( .A(i_data_FEalures[12]), .Q(n730) );
  INV3 U248 ( .A(i_data_FEalures[10]), .Q(n738) );
  INV3 U249 ( .A(i_data_FEalures[16]), .Q(n714) );
  NAND41 U250 ( .A(n1055), .B(n1054), .C(n1053), .D(n1052), .Q(
        alu_o_data_AluRes[30]) );
  OAI211 U251 ( .A(n962), .B(n920), .C(n919), .Q(alu_o_data_AluRes[20]) );
  OAI211 U252 ( .A(n962), .B(n958), .C(n957), .Q(alu_o_data_AluRes[23]) );
  OAI211 U253 ( .A(n962), .B(n908), .C(n907), .Q(alu_o_data_AluRes[19]) );
  OAI211 U254 ( .A(n962), .B(n945), .C(n944), .Q(alu_o_data_AluRes[22]) );
  INV2 U255 ( .A(n1070), .Q(n977) );
  OAI211 U256 ( .A(n962), .B(n933), .C(n932), .Q(alu_o_data_AluRes[21]) );
  OAI211 U257 ( .A(n962), .B(n896), .C(n895), .Q(alu_o_data_AluRes[18]) );
  NAND22 U258 ( .A(n1069), .B(u_alu_pre_subb[8]), .Q(n970) );
  INV2 U259 ( .A(u_alu_N173), .Q(n860) );
  NAND21 U260 ( .A(u_alu_pre_subb[15]), .B(n1069), .Q(n1074) );
  NOR23 U261 ( .A(n861), .B(u_alu_sub_x_2_n2), .Q(n1069) );
  INV1 U262 ( .A(n1068), .Q(n230) );
  NAND20 U263 ( .A(u_alu_N168), .B(n859), .Q(n821) );
  NAND20 U264 ( .A(u_alu_N167), .B(n859), .Q(n824) );
  IMUX21 U265 ( .A(n227), .B(u_alu_pre_suba[11]), .S(n216), .Q(
        u_alu_pre_subb[11]) );
  NAND20 U266 ( .A(u_alu_N166), .B(n859), .Q(n791) );
  OAI221 U267 ( .A(n1143), .B(n1160), .C(n1161), .D(n1162), .Q(n1157) );
  IMUX21 U268 ( .A(n226), .B(u_alu_pre_suba[9]), .S(n214), .Q(
        u_alu_pre_subb[9]) );
  OAI2111 U269 ( .A(compare_i_data_rs[2]), .B(n1121), .C(n1122), .D(n1123), 
        .Q(alu_o_data_AluRes[2]) );
  OAI2111 U270 ( .A(compare_i_data_rs[1]), .B(n1135), .C(n1136), .D(n1137), 
        .Q(alu_o_data_AluRes[1]) );
  INV2 U271 ( .A(u_alu_pre_sum_3b[8]), .Q(n960) );
  OAI2111 U272 ( .A(compare_i_data_rs[4]), .B(n1109), .C(n1110), .D(n1111), 
        .Q(alu_o_data_AluRes[4]) );
  NAND21 U273 ( .A(u_alu_half_sub_7_), .B(n826), .Q(n801) );
  OAI211 U274 ( .A(n196), .B(n195), .C(n194), .Q(n197) );
  NAND21 U275 ( .A(u_alu_half_sub_6_), .B(n826), .Q(n804) );
  INV2 U276 ( .A(u_alu_pre_sum_3a[8]), .Q(n961) );
  INV2 U277 ( .A(u_alu_pre_sum_3a[7]), .Q(n958) );
  NAND21 U278 ( .A(u_alu_N201), .B(n519), .Q(n797) );
  AOI220 U279 ( .A(n1077), .B(u_alu_N231), .C(u_alu_N199), .D(n519), .Q(n803)
         );
  NAND21 U280 ( .A(u_alu_N195), .B(n519), .Q(n816) );
  AOI220 U281 ( .A(n1077), .B(u_alu_N234), .C(u_alu_N202), .D(n519), .Q(n790)
         );
  AOI220 U282 ( .A(n1077), .B(u_alu_N235), .C(u_alu_N203), .D(n519), .Q(n823)
         );
  NAND21 U283 ( .A(u_alu_N194), .B(n519), .Q(n819) );
  AOI220 U284 ( .A(u_alu_N197), .B(n519), .C(u_alu_sum_1_4_), .D(n859), .Q(
        n810) );
  AOI220 U285 ( .A(n1077), .B(u_alu_N232), .C(u_alu_N200), .D(n519), .Q(n800)
         );
  AOI220 U286 ( .A(n1077), .B(u_alu_N236), .C(u_alu_N204), .D(n519), .Q(n820)
         );
  NAND21 U287 ( .A(u_alu_N196), .B(n519), .Q(n813) );
  NAND21 U288 ( .A(u_alu_half_sub_5_), .B(n826), .Q(n807) );
  INV2 U289 ( .A(u_alu_pre_sum_3a[6]), .Q(n945) );
  AOI220 U290 ( .A(n1077), .B(u_alu_N230), .C(u_alu_N198), .D(n519), .Q(n806)
         );
  OAI311 U291 ( .A(i_con_bop[0]), .B(n1275), .C(compare_i_data_rs[31]), .D(
        n1274), .Q(o_con_ifbranch) );
  NAND21 U292 ( .A(u_alu_N215), .B(n519), .Q(n941) );
  NAND21 U293 ( .A(u_alu_N221), .B(n519), .Q(n1022) );
  NAND21 U294 ( .A(u_alu_N212), .B(n519), .Q(n904) );
  NAND21 U295 ( .A(u_alu_N213), .B(n519), .Q(n916) );
  NAND21 U296 ( .A(u_alu_N224), .B(n519), .Q(n1065) );
  NAND21 U297 ( .A(u_alu_N222), .B(n519), .Q(n1037) );
  NAND21 U298 ( .A(u_alu_N214), .B(n519), .Q(n929) );
  NAND21 U299 ( .A(u_alu_N220), .B(n519), .Q(n1011) );
  NAND21 U300 ( .A(u_alu_N216), .B(n519), .Q(n953) );
  NAND21 U301 ( .A(n1077), .B(u_alu_N226), .Q(n817) );
  NAND21 U302 ( .A(u_alu_N218), .B(n519), .Q(n985) );
  AOI220 U303 ( .A(u_alu_N210), .B(n519), .C(u_alu_N242), .D(n1077), .Q(n877)
         );
  NAND21 U304 ( .A(u_alu_N223), .B(n519), .Q(n1049) );
  MUX22 U305 ( .A(n274), .B(n353), .S(n372), .Q(u_alu_N212) );
  INV2 U306 ( .A(n314), .Q(n370) );
  INV2 U307 ( .A(n358), .Q(n368) );
  INV2 U308 ( .A(n359), .Q(n369) );
  INV2 U309 ( .A(n320), .Q(n371) );
  NAND21 U310 ( .A(u_alu_N243), .B(n1077), .Q(n892) );
  INV2 U311 ( .A(n357), .Q(n367) );
  MUX22 U312 ( .A(n269), .B(n336), .S(n372), .Q(u_alu_N211) );
  MUX22 U313 ( .A(n290), .B(n356), .S(n372), .Q(u_alu_N215) );
  MUX22 U314 ( .A(n280), .B(n354), .S(n372), .Q(u_alu_N213) );
  INV2 U315 ( .A(n356), .Q(n366) );
  INV2 U316 ( .A(n354), .Q(n364) );
  MUX22 U317 ( .A(n315), .B(n314), .S(n372), .Q(u_alu_N219) );
  NAND21 U318 ( .A(n1077), .B(u_alu_N228), .Q(n811) );
  AOI220 U319 ( .A(n826), .B(u_alu_half_sub_3_), .C(n859), .D(u_alu_sum_1_3_), 
        .Q(n812) );
  INV2 U320 ( .A(n353), .Q(n363) );
  MUX22 U321 ( .A(n321), .B(n320), .S(n372), .Q(u_alu_N220) );
  INV2 U322 ( .A(n355), .Q(n365) );
  NAND21 U323 ( .A(n1077), .B(u_alu_N227), .Q(n814) );
  INV2 U324 ( .A(n336), .Q(n362) );
  INV2 U325 ( .A(n275), .Q(n361) );
  AOI210 U326 ( .A(n1077), .B(u_alu_N253), .C(n1019), .Q(n1020) );
  OAI2111 U327 ( .A(n829), .B(compare_i_data_rs[0]), .C(n828), .D(n827), .Q(
        n1158) );
  NAND21 U328 ( .A(u_alu_N249), .B(n1077), .Q(n971) );
  MUX22 U329 ( .A(n378), .B(n414), .S(i_data_immext[10]), .Q(u_alu_N225) );
  MUX22 U330 ( .A(n295), .B(n357), .S(n372), .Q(u_alu_N216) );
  MUX22 U331 ( .A(n302), .B(n358), .S(n372), .Q(u_alu_N217) );
  AOI210 U332 ( .A(n1077), .B(u_alu_N256), .C(n1059), .Q(n1066) );
  AOI2111 U333 ( .A(n1056), .B(n71), .C(n874), .D(n873), .Q(n879) );
  AOI220 U334 ( .A(n859), .B(u_alu_sum_1_2_), .C(n826), .D(u_alu_half_sub_2_), 
        .Q(n815) );
  IMUX21 U335 ( .A(n377), .B(n489), .S(u_alu_ashr_4_SH_3_), .Q(n378) );
  INV2 U336 ( .A(n414), .Q(n500) );
  AOI210 U337 ( .A(n1077), .B(u_alu_N255), .C(n1046), .Q(n1047) );
  AOI220 U338 ( .A(n859), .B(u_alu_sum_1_1_), .C(n826), .D(u_alu_half_sub_1_), 
        .Q(n818) );
  OAI211 U339 ( .A(i_con_bop[2]), .B(n1270), .C(n1269), .Q(n1273) );
  NAND21 U340 ( .A(i_con_bop[1]), .B(n1270), .Q(n1271) );
  INV2 U341 ( .A(n476), .Q(n503) );
  NAND20 U342 ( .A(n1056), .B(alu_i_data_B[15]), .Q(n1057) );
  AOI210 U343 ( .A(n1056), .B(alu_i_data_B[10]), .C(n990), .Q(n991) );
  AOI210 U344 ( .A(n1056), .B(alu_i_data_B[13]), .C(n1029), .Q(n1030) );
  INV2 U345 ( .A(n490), .Q(n499) );
  INV2 U346 ( .A(n454), .Q(n497) );
  AOI220 U347 ( .A(n859), .B(u_alu_sum_1_0_), .C(n826), .D(u_alu_half_sub_0_), 
        .Q(n827) );
  INV2 U348 ( .A(n428), .Q(n502) );
  INV1 U349 ( .A(u_alu_pre_suba[2]), .Q(n222) );
  INV2 U350 ( .A(n465), .Q(n506) );
  INV2 U351 ( .A(n494), .Q(n501) );
  NAND20 U352 ( .A(n1056), .B(alu_i_data_B[12]), .Q(n1018) );
  AOI210 U353 ( .A(n1056), .B(alu_i_data_B[11]), .C(n1003), .Q(n1004) );
  INV2 U354 ( .A(n444), .Q(n507) );
  OAI211 U355 ( .A(n170), .B(n169), .C(n178), .Q(n171) );
  INV2 U356 ( .A(n446), .Q(n504) );
  NAND20 U357 ( .A(n1056), .B(alu_i_data_B[14]), .Q(n1045) );
  INV2 U358 ( .A(u_alu_pre_sum_3a[1]), .Q(n883) );
  NOR20 U359 ( .A(n372), .B(n456), .Q(u_alu_N255) );
  MUX21 U360 ( .A(n395), .B(n394), .S(i_data_immext[8]), .Q(n432) );
  IMUX20 U361 ( .A(n262), .B(n261), .S(i_data_immext[8]), .Q(n308) );
  NOR40 U362 ( .A(n1264), .B(n1263), .C(n1262), .D(n1261), .Q(n1265) );
  INV2 U363 ( .A(u_alu_pre_subb[0]), .Q(n221) );
  ADD32 U364 ( .A(n74), .B(compare_i_data_rs[17]), .CI(
        u_alu_DP_OP_85J3_126_1427_n46), .CO(u_alu_DP_OP_85J3_126_1427_n45), 
        .S(u_alu_pre_suba[1]) );
  NOR20 U365 ( .A(i_data_immext[8]), .B(n498), .Q(n431) );
  IMUX20 U366 ( .A(n250), .B(n252), .S(i_data_immext[8]), .Q(n272) );
  NOR20 U367 ( .A(i_data_immext[8]), .B(n496), .Q(n436) );
  NOR20 U368 ( .A(i_data_immext[8]), .B(n505), .Q(n439) );
  NOR20 U369 ( .A(n372), .B(n457), .Q(u_alu_N256) );
  INV1 U370 ( .A(n188), .Q(n204) );
  IMUX21 U371 ( .A(n468), .B(n393), .S(i_data_immext[8]), .Q(n489) );
  INV2 U372 ( .A(n133), .Q(n205) );
  INV1 U373 ( .A(n430), .Q(n498) );
  INV2 U374 ( .A(n183), .Q(n203) );
  NOR21 U375 ( .A(i_data_immext[10]), .B(n360), .Q(u_alu_N193) );
  INV3 U376 ( .A(n71), .Q(n83) );
  INV2 U377 ( .A(n190), .Q(n206) );
  INV1 U378 ( .A(n435), .Q(n496) );
  INV1 U379 ( .A(n438), .Q(n505) );
  ADD22 U380 ( .A(compare_i_data_rs[16]), .B(alu_i_data_B[16]), .CO(
        u_alu_DP_OP_83J3_124_3384_n15), .S(u_alu_pre_sum_3a[0]) );
  NAND21 U381 ( .A(n793), .B(alu_i_con_AluCtrl[3]), .Q(n795) );
  INV2 U382 ( .A(n257), .Q(n360) );
  NAND21 U383 ( .A(alu_i_con_AluCtrl[3]), .B(n231), .Q(n783) );
  XNR20 U384 ( .A(compare_i_data_rs[27]), .B(alu_i_data_B[27]), .Q(n1005) );
  NOR20 U385 ( .A(n374), .B(n237), .Q(n238) );
  NOR20 U386 ( .A(compare_i_data_rs[28]), .B(alu_i_data_B[28]), .Q(n1017) );
  INV2 U387 ( .A(alu_i_data_B[31]), .Q(n1058) );
  NAND21 U388 ( .A(alu_i_data_B[31]), .B(n510), .Q(n404) );
  INV2 U389 ( .A(n229), .Q(n121) );
  NOR20 U390 ( .A(compare_i_data_rs[30]), .B(alu_i_data_B[30]), .Q(n1044) );
  INV3 U391 ( .A(alu_i_data_B[25]), .Q(n88) );
  INV3 U392 ( .A(alu_i_data_B[24]), .Q(n89) );
  INV3 U393 ( .A(alu_i_data_B[28]), .Q(n90) );
  INV1 U394 ( .A(compare_i_data_rs[7]), .Q(n844) );
  NAND21 U395 ( .A(compare_i_data_rt[18]), .B(n711), .Q(n706) );
  NAND21 U396 ( .A(compare_i_data_rt[25]), .B(n711), .Q(n671) );
  NAND21 U397 ( .A(compare_i_data_rt[24]), .B(n711), .Q(n676) );
  INV1 U398 ( .A(alu_i_con_AluCtrl[2]), .Q(n785) );
  NAND21 U399 ( .A(alu_i_data_B[0]), .B(n510), .Q(n237) );
  INV3 U400 ( .A(alu_i_data_B[11]), .Q(n91) );
  NAND31 U401 ( .A(i_con_bop[2]), .B(compare_i_data_rs[31]), .C(n1268), .Q(
        n1269) );
  INV2 U402 ( .A(alu_i_data_B[7]), .Q(n92) );
  INV2 U403 ( .A(compare_i_data_rs[21]), .Q(n924) );
  INV2 U404 ( .A(alu_i_data_B[4]), .Q(n93) );
  INV3 U405 ( .A(alu_i_data_B[12]), .Q(n94) );
  INV2 U406 ( .A(compare_i_data_rs[26]), .Q(n993) );
  INV2 U407 ( .A(compare_i_data_rs[27]), .Q(n1006) );
  INV2 U408 ( .A(alu_i_con_AluCtrl[3]), .Q(n784) );
  NAND21 U409 ( .A(compare_i_data_rt[19]), .B(n711), .Q(n701) );
  INV2 U410 ( .A(compare_i_data_rs[23]), .Q(n96) );
  INV3 U411 ( .A(compare_i_data_rs[4]), .Q(n841) );
  INV1 U412 ( .A(compare_i_data_rs[31]), .Q(n99) );
  INV2 U413 ( .A(compare_i_data_rs[12]), .Q(n853) );
  NAND21 U414 ( .A(compare_i_data_rt[28]), .B(n711), .Q(n656) );
  NAND21 U415 ( .A(compare_i_data_rt[29]), .B(n711), .Q(n651) );
  NAND21 U416 ( .A(compare_i_data_rt[27]), .B(n711), .Q(n661) );
  NAND21 U417 ( .A(compare_i_data_rt[26]), .B(n711), .Q(n666) );
  NAND21 U418 ( .A(compare_i_data_rt[30]), .B(n711), .Q(n646) );
  INV2 U419 ( .A(n1197), .Q(n1186) );
  OAI211 U420 ( .A(n517), .B(n1229), .C(n655), .Q(compare_i_data_rt[28]) );
  OAI211 U421 ( .A(n517), .B(n1231), .C(n645), .Q(compare_i_data_rt[30]) );
  OAI211 U422 ( .A(n517), .B(n1230), .C(n650), .Q(compare_i_data_rt[29]) );
  AOI211 U423 ( .A(n776), .B(i_data_rt[11]), .C(n735), .Q(n736) );
  AOI211 U424 ( .A(n776), .B(i_data_rt[13]), .C(n727), .Q(n728) );
  INV3 U425 ( .A(compare_i_data_rt[2]), .Q(n836) );
  OAI211 U426 ( .A(n517), .B(n1228), .C(n660), .Q(compare_i_data_rt[27]) );
  AOI211 U427 ( .A(n776), .B(i_data_rt[21]), .C(n689), .Q(n690) );
  INV3 U428 ( .A(compare_i_data_rt[3]), .Q(n843) );
  INV2 U429 ( .A(compare_i_data_rs[20]), .Q(n104) );
  INV2 U430 ( .A(compare_i_data_rs[6]), .Q(n105) );
  OAI211 U431 ( .A(n517), .B(n1232), .C(n640), .Q(compare_i_data_rt[31]) );
  AOI211 U432 ( .A(n776), .B(i_data_rt[15]), .C(n719), .Q(n720) );
  AOI221 U433 ( .A(n1185), .B(n1198), .C(i_con_Ealuop[0]), .D(i_con_Ealuop[5]), 
        .Q(n1197) );
  AOI211 U434 ( .A(n776), .B(i_data_rt[14]), .C(n723), .Q(n724) );
  INV2 U435 ( .A(compare_i_data_rs[8]), .Q(n107) );
  OAI211 U436 ( .A(n1200), .B(n1199), .C(n1198), .Q(n1201) );
  AOI211 U437 ( .A(n776), .B(i_data_rt[24]), .C(n674), .Q(n675) );
  INV3 U438 ( .A(compare_i_data_rs[10]), .Q(n108) );
  AOI211 U439 ( .A(n776), .B(i_data_rt[23]), .C(n679), .Q(n680) );
  AOI211 U440 ( .A(n776), .B(i_data_rt[22]), .C(n684), .Q(n685) );
  INV2 U441 ( .A(compare_i_data_rs[22]), .Q(n109) );
  INV2 U442 ( .A(compare_i_data_rs[24]), .Q(n110) );
  AOI211 U443 ( .A(n776), .B(i_data_rt[10]), .C(n739), .Q(n740) );
  OAI211 U444 ( .A(n517), .B(n1227), .C(n665), .Q(compare_i_data_rt[26]) );
  AOI211 U445 ( .A(n776), .B(i_data_rt[25]), .C(n669), .Q(n670) );
  AOI211 U446 ( .A(n776), .B(i_data_rt[12]), .C(n731), .Q(n732) );
  NAND31 U447 ( .A(n769), .B(n768), .C(n767), .Q(compare_i_data_rt[3]) );
  INV2 U448 ( .A(n1184), .Q(n1185) );
  NAND31 U449 ( .A(n781), .B(n780), .C(n779), .Q(compare_i_data_rt[0]) );
  NAND31 U450 ( .A(n772), .B(n771), .C(n770), .Q(compare_i_data_rt[2]) );
  AOI311 U451 ( .A(i_data_immext[5]), .B(n1209), .C(n1207), .D(n1183), .Q(
        n1192) );
  OAI211 U452 ( .A(n1195), .B(n1194), .C(n1198), .Q(n1196) );
  OAI211 U453 ( .A(n516), .B(n742), .C(n741), .Q(n743) );
  OAI211 U454 ( .A(n516), .B(n750), .C(n749), .Q(n751) );
  OAI211 U455 ( .A(n516), .B(n708), .C(n707), .Q(n709) );
  OAI211 U456 ( .A(n512), .B(n742), .C(n595), .Q(n596) );
  OAI211 U457 ( .A(n512), .B(n746), .C(n598), .Q(n599) );
  OAI211 U458 ( .A(n516), .B(n730), .C(n729), .Q(n731) );
  OAI211 U459 ( .A(n516), .B(n714), .C(n713), .Q(n715) );
  OAI211 U460 ( .A(n512), .B(n738), .C(n592), .Q(n593) );
  OAI211 U461 ( .A(n516), .B(n746), .C(n745), .Q(n747) );
  OAI212 U462 ( .A(n512), .B(n638), .C(n529), .Q(n530) );
  OAI211 U463 ( .A(n512), .B(n754), .C(n604), .Q(n605) );
  OAI211 U464 ( .A(n516), .B(n703), .C(n702), .Q(n704) );
  OAI211 U465 ( .A(n516), .B(n722), .C(n721), .Q(n723) );
  OAI211 U466 ( .A(n512), .B(n714), .C(n574), .Q(n575) );
  OAI211 U467 ( .A(n516), .B(n693), .C(n692), .Q(n694) );
  OAI211 U468 ( .A(n516), .B(n754), .C(n753), .Q(n755) );
  AOI221 U469 ( .A(n778), .B(i_data_FMmemout[1]), .C(n518), .D(
        i_data_FWmemout[1]), .Q(n773) );
  AOI221 U470 ( .A(n778), .B(i_data_FMmemout[0]), .C(n518), .D(
        i_data_FWmemout[0]), .Q(n779) );
  NAND21 U471 ( .A(n776), .B(i_data_rt[3]), .Q(n769) );
  AOI221 U472 ( .A(n778), .B(i_data_FMmemout[2]), .C(n518), .D(
        i_data_FWmemout[2]), .Q(n770) );
  OAI211 U473 ( .A(n516), .B(n718), .C(n717), .Q(n719) );
  OAI211 U474 ( .A(n512), .B(n730), .C(n586), .Q(n587) );
  OAI211 U475 ( .A(n516), .B(n758), .C(n757), .Q(n759) );
  OAI211 U476 ( .A(n516), .B(n688), .C(n687), .Q(n689) );
  OAI211 U477 ( .A(n512), .B(n758), .C(n607), .Q(n608) );
  OAI211 U478 ( .A(n516), .B(n738), .C(n737), .Q(n739) );
  OAI211 U479 ( .A(n512), .B(n762), .C(n610), .Q(n612) );
  OAI211 U480 ( .A(n516), .B(n678), .C(n677), .Q(n679) );
  OAI211 U481 ( .A(n516), .B(n673), .C(n672), .Q(n674) );
  OAI211 U482 ( .A(n516), .B(n683), .C(n682), .Q(n684) );
  OAI211 U483 ( .A(n516), .B(n734), .C(n733), .Q(n735) );
  OAI211 U484 ( .A(n516), .B(n726), .C(n725), .Q(n727) );
  OAI211 U485 ( .A(n516), .B(n762), .C(n761), .Q(n764) );
  OAI211 U486 ( .A(n512), .B(n734), .C(n589), .Q(n590) );
  INV3 U487 ( .A(n614), .Q(n515) );
  INV3 U488 ( .A(n766), .Q(n518) );
  AOI311 U489 ( .A(i_con_Ealuop[3]), .B(i_con_Ealuop[2]), .C(n1178), .D(n1189), 
        .Q(n1202) );
  INV2 U490 ( .A(n1173), .Q(n1174) );
  INV2 U491 ( .A(n1193), .Q(n1194) );
  INV2 U492 ( .A(n1167), .Q(n1168) );
  NAND21 U493 ( .A(n1172), .B(n1205), .Q(n1170) );
  IMUX21 U494 ( .A(n1167), .B(i_data_immext[5]), .S(n1207), .Q(n1175) );
  AOI211 U495 ( .A(i_con_Ealuop[1]), .B(n1177), .C(n1203), .Q(n1189) );
  OAI211 U496 ( .A(i_con_Ealuop[5]), .B(n1180), .C(i_con_Ealuop[0]), .Q(n1181)
         );
  NAND21 U497 ( .A(i_data_immext[0]), .B(n1172), .Q(n1193) );
  NOR21 U498 ( .A(i_con_Ealuop[2]), .B(n1179), .Q(n1180) );
  AOI2111 U499 ( .A(i_data_immext[2]), .B(n1210), .C(i_data_immext[3]), .D(
        n1206), .Q(n1195) );
  INV2 U500 ( .A(u_alu_ashr_4_SH_3_), .Q(n508) );
  NOR21 U501 ( .A(i_con_Ealuop[4]), .B(n1203), .Q(n1178) );
  NOR21 U502 ( .A(n1187), .B(i_con_Ealuop[0]), .Q(n1198) );
  NAND21 U503 ( .A(i_data_immext[5]), .B(n1165), .Q(n1167) );
  NAND21 U504 ( .A(n1210), .B(n1207), .Q(n1166) );
  INV2 U505 ( .A(i_data_FEalures[24]), .Q(n673) );
  INV3 U506 ( .A(i_data_FWmemout[8]), .Q(n1237) );
  INV2 U507 ( .A(i_data_FEalures[30]), .Q(n643) );
  INV2 U508 ( .A(i_data_FEalures[27]), .Q(n658) );
  INV3 U509 ( .A(i_data_FEalures[5]), .Q(n758) );
  INV2 U510 ( .A(i_data_FEalures[19]), .Q(n698) );
  INV2 U511 ( .A(i_data_FEalures[25]), .Q(n668) );
  INV3 U512 ( .A(i_data_FWmemout[19]), .Q(n1220) );
  INV3 U513 ( .A(i_data_FWmemout[18]), .Q(n1219) );
  INV3 U514 ( .A(i_con_Ealuop[1]), .Q(n1187) );
  INV3 U515 ( .A(i_data_FWmemout[20]), .Q(n1221) );
  INV3 U516 ( .A(i_data_FWmemout[17]), .Q(n1218) );
  INV2 U517 ( .A(i_data_FEalures[20]), .Q(n693) );
  INV3 U518 ( .A(i_data_FEalures[7]), .Q(n750) );
  INV2 U519 ( .A(i_con_Ealuop[3]), .Q(n1179) );
  INV3 U520 ( .A(i_data_FWmemout[27]), .Q(n1228) );
  INV3 U521 ( .A(i_data_FWmemout[24]), .Q(n1225) );
  INV3 U522 ( .A(i_data_FWmemout[31]), .Q(n1232) );
  INV3 U523 ( .A(i_con_Ealuop[0]), .Q(n1203) );
  INV2 U524 ( .A(i_data_FEalures[26]), .Q(n663) );
  INV1 U525 ( .A(i_con_Ealuop[2]), .Q(n1176) );
  INV3 U526 ( .A(i_data_FWmemout[9]), .Q(n1238) );
  INV3 U527 ( .A(i_data_FWmemout[10]), .Q(n1211) );
  INV3 U528 ( .A(i_data_FWmemout[25]), .Q(n1226) );
  INV3 U529 ( .A(i_data_FWmemout[12]), .Q(n1213) );
  INV2 U530 ( .A(i_data_FEalures[18]), .Q(n703) );
  INV3 U531 ( .A(i_data_FEalures[14]), .Q(n722) );
  INV3 U532 ( .A(i_data_FWmemout[14]), .Q(n1215) );
  INV3 U533 ( .A(i_data_FEalures[6]), .Q(n754) );
  INV2 U534 ( .A(i_con_Ealuop[4]), .Q(n1204) );
  INV3 U535 ( .A(i_data_FWmemout[6]), .Q(n1235) );
  INV3 U536 ( .A(i_data_FWmemout[7]), .Q(n1236) );
  INV3 U537 ( .A(i_data_FWmemout[16]), .Q(n1217) );
  INV3 U538 ( .A(i_data_FWmemout[26]), .Q(n1227) );
  INV3 U539 ( .A(i_data_FWmemout[23]), .Q(n1224) );
  INV3 U540 ( .A(i_data_FEalures[15]), .Q(n718) );
  INV3 U541 ( .A(i_con_Malupc8), .Q(n1244) );
  INV3 U542 ( .A(i_data_FEalures[11]), .Q(n734) );
  INV3 U543 ( .A(i_data_FWmemout[21]), .Q(n1222) );
  INV3 U544 ( .A(i_data_FEalures[13]), .Q(n726) );
  INV3 U545 ( .A(i_data_FWmemout[28]), .Q(n1229) );
  INV2 U546 ( .A(i_data_FEalures[29]), .Q(n648) );
  INV2 U547 ( .A(i_data_FEalures[21]), .Q(n688) );
  BUF6 U548 ( .A(i_data_immext[9]), .Q(u_alu_ashr_4_SH_3_) );
  INV3 U549 ( .A(i_data_FWmemout[22]), .Q(n1223) );
  INV3 U550 ( .A(i_data_FEalures[4]), .Q(n762) );
  INV2 U551 ( .A(i_data_FEalures[28]), .Q(n653) );
  INV3 U552 ( .A(i_data_FWmemout[13]), .Q(n1214) );
  INV3 U553 ( .A(i_data_FWmemout[29]), .Q(n1230) );
  INV3 U554 ( .A(i_data_FWmemout[5]), .Q(n1234) );
  INV3 U555 ( .A(i_data_FWmemout[30]), .Q(n1231) );
  INV3 U556 ( .A(i_data_FWmemout[11]), .Q(n1212) );
  INV1 U557 ( .A(i_con_bop[1]), .Q(n1268) );
  INV3 U558 ( .A(i_data_FWmemout[15]), .Q(n1216) );
  INV3 U559 ( .A(i_data_FWmemout[4]), .Q(n1233) );
  BUF6 U560 ( .A(i_data_immext[10]), .Q(n372) );
  INV3 U561 ( .A(DP_OP_77J3_127_5954_n10), .Q(n119) );
  INV3 U562 ( .A(DP_OP_77J3_127_5954_n11), .Q(n118) );
  INV3 U563 ( .A(DP_OP_77J3_127_5954_n12), .Q(n117) );
  INV3 U564 ( .A(DP_OP_77J3_127_5954_n13), .Q(n116) );
  INV3 U565 ( .A(DP_OP_77J3_127_5954_n14), .Q(n115) );
  INV3 U566 ( .A(DP_OP_77J3_127_5954_n15), .Q(n114) );
  INV3 U567 ( .A(DP_OP_77J3_127_5954_n16), .Q(n113) );
  INV3 U568 ( .A(DP_OP_77J3_127_5954_n17), .Q(n112) );
  ADD32 U569 ( .A(n118), .B(alu_i_data_B[14]), .CI(DP_OP_77J3_127_5954_n3), 
        .CO(DP_OP_77J3_127_5954_n2), .S(u_alu_N171) );
  ADD32 U570 ( .A(n119), .B(alu_i_data_B[15]), .CI(DP_OP_77J3_127_5954_n2), 
        .CO(DP_OP_77J3_127_5954_n1), .S(u_alu_N172) );
  ADD32 U571 ( .A(n116), .B(alu_i_data_B[12]), .CI(DP_OP_77J3_127_5954_n5), 
        .CO(DP_OP_77J3_127_5954_n4), .S(u_alu_N169) );
  ADD32 U572 ( .A(n117), .B(alu_i_data_B[13]), .CI(DP_OP_77J3_127_5954_n4), 
        .CO(DP_OP_77J3_127_5954_n3), .S(u_alu_N170) );
  ADD22 U573 ( .A(compare_i_data_rs[0]), .B(alu_i_data_B[0]), .CO(
        u_alu_add_x_1_n8), .S(u_alu_sum_1_0_) );
  ADD32 U574 ( .A(compare_i_data_rs[6]), .B(alu_i_data_B[6]), .CI(
        u_alu_add_x_1_n3), .CO(u_alu_add_x_1_n2), .S(u_alu_sum_1_6_) );
  ADD32 U575 ( .A(compare_i_data_rs[7]), .B(alu_i_data_B[7]), .CI(
        u_alu_add_x_1_n2), .CO(u_alu_sum_1_8_), .S(u_alu_sum_1_7_) );
  INV3 U576 ( .A(alu_i_data_B[14]), .Q(n127) );
  INV3 U577 ( .A(alu_i_data_B[13]), .Q(n126) );
  IMUX20 U578 ( .A(n128), .B(compare_i_data_rs[0]), .S(alu_i_data_B[0]), .Q(
        u_alu_half_sub_0_) );
  INV3 U579 ( .A(alu_i_data_B[10]), .Q(n125) );
  INV3 U580 ( .A(alu_i_data_B[9]), .Q(n124) );
  NAND22 U581 ( .A(alu_i_data_B[0]), .B(n128), .Q(u_alu_sub_x_2_n17) );
  ADD32 U582 ( .A(n92), .B(compare_i_data_rs[7]), .CI(u_alu_sub_x_2_n11), .CO(
        u_alu_sub_x_2_n10), .S(u_alu_half_sub_7_) );
  ADD32 U583 ( .A(n75), .B(compare_i_data_rs[8]), .CI(u_alu_sub_x_2_n10), .CO(
        u_alu_sub_x_2_n9), .S(u_alu_half_sub_8_) );
  ADD32 U584 ( .A(n125), .B(compare_i_data_rs[10]), .CI(u_alu_sub_x_2_n8), 
        .CO(u_alu_sub_x_2_n7), .S(u_alu_half_sub_10_) );
  ADD32 U585 ( .A(n91), .B(compare_i_data_rs[11]), .CI(u_alu_sub_x_2_n7), .CO(
        u_alu_sub_x_2_n6), .S(u_alu_half_sub_11_) );
  MAJ31 U586 ( .A(alu_i_data_B[25]), .B(n102), .C(n132), .Q(n135) );
  MAJ31 U587 ( .A(alu_i_data_B[31]), .B(n99), .C(n137), .Q(n138) );
  NOR20 U588 ( .A(alu_i_data_B[17]), .B(n98), .Q(n181) );
  OAI220 U589 ( .A(n96), .B(alu_i_data_B[23]), .C(n109), .D(alu_i_data_B[22]), 
        .Q(n188) );
  NOR20 U590 ( .A(alu_i_data_B[19]), .B(n103), .Q(n143) );
  OAI210 U591 ( .A(alu_i_data_B[16]), .B(n81), .C(n184), .Q(n180) );
  OAI220 U592 ( .A(alu_i_data_B[11]), .B(n97), .C(alu_i_data_B[10]), .D(n108), 
        .Q(n167) );
  AOI2110 U593 ( .A(compare_i_data_rs[8]), .B(n75), .C(n146), .D(n167), .Q(
        n177) );
  NAND20 U594 ( .A(compare_i_data_rs[7]), .B(n92), .Q(n147) );
  OAI210 U595 ( .A(alu_i_data_B[6]), .B(n105), .C(n147), .Q(n162) );
  NOR20 U596 ( .A(alu_i_data_B[5]), .B(n201), .Q(n155) );
  NOR20 U597 ( .A(n229), .B(n200), .Q(n148) );
  AOI210 U598 ( .A(compare_i_data_rs[2]), .B(n95), .C(n148), .Q(n153) );
  OAI210 U599 ( .A(n71), .B(n199), .C(alu_i_data_B[0]), .Q(n149) );
  OAI220 U600 ( .A(compare_i_data_rs[0]), .B(n149), .C(compare_i_data_rs[1]), 
        .D(n83), .Q(n152) );
  NOR20 U601 ( .A(compare_i_data_rs[2]), .B(n95), .Q(n150) );
  MAJ31 U602 ( .A(n229), .B(n200), .C(n150), .Q(n151) );
  AOI2110 U603 ( .A(compare_i_data_rs[4]), .B(n93), .C(n155), .D(n154), .Q(
        n158) );
  NOR20 U604 ( .A(compare_i_data_rs[4]), .B(n93), .Q(n156) );
  MAJ31 U605 ( .A(alu_i_data_B[5]), .B(n201), .C(n156), .Q(n157) );
  NAND20 U606 ( .A(alu_i_data_B[6]), .B(n105), .Q(n159) );
  MAJ31 U607 ( .A(compare_i_data_rs[7]), .B(n92), .C(n159), .Q(n160) );
  MAJ31 U608 ( .A(compare_i_data_rs[15]), .B(n80), .C(n164), .Q(n172) );
  IMAJ30 U609 ( .A(n91), .B(compare_i_data_rs[11]), .C(n165), .Q(n170) );
  NOR40 U610 ( .A(n181), .B(n185), .C(n180), .D(n179), .Q(n196) );
  NAND20 U611 ( .A(alu_i_data_B[20]), .B(n104), .Q(n182) );
  MAJ31 U612 ( .A(compare_i_data_rs[21]), .B(n72), .C(n182), .Q(n189) );
  NOR40 U613 ( .A(n193), .B(n192), .C(n191), .D(n206), .Q(n194) );
  INV0 U614 ( .A(compare_i_data_rs[9]), .Q(n202) );
  INV0 U615 ( .A(compare_i_data_rs[5]), .Q(n201) );
  INV0 U616 ( .A(compare_i_data_rs[3]), .Q(n200) );
  INV0 U617 ( .A(compare_i_data_rs[1]), .Q(n199) );
  AOI211 U618 ( .A(n190), .B(n135), .C(n134), .Q(n136) );
  NOR21 U619 ( .A(n191), .B(n136), .Q(n139) );
  AOI2111 U620 ( .A(n141), .B(n140), .C(n139), .D(n138), .Q(n198) );
  AOI211 U621 ( .A(n153), .B(n152), .C(n151), .Q(n154) );
  NOR21 U622 ( .A(n158), .B(n157), .Q(n161) );
  NOR21 U623 ( .A(n168), .B(n167), .Q(n169) );
  OAI2111 U624 ( .A(n174), .B(n173), .C(n172), .D(n171), .Q(n175) );
  AOI311 U625 ( .A(n178), .B(n177), .C(n176), .D(n175), .Q(n179) );
  OAI2111 U626 ( .A(n189), .B(n188), .C(n187), .D(n186), .Q(n195) );
  NAND22 U627 ( .A(n198), .B(n197), .Q(u_alu_N306) );
  AOI211 U628 ( .A(compare_i_data_rs[30]), .B(n77), .C(n129), .Q(n141) );
  OAI2111 U629 ( .A(alu_i_data_B[28]), .B(n101), .C(n141), .D(n131), .Q(n191)
         );
  AOI221 U630 ( .A(n76), .B(compare_i_data_rs[27]), .C(n78), .D(
        compare_i_data_rs[26]), .Q(n190) );
  OAI2111 U631 ( .A(alu_i_data_B[20]), .B(n104), .C(n204), .D(n142), .Q(n185)
         );
  AOI211 U632 ( .A(compare_i_data_rs[18]), .B(n73), .C(n143), .Q(n184) );
  IMAJ30 U633 ( .A(n79), .B(compare_i_data_rs[29]), .C(n130), .Q(n140) );
  NAND20 U634 ( .A(compare_i_data_rs[15]), .B(n80), .Q(n144) );
  AOI2110 U635 ( .A(compare_i_data_rs[12]), .B(n94), .C(n145), .D(n173), .Q(
        n178) );
  NOR20 U636 ( .A(alu_i_data_B[9]), .B(n202), .Q(n146) );
  NOR20 U637 ( .A(n94), .B(compare_i_data_rs[12]), .Q(n163) );
  NAND20 U638 ( .A(n108), .B(alu_i_data_B[10]), .Q(n165) );
  NOR20 U639 ( .A(n75), .B(compare_i_data_rs[8]), .Q(n166) );
  IMAJ30 U640 ( .A(n202), .B(alu_i_data_B[9]), .C(n166), .Q(n168) );
  NAND20 U641 ( .A(alu_i_data_B[22]), .B(n109), .Q(n183) );
  XOR21 U642 ( .A(u_alu_pre_sum_3a[8]), .B(u_alu_DP_OP_83J3_124_3384_n1), .Q(
        u_alu_pre_sum_3b[8]) );
  XOR31 U643 ( .A(alu_i_data_B[31]), .B(u_alu_DP_OP_84J3_125_2615_n9), .C(
        compare_i_data_rs[31]), .Q(u_alu_pre_sum_4a[7]) );
  OAI210 U644 ( .A(n220), .B(u_alu_pre_suba[14]), .C(u_alu_pre_suba[15]), .Q(
        n219) );
  XNR21 U645 ( .A(u_alu_pre_suba[14]), .B(n220), .Q(u_alu_pre_subb[14]) );
  XNR31 U646 ( .A(alu_i_data_B[31]), .B(u_alu_DP_OP_85J3_126_1427_n32), .C(
        compare_i_data_rs[31]), .Q(u_alu_pre_suba[15]) );
  XNR21 U647 ( .A(alu_i_data_B[16]), .B(compare_i_data_rs[16]), .Q(
        u_alu_pre_subb[0]) );
  XNR21 U648 ( .A(u_alu_pre_suba[10]), .B(n215), .Q(u_alu_pre_subb[10]) );
  XNR21 U649 ( .A(u_alu_pre_suba[12]), .B(n217), .Q(u_alu_pre_subb[12]) );
  XNR21 U650 ( .A(u_alu_pre_suba[8]), .B(n213), .Q(u_alu_pre_subb[8]) );
  XNR21 U651 ( .A(u_alu_pre_suba[6]), .B(n211), .Q(u_alu_pre_subb[6]) );
  XNR21 U652 ( .A(u_alu_pre_suba[4]), .B(n209), .Q(u_alu_pre_subb[4]) );
  NAND22 U653 ( .A(alu_i_data_B[16]), .B(n81), .Q(
        u_alu_DP_OP_85J3_126_1427_n46) );
  NOR31 U654 ( .A(u_alu_pre_suba[2]), .B(u_alu_pre_suba[1]), .C(n221), .Q(n208) );
  NAND22 U655 ( .A(n208), .B(n223), .Q(n209) );
  NOR21 U656 ( .A(u_alu_pre_suba[4]), .B(n209), .Q(n210) );
  INV3 U657 ( .A(u_alu_pre_suba[5]), .Q(n224) );
  NAND22 U658 ( .A(n210), .B(n224), .Q(n211) );
  NOR21 U659 ( .A(u_alu_pre_suba[6]), .B(n211), .Q(n212) );
  NAND22 U660 ( .A(n212), .B(n225), .Q(n213) );
  NOR21 U661 ( .A(u_alu_pre_suba[8]), .B(n213), .Q(n214) );
  NAND22 U662 ( .A(n214), .B(n226), .Q(n215) );
  NOR21 U663 ( .A(u_alu_pre_suba[10]), .B(n215), .Q(n216) );
  INV3 U664 ( .A(u_alu_pre_suba[11]), .Q(n227) );
  NAND22 U665 ( .A(n216), .B(n227), .Q(n217) );
  NOR21 U666 ( .A(u_alu_pre_suba[12]), .B(n217), .Q(n218) );
  INV3 U667 ( .A(u_alu_pre_suba[13]), .Q(n228) );
  NAND22 U668 ( .A(n218), .B(n228), .Q(n220) );
  OAI311 U669 ( .A(n220), .B(u_alu_pre_suba[14]), .C(u_alu_pre_suba[15]), .D(
        n219), .Q(u_alu_pre_subb[15]) );
  NOR21 U670 ( .A(u_alu_pre_suba[1]), .B(n221), .Q(n207) );
  IMUX21 U671 ( .A(n222), .B(u_alu_pre_suba[2]), .S(n207), .Q(
        u_alu_pre_subb[2]) );
  IMUX21 U672 ( .A(n224), .B(u_alu_pre_suba[5]), .S(n210), .Q(
        u_alu_pre_subb[5]) );
  IMUX21 U673 ( .A(n223), .B(u_alu_pre_suba[3]), .S(n208), .Q(
        u_alu_pre_subb[3]) );
  IMUX21 U674 ( .A(n225), .B(u_alu_pre_suba[7]), .S(n212), .Q(
        u_alu_pre_subb[7]) );
  IMUX21 U675 ( .A(n228), .B(u_alu_pre_suba[13]), .S(n218), .Q(
        u_alu_pre_subb[13]) );
  OAI2111 U676 ( .A(compare_i_data_rs[3]), .B(n1114), .C(n1115), .D(n1116), 
        .Q(alu_o_data_AluRes[3]) );
  AOI210 U677 ( .A(alu_i_con_AluCtrl[0]), .B(n1157), .C(n1158), .Q(n1156) );
  AOI220 U678 ( .A(n1077), .B(u_alu_N233), .C(n82), .D(alu_i_data_B[8]), .Q(
        n799) );
  IMUX21 U679 ( .A(n416), .B(n415), .S(i_data_immext[8]), .Q(n492) );
  IMUX21 U680 ( .A(n410), .B(n413), .S(i_data_immext[8]), .Q(n422) );
  OAI310 U681 ( .A(alu_i_data_B[23]), .B(compare_i_data_rs[23]), .C(n1060), 
        .D(n947), .Q(n950) );
  IMUX21 U682 ( .A(n440), .B(n439), .S(u_alu_ashr_4_SH_3_), .Q(n486) );
  IMUX21 U683 ( .A(n400), .B(n403), .S(n374), .Q(n413) );
  IMUX21 U684 ( .A(n406), .B(n409), .S(i_data_immext[8]), .Q(n420) );
  IMUX21 U685 ( .A(n432), .B(n431), .S(u_alu_ashr_4_SH_3_), .Q(n470) );
  IMUX21 U686 ( .A(n437), .B(n436), .S(u_alu_ashr_4_SH_3_), .Q(n481) );
  IMUX21 U687 ( .A(n386), .B(n385), .S(n374), .Q(n409) );
  IMUX21 U688 ( .A(n415), .B(n418), .S(i_data_immext[8]), .Q(n434) );
  IMUX21 U689 ( .A(n401), .B(n400), .S(n374), .Q(n415) );
  OAI310 U690 ( .A(alu_i_data_B[24]), .B(compare_i_data_rs[24]), .C(n1060), 
        .D(n967), .Q(n968) );
  AOI210 U691 ( .A(n521), .B(compare_i_data_rs[24]), .C(n82), .Q(n965) );
  IMUX21 U692 ( .A(n255), .B(n238), .S(i_data_immext[8]), .Q(n279) );
  IMUX21 U693 ( .A(n254), .B(n256), .S(i_data_immext[8]), .Q(n278) );
  IMUX21 U694 ( .A(n248), .B(n247), .S(i_data_immext[8]), .Q(n289) );
  IMUX21 U695 ( .A(n266), .B(n246), .S(i_data_immext[8]), .Q(n288) );
  IMUX21 U696 ( .A(n256), .B(n255), .S(i_data_immext[8]), .Q(n301) );
  IMUX21 U697 ( .A(n236), .B(n235), .S(n374), .Q(n255) );
  IMUX21 U698 ( .A(n234), .B(n233), .S(n374), .Q(n256) );
  IMUX21 U699 ( .A(n394), .B(n430), .S(i_data_immext[8]), .Q(n441) );
  IMUX21 U700 ( .A(n385), .B(n388), .S(n374), .Q(n394) );
  IMUX21 U701 ( .A(n392), .B(n395), .S(i_data_immext[8]), .Q(n488) );
  IMUX21 U702 ( .A(n408), .B(n435), .S(i_data_immext[8]), .Q(n419) );
  IMUX21 U703 ( .A(n388), .B(n387), .S(n374), .Q(n408) );
  OAI310 U704 ( .A(alu_i_data_B[26]), .B(compare_i_data_rs[26]), .C(n1060), 
        .D(n991), .Q(n995) );
  IMUX21 U705 ( .A(n235), .B(n237), .S(u_alu_ashr_4_SH_1_), .Q(n247) );
  IMUX21 U706 ( .A(n246), .B(n248), .S(i_data_immext[8]), .Q(n267) );
  IMUX21 U707 ( .A(n233), .B(n236), .S(n374), .Q(n248) );
  IMUX21 U708 ( .A(n232), .B(n234), .S(n374), .Q(n246) );
  NAND22 U709 ( .A(n1068), .B(u_alu_pre_suba[11]), .Q(n1010) );
  OAI310 U710 ( .A(alu_i_data_B[27]), .B(compare_i_data_rs[27]), .C(n1060), 
        .D(n1004), .Q(n1008) );
  IMUX21 U711 ( .A(n412), .B(n438), .S(i_data_immext[8]), .Q(n421) );
  IMUX21 U712 ( .A(n402), .B(n405), .S(n374), .Q(n412) );
  NAND22 U713 ( .A(n1068), .B(u_alu_pre_suba[13]), .Q(n1036) );
  IMUX21 U714 ( .A(n261), .B(n263), .S(i_data_immext[8]), .Q(n284) );
  IMUX21 U715 ( .A(n260), .B(n262), .S(i_data_immext[8]), .Q(n283) );
  OAI310 U716 ( .A(alu_i_data_B[29]), .B(compare_i_data_rs[29]), .C(n1060), 
        .D(n1030), .Q(n1034) );
  IMUX21 U717 ( .A(n241), .B(n240), .S(n374), .Q(n262) );
  OAI310 U718 ( .A(alu_i_data_B[25]), .B(compare_i_data_rs[25]), .C(n1060), 
        .D(n979), .Q(n982) );
  AOI210 U719 ( .A(n1056), .B(alu_i_data_B[9]), .C(n978), .Q(n979) );
  IMUX21 U720 ( .A(n418), .B(n417), .S(i_data_immext[8]), .Q(n442) );
  IMUX21 U721 ( .A(n405), .B(n404), .S(u_alu_ashr_4_SH_1_), .Q(n417) );
  IMUX21 U722 ( .A(n403), .B(n402), .S(n374), .Q(n418) );
  NOR22 U723 ( .A(n783), .B(n794), .Q(n1079) );
  IMUX21 U724 ( .A(n252), .B(n251), .S(i_data_immext[8]), .Q(n294) );
  IMUX21 U725 ( .A(n271), .B(n250), .S(i_data_immext[8]), .Q(n293) );
  IMUX21 U726 ( .A(n239), .B(n241), .S(n374), .Q(n250) );
  AOI221 U727 ( .A(n626), .B(i_data_FMmemout[0]), .C(n515), .D(
        i_data_FWmemout[0]), .Q(n627) );
  IMUX23 U728 ( .A(n852), .B(n1205), .S(n70), .Q(alu_i_data_B[0]) );
  AOI221 U729 ( .A(n625), .B(i_data_FMalures[3]), .C(n513), .D(
        i_data_FEalures[3]), .Q(n616) );
  AOI211 U730 ( .A(n624), .B(i_data_rs[6]), .C(n605), .Q(n606) );
  AOI211 U731 ( .A(n776), .B(i_data_rt[8]), .C(n747), .Q(n748) );
  AOI211 U732 ( .A(n776), .B(i_data_rt[9]), .C(n743), .Q(n744) );
  MUX22 U733 ( .A(compare_i_data_rt[12]), .B(i_data_immext[12]), .S(n70), .Q(
        alu_i_data_B[12]) );
  AOI211 U734 ( .A(n624), .B(i_data_rs[13]), .C(n584), .Q(n585) );
  MUX22 U735 ( .A(compare_i_data_rt[13]), .B(i_data_immext[13]), .S(n70), .Q(
        alu_i_data_B[13]) );
  MUX22 U736 ( .A(compare_i_data_rt[14]), .B(i_data_immext[14]), .S(n70), .Q(
        alu_i_data_B[14]) );
  OAI212 U737 ( .A(n517), .B(n1215), .C(n724), .Q(compare_i_data_rt[14]) );
  MUX22 U738 ( .A(compare_i_data_rt[15]), .B(i_data_immext[15]), .S(n70), .Q(
        alu_i_data_B[15]) );
  OAI212 U739 ( .A(n517), .B(n1216), .C(n720), .Q(compare_i_data_rt[15]) );
  AOI2111 U740 ( .A(i_data_immext[0]), .B(n1175), .C(n1199), .D(n1183), .Q(
        n1182) );
  AOI210 U741 ( .A(n624), .B(i_data_rs[16]), .C(n575), .Q(n576) );
  AOI211 U742 ( .A(n624), .B(i_data_rs[19]), .C(n566), .Q(n567) );
  AOI211 U743 ( .A(n776), .B(i_data_rt[20]), .C(n694), .Q(n695) );
  IMUX21 U744 ( .A(n492), .B(n442), .S(u_alu_ashr_4_SH_3_), .Q(n428) );
  IMUX21 U745 ( .A(n422), .B(n421), .S(u_alu_ashr_4_SH_3_), .Q(n465) );
  IMUX21 U746 ( .A(n420), .B(n419), .S(u_alu_ashr_4_SH_3_), .Q(n454) );
  IMUX21 U747 ( .A(n434), .B(n433), .S(u_alu_ashr_4_SH_3_), .Q(n476) );
  IMUX21 U748 ( .A(n301), .B(n300), .S(u_alu_ashr_4_SH_3_), .Q(n358) );
  IMUX21 U749 ( .A(n278), .B(n279), .S(u_alu_ashr_4_SH_3_), .Q(n327) );
  IMUX21 U750 ( .A(n288), .B(n289), .S(u_alu_ashr_4_SH_3_), .Q(n343) );
  IMUX21 U751 ( .A(n488), .B(n441), .S(u_alu_ashr_4_SH_3_), .Q(n414) );
  IMUX21 U752 ( .A(n267), .B(n268), .S(u_alu_ashr_4_SH_3_), .Q(n314) );
  IMUX21 U753 ( .A(n272), .B(n273), .S(u_alu_ashr_4_SH_3_), .Q(n320) );
  IMUX21 U754 ( .A(n283), .B(n284), .S(u_alu_ashr_4_SH_3_), .Q(n334) );
  IMUX21 U755 ( .A(n308), .B(n307), .S(u_alu_ashr_4_SH_3_), .Q(n359) );
  IMUX21 U756 ( .A(n293), .B(n294), .S(u_alu_ashr_4_SH_3_), .Q(n351) );
  IMUX20 U757 ( .A(n382), .B(n381), .S(n374), .Q(n407) );
  IMUX20 U758 ( .A(n460), .B(n425), .S(n374), .Q(n472) );
  IMUX20 U759 ( .A(n396), .B(n399), .S(n374), .Q(n411) );
  IMUX20 U760 ( .A(n265), .B(n253), .S(n374), .Q(n277) );
  IMUX20 U761 ( .A(n296), .B(n286), .S(n374), .Q(n311) );
  IMUX20 U762 ( .A(n270), .B(n259), .S(n374), .Q(n282) );
  IMUX21 U763 ( .A(n242), .B(n244), .S(n374), .Q(n251) );
  IMUX20 U764 ( .A(n303), .B(n291), .S(n374), .Q(n317) );
  MUX22 U765 ( .A(compare_i_data_rt[6]), .B(i_data_immext[6]), .S(n70), .Q(
        alu_i_data_B[6]) );
  BUF2 U766 ( .A(alu_i_con_AluCtrl[0]), .Q(n231) );
  NOR20 U767 ( .A(i_data_immext[3]), .B(i_data_immext[1]), .Q(n1165) );
  NOR21 U768 ( .A(i_con_Efamux[1]), .B(n525), .Q(n526) );
  IMUX20 U769 ( .A(n426), .B(n416), .S(i_data_immext[8]), .Q(n474) );
  IMUX20 U770 ( .A(n484), .B(n411), .S(i_data_immext[8]), .Q(n463) );
  AOI210 U771 ( .A(alu_i_data_B[6]), .B(n82), .C(n1103), .Q(n1100) );
  IMUX20 U772 ( .A(n479), .B(n407), .S(i_data_immext[8]), .Q(n452) );
  IMUX20 U773 ( .A(n472), .B(n426), .S(i_data_immext[8]), .Q(n493) );
  NOR40 U774 ( .A(n857), .B(n856), .C(n855), .D(n854), .Q(n1266) );
  IMUX20 U775 ( .A(n297), .B(n277), .S(i_data_immext[8]), .Q(n325) );
  IMUX20 U776 ( .A(n311), .B(n287), .S(i_data_immext[8]), .Q(n341) );
  IMUX20 U777 ( .A(n277), .B(n254), .S(i_data_immext[8]), .Q(n298) );
  IMUX20 U778 ( .A(alu_i_data_B[30]), .B(alu_i_data_B[31]), .S(n511), .Q(n389)
         );
  IMUX20 U779 ( .A(n287), .B(n266), .S(i_data_immext[8]), .Q(n312) );
  IMUX20 U780 ( .A(n292), .B(n271), .S(i_data_immext[8]), .Q(n318) );
  IMUX20 U781 ( .A(n304), .B(n282), .S(i_data_immext[8]), .Q(n332) );
  IMUX20 U782 ( .A(n282), .B(n260), .S(i_data_immext[8]), .Q(n305) );
  INV3 U783 ( .A(n964), .Q(n859) );
  NOR21 U784 ( .A(n795), .B(n794), .Q(n1076) );
  IMUX20 U785 ( .A(n317), .B(n292), .S(i_data_immext[8]), .Q(n349) );
  AOI221 U786 ( .A(n625), .B(i_data_FMalures[0]), .C(n513), .D(
        i_data_FEalures[0]), .Q(n628) );
  AOI221 U787 ( .A(n777), .B(i_data_FMalures[0]), .C(n111), .D(
        i_data_FEalures[0]), .Q(n780) );
  NAND22 U788 ( .A(n776), .B(i_data_rt[0]), .Q(n781) );
  NAND33 U789 ( .A(n775), .B(n774), .C(n773), .Q(compare_i_data_rt[1]) );
  AOI220 U790 ( .A(n626), .B(i_data_FMmemout[4]), .C(n625), .D(
        i_data_FMalures[4]), .Q(n610) );
  INV3 U791 ( .A(compare_i_data_rt[5]), .Q(n842) );
  AOI220 U792 ( .A(n778), .B(i_data_FMmemout[6]), .C(n777), .D(
        i_data_FMalures[6]), .Q(n753) );
  MUX22 U793 ( .A(compare_i_data_rt[7]), .B(u_alu_ashr_4_SH_1_), .S(n70), .Q(
        alu_i_data_B[7]) );
  NOR40 U794 ( .A(i_data_immext[2]), .B(n1209), .C(n1210), .D(n1206), .Q(n1172) );
  IMUX20 U795 ( .A(n450), .B(n449), .S(u_alu_ashr_4_SH_1_), .Q(n480) );
  IMUX20 U796 ( .A(n380), .B(n379), .S(u_alu_ashr_4_SH_1_), .Q(n479) );
  IMUX20 U797 ( .A(n397), .B(n396), .S(u_alu_ashr_4_SH_1_), .Q(n426) );
  IMUX20 U798 ( .A(n425), .B(n397), .S(u_alu_ashr_4_SH_1_), .Q(n484) );
  IMUX20 U799 ( .A(n461), .B(n460), .S(u_alu_ashr_4_SH_1_), .Q(n485) );
  NOR40 U800 ( .A(n1248), .B(n1247), .C(n1246), .D(n1245), .Q(n1267) );
  IMUX20 U801 ( .A(n447), .B(n450), .S(u_alu_ashr_4_SH_1_), .Q(n469) );
  IMUX20 U802 ( .A(n379), .B(n382), .S(u_alu_ashr_4_SH_1_), .Q(n393) );
  IMUX20 U803 ( .A(n449), .B(n380), .S(u_alu_ashr_4_SH_1_), .Q(n468) );
  IMUX20 U804 ( .A(n399), .B(n398), .S(u_alu_ashr_4_SH_1_), .Q(n416) );
  IMUX20 U805 ( .A(n398), .B(n401), .S(u_alu_ashr_4_SH_1_), .Q(n410) );
  IMUX20 U806 ( .A(n384), .B(n383), .S(u_alu_ashr_4_SH_1_), .Q(n406) );
  AOI221 U807 ( .A(n519), .B(u_alu_N217), .C(n966), .D(alu_i_data_B[24]), .Q(
        n973) );
  IMUX20 U808 ( .A(n286), .B(n276), .S(u_alu_ashr_4_SH_1_), .Q(n297) );
  IMUX20 U809 ( .A(n245), .B(n232), .S(u_alu_ashr_4_SH_1_), .Q(n254) );
  IMUX20 U810 ( .A(n383), .B(n386), .S(u_alu_ashr_4_SH_1_), .Q(n395) );
  IMUX20 U811 ( .A(n381), .B(n384), .S(u_alu_ashr_4_SH_1_), .Q(n392) );
  IMUX20 U812 ( .A(n253), .B(n245), .S(u_alu_ashr_4_SH_1_), .Q(n266) );
  IMUX20 U813 ( .A(n276), .B(n265), .S(u_alu_ashr_4_SH_1_), .Q(n287) );
  IMUX20 U814 ( .A(n249), .B(n239), .S(u_alu_ashr_4_SH_1_), .Q(n260) );
  IMUX20 U815 ( .A(n291), .B(n281), .S(u_alu_ashr_4_SH_1_), .Q(n304) );
  INV3 U816 ( .A(n1080), .Q(n520) );
  IMUX20 U817 ( .A(n259), .B(n249), .S(u_alu_ashr_4_SH_1_), .Q(n271) );
  IMUX20 U818 ( .A(n281), .B(n270), .S(u_alu_ashr_4_SH_1_), .Q(n292) );
  INV3 U819 ( .A(n510), .Q(n511) );
  NAND22 U820 ( .A(n1081), .B(n782), .Q(n1087) );
  AOI221 U821 ( .A(n625), .B(i_data_FMalures[1]), .C(n513), .D(
        i_data_FEalures[1]), .Q(n622) );
  AOI221 U822 ( .A(n777), .B(i_data_FMalures[1]), .C(n111), .D(
        i_data_FEalures[1]), .Q(n774) );
  AOI220 U823 ( .A(n626), .B(i_data_FMmemout[5]), .C(n625), .D(
        i_data_FMalures[5]), .Q(n607) );
  AOI220 U824 ( .A(n778), .B(i_data_FMmemout[7]), .C(n777), .D(
        i_data_FMalures[7]), .Q(n749) );
  OAI2111 U825 ( .A(n1182), .B(n1191), .C(n1202), .D(n1181), .Q(
        alu_i_con_AluCtrl[0]) );
  NOR21 U826 ( .A(i_con_Efamux[2]), .B(i_con_Efamux[0]), .Q(n525) );
  AOI210 U827 ( .A(u_alu_lt_x_11_B_2_), .B(n82), .C(n1125), .Q(n1122) );
  AOI210 U828 ( .A(n229), .B(n82), .C(n1118), .Q(n1115) );
  AOI210 U829 ( .A(alu_i_data_B[4]), .B(n82), .C(n1113), .Q(n1110) );
  AOI210 U830 ( .A(n71), .B(n82), .C(n1139), .Q(n1136) );
  AOI210 U831 ( .A(alu_i_data_B[5]), .B(n82), .C(n1108), .Q(n1105) );
  INV3 U832 ( .A(n1079), .Q(n1086) );
  NOR21 U833 ( .A(n793), .B(n1087), .Q(n1080) );
  NAND33 U834 ( .A(n623), .B(n622), .C(n621), .Q(compare_i_data_rs[1]) );
  AOI221 U835 ( .A(n626), .B(i_data_FMmemout[1]), .C(n515), .D(
        i_data_FWmemout[1]), .Q(n621) );
  NAND22 U836 ( .A(n776), .B(i_data_rt[1]), .Q(n775) );
  AOI221 U837 ( .A(n626), .B(i_data_FMmemout[2]), .C(n515), .D(
        i_data_FWmemout[2]), .Q(n618) );
  AOI221 U838 ( .A(n625), .B(i_data_FMalures[2]), .C(n513), .D(
        i_data_FEalures[2]), .Q(n619) );
  AOI221 U839 ( .A(n777), .B(i_data_FMalures[2]), .C(n111), .D(
        i_data_FEalures[2]), .Q(n771) );
  AOI221 U840 ( .A(n626), .B(i_data_FMmemout[3]), .C(n515), .D(
        i_data_FWmemout[3]), .Q(n615) );
  AOI220 U841 ( .A(n626), .B(i_data_FMmemout[6]), .C(n625), .D(
        i_data_FMalures[6]), .Q(n604) );
  AOI220 U842 ( .A(n626), .B(i_data_FMmemout[7]), .C(n625), .D(
        i_data_FMalures[7]), .Q(n601) );
  BUF2 U843 ( .A(i_data_immext[7]), .Q(u_alu_ashr_4_SH_1_) );
  NAND31 U844 ( .A(n1197), .B(n1202), .C(n1196), .Q(alu_i_con_AluCtrl[2]) );
  OAI2111 U845 ( .A(n1204), .B(n1203), .C(n1202), .D(n1201), .Q(
        alu_i_con_AluCtrl[3]) );
  NOR40 U846 ( .A(i_data_immext[0]), .B(i_data_immext[3]), .C(i_data_immext[1]), .D(n1166), .Q(n1173) );
  OAI212 U847 ( .A(n70), .B(n830), .C(n1208), .Q(alu_i_data_B[16]) );
  OAI210 U848 ( .A(n82), .B(n1147), .C(alu_i_data_B[11]), .Q(n1146) );
  OAI210 U849 ( .A(n82), .B(n1152), .C(alu_i_data_B[10]), .Q(n1151) );
  NOR22 U850 ( .A(alu_i_con_AluCtrl[3]), .B(n794), .Q(n1077) );
  NAND22 U851 ( .A(n624), .B(i_data_rs[1]), .Q(n623) );
  NAND22 U852 ( .A(n624), .B(i_data_rs[2]), .Q(n620) );
  AOI221 U853 ( .A(n778), .B(i_data_FMmemout[3]), .C(n518), .D(
        i_data_FWmemout[3]), .Q(n767) );
  NOR40 U854 ( .A(n1210), .B(n1207), .C(n1206), .D(i_data_immext[3]), .Q(n1200) );
  AOI210 U855 ( .A(n624), .B(i_data_rs[22]), .C(n557), .Q(n558) );
  NAND22 U856 ( .A(n524), .B(n523), .Q(n614) );
  INV3 U857 ( .A(n70), .Q(n711) );
  OAI210 U858 ( .A(n82), .B(n1124), .C(compare_i_data_rs[2]), .Q(n1123) );
  OAI210 U859 ( .A(n82), .B(n1117), .C(compare_i_data_rs[3]), .Q(n1116) );
  OAI210 U860 ( .A(n82), .B(n1138), .C(compare_i_data_rs[1]), .Q(n1137) );
  OAI210 U861 ( .A(n82), .B(n1085), .C(compare_i_data_rs[9]), .Q(n1084) );
  NAND22 U862 ( .A(n1068), .B(u_alu_pre_suba[1]), .Q(n876) );
  NAND22 U863 ( .A(n1068), .B(u_alu_pre_suba[7]), .Q(n952) );
  AOI211 U864 ( .A(n969), .B(compare_i_data_rs[24]), .C(n968), .Q(n972) );
  MUX22 U865 ( .A(u_alu_pre_sum_3a[8]), .B(u_alu_pre_sum_3b[8]), .S(u_alu_N173), .Q(n963) );
  AOI210 U866 ( .A(n624), .B(i_data_rs[20]), .C(n563), .Q(n564) );
  AOI210 U867 ( .A(n624), .B(i_data_rs[24]), .C(n551), .Q(n552) );
  AOI210 U868 ( .A(n776), .B(i_data_rt[26]), .C(n664), .Q(n665) );
  AOI210 U869 ( .A(n776), .B(i_data_rt[27]), .C(n659), .Q(n660) );
  AOI210 U870 ( .A(n776), .B(i_data_rt[28]), .C(n654), .Q(n655) );
  AOI210 U871 ( .A(n776), .B(i_data_rt[29]), .C(n649), .Q(n650) );
  NAND22 U872 ( .A(n70), .B(i_data_immext[16]), .Q(n1208) );
  AOI210 U873 ( .A(n776), .B(i_data_rt[31]), .C(n639), .Q(n640) );
  OAI210 U874 ( .A(n82), .B(n1107), .C(compare_i_data_rs[5]), .Q(n1106) );
  OAI210 U875 ( .A(n82), .B(n1102), .C(compare_i_data_rs[6]), .Q(n1101) );
  OAI210 U876 ( .A(n82), .B(n1097), .C(compare_i_data_rs[7]), .Q(n1096) );
  NAND22 U877 ( .A(n1069), .B(u_alu_pre_subb[3]), .Q(n902) );
  NAND22 U878 ( .A(n1068), .B(u_alu_pre_suba[3]), .Q(n903) );
  NAND22 U879 ( .A(n1069), .B(u_alu_pre_subb[7]), .Q(n951) );
  NAND22 U880 ( .A(n1069), .B(u_alu_pre_subb[2]), .Q(n890) );
  NAND22 U881 ( .A(n1068), .B(u_alu_pre_suba[2]), .Q(n891) );
  NAND22 U882 ( .A(n1069), .B(u_alu_pre_subb[4]), .Q(n914) );
  NAND22 U883 ( .A(n1068), .B(u_alu_pre_suba[4]), .Q(n915) );
  NAND22 U884 ( .A(n1069), .B(u_alu_pre_subb[6]), .Q(n939) );
  NAND22 U885 ( .A(n1068), .B(u_alu_pre_suba[6]), .Q(n940) );
  NAND22 U886 ( .A(n1069), .B(u_alu_pre_subb[5]), .Q(n927) );
  NAND22 U887 ( .A(n1068), .B(u_alu_pre_suba[5]), .Q(n928) );
  OAI2111 U888 ( .A(n868), .B(n1154), .C(n867), .D(n866), .Q(n869) );
  IMUX21 U889 ( .A(n387), .B(n389), .S(n374), .Q(n430) );
  NAND22 U890 ( .A(n1068), .B(u_alu_pre_suba[10]), .Q(n997) );
  NAND22 U891 ( .A(n1068), .B(u_alu_pre_suba[9]), .Q(n984) );
  INV3 U892 ( .A(n231), .Q(n793) );
  NAND22 U893 ( .A(n1244), .B(n1239), .Q(o_addr_Erd[0]) );
  NAND22 U894 ( .A(n1244), .B(n1241), .Q(o_addr_Erd[2]) );
  NAND22 U895 ( .A(n1244), .B(n1243), .Q(o_addr_Erd[4]) );
  NAND22 U896 ( .A(n1244), .B(n1242), .Q(o_addr_Erd[3]) );
  NAND22 U897 ( .A(n1244), .B(n1240), .Q(o_addr_Erd[1]) );
  IMUX20 U898 ( .A(n1086), .B(n1087), .S(u_alu_lt_x_11_B_2_), .Q(n1124) );
  NAND31 U899 ( .A(n816), .B(n815), .C(n814), .Q(n1125) );
  IMUX20 U900 ( .A(n453), .B(n452), .S(u_alu_ashr_4_SH_3_), .Q(n455) );
  NOR21 U901 ( .A(n372), .B(n362), .Q(u_alu_N195) );
  IMUX20 U902 ( .A(n1076), .B(n1079), .S(u_alu_lt_x_11_B_2_), .Q(n1121) );
  IMUX20 U903 ( .A(n1086), .B(n1087), .S(n229), .Q(n1117) );
  NAND31 U904 ( .A(n813), .B(n812), .C(n811), .Q(n1118) );
  IMUX20 U905 ( .A(n464), .B(n463), .S(u_alu_ashr_4_SH_3_), .Q(n466) );
  NOR21 U906 ( .A(n372), .B(n363), .Q(u_alu_N196) );
  IMUX20 U907 ( .A(n1076), .B(n1079), .S(n229), .Q(n1114) );
  IMUX20 U908 ( .A(n1086), .B(n1087), .S(alu_i_data_B[4]), .Q(n1112) );
  NAND22 U909 ( .A(n810), .B(n809), .Q(n1113) );
  NOR21 U910 ( .A(n372), .B(n364), .Q(u_alu_N197) );
  IMUX20 U911 ( .A(n1076), .B(n1079), .S(alu_i_data_B[4]), .Q(n1109) );
  MUX21 U912 ( .A(n393), .B(n392), .S(i_data_immext[8]), .Q(n467) );
  IMUX20 U913 ( .A(n1086), .B(n1087), .S(n71), .Q(n1138) );
  NAND31 U914 ( .A(n819), .B(n818), .C(n817), .Q(n1139) );
  IMUX20 U915 ( .A(n427), .B(n493), .S(u_alu_ashr_4_SH_3_), .Q(n429) );
  IMUX20 U916 ( .A(n229), .B(alu_i_data_B[4]), .S(n511), .Q(n459) );
  IMUX20 U917 ( .A(n71), .B(u_alu_lt_x_11_B_2_), .S(i_data_immext[6]), .Q(n423) );
  NOR21 U918 ( .A(n372), .B(n361), .Q(u_alu_N194) );
  IMUX20 U919 ( .A(n1076), .B(n1079), .S(n71), .Q(n1135) );
  OAI2111 U920 ( .A(compare_i_data_rs[5]), .B(n1104), .C(n1105), .D(n1106), 
        .Q(alu_o_data_AluRes[5]) );
  IMUX20 U921 ( .A(n1086), .B(n1087), .S(alu_i_data_B[5]), .Q(n1107) );
  NAND31 U922 ( .A(n808), .B(n807), .C(n806), .Q(n1108) );
  NOR21 U923 ( .A(n372), .B(n365), .Q(u_alu_N198) );
  IMUX20 U924 ( .A(n475), .B(n474), .S(u_alu_ashr_4_SH_3_), .Q(n477) );
  IMUX20 U925 ( .A(n458), .B(n461), .S(n374), .Q(n473) );
  IMUX20 U926 ( .A(alu_i_data_B[5]), .B(alu_i_data_B[6]), .S(n511), .Q(n458)
         );
  IMUX20 U927 ( .A(n1076), .B(n1079), .S(alu_i_data_B[5]), .Q(n1104) );
  OAI2111 U928 ( .A(alu_i_data_B[11]), .B(n1144), .C(n1145), .D(n1146), .Q(
        alu_o_data_AluRes[11]) );
  IMUX20 U929 ( .A(n1086), .B(n1087), .S(compare_i_data_rs[11]), .Q(n1147) );
  OAI2111 U930 ( .A(n861), .B(n822), .C(n821), .D(n820), .Q(n1148) );
  IMUX20 U931 ( .A(n463), .B(n422), .S(u_alu_ashr_4_SH_3_), .Q(n391) );
  INV3 U932 ( .A(u_alu_half_sub_11_), .Q(n822) );
  IMUX20 U933 ( .A(n1076), .B(n1079), .S(compare_i_data_rs[11]), .Q(n1144) );
  OAI2111 U934 ( .A(compare_i_data_rs[6]), .B(n1099), .C(n1100), .D(n1101), 
        .Q(alu_o_data_AluRes[6]) );
  IMUX20 U935 ( .A(n1086), .B(n1087), .S(alu_i_data_B[6]), .Q(n1102) );
  NAND31 U936 ( .A(n805), .B(n804), .C(n803), .Q(n1103) );
  NOR21 U937 ( .A(n372), .B(n366), .Q(u_alu_N199) );
  IMUX20 U938 ( .A(n1076), .B(n1079), .S(alu_i_data_B[6]), .Q(n1099) );
  OAI2111 U939 ( .A(alu_i_data_B[10]), .B(n1149), .C(n1150), .D(n1151), .Q(
        alu_o_data_AluRes[10]) );
  IMUX20 U940 ( .A(n1086), .B(n1087), .S(compare_i_data_rs[10]), .Q(n1152) );
  OAI2111 U941 ( .A(n861), .B(n825), .C(n824), .D(n823), .Q(n1153) );
  IMUX20 U942 ( .A(n452), .B(n420), .S(u_alu_ashr_4_SH_3_), .Q(n390) );
  INV3 U943 ( .A(u_alu_half_sub_10_), .Q(n825) );
  IMUX20 U944 ( .A(n1076), .B(n1079), .S(compare_i_data_rs[10]), .Q(n1149) );
  OAI2111 U945 ( .A(compare_i_data_rs[9]), .B(n1082), .C(n1083), .D(n1084), 
        .Q(alu_o_data_AluRes[9]) );
  IMUX20 U946 ( .A(n1086), .B(n1087), .S(alu_i_data_B[9]), .Q(n1085) );
  OAI2111 U947 ( .A(n861), .B(n792), .C(n791), .D(n790), .Q(n1088) );
  NOR21 U948 ( .A(n372), .B(n369), .Q(u_alu_N202) );
  IMUX20 U949 ( .A(n493), .B(n492), .S(u_alu_ashr_4_SH_3_), .Q(n495) );
  INV3 U950 ( .A(u_alu_half_sub_9_), .Q(n792) );
  IMUX20 U951 ( .A(n1076), .B(n1079), .S(alu_i_data_B[9]), .Q(n1082) );
  OAI2111 U952 ( .A(compare_i_data_rs[7]), .B(n1094), .C(n1095), .D(n1096), 
        .Q(alu_o_data_AluRes[7]) );
  IMUX20 U953 ( .A(n1086), .B(n1087), .S(alu_i_data_B[7]), .Q(n1097) );
  NAND31 U954 ( .A(n802), .B(n801), .C(n800), .Q(n1098) );
  NOR21 U955 ( .A(n372), .B(n367), .Q(u_alu_N200) );
  IMUX20 U956 ( .A(alu_i_data_B[13]), .B(alu_i_data_B[14]), .S(n511), .Q(n397)
         );
  IMUX20 U957 ( .A(alu_i_data_B[11]), .B(alu_i_data_B[12]), .S(n511), .Q(n425)
         );
  IMUX20 U958 ( .A(alu_i_data_B[9]), .B(alu_i_data_B[10]), .S(n511), .Q(n460)
         );
  IMUX20 U959 ( .A(alu_i_data_B[7]), .B(alu_i_data_B[8]), .S(n511), .Q(n461)
         );
  IMUX20 U960 ( .A(n1076), .B(n1079), .S(alu_i_data_B[7]), .Q(n1094) );
  AOI221 U961 ( .A(n1273), .B(i_con_bop[0]), .C(n1272), .D(
        compare_i_data_rs[31]), .Q(n1274) );
  NOR21 U962 ( .A(i_con_bop[2]), .B(n1271), .Q(n1272) );
  IMAJ31 U963 ( .A(i_con_bop[2]), .B(i_con_bop[1]), .C(n1270), .Q(n1275) );
  NAND41 U964 ( .A(n1260), .B(n1259), .C(n1258), .D(n1257), .Q(n1261) );
  NAND31 U965 ( .A(n851), .B(n850), .C(n849), .Q(n1262) );
  OAI2111 U966 ( .A(n520), .B(n1154), .C(n1155), .D(n1156), .Q(
        alu_o_data_AluRes[0]) );
  IMUX20 U967 ( .A(n1087), .B(n1086), .S(n1154), .Q(n1159) );
  INV3 U968 ( .A(u_alu_N306), .Q(n1161) );
  AOI221 U969 ( .A(n519), .B(u_alu_N193), .C(n1077), .D(u_alu_N225), .Q(n1155)
         );
  IMUX20 U970 ( .A(n376), .B(n469), .S(i_data_immext[8]), .Q(n377) );
  IMUX20 U971 ( .A(alu_i_data_B[6]), .B(alu_i_data_B[7]), .S(n511), .Q(n450)
         );
  IMUX20 U972 ( .A(alu_i_data_B[4]), .B(alu_i_data_B[5]), .S(n511), .Q(n447)
         );
  IMUX20 U973 ( .A(u_alu_lt_x_11_B_2_), .B(n229), .S(n511), .Q(n448) );
  IMUX20 U974 ( .A(alu_i_data_B[0]), .B(n71), .S(i_data_immext[6]), .Q(n375)
         );
  AOI211 U975 ( .A(compare_i_data_rs[8]), .B(n1091), .C(n1092), .Q(n1090) );
  NAND41 U976 ( .A(n799), .B(n798), .C(n797), .D(n796), .Q(n1092) );
  IMUX20 U977 ( .A(n489), .B(n488), .S(u_alu_ashr_4_SH_3_), .Q(n491) );
  IMUX20 U978 ( .A(alu_i_data_B[14]), .B(alu_i_data_B[15]), .S(n511), .Q(n382)
         );
  IMUX20 U979 ( .A(alu_i_data_B[12]), .B(alu_i_data_B[13]), .S(n511), .Q(n379)
         );
  IMUX20 U980 ( .A(alu_i_data_B[10]), .B(alu_i_data_B[11]), .S(n511), .Q(n380)
         );
  IMUX20 U981 ( .A(alu_i_data_B[8]), .B(alu_i_data_B[9]), .S(n511), .Q(n449)
         );
  OAI2111 U982 ( .A(n883), .B(n962), .C(n882), .D(n881), .Q(
        alu_o_data_AluRes[17]) );
  AOI211 U983 ( .A(n1069), .B(u_alu_pre_subb[1]), .C(n880), .Q(n881) );
  NAND41 U984 ( .A(n879), .B(n878), .C(n877), .D(n876), .Q(n880) );
  NOR21 U985 ( .A(n372), .B(n502), .Q(u_alu_N242) );
  NOR21 U986 ( .A(u_alu_ashr_4_SH_3_), .B(n307), .Q(n275) );
  IMUX20 U987 ( .A(n305), .B(n308), .S(u_alu_ashr_4_SH_3_), .Q(n264) );
  NAND22 U988 ( .A(n956), .B(u_alu_pre_sum_3b[1]), .Q(n882) );
  IMUX20 U989 ( .A(alu_i_data_B[17]), .B(alu_i_data_B[18]), .S(n511), .Q(n399)
         );
  IMUX20 U990 ( .A(alu_i_data_B[15]), .B(alu_i_data_B[16]), .S(n511), .Q(n396)
         );
  AOI211 U991 ( .A(n956), .B(u_alu_pre_sum_3b[3]), .C(n906), .Q(n907) );
  NAND41 U992 ( .A(n905), .B(n904), .C(n903), .D(n902), .Q(n906) );
  NOR21 U993 ( .A(u_alu_ashr_4_SH_3_), .B(n273), .Q(n353) );
  IMUX20 U994 ( .A(n318), .B(n272), .S(u_alu_ashr_4_SH_3_), .Q(n274) );
  IMUX20 U995 ( .A(alu_i_data_B[19]), .B(alu_i_data_B[20]), .S(n511), .Q(n398)
         );
  AOI211 U996 ( .A(n956), .B(u_alu_pre_sum_3b[7]), .C(n955), .Q(n957) );
  NAND41 U997 ( .A(n954), .B(n953), .C(n952), .D(n951), .Q(n955) );
  NOR21 U998 ( .A(u_alu_ashr_4_SH_3_), .B(n294), .Q(n357) );
  IMUX20 U999 ( .A(n349), .B(n293), .S(u_alu_ashr_4_SH_3_), .Q(n295) );
  NOR21 U1000 ( .A(n372), .B(n486), .Q(u_alu_N248) );
  AOI211 U1001 ( .A(n956), .B(u_alu_pre_sum_3b[2]), .C(n894), .Q(n895) );
  NAND41 U1002 ( .A(n893), .B(n892), .C(n891), .D(n890), .Q(n894) );
  NOR21 U1003 ( .A(n372), .B(n497), .Q(u_alu_N243) );
  AOI2111 U1004 ( .A(n519), .B(u_alu_N211), .C(n889), .D(n888), .Q(n893) );
  NOR21 U1005 ( .A(u_alu_ashr_4_SH_3_), .B(n268), .Q(n336) );
  IMUX20 U1006 ( .A(n312), .B(n267), .S(u_alu_ashr_4_SH_3_), .Q(n269) );
  AOI211 U1007 ( .A(n956), .B(u_alu_pre_sum_3b[4]), .C(n918), .Q(n919) );
  NAND41 U1008 ( .A(n917), .B(n916), .C(n915), .D(n914), .Q(n918) );
  NOR21 U1009 ( .A(u_alu_ashr_4_SH_3_), .B(n279), .Q(n354) );
  IMUX20 U1010 ( .A(n325), .B(n278), .S(u_alu_ashr_4_SH_3_), .Q(n280) );
  AOI211 U1011 ( .A(n956), .B(u_alu_pre_sum_3b[6]), .C(n943), .Q(n944) );
  NAND41 U1012 ( .A(n942), .B(n941), .C(n940), .D(n939), .Q(n943) );
  NOR21 U1013 ( .A(u_alu_ashr_4_SH_3_), .B(n289), .Q(n356) );
  IMUX20 U1014 ( .A(n341), .B(n288), .S(u_alu_ashr_4_SH_3_), .Q(n290) );
  NOR21 U1015 ( .A(n372), .B(n481), .Q(u_alu_N247) );
  AOI211 U1016 ( .A(n956), .B(u_alu_pre_sum_3b[5]), .C(n931), .Q(n932) );
  NAND41 U1017 ( .A(n930), .B(n929), .C(n928), .D(n927), .Q(n931) );
  NOR21 U1018 ( .A(u_alu_ashr_4_SH_3_), .B(n284), .Q(n355) );
  IMUX20 U1019 ( .A(n332), .B(n283), .S(u_alu_ashr_4_SH_3_), .Q(n285) );
  NOR21 U1020 ( .A(n372), .B(n503), .Q(u_alu_N246) );
  IMUX20 U1021 ( .A(alu_i_data_B[23]), .B(alu_i_data_B[24]), .S(n511), .Q(n400) );
  IMUX20 U1022 ( .A(alu_i_data_B[21]), .B(alu_i_data_B[22]), .S(n511), .Q(n401) );
  OAI2111 U1023 ( .A(n977), .B(u_alu_pre_sum_4a[0]), .C(n976), .D(n975), .Q(
        alu_o_data_AluRes[24]) );
  AOI211 U1024 ( .A(n1068), .B(u_alu_pre_suba[8]), .C(n974), .Q(n975) );
  NOR21 U1025 ( .A(n372), .B(n499), .Q(u_alu_N249) );
  NOR21 U1026 ( .A(u_alu_ashr_4_SH_3_), .B(n441), .Q(n490) );
  IMUX20 U1027 ( .A(n299), .B(n298), .S(u_alu_ashr_4_SH_3_), .Q(n302) );
  NAND22 U1028 ( .A(n1071), .B(u_alu_pre_sum_4a[0]), .Q(n976) );
  NAND22 U1029 ( .A(n1071), .B(u_alu_pre_sum_4a[4]), .Q(n1025) );
  NAND22 U1030 ( .A(n1070), .B(u_alu_pre_sum_4b[4]), .Q(n1026) );
  NAND22 U1031 ( .A(n1069), .B(u_alu_pre_subb[12]), .Q(n1027) );
  AOI211 U1032 ( .A(n1068), .B(u_alu_pre_suba[12]), .C(n1024), .Q(n1028) );
  NAND41 U1033 ( .A(n1023), .B(n1022), .C(n1021), .D(n1020), .Q(n1024) );
  NAND31 U1034 ( .A(n508), .B(n509), .C(n430), .Q(n445) );
  IMUX20 U1035 ( .A(n326), .B(n325), .S(u_alu_ashr_4_SH_3_), .Q(n328) );
  IMUX20 U1036 ( .A(n310), .B(n296), .S(n374), .Q(n323) );
  IMUX20 U1037 ( .A(n337), .B(n322), .S(n374), .Q(n324) );
  NAND22 U1038 ( .A(n1071), .B(u_alu_pre_sum_4a[6]), .Q(n1052) );
  NAND22 U1039 ( .A(n1070), .B(u_alu_pre_sum_4b[6]), .Q(n1053) );
  AOI211 U1040 ( .A(n1068), .B(u_alu_pre_suba[14]), .C(n1051), .Q(n1055) );
  NAND41 U1041 ( .A(n1050), .B(n1049), .C(n1048), .D(n1047), .Q(n1051) );
  NAND31 U1042 ( .A(n435), .B(n508), .C(n509), .Q(n456) );
  IMUX20 U1043 ( .A(n342), .B(n341), .S(u_alu_ashr_4_SH_3_), .Q(n344) );
  IMUX20 U1044 ( .A(n338), .B(n337), .S(n374), .Q(n340) );
  IMUX20 U1045 ( .A(alu_i_data_B[30]), .B(alu_i_data_B[29]), .S(
        i_data_immext[6]), .Q(n338) );
  OAI2111 U1046 ( .A(u_alu_pre_subb[0]), .B(n230), .C(n871), .D(n870), .Q(n872) );
  AOI211 U1047 ( .A(n1077), .B(u_alu_N241), .C(n869), .Q(n870) );
  IMUX20 U1048 ( .A(n298), .B(n301), .S(u_alu_ashr_4_SH_3_), .Q(n258) );
  NOR21 U1049 ( .A(n372), .B(n500), .Q(u_alu_N241) );
  IMUX20 U1050 ( .A(alu_i_data_B[24]), .B(alu_i_data_B[25]), .S(n511), .Q(n385) );
  IMUX20 U1051 ( .A(alu_i_data_B[22]), .B(alu_i_data_B[23]), .S(n511), .Q(n386) );
  IMUX20 U1052 ( .A(alu_i_data_B[20]), .B(alu_i_data_B[21]), .S(n511), .Q(n383) );
  IMUX20 U1053 ( .A(alu_i_data_B[18]), .B(alu_i_data_B[19]), .S(n511), .Q(n384) );
  IMUX20 U1054 ( .A(alu_i_data_B[16]), .B(alu_i_data_B[17]), .S(n511), .Q(n381) );
  NAND22 U1055 ( .A(n1002), .B(n1001), .Q(alu_o_data_AluRes[26]) );
  NAND22 U1056 ( .A(n1071), .B(u_alu_pre_sum_4a[2]), .Q(n1001) );
  AOI211 U1057 ( .A(n1070), .B(u_alu_pre_sum_4b[2]), .C(n1000), .Q(n1002) );
  NAND41 U1058 ( .A(n999), .B(n998), .C(n997), .D(n996), .Q(n1000) );
  NAND22 U1059 ( .A(n1069), .B(u_alu_pre_subb[10]), .Q(n996) );
  NOR21 U1060 ( .A(u_alu_ashr_4_SH_3_), .B(n419), .Q(n443) );
  NOR21 U1061 ( .A(u_alu_ashr_4_SH_1_), .B(n389), .Q(n435) );
  IMUX20 U1062 ( .A(alu_i_data_B[28]), .B(alu_i_data_B[29]), .S(n511), .Q(n387) );
  IMUX20 U1063 ( .A(alu_i_data_B[26]), .B(alu_i_data_B[27]), .S(n511), .Q(n388) );
  AOI2111 U1064 ( .A(n519), .B(u_alu_N219), .C(n995), .D(n994), .Q(n999) );
  NAND22 U1065 ( .A(n509), .B(n247), .Q(n268) );
  IMUX20 U1066 ( .A(u_alu_lt_x_11_B_2_), .B(n71), .S(n511), .Q(n235) );
  IMUX20 U1067 ( .A(alu_i_data_B[4]), .B(n229), .S(n511), .Q(n236) );
  IMUX20 U1068 ( .A(alu_i_data_B[6]), .B(alu_i_data_B[5]), .S(n511), .Q(n233)
         );
  IMUX20 U1069 ( .A(alu_i_data_B[8]), .B(alu_i_data_B[7]), .S(n511), .Q(n234)
         );
  IMUX20 U1070 ( .A(alu_i_data_B[10]), .B(alu_i_data_B[9]), .S(n511), .Q(n232)
         );
  IMUX20 U1071 ( .A(n313), .B(n312), .S(u_alu_ashr_4_SH_3_), .Q(n315) );
  IMUX20 U1072 ( .A(alu_i_data_B[12]), .B(alu_i_data_B[11]), .S(n511), .Q(n245) );
  IMUX20 U1073 ( .A(alu_i_data_B[14]), .B(alu_i_data_B[13]), .S(n511), .Q(n253) );
  IMUX20 U1074 ( .A(alu_i_data_B[16]), .B(alu_i_data_B[15]), .S(n511), .Q(n265) );
  IMUX20 U1075 ( .A(alu_i_data_B[18]), .B(alu_i_data_B[17]), .S(n511), .Q(n276) );
  IMUX20 U1076 ( .A(alu_i_data_B[22]), .B(alu_i_data_B[21]), .S(n511), .Q(n296) );
  IMUX20 U1077 ( .A(n322), .B(n310), .S(n374), .Q(n339) );
  NAND22 U1078 ( .A(n1015), .B(n1014), .Q(alu_o_data_AluRes[27]) );
  NAND22 U1079 ( .A(n1071), .B(u_alu_pre_sum_4a[3]), .Q(n1014) );
  AOI211 U1080 ( .A(n1070), .B(u_alu_pre_sum_4b[3]), .C(n1013), .Q(n1015) );
  NAND41 U1081 ( .A(n1012), .B(n1011), .C(n1010), .D(n1009), .Q(n1013) );
  NAND22 U1082 ( .A(n1069), .B(u_alu_pre_subb[11]), .Q(n1009) );
  NAND22 U1083 ( .A(n509), .B(n251), .Q(n273) );
  IMUX20 U1084 ( .A(n319), .B(n318), .S(u_alu_ashr_4_SH_3_), .Q(n321) );
  NOR21 U1085 ( .A(n372), .B(n507), .Q(u_alu_N252) );
  NOR21 U1086 ( .A(u_alu_ashr_4_SH_3_), .B(n421), .Q(n444) );
  NAND22 U1087 ( .A(n1041), .B(n1040), .Q(alu_o_data_AluRes[29]) );
  NAND22 U1088 ( .A(n1071), .B(u_alu_pre_sum_4a[5]), .Q(n1040) );
  AOI211 U1089 ( .A(n1070), .B(u_alu_pre_sum_4b[5]), .C(n1039), .Q(n1041) );
  NAND41 U1090 ( .A(n1038), .B(n1037), .C(n1036), .D(n1035), .Q(n1039) );
  NAND22 U1091 ( .A(n1069), .B(u_alu_pre_subb[13]), .Q(n1035) );
  IMUX20 U1092 ( .A(n333), .B(n332), .S(u_alu_ashr_4_SH_3_), .Q(n335) );
  IMUX20 U1093 ( .A(n345), .B(n329), .S(n374), .Q(n331) );
  NOR21 U1094 ( .A(n372), .B(n504), .Q(u_alu_N254) );
  NOR21 U1095 ( .A(u_alu_ashr_4_SH_3_), .B(n433), .Q(n446) );
  NAND22 U1096 ( .A(n509), .B(n417), .Q(n433) );
  NAND22 U1097 ( .A(n989), .B(n988), .Q(alu_o_data_AluRes[25]) );
  NAND22 U1098 ( .A(n1071), .B(u_alu_pre_sum_4a[1]), .Q(n988) );
  AOI211 U1099 ( .A(n1070), .B(u_alu_pre_sum_4b[1]), .C(n987), .Q(n989) );
  NAND41 U1100 ( .A(n986), .B(n985), .C(n984), .D(n983), .Q(n987) );
  NAND22 U1101 ( .A(n1069), .B(u_alu_pre_subb[9]), .Q(n983) );
  NAND22 U1102 ( .A(n263), .B(n509), .Q(n307) );
  NOR21 U1103 ( .A(u_alu_ashr_4_SH_1_), .B(n244), .Q(n263) );
  IMUX20 U1104 ( .A(n306), .B(n305), .S(u_alu_ashr_4_SH_3_), .Q(n309) );
  IMUX20 U1105 ( .A(n316), .B(n303), .S(n374), .Q(n330) );
  NOR21 U1106 ( .A(n372), .B(n501), .Q(u_alu_N250) );
  NOR21 U1107 ( .A(u_alu_ashr_4_SH_3_), .B(n442), .Q(n494) );
  IMUX20 U1108 ( .A(alu_i_data_B[29]), .B(alu_i_data_B[30]), .S(n511), .Q(n405) );
  IMUX20 U1109 ( .A(alu_i_data_B[27]), .B(alu_i_data_B[28]), .S(n511), .Q(n402) );
  IMUX20 U1110 ( .A(alu_i_data_B[25]), .B(alu_i_data_B[26]), .S(n511), .Q(n403) );
  NAND41 U1111 ( .A(n1075), .B(n1074), .C(n1073), .D(n1072), .Q(
        alu_o_data_AluRes[31]) );
  NAND22 U1112 ( .A(n1071), .B(u_alu_pre_sum_4a[7]), .Q(n1072) );
  OAI222 U1113 ( .A(n962), .B(n961), .C(n960), .D(n959), .Q(n1070) );
  AOI211 U1114 ( .A(u_alu_pre_suba[15]), .B(n1068), .C(n1067), .Q(n1075) );
  NAND41 U1115 ( .A(n1066), .B(n1065), .C(n1064), .D(n1063), .Q(n1067) );
  INV3 U1116 ( .A(n1076), .Q(n1060) );
  NOR31 U1117 ( .A(alu_i_con_AluCtrl[2]), .B(n793), .C(n789), .Q(n1078) );
  IMUX20 U1118 ( .A(n71), .B(alu_i_data_B[0]), .S(n511), .Q(n244) );
  IMUX20 U1119 ( .A(n229), .B(u_alu_lt_x_11_B_2_), .S(n511), .Q(n242) );
  IMUX20 U1120 ( .A(alu_i_data_B[5]), .B(alu_i_data_B[4]), .S(n511), .Q(n243)
         );
  IMUX20 U1121 ( .A(alu_i_data_B[7]), .B(alu_i_data_B[6]), .S(n511), .Q(n240)
         );
  IMUX20 U1122 ( .A(alu_i_data_B[9]), .B(alu_i_data_B[8]), .S(n511), .Q(n241)
         );
  IMUX20 U1123 ( .A(alu_i_data_B[11]), .B(alu_i_data_B[10]), .S(n511), .Q(n239) );
  IMUX20 U1124 ( .A(alu_i_data_B[13]), .B(alu_i_data_B[12]), .S(n511), .Q(n249) );
  IMUX20 U1125 ( .A(alu_i_data_B[15]), .B(alu_i_data_B[14]), .S(n511), .Q(n259) );
  IMUX20 U1126 ( .A(n350), .B(n349), .S(u_alu_ashr_4_SH_3_), .Q(n352) );
  IMUX20 U1127 ( .A(alu_i_data_B[17]), .B(alu_i_data_B[16]), .S(n511), .Q(n270) );
  IMUX20 U1128 ( .A(alu_i_data_B[23]), .B(alu_i_data_B[22]), .S(n511), .Q(n303) );
  IMUX20 U1129 ( .A(n329), .B(n316), .S(n374), .Q(n347) );
  IMUX20 U1130 ( .A(n346), .B(n345), .S(n374), .Q(n348) );
  INV3 U1131 ( .A(n373), .Q(n374) );
  IMUX20 U1132 ( .A(alu_i_data_B[31]), .B(alu_i_data_B[30]), .S(
        i_data_immext[6]), .Q(n346) );
  NOR21 U1133 ( .A(alu_i_con_AluCtrl[2]), .B(alu_i_con_AluCtrl[3]), .Q(n782)
         );
  NAND31 U1134 ( .A(n438), .B(n508), .C(n509), .Q(n457) );
  NOR21 U1135 ( .A(u_alu_ashr_4_SH_1_), .B(n404), .Q(n438) );
  INV3 U1136 ( .A(i_data_immext[6]), .Q(n510) );
  NAND22 U1137 ( .A(n624), .B(i_data_rs[3]), .Q(n617) );
  OAI212 U1138 ( .A(n514), .B(n1233), .C(n613), .Q(compare_i_data_rs[4]) );
  OAI212 U1139 ( .A(n517), .B(n1233), .C(n765), .Q(compare_i_data_rt[4]) );
  AOI211 U1140 ( .A(n776), .B(i_data_rt[4]), .C(n764), .Q(n765) );
  OAI212 U1141 ( .A(n514), .B(n1234), .C(n609), .Q(compare_i_data_rs[5]) );
  AOI211 U1142 ( .A(n624), .B(i_data_rs[5]), .C(n608), .Q(n609) );
  OAI212 U1143 ( .A(n517), .B(n1234), .C(n760), .Q(compare_i_data_rt[5]) );
  AOI211 U1144 ( .A(n776), .B(i_data_rt[5]), .C(n759), .Q(n760) );
  OAI212 U1145 ( .A(n514), .B(n1235), .C(n606), .Q(compare_i_data_rs[6]) );
  OAI212 U1146 ( .A(n517), .B(n1235), .C(n756), .Q(compare_i_data_rt[6]) );
  AOI211 U1147 ( .A(n776), .B(i_data_rt[6]), .C(n755), .Q(n756) );
  OAI212 U1148 ( .A(n514), .B(n1236), .C(n603), .Q(compare_i_data_rs[7]) );
  AOI211 U1149 ( .A(n624), .B(i_data_rs[7]), .C(n602), .Q(n603) );
  OAI212 U1150 ( .A(n517), .B(n1236), .C(n752), .Q(compare_i_data_rt[7]) );
  AOI211 U1151 ( .A(n776), .B(i_data_rt[7]), .C(n751), .Q(n752) );
  OAI212 U1152 ( .A(n514), .B(n1237), .C(n600), .Q(compare_i_data_rs[8]) );
  MUX22 U1153 ( .A(compare_i_data_rt[8]), .B(i_data_immext[8]), .S(n70), .Q(
        alu_i_data_B[8]) );
  OAI212 U1154 ( .A(n514), .B(n1238), .C(n597), .Q(compare_i_data_rs[9]) );
  AOI211 U1155 ( .A(n624), .B(i_data_rs[9]), .C(n596), .Q(n597) );
  MUX22 U1156 ( .A(compare_i_data_rt[9]), .B(u_alu_ashr_4_SH_3_), .S(n70), .Q(
        alu_i_data_B[9]) );
  OAI212 U1157 ( .A(n517), .B(n1238), .C(n744), .Q(compare_i_data_rt[9]) );
  OAI212 U1158 ( .A(n514), .B(n1211), .C(n594), .Q(compare_i_data_rs[10]) );
  MUX22 U1159 ( .A(compare_i_data_rt[10]), .B(i_data_immext[10]), .S(n70), .Q(
        alu_i_data_B[10]) );
  OAI212 U1160 ( .A(n517), .B(n1211), .C(n740), .Q(compare_i_data_rt[10]) );
  OAI212 U1161 ( .A(n514), .B(n1212), .C(n591), .Q(compare_i_data_rs[11]) );
  AOI211 U1162 ( .A(n624), .B(i_data_rs[11]), .C(n590), .Q(n591) );
  MUX22 U1163 ( .A(compare_i_data_rt[11]), .B(i_data_immext[11]), .S(n70), .Q(
        alu_i_data_B[11]) );
  OAI212 U1164 ( .A(n517), .B(n1212), .C(n736), .Q(compare_i_data_rt[11]) );
  OAI212 U1165 ( .A(n514), .B(n1213), .C(n588), .Q(compare_i_data_rs[12]) );
  OAI212 U1166 ( .A(n517), .B(n1213), .C(n732), .Q(compare_i_data_rt[12]) );
  OAI212 U1167 ( .A(n514), .B(n1214), .C(n585), .Q(compare_i_data_rs[13]) );
  OAI212 U1168 ( .A(n517), .B(n1214), .C(n728), .Q(compare_i_data_rt[13]) );
  OAI212 U1169 ( .A(n514), .B(n1215), .C(n582), .Q(compare_i_data_rs[14]) );
  OAI212 U1170 ( .A(n514), .B(n1216), .C(n579), .Q(compare_i_data_rs[15]) );
  NOR21 U1171 ( .A(n785), .B(n231), .Q(n786) );
  OAI2111 U1172 ( .A(i_data_immext[0]), .B(n1171), .C(n1184), .D(n1170), .Q(
        n1199) );
  NOR21 U1173 ( .A(i_data_immext[4]), .B(n1169), .Q(n1184) );
  NAND22 U1174 ( .A(n1193), .B(n1174), .Q(n1183) );
  OAI212 U1175 ( .A(n614), .B(n1232), .C(n531), .Q(compare_i_data_rs[31]) );
  AOI211 U1176 ( .A(n624), .B(i_data_rs[31]), .C(n530), .Q(n531) );
  OAI212 U1177 ( .A(n514), .B(n1217), .C(n576), .Q(compare_i_data_rs[16]) );
  INV3 U1178 ( .A(compare_i_data_rt[16]), .Q(n830) );
  OAI212 U1179 ( .A(n517), .B(n1217), .C(n716), .Q(compare_i_data_rt[16]) );
  AOI211 U1180 ( .A(n776), .B(i_data_rt[16]), .C(n715), .Q(n716) );
  OAI212 U1181 ( .A(n514), .B(n1218), .C(n573), .Q(compare_i_data_rs[17]) );
  AOI211 U1182 ( .A(n624), .B(i_data_rs[17]), .C(n572), .Q(n573) );
  NAND22 U1183 ( .A(n712), .B(n1208), .Q(alu_i_data_B[17]) );
  OAI212 U1184 ( .A(n517), .B(n1218), .C(n710), .Q(compare_i_data_rt[17]) );
  AOI211 U1185 ( .A(n776), .B(i_data_rt[17]), .C(n709), .Q(n710) );
  OAI212 U1186 ( .A(n514), .B(n1219), .C(n570), .Q(compare_i_data_rs[18]) );
  AOI211 U1187 ( .A(n624), .B(i_data_rs[18]), .C(n569), .Q(n570) );
  NAND22 U1188 ( .A(n706), .B(n1208), .Q(alu_i_data_B[18]) );
  OAI212 U1189 ( .A(n517), .B(n1219), .C(n705), .Q(compare_i_data_rt[18]) );
  AOI211 U1190 ( .A(n776), .B(i_data_rt[18]), .C(n704), .Q(n705) );
  OAI212 U1191 ( .A(n514), .B(n1220), .C(n567), .Q(compare_i_data_rs[19]) );
  NAND22 U1192 ( .A(n701), .B(n1208), .Q(alu_i_data_B[19]) );
  OAI212 U1193 ( .A(n517), .B(n1220), .C(n700), .Q(compare_i_data_rt[19]) );
  AOI211 U1194 ( .A(n776), .B(i_data_rt[19]), .C(n699), .Q(n700) );
  OAI212 U1195 ( .A(n514), .B(n1221), .C(n564), .Q(compare_i_data_rs[20]) );
  NAND22 U1196 ( .A(n696), .B(n1208), .Q(alu_i_data_B[20]) );
  OAI212 U1197 ( .A(n517), .B(n1221), .C(n695), .Q(compare_i_data_rt[20]) );
  OAI212 U1198 ( .A(n514), .B(n1222), .C(n561), .Q(compare_i_data_rs[21]) );
  NAND22 U1199 ( .A(n691), .B(n1208), .Q(alu_i_data_B[21]) );
  NAND22 U1200 ( .A(compare_i_data_rt[21]), .B(n711), .Q(n691) );
  OAI212 U1201 ( .A(n517), .B(n1222), .C(n690), .Q(compare_i_data_rt[21]) );
  OAI212 U1202 ( .A(n514), .B(n1223), .C(n558), .Q(compare_i_data_rs[22]) );
  NAND22 U1203 ( .A(n686), .B(n1208), .Q(alu_i_data_B[22]) );
  NAND22 U1204 ( .A(compare_i_data_rt[22]), .B(n711), .Q(n686) );
  OAI212 U1205 ( .A(n517), .B(n1223), .C(n685), .Q(compare_i_data_rt[22]) );
  OAI212 U1206 ( .A(n514), .B(n1224), .C(n555), .Q(compare_i_data_rs[23]) );
  NAND22 U1207 ( .A(n681), .B(n1208), .Q(alu_i_data_B[23]) );
  NAND22 U1208 ( .A(compare_i_data_rt[23]), .B(n711), .Q(n681) );
  OAI212 U1209 ( .A(n517), .B(n1224), .C(n680), .Q(compare_i_data_rt[23]) );
  OAI212 U1210 ( .A(n514), .B(n1225), .C(n552), .Q(compare_i_data_rs[24]) );
  NAND22 U1211 ( .A(n676), .B(n1208), .Q(alu_i_data_B[24]) );
  OAI212 U1212 ( .A(n514), .B(n1226), .C(n549), .Q(compare_i_data_rs[25]) );
  NAND22 U1213 ( .A(n671), .B(n1208), .Q(alu_i_data_B[25]) );
  OAI212 U1214 ( .A(n514), .B(n1227), .C(n546), .Q(compare_i_data_rs[26]) );
  NAND22 U1215 ( .A(n666), .B(n1208), .Q(alu_i_data_B[26]) );
  OAI212 U1216 ( .A(n514), .B(n1228), .C(n543), .Q(compare_i_data_rs[27]) );
  NAND22 U1217 ( .A(n661), .B(n1208), .Q(alu_i_data_B[27]) );
  OAI212 U1218 ( .A(n514), .B(n1229), .C(n540), .Q(compare_i_data_rs[28]) );
  NAND22 U1219 ( .A(n656), .B(n1208), .Q(alu_i_data_B[28]) );
  OAI212 U1220 ( .A(n514), .B(n1230), .C(n537), .Q(compare_i_data_rs[29]) );
  NAND22 U1221 ( .A(n651), .B(n1208), .Q(alu_i_data_B[29]) );
  OAI212 U1222 ( .A(n514), .B(n1231), .C(n534), .Q(compare_i_data_rs[30]) );
  NAND22 U1223 ( .A(n646), .B(n1208), .Q(alu_i_data_B[30]) );
  NAND22 U1224 ( .A(n641), .B(n1208), .Q(alu_i_data_B[31]) );
  NAND22 U1225 ( .A(i_con_Efbmux[2]), .B(i_con_Efbmux[0]), .Q(n630) );
  IMUX20 U1226 ( .A(n448), .B(n447), .S(n374), .Q(n451) );
  IMUX20 U1227 ( .A(n459), .B(n458), .S(n374), .Q(n462) );
  IMUX20 U1228 ( .A(n423), .B(n459), .S(u_alu_ashr_4_SH_1_), .Q(n424) );
  IMUX20 U1229 ( .A(n375), .B(n448), .S(u_alu_ashr_4_SH_1_), .Q(n376) );
  MUX21 U1230 ( .A(n264), .B(n275), .S(n372), .Q(u_alu_N210) );
  MUX21 U1231 ( .A(n328), .B(n327), .S(n372), .Q(u_alu_N221) );
  MUX21 U1232 ( .A(n344), .B(n343), .S(n372), .Q(u_alu_N223) );
  IMUX20 U1233 ( .A(alu_i_data_B[28]), .B(alu_i_data_B[27]), .S(
        i_data_immext[6]), .Q(n337) );
  MUX21 U1234 ( .A(n258), .B(n257), .S(n372), .Q(u_alu_N209) );
  IMUX20 U1235 ( .A(alu_i_data_B[20]), .B(alu_i_data_B[19]), .S(
        i_data_immext[6]), .Q(n286) );
  IMUX20 U1236 ( .A(alu_i_data_B[24]), .B(alu_i_data_B[23]), .S(
        i_data_immext[6]), .Q(n310) );
  IMUX20 U1237 ( .A(alu_i_data_B[26]), .B(alu_i_data_B[25]), .S(
        i_data_immext[6]), .Q(n322) );
  IMUX20 U1238 ( .A(n243), .B(n242), .S(u_alu_ashr_4_SH_1_), .Q(n261) );
  NAND22 U1239 ( .A(u_alu_N173), .B(n859), .Q(n959) );
  NAND22 U1240 ( .A(n788), .B(n787), .Q(n964) );
  NOR21 U1241 ( .A(alu_i_con_AluCtrl[2]), .B(n231), .Q(n787) );
  MUX21 U1242 ( .A(n352), .B(n351), .S(n372), .Q(u_alu_N224) );
  IMUX20 U1243 ( .A(n240), .B(n243), .S(u_alu_ashr_4_SH_1_), .Q(n252) );
  IMUX20 U1244 ( .A(alu_i_data_B[19]), .B(alu_i_data_B[18]), .S(
        i_data_immext[6]), .Q(n281) );
  IMUX20 U1245 ( .A(alu_i_data_B[21]), .B(alu_i_data_B[20]), .S(
        i_data_immext[6]), .Q(n291) );
  IMUX20 U1246 ( .A(alu_i_data_B[25]), .B(alu_i_data_B[24]), .S(
        i_data_immext[6]), .Q(n316) );
  IMUX20 U1247 ( .A(alu_i_data_B[27]), .B(alu_i_data_B[26]), .S(
        i_data_immext[6]), .Q(n329) );
  IMUX20 U1248 ( .A(alu_i_data_B[29]), .B(alu_i_data_B[28]), .S(
        i_data_immext[6]), .Q(n345) );
  NAND22 U1249 ( .A(n1081), .B(alu_i_con_AluCtrl[2]), .Q(n794) );
  NAND22 U1250 ( .A(n788), .B(n786), .Q(n861) );
  NAND22 U1251 ( .A(alu_i_con_AluCtrl[1]), .B(n784), .Q(n789) );
  INV3 U1252 ( .A(n1198), .Q(n1191) );
  NAND22 U1253 ( .A(n525), .B(i_con_Efamux[1]), .Q(n611) );
  NAND22 U1254 ( .A(i_con_Efamux[2]), .B(i_con_Efamux[0]), .Q(n522) );
  XNR21 U1255 ( .A(compare_i_data_rt[27]), .B(n1006), .Q(n1253) );
  XNR21 U1256 ( .A(compare_i_data_rt[26]), .B(n993), .Q(n1254) );
  XNR21 U1257 ( .A(compare_i_data_rt[25]), .B(n102), .Q(n1255) );
  XNR21 U1258 ( .A(compare_i_data_rt[24]), .B(n110), .Q(n1256) );
  NOR40 U1259 ( .A(n840), .B(n839), .C(n838), .D(n837), .Q(n1258) );
  XNR21 U1260 ( .A(compare_i_data_rt[30]), .B(n1042), .Q(n837) );
  XNR21 U1261 ( .A(compare_i_data_rt[28]), .B(n101), .Q(n838) );
  XNR21 U1262 ( .A(compare_i_data_rt[29]), .B(n1032), .Q(n839) );
  XNR21 U1263 ( .A(compare_i_data_rs[2]), .B(n836), .Q(n840) );
  NOR40 U1264 ( .A(n835), .B(n834), .C(n833), .D(n832), .Q(n1259) );
  XNR21 U1265 ( .A(compare_i_data_rt[19]), .B(n103), .Q(n832) );
  XNR21 U1266 ( .A(compare_i_data_rt[17]), .B(n98), .Q(n833) );
  XNR21 U1267 ( .A(compare_i_data_rt[18]), .B(n887), .Q(n834) );
  XNR21 U1268 ( .A(compare_i_data_rs[1]), .B(n831), .Q(n835) );
  XNR21 U1269 ( .A(compare_i_data_rt[23]), .B(n96), .Q(n1249) );
  XNR21 U1270 ( .A(compare_i_data_rt[22]), .B(n109), .Q(n1250) );
  XNR21 U1271 ( .A(compare_i_data_rt[21]), .B(n924), .Q(n1251) );
  XNR21 U1272 ( .A(compare_i_data_rt[20]), .B(n104), .Q(n1252) );
  XNR21 U1273 ( .A(compare_i_data_rt[31]), .B(compare_i_data_rs[31]), .Q(n849)
         );
  XNR21 U1274 ( .A(compare_i_data_rt[9]), .B(compare_i_data_rs[9]), .Q(n850)
         );
  NOR40 U1275 ( .A(n848), .B(n847), .C(n846), .D(n845), .Q(n851) );
  XNR21 U1276 ( .A(compare_i_data_rt[7]), .B(n844), .Q(n845) );
  XNR21 U1277 ( .A(compare_i_data_rt[8]), .B(n107), .Q(n846) );
  XNR21 U1278 ( .A(compare_i_data_rt[6]), .B(n105), .Q(n847) );
  XNR21 U1279 ( .A(compare_i_data_rs[3]), .B(n843), .Q(n848) );
  XNR21 U1280 ( .A(compare_i_data_rs[5]), .B(n842), .Q(n1263) );
  XNR21 U1281 ( .A(compare_i_data_rt[4]), .B(n841), .Q(n1264) );
  XNR21 U1282 ( .A(compare_i_data_rt[11]), .B(n97), .Q(n854) );
  XNR21 U1283 ( .A(compare_i_data_rt[12]), .B(n853), .Q(n855) );
  XNR21 U1284 ( .A(compare_i_data_rt[10]), .B(n108), .Q(n856) );
  XNR21 U1285 ( .A(compare_i_data_rs[0]), .B(n852), .Q(n857) );
  XNR21 U1286 ( .A(compare_i_data_rt[15]), .B(n858), .Q(n1246) );
  XNR21 U1287 ( .A(compare_i_data_rt[14]), .B(n106), .Q(n1247) );
  XNR21 U1288 ( .A(compare_i_data_rt[13]), .B(n100), .Q(n1248) );
  OAI210 U1289 ( .A(n1159), .B(n82), .C(compare_i_data_rs[0]), .Q(n828) );
  IMUX20 U1290 ( .A(n1079), .B(n1076), .S(n1154), .Q(n829) );
  AOI220 U1291 ( .A(n1079), .B(n875), .C(n82), .D(compare_i_data_rs[17]), .Q(
        n878) );
  XNR21 U1292 ( .A(n98), .B(alu_i_data_B[17]), .Q(n875) );
  NOR30 U1293 ( .A(alu_i_data_B[17]), .B(compare_i_data_rs[17]), .C(n1060), 
        .Q(n873) );
  NOR30 U1294 ( .A(n74), .B(n1142), .C(n1087), .Q(n874) );
  OAI220 U1295 ( .A(n103), .B(n520), .C(n1086), .D(n899), .Q(n900) );
  XNR21 U1296 ( .A(compare_i_data_rs[19]), .B(alu_i_data_B[19]), .Q(n899) );
  OAI310 U1297 ( .A(alu_i_data_B[19]), .B(compare_i_data_rs[19]), .C(n1060), 
        .D(n898), .Q(n901) );
  AOI210 U1298 ( .A(n1056), .B(n229), .C(n897), .Q(n898) );
  NOR30 U1299 ( .A(n86), .B(n1140), .C(n1087), .Q(n897) );
  OAI220 U1300 ( .A(n96), .B(n520), .C(n1086), .D(n948), .Q(n949) );
  XNR21 U1301 ( .A(compare_i_data_rs[23]), .B(alu_i_data_B[23]), .Q(n948) );
  AOI210 U1302 ( .A(n1056), .B(alu_i_data_B[7]), .C(n946), .Q(n947) );
  NOR30 U1303 ( .A(n84), .B(n1131), .C(n1087), .Q(n946) );
  OAI220 U1304 ( .A(n887), .B(n520), .C(n1086), .D(n886), .Q(n888) );
  XNR21 U1305 ( .A(compare_i_data_rs[18]), .B(alu_i_data_B[18]), .Q(n886) );
  OAI310 U1306 ( .A(alu_i_data_B[18]), .B(compare_i_data_rs[18]), .C(n1060), 
        .D(n885), .Q(n889) );
  AOI210 U1307 ( .A(n1056), .B(u_alu_lt_x_11_B_2_), .C(n884), .Q(n885) );
  NOR30 U1308 ( .A(n73), .B(n1141), .C(n1087), .Q(n884) );
  OAI220 U1309 ( .A(n104), .B(n520), .C(n1086), .D(n911), .Q(n912) );
  XNR21 U1310 ( .A(compare_i_data_rs[20]), .B(alu_i_data_B[20]), .Q(n911) );
  OAI310 U1311 ( .A(alu_i_data_B[20]), .B(compare_i_data_rs[20]), .C(n1060), 
        .D(n910), .Q(n913) );
  AOI210 U1312 ( .A(n1056), .B(alu_i_data_B[4]), .C(n909), .Q(n910) );
  NOR30 U1313 ( .A(n87), .B(n1134), .C(n1087), .Q(n909) );
  OAI220 U1314 ( .A(n109), .B(n520), .C(n1086), .D(n936), .Q(n937) );
  XNR21 U1315 ( .A(compare_i_data_rs[22]), .B(alu_i_data_B[22]), .Q(n936) );
  OAI310 U1316 ( .A(alu_i_data_B[22]), .B(compare_i_data_rs[22]), .C(n1060), 
        .D(n935), .Q(n938) );
  AOI210 U1317 ( .A(n1056), .B(alu_i_data_B[6]), .C(n934), .Q(n935) );
  NOR30 U1318 ( .A(n85), .B(n1132), .C(n1087), .Q(n934) );
  OAI220 U1319 ( .A(n924), .B(n520), .C(n1086), .D(n923), .Q(n925) );
  XNR21 U1320 ( .A(compare_i_data_rs[21]), .B(alu_i_data_B[21]), .Q(n923) );
  OAI310 U1321 ( .A(alu_i_data_B[21]), .B(compare_i_data_rs[21]), .C(n1060), 
        .D(n922), .Q(n926) );
  AOI210 U1322 ( .A(n1056), .B(alu_i_data_B[5]), .C(n921), .Q(n922) );
  NOR30 U1323 ( .A(n72), .B(n1133), .C(n1087), .Q(n921) );
  NAND20 U1324 ( .A(n1056), .B(alu_i_data_B[8]), .Q(n967) );
  OAI210 U1325 ( .A(alu_i_data_B[24]), .B(n1086), .C(n520), .Q(n969) );
  OAI210 U1326 ( .A(compare_i_data_rs[24]), .B(n1086), .C(n965), .Q(n966) );
  OAI310 U1327 ( .A(n90), .B(n1127), .C(n1087), .D(n1018), .Q(n1019) );
  AOI220 U1328 ( .A(n1076), .B(n1017), .C(n1079), .D(n1016), .Q(n1021) );
  XNR21 U1329 ( .A(n101), .B(alu_i_data_B[28]), .Q(n1016) );
  NAND20 U1330 ( .A(n82), .B(compare_i_data_rs[28]), .Q(n1023) );
  OAI310 U1331 ( .A(n77), .B(n1120), .C(n1087), .D(n1045), .Q(n1046) );
  AOI220 U1332 ( .A(n1076), .B(n1044), .C(n1079), .D(n1043), .Q(n1048) );
  XNR21 U1333 ( .A(n1042), .B(alu_i_data_B[30]), .Q(n1043) );
  NAND20 U1334 ( .A(n82), .B(compare_i_data_rs[30]), .Q(n1050) );
  OAI210 U1335 ( .A(alu_i_data_B[16]), .B(n1086), .C(n520), .Q(n864) );
  OAI220 U1336 ( .A(n993), .B(n520), .C(n1086), .D(n992), .Q(n994) );
  NOR30 U1337 ( .A(n78), .B(n1129), .C(n1087), .Q(n990) );
  OAI220 U1338 ( .A(n1006), .B(n520), .C(n1086), .D(n1005), .Q(n1007) );
  NOR30 U1339 ( .A(n76), .B(n1128), .C(n1087), .Q(n1003) );
  OAI220 U1340 ( .A(n1032), .B(n520), .C(n1086), .D(n1031), .Q(n1033) );
  XNR21 U1341 ( .A(compare_i_data_rs[29]), .B(alu_i_data_B[29]), .Q(n1031) );
  NOR30 U1342 ( .A(n79), .B(n1126), .C(n1087), .Q(n1029) );
  OAI220 U1343 ( .A(n102), .B(n520), .C(n1086), .D(n980), .Q(n981) );
  XNR21 U1344 ( .A(compare_i_data_rs[25]), .B(alu_i_data_B[25]), .Q(n980) );
  NOR30 U1345 ( .A(n88), .B(n1130), .C(n1087), .Q(n978) );
  AOI210 U1346 ( .A(n1079), .B(n1062), .C(n1061), .Q(n1063) );
  NOR30 U1347 ( .A(alu_i_data_B[31]), .B(compare_i_data_rs[31]), .C(n1060), 
        .Q(n1061) );
  XNR21 U1348 ( .A(n99), .B(alu_i_data_B[31]), .Q(n1062) );
  NAND20 U1349 ( .A(n82), .B(compare_i_data_rs[31]), .Q(n1064) );
  OAI310 U1350 ( .A(n1058), .B(n1119), .C(n1087), .D(n1057), .Q(n1059) );
  NAND20 U1351 ( .A(alu_i_con_AluCtrl[3]), .B(n1164), .Q(n1143) );
  INV3 U1352 ( .A(alu_i_con_AluCtrl[1]), .Q(n1081) );
  AOI220 U1353 ( .A(n626), .B(i_data_FMmemout[8]), .C(n625), .D(
        i_data_FMalures[8]), .Q(n598) );
  AOI220 U1354 ( .A(n778), .B(i_data_FMmemout[8]), .C(n777), .D(
        i_data_FMalures[8]), .Q(n745) );
  AOI220 U1355 ( .A(n626), .B(i_data_FMmemout[9]), .C(n625), .D(
        i_data_FMalures[9]), .Q(n595) );
  AOI220 U1356 ( .A(n778), .B(i_data_FMmemout[9]), .C(n777), .D(
        i_data_FMalures[9]), .Q(n741) );
  AOI220 U1357 ( .A(n626), .B(i_data_FMmemout[10]), .C(n625), .D(
        i_data_FMalures[10]), .Q(n592) );
  AOI220 U1358 ( .A(n778), .B(i_data_FMmemout[10]), .C(n777), .D(
        i_data_FMalures[10]), .Q(n737) );
  AOI220 U1359 ( .A(n626), .B(i_data_FMmemout[11]), .C(n625), .D(
        i_data_FMalures[11]), .Q(n589) );
  AOI220 U1360 ( .A(n778), .B(i_data_FMmemout[11]), .C(n777), .D(
        i_data_FMalures[11]), .Q(n733) );
  AOI220 U1361 ( .A(n626), .B(i_data_FMmemout[12]), .C(n625), .D(
        i_data_FMalures[12]), .Q(n586) );
  AOI220 U1362 ( .A(n778), .B(i_data_FMmemout[12]), .C(n777), .D(
        i_data_FMalures[12]), .Q(n729) );
  AOI220 U1363 ( .A(n626), .B(i_data_FMmemout[13]), .C(n625), .D(
        i_data_FMalures[13]), .Q(n583) );
  AOI220 U1364 ( .A(n778), .B(i_data_FMmemout[13]), .C(n777), .D(
        i_data_FMalures[13]), .Q(n725) );
  AOI220 U1365 ( .A(n626), .B(i_data_FMmemout[14]), .C(n625), .D(
        i_data_FMalures[14]), .Q(n580) );
  AOI220 U1366 ( .A(n778), .B(i_data_FMmemout[14]), .C(n777), .D(
        i_data_FMalures[14]), .Q(n721) );
  AOI220 U1367 ( .A(n626), .B(i_data_FMmemout[15]), .C(n625), .D(
        i_data_FMalures[15]), .Q(n577) );
  AOI220 U1368 ( .A(n778), .B(i_data_FMmemout[15]), .C(n777), .D(
        i_data_FMalures[15]), .Q(n717) );
  INV3 U1369 ( .A(n789), .Q(n788) );
  OAI212 U1370 ( .A(n1192), .B(n1191), .C(n1190), .Q(alu_i_con_AluCtrl[1]) );
  INV3 U1371 ( .A(i_data_immext[1]), .Q(n1206) );
  INV3 U1372 ( .A(i_data_immext[5]), .Q(n1210) );
  INV3 U1373 ( .A(i_data_immext[2]), .Q(n1207) );
  INV3 U1374 ( .A(i_data_immext[3]), .Q(n1209) );
  AOI220 U1375 ( .A(n626), .B(i_data_FMmemout[16]), .C(n625), .D(
        i_data_FMalures[16]), .Q(n574) );
  AOI220 U1376 ( .A(n778), .B(i_data_FMmemout[16]), .C(n777), .D(
        i_data_FMalures[16]), .Q(n713) );
  OAI210 U1377 ( .A(n512), .B(n708), .C(n571), .Q(n572) );
  AOI220 U1378 ( .A(n626), .B(i_data_FMmemout[17]), .C(n625), .D(
        i_data_FMalures[17]), .Q(n571) );
  AOI220 U1379 ( .A(n778), .B(i_data_FMmemout[17]), .C(n777), .D(
        i_data_FMalures[17]), .Q(n707) );
  OAI210 U1380 ( .A(n512), .B(n703), .C(n568), .Q(n569) );
  AOI220 U1381 ( .A(n626), .B(i_data_FMmemout[18]), .C(n625), .D(
        i_data_FMalures[18]), .Q(n568) );
  AOI220 U1382 ( .A(n778), .B(i_data_FMmemout[18]), .C(n777), .D(
        i_data_FMalures[18]), .Q(n702) );
  OAI210 U1383 ( .A(n512), .B(n698), .C(n565), .Q(n566) );
  AOI220 U1384 ( .A(n626), .B(i_data_FMmemout[19]), .C(n625), .D(
        i_data_FMalures[19]), .Q(n565) );
  AOI220 U1385 ( .A(n778), .B(i_data_FMmemout[19]), .C(n777), .D(
        i_data_FMalures[19]), .Q(n697) );
  AOI220 U1386 ( .A(n626), .B(i_data_FMmemout[20]), .C(n625), .D(
        i_data_FMalures[20]), .Q(n562) );
  AOI220 U1387 ( .A(n778), .B(i_data_FMmemout[20]), .C(n777), .D(
        i_data_FMalures[20]), .Q(n692) );
  AOI220 U1388 ( .A(n626), .B(i_data_FMmemout[21]), .C(n625), .D(
        i_data_FMalures[21]), .Q(n559) );
  AOI220 U1389 ( .A(n778), .B(i_data_FMmemout[21]), .C(n777), .D(
        i_data_FMalures[21]), .Q(n687) );
  OAI210 U1390 ( .A(n611), .B(n683), .C(n556), .Q(n557) );
  AOI220 U1391 ( .A(n626), .B(i_data_FMmemout[22]), .C(n625), .D(
        i_data_FMalures[22]), .Q(n556) );
  AOI220 U1392 ( .A(n778), .B(i_data_FMmemout[22]), .C(n777), .D(
        i_data_FMalures[22]), .Q(n682) );
  OAI210 U1393 ( .A(n611), .B(n678), .C(n553), .Q(n554) );
  AOI220 U1394 ( .A(n626), .B(i_data_FMmemout[23]), .C(n625), .D(
        i_data_FMalures[23]), .Q(n553) );
  AOI220 U1395 ( .A(n778), .B(i_data_FMmemout[23]), .C(n777), .D(
        i_data_FMalures[23]), .Q(n677) );
  OAI210 U1396 ( .A(n512), .B(n673), .C(n550), .Q(n551) );
  AOI220 U1397 ( .A(n626), .B(i_data_FMmemout[24]), .C(n625), .D(
        i_data_FMalures[24]), .Q(n550) );
  AOI220 U1398 ( .A(n778), .B(i_data_FMmemout[24]), .C(n777), .D(
        i_data_FMalures[24]), .Q(n672) );
  OAI210 U1399 ( .A(n668), .B(n512), .C(n547), .Q(n548) );
  AOI220 U1400 ( .A(n626), .B(i_data_FMmemout[25]), .C(i_data_FMalures[25]), 
        .D(n625), .Q(n547) );
  AOI220 U1401 ( .A(n778), .B(i_data_FMmemout[25]), .C(n777), .D(
        i_data_FMalures[25]), .Q(n667) );
  OAI210 U1402 ( .A(n512), .B(n663), .C(n544), .Q(n545) );
  AOI220 U1403 ( .A(n626), .B(i_data_FMmemout[26]), .C(n625), .D(
        i_data_FMalures[26]), .Q(n544) );
  AOI220 U1404 ( .A(n778), .B(i_data_FMmemout[26]), .C(n777), .D(
        i_data_FMalures[26]), .Q(n662) );
  OAI210 U1405 ( .A(n512), .B(n658), .C(n541), .Q(n542) );
  AOI220 U1406 ( .A(n626), .B(i_data_FMmemout[27]), .C(n625), .D(
        i_data_FMalures[27]), .Q(n541) );
  AOI220 U1407 ( .A(n778), .B(i_data_FMmemout[27]), .C(n777), .D(
        i_data_FMalures[27]), .Q(n657) );
  OAI210 U1408 ( .A(n512), .B(n653), .C(n538), .Q(n539) );
  AOI220 U1409 ( .A(n626), .B(i_data_FMmemout[28]), .C(n625), .D(
        i_data_FMalures[28]), .Q(n538) );
  OAI210 U1410 ( .A(n763), .B(n653), .C(n652), .Q(n654) );
  AOI220 U1411 ( .A(n778), .B(i_data_FMmemout[28]), .C(n777), .D(
        i_data_FMalures[28]), .Q(n652) );
  OAI210 U1412 ( .A(n512), .B(n648), .C(n535), .Q(n536) );
  AOI220 U1413 ( .A(n626), .B(i_data_FMmemout[29]), .C(n625), .D(
        i_data_FMalures[29]), .Q(n535) );
  AOI220 U1414 ( .A(n778), .B(i_data_FMmemout[29]), .C(n777), .D(
        i_data_FMalures[29]), .Q(n647) );
  OAI210 U1415 ( .A(n611), .B(n643), .C(n532), .Q(n533) );
  AOI220 U1416 ( .A(n626), .B(i_data_FMmemout[30]), .C(n625), .D(
        i_data_FMalures[30]), .Q(n532) );
  INV3 U1417 ( .A(n522), .Q(n523) );
  AOI210 U1418 ( .A(n776), .B(i_data_rt[30]), .C(n644), .Q(n645) );
  OAI210 U1419 ( .A(n763), .B(n643), .C(n642), .Q(n644) );
  AOI220 U1420 ( .A(n778), .B(i_data_FMmemout[30]), .C(n777), .D(
        i_data_FMalures[30]), .Q(n642) );
  OAI210 U1421 ( .A(n763), .B(n638), .C(n637), .Q(n639) );
  AOI220 U1422 ( .A(n778), .B(i_data_FMmemout[31]), .C(n777), .D(
        i_data_FMalures[31]), .Q(n637) );
  INV3 U1423 ( .A(n630), .Q(n631) );
  NAND22 U1424 ( .A(n632), .B(n631), .Q(n766) );
  AOI220 U1425 ( .A(n864), .B(compare_i_data_rs[16]), .C(alu_i_data_B[16]), 
        .D(n863), .Q(n871) );
  OAI210 U1426 ( .A(compare_i_data_rs[16]), .B(n1086), .C(n862), .Q(n863) );
  AOI210 U1427 ( .A(n521), .B(compare_i_data_rs[16]), .C(n82), .Q(n862) );
  XNR21 U1428 ( .A(compare_i_data_rs[16]), .B(n830), .Q(n1245) );
  NOR40 U1429 ( .A(u_alu_ashr_4_SH_3_), .B(i_data_immext[8]), .C(n374), .D(
        n237), .Q(n257) );
  NOR20 U1430 ( .A(i_data_immext[10]), .B(n370), .Q(u_alu_N203) );
  NOR20 U1431 ( .A(i_data_immext[10]), .B(n371), .Q(u_alu_N204) );
  MUX21 U1432 ( .A(n285), .B(n355), .S(i_data_immext[10]), .Q(u_alu_N214) );
  IMUX20 U1433 ( .A(n323), .B(n297), .S(i_data_immext[8]), .Q(n299) );
  NAND40 U1434 ( .A(alu_i_data_B[0]), .B(n509), .C(n373), .D(n510), .Q(n300)
         );
  IMUX20 U1435 ( .A(n330), .B(n304), .S(i_data_immext[8]), .Q(n306) );
  MUX21 U1436 ( .A(n309), .B(n359), .S(i_data_immext[10]), .Q(u_alu_N218) );
  IMUX20 U1437 ( .A(n339), .B(n311), .S(i_data_immext[8]), .Q(n313) );
  IMUX20 U1438 ( .A(n347), .B(n317), .S(i_data_immext[8]), .Q(n319) );
  IMUX20 U1439 ( .A(n324), .B(n323), .S(i_data_immext[8]), .Q(n326) );
  IMUX20 U1440 ( .A(n331), .B(n330), .S(i_data_immext[8]), .Q(n333) );
  MUX21 U1441 ( .A(n335), .B(n334), .S(i_data_immext[10]), .Q(u_alu_N222) );
  IMUX20 U1442 ( .A(n340), .B(n339), .S(i_data_immext[8]), .Q(n342) );
  IMUX20 U1443 ( .A(n348), .B(n347), .S(i_data_immext[8]), .Q(n350) );
  NOR20 U1444 ( .A(i_data_immext[10]), .B(n368), .Q(u_alu_N201) );
  MUX21 U1445 ( .A(n390), .B(n443), .S(i_data_immext[10]), .Q(u_alu_N235) );
  MUX21 U1446 ( .A(n391), .B(n444), .S(i_data_immext[10]), .Q(u_alu_N236) );
  MUX21 U1447 ( .A(n407), .B(n406), .S(i_data_immext[8]), .Q(n478) );
  MUX21 U1448 ( .A(n411), .B(n410), .S(i_data_immext[8]), .Q(n483) );
  IMUX20 U1449 ( .A(n424), .B(n473), .S(i_data_immext[8]), .Q(n427) );
  MUX21 U1450 ( .A(n429), .B(n428), .S(i_data_immext[10]), .Q(u_alu_N226) );
  NOR20 U1451 ( .A(i_data_immext[10]), .B(n470), .Q(u_alu_N245) );
  IMUX20 U1452 ( .A(n451), .B(n480), .S(i_data_immext[8]), .Q(n453) );
  MUX21 U1453 ( .A(n455), .B(n454), .S(i_data_immext[10]), .Q(u_alu_N227) );
  IMUX20 U1454 ( .A(n462), .B(n485), .S(i_data_immext[8]), .Q(n464) );
  MUX21 U1455 ( .A(n466), .B(n465), .S(i_data_immext[10]), .Q(u_alu_N228) );
  IMUX30 U1456 ( .A(n469), .B(n468), .C(n467), .S0(i_data_immext[8]), .S1(
        u_alu_ashr_4_SH_3_), .Q(n471) );
  IMUX20 U1457 ( .A(n471), .B(n470), .S(i_data_immext[10]), .Q(u_alu_N229) );
  IMUX20 U1458 ( .A(n473), .B(n472), .S(i_data_immext[8]), .Q(n475) );
  MUX21 U1459 ( .A(n477), .B(n476), .S(i_data_immext[10]), .Q(u_alu_N230) );
  IMUX30 U1460 ( .A(n480), .B(n479), .C(n478), .S0(i_data_immext[8]), .S1(
        u_alu_ashr_4_SH_3_), .Q(n482) );
  IMUX20 U1461 ( .A(n482), .B(n481), .S(i_data_immext[10]), .Q(u_alu_N231) );
  IMUX30 U1462 ( .A(n485), .B(n484), .C(n483), .S0(i_data_immext[8]), .S1(
        u_alu_ashr_4_SH_3_), .Q(n487) );
  IMUX20 U1463 ( .A(n487), .B(n486), .S(i_data_immext[10]), .Q(u_alu_N232) );
  MUX21 U1464 ( .A(n491), .B(n490), .S(i_data_immext[10]), .Q(u_alu_N233) );
  MUX21 U1465 ( .A(n495), .B(n494), .S(i_data_immext[10]), .Q(u_alu_N234) );
  OAI220 U1466 ( .A(n1087), .B(n1093), .C(alu_i_data_B[8]), .D(n1086), .Q(
        n1091) );
  NOR20 U1467 ( .A(n231), .B(alu_i_data_B[8]), .Q(n1093) );
  IMUX20 U1468 ( .A(n1079), .B(n1076), .S(n75), .Q(n1089) );
  OAI210 U1469 ( .A(n82), .B(n1112), .C(compare_i_data_rs[4]), .Q(n1111) );
  NOR20 U1470 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[31]), .Q(n1119)
         );
  NOR20 U1471 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[30]), .Q(n1120)
         );
  NOR20 U1472 ( .A(n231), .B(compare_i_data_rs[29]), .Q(n1126) );
  NOR20 U1473 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[28]), .Q(n1127)
         );
  NOR20 U1474 ( .A(n231), .B(compare_i_data_rs[27]), .Q(n1128) );
  NOR20 U1475 ( .A(n231), .B(compare_i_data_rs[26]), .Q(n1129) );
  NOR20 U1476 ( .A(n231), .B(compare_i_data_rs[25]), .Q(n1130) );
  NOR20 U1477 ( .A(n231), .B(compare_i_data_rs[23]), .Q(n1131) );
  NOR20 U1478 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[22]), .Q(n1132)
         );
  NOR20 U1479 ( .A(n231), .B(compare_i_data_rs[21]), .Q(n1133) );
  NOR20 U1480 ( .A(n231), .B(compare_i_data_rs[20]), .Q(n1134) );
  NOR20 U1481 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[19]), .Q(n1140)
         );
  NOR20 U1482 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[18]), .Q(n1141)
         );
  NOR20 U1483 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[17]), .Q(n1142)
         );
  NAND20 U1484 ( .A(alu_i_con_AluCtrl[2]), .B(n1163), .Q(n1162) );
  NOR20 U1485 ( .A(alu_i_con_AluCtrl[3]), .B(n1081), .Q(n1163) );
  IMAJ30 U1486 ( .A(compare_i_data_rs[31]), .B(u_alu_N306), .C(n1058), .Q(
        n1160) );
  NOR20 U1487 ( .A(alu_i_con_AluCtrl[1]), .B(alu_i_con_AluCtrl[2]), .Q(n1164)
         );
  NOR40 U1488 ( .A(n1172), .B(n1195), .C(n1173), .D(n1168), .Q(n1169) );
  NOR30 U1489 ( .A(i_con_Ealuop[2]), .B(i_con_Ealuop[3]), .C(n1203), .Q(n1188)
         );
  NOR40 U1490 ( .A(n1189), .B(n1188), .C(n1187), .D(n1186), .Q(n1190) );
  IMUX20 U1491 ( .A(i_addr_rt[0]), .B(i_data_immext[11]), .S(i_con_Eregdst), 
        .Q(n1239) );
  IMUX20 U1492 ( .A(i_addr_rt[1]), .B(i_data_immext[12]), .S(i_con_Eregdst), 
        .Q(n1240) );
  IMUX20 U1493 ( .A(i_addr_rt[2]), .B(i_data_immext[13]), .S(i_con_Eregdst), 
        .Q(n1241) );
  IMUX20 U1494 ( .A(i_addr_rt[3]), .B(i_data_immext[14]), .S(i_con_Eregdst), 
        .Q(n1242) );
  IMUX20 U1495 ( .A(i_addr_rt[4]), .B(i_data_immext[15]), .S(i_con_Eregdst), 
        .Q(n1243) );
  NOR40 U1496 ( .A(n1252), .B(n1251), .C(n1250), .D(n1249), .Q(n1260) );
  NOR40 U1497 ( .A(n1256), .B(n1255), .C(n1254), .D(n1253), .Q(n1257) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Mmemread, ex_con_Mmemwrite, ex_con_Malupc8, ex_con_Wmemtoreg,
         mem_con_Malupc8, mem_con_Wmemtoreg, wb_con_Wmemtoreg,
         u_fetch_jmux_i_addr_pc4_3_, u_fetch_jmux_i_addr_pc4_4_,
         u_fetch_jmux_i_addr_pc4_5_, u_fetch_jmux_i_addr_pc4_6_,
         u_fetch_jmux_i_addr_pc4_7_, u_fetch_jmux_i_addr_pc4_8_,
         u_fetch_jmux_i_addr_pc4_9_, u_fetch_jmux_i_addr_pc4_10_,
         u_fetch_jmux_i_addr_pc4_11_, u_fetch_jmux_i_addr_pc4_12_,
         u_fetch_jmux_i_addr_pc4_13_, u_fetch_jmux_i_addr_pc4_14_,
         u_fetch_jmux_i_addr_pc4_15_, u_fetch_jmux_i_addr_pc4_16_,
         u_fetch_jmux_i_addr_pc4_17_, u_fetch_jmux_i_addr_pc4_18_,
         u_fetch_jmux_i_addr_pc4_19_, u_fetch_jmux_i_addr_pc4_20_,
         u_fetch_jmux_i_addr_pc4_21_, u_fetch_jmux_i_addr_pc4_22_,
         u_fetch_jmux_i_addr_pc4_23_, u_fetch_jmux_i_addr_pc4_24_,
         u_fetch_jmux_i_addr_pc4_25_, u_fetch_jmux_i_addr_pc4_26_,
         u_fetch_jmux_i_addr_pc4_27_, u_fetch_jmux_i_addr_pc4_28_,
         u_fetch_jmux_i_addr_pc4_29_, u_fetch_jmux_i_addr_pc4_30_,
         u_fetch_jmux_i_addr_pc4_31_, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, add_x_4_n28, add_x_4_n27, add_x_4_n26, add_x_4_n25,
         add_x_4_n24, add_x_4_n23, add_x_4_n22, add_x_4_n21, add_x_4_n20,
         add_x_4_n19, add_x_4_n18, add_x_4_n17, add_x_4_n16, add_x_4_n15,
         add_x_4_n14, add_x_4_n13, add_x_4_n12, add_x_4_n11, add_x_4_n10,
         add_x_4_n9, add_x_4_n8, add_x_4_n7, add_x_4_n6, add_x_4_n5,
         add_x_4_n4, add_x_4_n3, add_x_4_n2, add_x_4_n1, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20;
  wire   [31:0] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [31:0] id_addr_pc4;
  wire   [31:0] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] wb_data_memout;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [16:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] mem_data_alures;
  wire   [31:2] mem_data_pc4;
  wire   [31:0] u_mem_resmux_o_data_alu;
  wire   [1:0] u_mem_pc8;

  decode u_decode ( .i_clk(clk), .i_nrst(rst_n), .i_addr_pc4(id_addr_pc4), 
        .i_con_Wregwrite(id_con_Wregwrite), .i_data_Wregwrite(
        id_data_Wregwrite), .i_addr_Wregwrite(id_addr_Wregwrite), .i_addr_Erd(
        for_o_addr_Erd), .i_addr_Mrd(mem_addr_regdst), .i_con_Eregwrite(
        ex_con_Wregwrite), .i_con_Mregwrite(mem_con_Wregwrite), .i_addr_rtM(
        for_addr_rtM), .i_addr_rtW(for_addr_rtW), .i_con_memreadM(mem_read), 
        .i_con_memreadW(for_FWmemread), .i_data_Wmemout(wb_data_memout), 
        .o_data_rs(id_data_rs), .o_data_rt(ex_data_rt), .o_addr_rd({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5}), .o_addr_rt(
        ex_addr_rt), .o_data_jr(id_data_jr), .o_con_jump(if_con_j), 
        .o_addr_pc4(ex_data_pc4), .o_addr_branch(if_addr_b), .o_con_Ealuop(
        ex_con_Ealuop), .o_con_Eregdst(ex_con_Eregdst), .o_con_Mmemread(
        ex_con_Mmemread), .o_con_Mmemwrite(ex_con_Mmemwrite), .o_con_Malupc8(
        ex_con_Malupc8), .o_con_Wmemtoreg(ex_con_Wmemtoreg), .o_con_Wregwrite(
        ex_con_Wregwrite), .o_con_ifstall(if_con_ifstall), .o_con_Ebop(
        ex_con_bop), .o_data_signext({SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, ex_data_immext}), .o_con_Efamux(
        for_o_con_Efamux), .o_con_Efbmux(for_o_con_Efbmux), .o_data_Fmemout(
        for_memout), .o_addr_jump_31_(if_addr_j[31]), .o_addr_jump_30_(
        if_addr_j[30]), .o_addr_jump_29_(if_addr_j[29]), .o_addr_jump_28_(
        if_addr_j[28]), .o_addr_jump_27_(if_addr_j[27]), .o_addr_jump_26_(
        if_addr_j[26]), .o_addr_jump_25_(if_addr_j[25]), .o_addr_jump_24_(
        if_addr_j[24]), .o_addr_jump_23_(if_addr_j[23]), .o_addr_jump_22_(
        if_addr_j[22]), .o_addr_jump_21_(if_addr_j[21]), .o_addr_jump_20_(
        if_addr_j[20]), .o_addr_jump_19_(if_addr_j[19]), .o_addr_jump_17_(
        if_addr_j[17]), .o_addr_jump_16_(if_addr_j[16]), .o_addr_jump_15_(
        if_addr_j[15]), .o_addr_jump_14_(if_addr_j[14]), .o_addr_jump_13_(
        if_addr_j[13]), .o_addr_jump_12_(if_addr_j[12]), .o_addr_jump_11_(
        if_addr_j[11]), .o_addr_jump_10_(if_addr_j[10]), .o_addr_jump_9_(
        if_addr_j[9]), .o_addr_jump_8_(if_addr_j[8]), .o_addr_jump_7_(
        if_addr_j[7]), .o_addr_jump_6_(if_addr_j[6]), .o_addr_jump_5_(
        if_addr_j[5]), .o_addr_jump_4_(if_addr_j[4]), .o_addr_jump_3_(
        if_addr_j[3]), .o_addr_jump_2_(if_addr_j[2]), .i_data_instr_31_(
        id_data_instr[31]), .i_data_instr_30_(id_data_instr[30]), 
        .i_data_instr_29_(id_data_instr[29]), .i_data_instr_28_(
        id_data_instr[28]), .i_data_instr_27_(id_data_instr[27]), 
        .i_data_instr_26_(id_data_instr[26]), .i_data_instr_25_(
        id_data_instr[25]), .i_data_instr_24_(id_data_instr[24]), 
        .i_data_instr_23_(id_data_instr[23]), .i_data_instr_22_(
        id_data_instr[22]), .i_data_instr_21_(id_data_instr[21]), 
        .i_data_instr_20_(id_data_instr[20]), .i_data_instr_19_(
        id_data_instr[19]), .i_data_instr_18_(id_data_instr[18]), 
        .i_data_instr_17_(id_data_instr[17]), .i_data_instr_14_(
        id_data_instr[14]), .i_data_instr_13_(id_data_instr[13]), 
        .i_data_instr_12_(id_data_instr[12]), .i_data_instr_11_(
        id_data_instr[11]), .i_data_instr_10_(id_data_instr[10]), 
        .i_data_instr_9_(id_data_instr[9]), .i_data_instr_8_(id_data_instr[8]), 
        .i_data_instr_7_(id_data_instr[7]), .i_data_instr_6_(id_data_instr[6]), 
        .i_data_instr_5_(id_data_instr[5]), .i_data_instr_4_(id_data_instr[4]), 
        .i_data_instr_3_(id_data_instr[3]), .i_data_instr_2_(id_data_instr[2]), 
        .i_data_instr_1_(id_data_instr[1]), .i_data_instr_0_(id_data_instr[0]), 
        .o_addr_jump_18_(if_addr_j[18]), .i_data_instr_16_(id_data_instr[16]), 
        .i_data_instr_15__BAR(n142), .o_con_Ealusrc_BAR(ex_con_Ealusrc) );
  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext({n146, 
        n146, n146, n146, n146, n146, n146, n146, n146, n146, n146, n146, n146, 
        n146, n146, ex_data_immext}), .i_addr_rt(ex_addr_rt), .i_addr_rd({n146, 
        n146, n146, n146, n146}), .i_data_FEalures(data_address), 
        .i_data_FMalures(mem_data_alures), .i_data_FMmemout(wb_data_memout), 
        .i_data_FWmemout(for_memout), .i_con_Efamux(for_o_con_Efamux), 
        .i_con_Efbmux(for_o_con_Efbmux), .i_con_Ealuop(ex_con_Ealuop), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), 
        .i_con_Mmemwrite(ex_con_Mmemwrite), .i_con_Malupc8(ex_con_Malupc8), 
        .i_con_Wmemtoreg(ex_con_Wmemtoreg), .i_con_Wregwrite(ex_con_Wregwrite), 
        .i_con_bop(ex_con_bop), .o_data_alures(data_address), .o_data_rt(
        write_data), .o_addr_regdst(mem_addr_regdst), .o_con_Mmemread(mem_read), .o_con_Mmemwrite(mem_write), .o_con_Malupc8(mem_con_Malupc8), 
        .o_con_Wmemtoreg(mem_con_Wmemtoreg), .o_con_Wregwrite(
        mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), .o_addr_Mrt(
        for_addr_rtM), .o_con_ifbranch(if_con_b), .i_con_Ealusrc_BAR(
        ex_con_Ealusrc), .o_data_pc4_31_(mem_data_pc4[31]), .o_data_pc4_30_(
        mem_data_pc4[30]), .o_data_pc4_29__BAR(mem_data_pc4[29]), 
        .o_data_pc4_28_(mem_data_pc4[28]), .o_data_pc4_26_(mem_data_pc4[26]), 
        .o_data_pc4_24_(mem_data_pc4[24]), .o_data_pc4_22_(mem_data_pc4[22]), 
        .o_data_pc4_20_(mem_data_pc4[20]), .o_data_pc4_18_(mem_data_pc4[18]), 
        .o_data_pc4_16_(mem_data_pc4[16]), .o_data_pc4_14_(mem_data_pc4[14]), 
        .o_data_pc4_12_(mem_data_pc4[12]), .o_data_pc4_10_(mem_data_pc4[10]), 
        .o_data_pc4_8_(mem_data_pc4[8]), .o_data_pc4_6_(mem_data_pc4[6]), 
        .o_data_pc4_4_(mem_data_pc4[4]), .o_data_pc4_3_(mem_data_pc4[3]), 
        .o_data_pc4_2_(mem_data_pc4[2]), .o_data_pc4_1_(u_mem_pc8[1]), 
        .o_data_pc4_0_(u_mem_pc8[0]), .o_data_pc4_27__BAR(mem_data_pc4[27]), 
        .o_data_pc4_25__BAR(mem_data_pc4[25]), .o_data_pc4_23__BAR(
        mem_data_pc4[23]), .o_data_pc4_21__BAR(mem_data_pc4[21]), 
        .o_data_pc4_19__BAR(mem_data_pc4[19]), .o_data_pc4_17__BAR(
        mem_data_pc4[17]), .o_data_pc4_15__BAR(mem_data_pc4[15]), 
        .o_data_pc4_13__BAR(mem_data_pc4[13]), .o_data_pc4_11__BAR(
        mem_data_pc4[11]), .o_data_pc4_9__BAR(mem_data_pc4[9]), 
        .o_data_pc4_7__BAR(mem_data_pc4[7]), .o_data_pc4_5__BAR(
        mem_data_pc4[5]) );
  DFC1 u_fetch_pipe_pc4_reg_0_ ( .D(instruction_address[0]), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[0]) );
  DFC1 u_fetch_pipe_pc4_reg_1_ ( .D(instruction_address[1]), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[1]) );
  DFC1 u_fetch_pipe_pc4_reg_2_ ( .D(n145), .C(clk), .RN(rst_n), .Q(
        id_addr_pc4[2]) );
  DFC1 u_fetch_pipe_pc4_reg_3_ ( .D(u_fetch_jmux_i_addr_pc4_3_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[3]) );
  DFC1 u_fetch_pipe_pc4_reg_4_ ( .D(u_fetch_jmux_i_addr_pc4_4_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[4]) );
  DFC1 u_fetch_pipe_pc4_reg_5_ ( .D(u_fetch_jmux_i_addr_pc4_5_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[5]) );
  DFC1 u_fetch_pipe_pc4_reg_6_ ( .D(u_fetch_jmux_i_addr_pc4_6_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[6]) );
  DFC1 u_fetch_pipe_pc4_reg_7_ ( .D(u_fetch_jmux_i_addr_pc4_7_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[7]) );
  DFC1 u_fetch_pipe_pc4_reg_8_ ( .D(u_fetch_jmux_i_addr_pc4_8_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[8]) );
  DFC1 u_fetch_pipe_pc4_reg_9_ ( .D(u_fetch_jmux_i_addr_pc4_9_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[9]) );
  DFC1 u_fetch_pipe_pc4_reg_10_ ( .D(u_fetch_jmux_i_addr_pc4_10_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[10]) );
  DFC1 u_fetch_pipe_pc4_reg_11_ ( .D(u_fetch_jmux_i_addr_pc4_11_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[11]) );
  DFC1 u_fetch_pipe_pc4_reg_12_ ( .D(u_fetch_jmux_i_addr_pc4_12_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[12]) );
  DFC1 u_fetch_pipe_pc4_reg_13_ ( .D(u_fetch_jmux_i_addr_pc4_13_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[13]) );
  DFC1 u_fetch_pipe_pc4_reg_14_ ( .D(u_fetch_jmux_i_addr_pc4_14_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[14]) );
  DFC1 u_fetch_pipe_pc4_reg_15_ ( .D(u_fetch_jmux_i_addr_pc4_15_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[15]) );
  DFC1 u_fetch_pipe_pc4_reg_16_ ( .D(u_fetch_jmux_i_addr_pc4_16_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[16]) );
  DFC1 u_fetch_pipe_pc4_reg_17_ ( .D(u_fetch_jmux_i_addr_pc4_17_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[17]) );
  DFC1 u_fetch_pipe_pc4_reg_18_ ( .D(u_fetch_jmux_i_addr_pc4_18_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[18]) );
  DFC1 u_fetch_pipe_pc4_reg_19_ ( .D(u_fetch_jmux_i_addr_pc4_19_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[19]) );
  DFC1 u_fetch_pipe_pc4_reg_20_ ( .D(u_fetch_jmux_i_addr_pc4_20_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[20]) );
  DFC1 u_fetch_pipe_pc4_reg_21_ ( .D(u_fetch_jmux_i_addr_pc4_21_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[21]) );
  DFC1 u_fetch_pipe_pc4_reg_22_ ( .D(u_fetch_jmux_i_addr_pc4_22_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[22]) );
  DFC1 u_fetch_pipe_pc4_reg_23_ ( .D(u_fetch_jmux_i_addr_pc4_23_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[23]) );
  DFC1 u_fetch_pipe_pc4_reg_24_ ( .D(u_fetch_jmux_i_addr_pc4_24_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[24]) );
  DFC1 u_fetch_pipe_pc4_reg_25_ ( .D(u_fetch_jmux_i_addr_pc4_25_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[25]) );
  DFC1 u_fetch_pipe_pc4_reg_26_ ( .D(u_fetch_jmux_i_addr_pc4_26_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[26]) );
  DFC1 u_fetch_pipe_pc4_reg_27_ ( .D(u_fetch_jmux_i_addr_pc4_27_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[27]) );
  DFC1 u_fetch_pipe_pc4_reg_28_ ( .D(u_fetch_jmux_i_addr_pc4_28_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[28]) );
  DFC1 u_fetch_pipe_pc4_reg_29_ ( .D(u_fetch_jmux_i_addr_pc4_29_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[29]) );
  DFC1 u_fetch_pipe_pc4_reg_30_ ( .D(u_fetch_jmux_i_addr_pc4_30_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[30]) );
  DFC1 u_fetch_pipe_pc4_reg_31_ ( .D(u_fetch_jmux_i_addr_pc4_31_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[31]) );
  DFC1 u_fetch_pipe_instr_reg_1_ ( .D(read_instruction[1]), .C(clk), .RN(rst_n), .Q(id_data_instr[1]) );
  DFC1 u_fetch_pipe_instr_reg_2_ ( .D(read_instruction[2]), .C(clk), .RN(rst_n), .Q(id_data_instr[2]) );
  DFC1 u_fetch_pipe_instr_reg_3_ ( .D(read_instruction[3]), .C(clk), .RN(rst_n), .Q(id_data_instr[3]) );
  DFC1 u_fetch_pipe_instr_reg_4_ ( .D(read_instruction[4]), .C(clk), .RN(rst_n), .Q(id_data_instr[4]) );
  DFC1 u_fetch_pipe_instr_reg_5_ ( .D(read_instruction[5]), .C(clk), .RN(rst_n), .Q(id_data_instr[5]) );
  DFC1 u_fetch_pipe_instr_reg_6_ ( .D(read_instruction[6]), .C(clk), .RN(rst_n), .Q(id_data_instr[6]) );
  DFC1 u_fetch_pipe_instr_reg_7_ ( .D(read_instruction[7]), .C(clk), .RN(rst_n), .Q(id_data_instr[7]) );
  DFC1 u_fetch_pipe_instr_reg_8_ ( .D(read_instruction[8]), .C(clk), .RN(rst_n), .Q(id_data_instr[8]) );
  DFC1 u_fetch_pipe_instr_reg_9_ ( .D(read_instruction[9]), .C(clk), .RN(rst_n), .Q(id_data_instr[9]) );
  DFC1 u_fetch_pipe_instr_reg_10_ ( .D(read_instruction[10]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[10]) );
  DFC1 u_fetch_pipe_instr_reg_11_ ( .D(read_instruction[11]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[11]) );
  DFC1 u_fetch_pipe_instr_reg_12_ ( .D(read_instruction[12]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[12]) );
  DFC1 u_fetch_pipe_instr_reg_13_ ( .D(read_instruction[13]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[13]) );
  DFC1 u_fetch_pipe_instr_reg_14_ ( .D(read_instruction[14]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[14]) );
  DFC1 u_fetch_pipe_instr_reg_15_ ( .D(read_instruction[15]), .C(clk), .RN(
        rst_n), .QN(n142) );
  DFC1 u_fetch_pipe_instr_reg_16_ ( .D(read_instruction[16]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[16]) );
  DFC1 u_fetch_pipe_instr_reg_17_ ( .D(read_instruction[17]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[17]) );
  DFC1 u_fetch_pipe_instr_reg_18_ ( .D(read_instruction[18]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[18]) );
  DFC1 u_fetch_pipe_instr_reg_20_ ( .D(read_instruction[20]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[20]) );
  DFC1 u_fetch_pipe_instr_reg_21_ ( .D(read_instruction[21]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[21]) );
  DFC1 u_fetch_pipe_instr_reg_22_ ( .D(read_instruction[22]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[22]) );
  DFC1 u_fetch_pipe_instr_reg_23_ ( .D(read_instruction[23]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[23]) );
  DFC1 u_fetch_pipe_instr_reg_24_ ( .D(read_instruction[24]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[24]) );
  DFC1 u_fetch_pipe_instr_reg_26_ ( .D(read_instruction[26]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[26]) );
  DFC1 u_fetch_pipe_instr_reg_27_ ( .D(read_instruction[27]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[27]) );
  DFC1 u_fetch_pipe_instr_reg_28_ ( .D(read_instruction[28]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[28]) );
  DFC1 u_fetch_pipe_instr_reg_29_ ( .D(read_instruction[29]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[29]) );
  DFC1 u_fetch_pipe_instr_reg_30_ ( .D(read_instruction[30]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[30]) );
  DFC1 u_fetch_pipe_instr_reg_31_ ( .D(read_instruction[31]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[31]) );
  DFC1 u_mem_pipe_data_memout_reg_0_ ( .D(read_data[0]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[0]) );
  DFC1 u_mem_pipe_data_memout_reg_1_ ( .D(read_data[1]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[1]) );
  DFC1 u_mem_pipe_data_memout_reg_2_ ( .D(read_data[2]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[2]) );
  DFC1 u_mem_pipe_data_memout_reg_3_ ( .D(read_data[3]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[3]) );
  DFC1 u_mem_pipe_data_memout_reg_4_ ( .D(read_data[4]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[4]) );
  DFC1 u_mem_pipe_data_memout_reg_5_ ( .D(read_data[5]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[5]) );
  DFC1 u_mem_pipe_data_memout_reg_6_ ( .D(read_data[6]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[6]) );
  DFC1 u_mem_pipe_data_memout_reg_7_ ( .D(read_data[7]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[7]) );
  DFC1 u_mem_pipe_data_memout_reg_8_ ( .D(read_data[8]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[8]) );
  DFC1 u_mem_pipe_data_memout_reg_9_ ( .D(read_data[9]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[9]) );
  DFC1 u_mem_pipe_data_memout_reg_10_ ( .D(read_data[10]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[10]) );
  DFC1 u_mem_pipe_data_memout_reg_11_ ( .D(read_data[11]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[11]) );
  DFC1 u_mem_pipe_data_memout_reg_12_ ( .D(read_data[12]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[12]) );
  DFC1 u_mem_pipe_data_memout_reg_13_ ( .D(read_data[13]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[13]) );
  DFC1 u_mem_pipe_data_memout_reg_14_ ( .D(read_data[14]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[14]) );
  DFC1 u_mem_pipe_data_memout_reg_15_ ( .D(read_data[15]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[15]) );
  DFC1 u_mem_pipe_data_memout_reg_16_ ( .D(read_data[16]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[16]) );
  DFC1 u_mem_pipe_data_memout_reg_17_ ( .D(read_data[17]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[17]) );
  DFC1 u_mem_pipe_data_memout_reg_18_ ( .D(read_data[18]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[18]) );
  DFC1 u_mem_pipe_data_memout_reg_19_ ( .D(read_data[19]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[19]) );
  DFC1 u_mem_pipe_data_memout_reg_20_ ( .D(read_data[20]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[20]) );
  DFC1 u_mem_pipe_data_memout_reg_21_ ( .D(read_data[21]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[21]) );
  DFC1 u_mem_pipe_data_memout_reg_22_ ( .D(read_data[22]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[22]) );
  DFC1 u_mem_pipe_data_memout_reg_23_ ( .D(read_data[23]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[23]) );
  DFC1 u_mem_pipe_data_memout_reg_24_ ( .D(read_data[24]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[24]) );
  DFC1 u_mem_pipe_data_memout_reg_25_ ( .D(read_data[25]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[25]) );
  DFC1 u_mem_pipe_data_memout_reg_26_ ( .D(read_data[26]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[26]) );
  DFC1 u_mem_pipe_data_memout_reg_27_ ( .D(read_data[27]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[27]) );
  DFC1 u_mem_pipe_data_memout_reg_28_ ( .D(read_data[28]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[28]) );
  DFC1 u_mem_pipe_data_memout_reg_29_ ( .D(read_data[29]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[29]) );
  DFC1 u_mem_pipe_data_memout_reg_30_ ( .D(read_data[30]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[30]) );
  DFC1 u_mem_pipe_data_memout_reg_31_ ( .D(read_data[31]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[31]) );
  DFC1 u_mem_pipe_rt_reg_4_ ( .D(for_addr_rtM[4]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[4]) );
  DFC1 u_mem_pipe_con_FWmemread_reg ( .D(ex_con_Mmemread), .C(clk), .RN(rst_n), 
        .Q(for_FWmemread) );
  DFC1 u_mem_pipe_rt_reg_0_ ( .D(for_addr_rtM[0]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[0]) );
  DFC1 u_mem_pipe_rt_reg_1_ ( .D(for_addr_rtM[1]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[1]) );
  DFC1 u_mem_pipe_rt_reg_2_ ( .D(for_addr_rtM[2]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[2]) );
  DFC1 u_mem_pipe_rt_reg_3_ ( .D(for_addr_rtM[3]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[3]) );
  DFC1 u_mem_pipe_con_Wregwrite_reg ( .D(mem_con_Wregwrite), .C(clk), .RN(
        rst_n), .Q(id_con_Wregwrite) );
  DFC1 u_mem_pipe_addr_regdst_reg_1_ ( .D(mem_addr_regdst[1]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[1]) );
  DFC1 u_mem_pipe_addr_regdst_reg_2_ ( .D(mem_addr_regdst[2]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[2]) );
  DFC1 u_mem_pipe_addr_regdst_reg_4_ ( .D(mem_addr_regdst[4]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[4]) );
  DFC1 u_mem_pipe_data_alures_reg_0_ ( .D(u_mem_resmux_o_data_alu[0]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[0]) );
  DFC1 u_mem_pipe_data_alures_reg_1_ ( .D(u_mem_resmux_o_data_alu[1]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[1]) );
  DFC1 u_mem_pipe_data_alures_reg_2_ ( .D(u_mem_resmux_o_data_alu[2]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[2]) );
  DFC1 u_mem_pipe_data_alures_reg_3_ ( .D(u_mem_resmux_o_data_alu[3]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[3]) );
  DFC1 u_mem_pipe_data_alures_reg_4_ ( .D(u_mem_resmux_o_data_alu[4]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[4]) );
  DFC1 u_mem_pipe_data_alures_reg_5_ ( .D(u_mem_resmux_o_data_alu[5]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[5]) );
  DFC1 u_mem_pipe_data_alures_reg_6_ ( .D(u_mem_resmux_o_data_alu[6]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[6]) );
  DFC1 u_mem_pipe_data_alures_reg_7_ ( .D(u_mem_resmux_o_data_alu[7]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[7]) );
  DFC1 u_mem_pipe_data_alures_reg_8_ ( .D(u_mem_resmux_o_data_alu[8]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[8]) );
  DFC1 u_mem_pipe_data_alures_reg_9_ ( .D(u_mem_resmux_o_data_alu[9]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[9]) );
  DFC1 u_mem_pipe_data_alures_reg_10_ ( .D(u_mem_resmux_o_data_alu[10]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[10]) );
  DFC1 u_mem_pipe_data_alures_reg_11_ ( .D(u_mem_resmux_o_data_alu[11]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[11]) );
  DFC1 u_mem_pipe_data_alures_reg_12_ ( .D(u_mem_resmux_o_data_alu[12]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[12]) );
  DFC1 u_mem_pipe_data_alures_reg_13_ ( .D(u_mem_resmux_o_data_alu[13]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[13]) );
  DFC1 u_mem_pipe_data_alures_reg_14_ ( .D(u_mem_resmux_o_data_alu[14]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[14]) );
  DFC1 u_mem_pipe_data_alures_reg_15_ ( .D(u_mem_resmux_o_data_alu[15]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[15]) );
  DFC1 u_mem_pipe_data_alures_reg_16_ ( .D(u_mem_resmux_o_data_alu[16]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[16]) );
  DFC1 u_mem_pipe_data_alures_reg_17_ ( .D(u_mem_resmux_o_data_alu[17]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[17]) );
  DFC1 u_mem_pipe_data_alures_reg_18_ ( .D(u_mem_resmux_o_data_alu[18]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[18]) );
  DFC1 u_mem_pipe_data_alures_reg_19_ ( .D(u_mem_resmux_o_data_alu[19]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[19]) );
  DFC1 u_mem_pipe_data_alures_reg_20_ ( .D(u_mem_resmux_o_data_alu[20]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[20]) );
  DFC1 u_mem_pipe_data_alures_reg_21_ ( .D(u_mem_resmux_o_data_alu[21]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[21]) );
  DFC1 u_mem_pipe_data_alures_reg_22_ ( .D(u_mem_resmux_o_data_alu[22]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[22]) );
  DFC1 u_mem_pipe_data_alures_reg_23_ ( .D(u_mem_resmux_o_data_alu[23]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[23]) );
  DFC1 u_mem_pipe_data_alures_reg_24_ ( .D(u_mem_resmux_o_data_alu[24]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[24]) );
  DFC1 u_mem_pipe_data_alures_reg_25_ ( .D(u_mem_resmux_o_data_alu[25]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[25]) );
  DFC1 u_mem_pipe_data_alures_reg_26_ ( .D(u_mem_resmux_o_data_alu[26]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[26]) );
  DFC1 u_mem_pipe_data_alures_reg_27_ ( .D(u_mem_resmux_o_data_alu[27]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[27]) );
  DFC1 u_mem_pipe_data_alures_reg_28_ ( .D(u_mem_resmux_o_data_alu[28]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[28]) );
  DFC1 u_mem_pipe_data_alures_reg_29_ ( .D(u_mem_resmux_o_data_alu[29]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[29]) );
  DFC1 u_mem_pipe_data_alures_reg_30_ ( .D(u_mem_resmux_o_data_alu[30]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[30]) );
  DFC1 u_mem_pipe_data_alures_reg_31_ ( .D(u_mem_resmux_o_data_alu[31]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[31]) );
  DFC1 u_fetch_u_pc_program_counter_reg_0_ ( .D(n137), .C(clk), .RN(rst_n), 
        .Q(instruction_address[0]), .QN(n143) );
  DFC1 u_fetch_u_pc_program_counter_reg_1_ ( .D(n136), .C(clk), .RN(rst_n), 
        .Q(instruction_address[1]), .QN(n144) );
  DFC1 u_fetch_u_pc_program_counter_reg_4_ ( .D(n133), .C(clk), .RN(rst_n), 
        .Q(instruction_address[4]) );
  DFC1 u_fetch_u_pc_program_counter_reg_5_ ( .D(n132), .C(clk), .RN(rst_n), 
        .Q(instruction_address[5]) );
  DFC1 u_fetch_u_pc_program_counter_reg_6_ ( .D(n131), .C(clk), .RN(rst_n), 
        .Q(instruction_address[6]) );
  DFC1 u_fetch_u_pc_program_counter_reg_7_ ( .D(n130), .C(clk), .RN(rst_n), 
        .Q(instruction_address[7]) );
  DFC1 u_fetch_u_pc_program_counter_reg_8_ ( .D(n129), .C(clk), .RN(rst_n), 
        .Q(instruction_address[8]) );
  DFC1 u_fetch_u_pc_program_counter_reg_9_ ( .D(n128), .C(clk), .RN(rst_n), 
        .Q(instruction_address[9]) );
  DFC1 u_fetch_u_pc_program_counter_reg_10_ ( .D(n127), .C(clk), .RN(rst_n), 
        .Q(instruction_address[10]) );
  DFC1 u_fetch_u_pc_program_counter_reg_11_ ( .D(n126), .C(clk), .RN(rst_n), 
        .Q(instruction_address[11]) );
  DFC1 u_fetch_u_pc_program_counter_reg_12_ ( .D(n125), .C(clk), .RN(rst_n), 
        .Q(instruction_address[12]) );
  DFC1 u_fetch_u_pc_program_counter_reg_13_ ( .D(n124), .C(clk), .RN(rst_n), 
        .Q(instruction_address[13]) );
  DFC1 u_fetch_u_pc_program_counter_reg_14_ ( .D(n123), .C(clk), .RN(rst_n), 
        .Q(instruction_address[14]) );
  DFC1 u_fetch_u_pc_program_counter_reg_15_ ( .D(n122), .C(clk), .RN(rst_n), 
        .Q(instruction_address[15]) );
  DFC1 u_fetch_u_pc_program_counter_reg_16_ ( .D(n121), .C(clk), .RN(rst_n), 
        .Q(instruction_address[16]) );
  DFC1 u_fetch_u_pc_program_counter_reg_17_ ( .D(n120), .C(clk), .RN(rst_n), 
        .Q(instruction_address[17]) );
  DFC1 u_fetch_u_pc_program_counter_reg_18_ ( .D(n119), .C(clk), .RN(rst_n), 
        .Q(instruction_address[18]) );
  DFC1 u_fetch_u_pc_program_counter_reg_19_ ( .D(n118), .C(clk), .RN(rst_n), 
        .Q(instruction_address[19]) );
  DFC1 u_fetch_u_pc_program_counter_reg_20_ ( .D(n117), .C(clk), .RN(rst_n), 
        .Q(instruction_address[20]) );
  DFC1 u_fetch_u_pc_program_counter_reg_21_ ( .D(n116), .C(clk), .RN(rst_n), 
        .Q(instruction_address[21]) );
  DFC1 u_fetch_u_pc_program_counter_reg_22_ ( .D(n115), .C(clk), .RN(rst_n), 
        .Q(instruction_address[22]) );
  DFC1 u_fetch_u_pc_program_counter_reg_23_ ( .D(n114), .C(clk), .RN(rst_n), 
        .Q(instruction_address[23]) );
  DFC1 u_fetch_u_pc_program_counter_reg_24_ ( .D(n113), .C(clk), .RN(rst_n), 
        .Q(instruction_address[24]) );
  DFC1 u_fetch_u_pc_program_counter_reg_25_ ( .D(n112), .C(clk), .RN(rst_n), 
        .Q(instruction_address[25]) );
  DFC1 u_fetch_u_pc_program_counter_reg_26_ ( .D(n111), .C(clk), .RN(rst_n), 
        .Q(instruction_address[26]) );
  DFC1 u_fetch_u_pc_program_counter_reg_27_ ( .D(n110), .C(clk), .RN(rst_n), 
        .Q(instruction_address[27]) );
  DFC1 u_fetch_u_pc_program_counter_reg_28_ ( .D(n109), .C(clk), .RN(rst_n), 
        .Q(instruction_address[28]) );
  DFC1 u_fetch_u_pc_program_counter_reg_29_ ( .D(n108), .C(clk), .RN(rst_n), 
        .Q(instruction_address[29]) );
  DFC1 u_fetch_u_pc_program_counter_reg_30_ ( .D(n107), .C(clk), .RN(rst_n), 
        .Q(instruction_address[30]) );
  DFC1 u_fetch_u_pc_program_counter_reg_31_ ( .D(n138), .C(clk), .RN(rst_n), 
        .Q(instruction_address[31]) );
  DFC3 u_fetch_pipe_instr_reg_0_ ( .D(read_instruction[0]), .C(clk), .RN(rst_n), .Q(id_data_instr[0]) );
  DFC3 u_mem_pipe_con_Wmemtoreg_reg ( .D(mem_con_Wmemtoreg), .C(clk), .RN(
        rst_n), .Q(wb_con_Wmemtoreg) );
  ADD22 add_x_4_U3 ( .A(add_x_4_n3), .B(instruction_address[29]), .CO(
        add_x_4_n2), .S(u_fetch_jmux_i_addr_pc4_29_) );
  ADD22 add_x_4_U2 ( .A(add_x_4_n2), .B(instruction_address[30]), .CO(
        add_x_4_n1), .S(u_fetch_jmux_i_addr_pc4_30_) );
  ADD22 add_x_4_U8 ( .A(add_x_4_n8), .B(instruction_address[24]), .CO(
        add_x_4_n7), .S(u_fetch_jmux_i_addr_pc4_24_) );
  ADD22 add_x_4_U7 ( .A(add_x_4_n7), .B(instruction_address[25]), .CO(
        add_x_4_n6), .S(u_fetch_jmux_i_addr_pc4_25_) );
  ADD22 add_x_4_U5 ( .A(add_x_4_n5), .B(instruction_address[27]), .CO(
        add_x_4_n4), .S(u_fetch_jmux_i_addr_pc4_27_) );
  ADD22 add_x_4_U4 ( .A(add_x_4_n4), .B(instruction_address[28]), .CO(
        add_x_4_n3), .S(u_fetch_jmux_i_addr_pc4_28_) );
  DFC3 u_fetch_u_pc_program_counter_reg_2_ ( .D(n135), .C(clk), .RN(rst_n), 
        .Q(instruction_address[2]), .QN(n145) );
  DFC3 u_fetch_u_pc_program_counter_reg_3_ ( .D(n134), .C(clk), .RN(rst_n), 
        .Q(instruction_address[3]) );
  DFC3 u_fetch_pipe_instr_reg_19_ ( .D(read_instruction[19]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[19]) );
  DFC3 u_fetch_pipe_instr_reg_25_ ( .D(read_instruction[25]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[25]) );
  DFC3 u_mem_pipe_addr_regdst_reg_0_ ( .D(mem_addr_regdst[0]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[0]) );
  DFC3 u_mem_pipe_addr_regdst_reg_3_ ( .D(mem_addr_regdst[3]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[3]) );
  ADD22 add_x_4_U28 ( .A(add_x_4_n28), .B(instruction_address[4]), .CO(
        add_x_4_n27), .S(u_fetch_jmux_i_addr_pc4_4_) );
  ADD22 add_x_4_U27 ( .A(add_x_4_n27), .B(instruction_address[5]), .CO(
        add_x_4_n26), .S(u_fetch_jmux_i_addr_pc4_5_) );
  ADD22 add_x_4_U26 ( .A(add_x_4_n26), .B(instruction_address[6]), .CO(
        add_x_4_n25), .S(u_fetch_jmux_i_addr_pc4_6_) );
  ADD22 add_x_4_U25 ( .A(add_x_4_n25), .B(instruction_address[7]), .CO(
        add_x_4_n24), .S(u_fetch_jmux_i_addr_pc4_7_) );
  ADD22 add_x_4_U24 ( .A(add_x_4_n24), .B(instruction_address[8]), .CO(
        add_x_4_n23), .S(u_fetch_jmux_i_addr_pc4_8_) );
  ADD22 add_x_4_U23 ( .A(add_x_4_n23), .B(instruction_address[9]), .CO(
        add_x_4_n22), .S(u_fetch_jmux_i_addr_pc4_9_) );
  ADD22 add_x_4_U22 ( .A(add_x_4_n22), .B(instruction_address[10]), .CO(
        add_x_4_n21), .S(u_fetch_jmux_i_addr_pc4_10_) );
  ADD22 add_x_4_U21 ( .A(add_x_4_n21), .B(instruction_address[11]), .CO(
        add_x_4_n20), .S(u_fetch_jmux_i_addr_pc4_11_) );
  ADD22 add_x_4_U20 ( .A(add_x_4_n20), .B(instruction_address[12]), .CO(
        add_x_4_n19), .S(u_fetch_jmux_i_addr_pc4_12_) );
  ADD22 add_x_4_U17 ( .A(add_x_4_n17), .B(instruction_address[15]), .CO(
        add_x_4_n16), .S(u_fetch_jmux_i_addr_pc4_15_) );
  ADD22 add_x_4_U16 ( .A(add_x_4_n16), .B(instruction_address[16]), .CO(
        add_x_4_n15), .S(u_fetch_jmux_i_addr_pc4_16_) );
  ADD22 add_x_4_U15 ( .A(add_x_4_n15), .B(instruction_address[17]), .CO(
        add_x_4_n14), .S(u_fetch_jmux_i_addr_pc4_17_) );
  ADD22 add_x_4_U14 ( .A(add_x_4_n14), .B(instruction_address[18]), .CO(
        add_x_4_n13), .S(u_fetch_jmux_i_addr_pc4_18_) );
  ADD22 add_x_4_U13 ( .A(add_x_4_n13), .B(instruction_address[19]), .CO(
        add_x_4_n12), .S(u_fetch_jmux_i_addr_pc4_19_) );
  ADD22 add_x_4_U12 ( .A(add_x_4_n12), .B(instruction_address[20]), .CO(
        add_x_4_n11), .S(u_fetch_jmux_i_addr_pc4_20_) );
  ADD22 add_x_4_U11 ( .A(add_x_4_n11), .B(instruction_address[21]), .CO(
        add_x_4_n10), .S(u_fetch_jmux_i_addr_pc4_21_) );
  ADD22 add_x_4_U6 ( .A(add_x_4_n6), .B(instruction_address[26]), .CO(
        add_x_4_n5), .S(u_fetch_jmux_i_addr_pc4_26_) );
  BUF2 U204 ( .A(n245), .Q(n148) );
  BUF2 U205 ( .A(n244), .Q(n147) );
  OAI220 U206 ( .A(if_con_j[0]), .B(n149), .C(if_con_j[1]), .D(n155), .Q(n140)
         );
  NOR30 U207 ( .A(if_con_b), .B(n242), .C(n140), .Q(n154) );
  XNR20 U208 ( .A(mem_data_pc4[31]), .B(n303), .Q(n141) );
  MUX21 U209 ( .A(data_address[31]), .B(n141), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[31]) );
  AOI221 U210 ( .A(n148), .B(id_data_jr[27]), .C(n147), .D(if_addr_j[27]), .Q(
        n233) );
  AOI221 U211 ( .A(n148), .B(id_data_jr[19]), .C(n147), .D(if_addr_j[19]), .Q(
        n209) );
  AOI220 U212 ( .A(n148), .B(id_data_jr[15]), .C(n147), .D(if_addr_j[15]), .Q(
        n197) );
  AOI221 U213 ( .A(n148), .B(id_data_jr[18]), .C(n147), .D(if_addr_j[18]), .Q(
        n206) );
  IMUX21 U214 ( .A(n281), .B(n280), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[22]) );
  AOI220 U215 ( .A(n148), .B(id_data_jr[12]), .C(n147), .D(if_addr_j[12]), .Q(
        n188) );
  AOI220 U216 ( .A(n148), .B(id_data_jr[11]), .C(n147), .D(if_addr_j[11]), .Q(
        n185) );
  OAI210 U217 ( .A(n307), .B(mem_data_pc4[4]), .C(n310), .Q(n308) );
  INV1 U218 ( .A(data_address[22]), .Q(n281) );
  INV1 U219 ( .A(data_address[2]), .Q(n299) );
  INV1 U220 ( .A(data_address[16]), .Q(n266) );
  MUX22 U221 ( .A(data_address[27]), .B(n293), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[27]) );
  MUX22 U222 ( .A(data_address[25]), .B(n288), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[25]) );
  IMUX21 U223 ( .A(n286), .B(n285), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[24]) );
  AOI220 U224 ( .A(n148), .B(id_data_jr[14]), .C(n147), .D(if_addr_j[14]), .Q(
        n194) );
  AOI220 U225 ( .A(n148), .B(id_data_jr[13]), .C(n147), .D(if_addr_j[13]), .Q(
        n191) );
  AOI221 U226 ( .A(n148), .B(id_data_jr[21]), .C(n147), .D(if_addr_j[21]), .Q(
        n215) );
  INV1 U227 ( .A(data_address[3]), .Q(n305) );
  INV1 U228 ( .A(data_address[8]), .Q(n319) );
  NAND21 U229 ( .A(mem_data_pc4[2]), .B(mem_data_pc4[3]), .Q(n304) );
  OAI2111 U230 ( .A(n249), .B(n158), .C(n157), .D(n156), .Q(n138) );
  INV2 U231 ( .A(u_fetch_jmux_i_addr_pc4_31_), .Q(n158) );
  IMUX21 U232 ( .A(n302), .B(n301), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[30]) );
  XOR21 U233 ( .A(add_x_4_n1), .B(instruction_address[31]), .Q(
        u_fetch_jmux_i_addr_pc4_31_) );
  INV2 U234 ( .A(u_fetch_jmux_i_addr_pc4_30_), .Q(n248) );
  INV2 U235 ( .A(u_fetch_jmux_i_addr_pc4_29_), .Q(n241) );
  MUX22 U236 ( .A(data_address[29]), .B(n298), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[29]) );
  OAI211 U237 ( .A(n300), .B(mem_data_pc4[30]), .C(n303), .Q(n301) );
  IMUX21 U238 ( .A(n296), .B(n295), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[28]) );
  INV2 U239 ( .A(u_fetch_jmux_i_addr_pc4_28_), .Q(n238) );
  INV2 U240 ( .A(u_fetch_jmux_i_addr_pc4_27_), .Q(n235) );
  INV2 U241 ( .A(u_fetch_jmux_i_addr_pc4_26_), .Q(n232) );
  IMUX21 U242 ( .A(n291), .B(n290), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[26]) );
  INV2 U243 ( .A(u_fetch_jmux_i_addr_pc4_25_), .Q(n229) );
  INV2 U244 ( .A(u_fetch_jmux_i_addr_pc4_24_), .Q(n226) );
  OAI2111 U245 ( .A(instruction_address[2]), .B(n249), .C(n160), .D(n159), .Q(
        n135) );
  OAI211 U246 ( .A(n153), .B(n143), .C(n151), .Q(n137) );
  OAI211 U247 ( .A(n153), .B(n144), .C(n152), .Q(n136) );
  INV2 U248 ( .A(u_fetch_jmux_i_addr_pc4_23_), .Q(n223) );
  AOI220 U249 ( .A(n148), .B(id_data_jr[17]), .C(n147), .D(if_addr_j[17]), .Q(
        n203) );
  AOI221 U250 ( .A(n148), .B(id_data_jr[30]), .C(n147), .D(if_addr_j[30]), .Q(
        n246) );
  AOI221 U251 ( .A(n148), .B(id_data_jr[9]), .C(n147), .D(if_addr_j[9]), .Q(
        n179) );
  AOI221 U252 ( .A(n148), .B(id_data_jr[29]), .C(n147), .D(if_addr_j[29]), .Q(
        n239) );
  INV2 U253 ( .A(u_fetch_jmux_i_addr_pc4_22_), .Q(n220) );
  AOI221 U254 ( .A(n148), .B(id_data_jr[10]), .C(n147), .D(if_addr_j[10]), .Q(
        n182) );
  AOI221 U255 ( .A(n148), .B(id_data_jr[31]), .C(n147), .D(if_addr_j[31]), .Q(
        n156) );
  NOR20 U256 ( .A(n154), .B(n242), .Q(n153) );
  INV2 U257 ( .A(u_fetch_jmux_i_addr_pc4_21_), .Q(n217) );
  INV3 U258 ( .A(n150), .Q(n243) );
  INV3 U259 ( .A(n154), .Q(n249) );
  INV2 U260 ( .A(u_fetch_jmux_i_addr_pc4_20_), .Q(n214) );
  INV2 U261 ( .A(u_fetch_jmux_i_addr_pc4_19_), .Q(n211) );
  INV2 U262 ( .A(u_fetch_jmux_i_addr_pc4_18_), .Q(n208) );
  INV2 U263 ( .A(u_fetch_jmux_i_addr_pc4_17_), .Q(n205) );
  INV2 U264 ( .A(u_fetch_jmux_i_addr_pc4_16_), .Q(n202) );
  INV2 U265 ( .A(u_fetch_jmux_i_addr_pc4_15_), .Q(n199) );
  INV2 U266 ( .A(u_fetch_jmux_i_addr_pc4_14_), .Q(n196) );
  INV2 U267 ( .A(u_fetch_jmux_i_addr_pc4_13_), .Q(n193) );
  INV2 U268 ( .A(u_fetch_jmux_i_addr_pc4_12_), .Q(n190) );
  INV2 U269 ( .A(u_fetch_jmux_i_addr_pc4_11_), .Q(n187) );
  INV2 U270 ( .A(u_fetch_jmux_i_addr_pc4_10_), .Q(n184) );
  INV2 U271 ( .A(u_fetch_jmux_i_addr_pc4_9_), .Q(n181) );
  INV2 U272 ( .A(u_fetch_jmux_i_addr_pc4_8_), .Q(n178) );
  INV2 U273 ( .A(u_fetch_jmux_i_addr_pc4_7_), .Q(n175) );
  INV2 U274 ( .A(u_fetch_jmux_i_addr_pc4_6_), .Q(n172) );
  INV2 U275 ( .A(u_fetch_jmux_i_addr_pc4_5_), .Q(n169) );
  INV2 U276 ( .A(u_fetch_jmux_i_addr_pc4_4_), .Q(n166) );
  INV2 U277 ( .A(u_fetch_jmux_i_addr_pc4_3_), .Q(n163) );
  INV1 U278 ( .A(data_address[6]), .Q(n314) );
  INV1 U279 ( .A(data_address[4]), .Q(n309) );
  INV2 U280 ( .A(data_address[26]), .Q(n291) );
  INV1 U281 ( .A(data_address[12]), .Q(n256) );
  MUX22 U282 ( .A(mem_data_alures[27]), .B(wb_data_memout[27]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[27]) );
  MUX22 U283 ( .A(mem_data_alures[28]), .B(wb_data_memout[28]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[28]) );
  INV2 U284 ( .A(data_address[18]), .Q(n271) );
  MUX22 U285 ( .A(mem_data_alures[17]), .B(wb_data_memout[17]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[17]) );
  MUX22 U286 ( .A(mem_data_alures[18]), .B(wb_data_memout[18]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[18]) );
  MUX22 U287 ( .A(mem_data_alures[5]), .B(wb_data_memout[5]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[5]) );
  MUX22 U288 ( .A(mem_data_alures[30]), .B(wb_data_memout[30]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[30]) );
  MUX22 U289 ( .A(mem_data_alures[1]), .B(wb_data_memout[1]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[1]) );
  MUX22 U290 ( .A(mem_data_alures[20]), .B(wb_data_memout[20]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[20]) );
  MUX22 U291 ( .A(mem_data_alures[6]), .B(wb_data_memout[6]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[6]) );
  MUX22 U292 ( .A(mem_data_alures[7]), .B(wb_data_memout[7]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[7]) );
  MUX22 U293 ( .A(mem_data_alures[29]), .B(wb_data_memout[29]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[29]) );
  MUX22 U294 ( .A(mem_data_alures[26]), .B(wb_data_memout[26]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[26]) );
  INV1 U295 ( .A(data_address[10]), .Q(n251) );
  MUX22 U296 ( .A(mem_data_alures[19]), .B(wb_data_memout[19]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[19]) );
  MUX22 U297 ( .A(mem_data_alures[31]), .B(wb_data_memout[31]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[31]) );
  MUX22 U298 ( .A(mem_data_alures[8]), .B(wb_data_memout[8]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[8]) );
  MUX22 U299 ( .A(mem_data_alures[9]), .B(wb_data_memout[9]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[9]) );
  MUX22 U300 ( .A(mem_data_alures[14]), .B(wb_data_memout[14]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[14]) );
  MUX22 U301 ( .A(mem_data_alures[13]), .B(wb_data_memout[13]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[13]) );
  MUX22 U302 ( .A(mem_data_alures[15]), .B(wb_data_memout[15]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[15]) );
  MUX22 U303 ( .A(mem_data_alures[24]), .B(wb_data_memout[24]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[24]) );
  MUX22 U304 ( .A(mem_data_alures[10]), .B(wb_data_memout[10]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[10]) );
  MUX22 U305 ( .A(mem_data_alures[0]), .B(wb_data_memout[0]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[0]) );
  MUX22 U306 ( .A(mem_data_alures[3]), .B(wb_data_memout[3]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[3]) );
  MUX22 U307 ( .A(mem_data_alures[21]), .B(wb_data_memout[21]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[21]) );
  MUX22 U308 ( .A(mem_data_alures[23]), .B(wb_data_memout[23]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[23]) );
  MUX22 U309 ( .A(mem_data_alures[25]), .B(wb_data_memout[25]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[25]) );
  MUX22 U310 ( .A(mem_data_alures[2]), .B(wb_data_memout[2]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[2]) );
  MUX22 U311 ( .A(mem_data_alures[11]), .B(wb_data_memout[11]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[11]) );
  MUX22 U312 ( .A(mem_data_alures[4]), .B(wb_data_memout[4]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[4]) );
  MUX22 U313 ( .A(mem_data_alures[22]), .B(wb_data_memout[22]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[22]) );
  MUX22 U314 ( .A(mem_data_alures[16]), .B(wb_data_memout[16]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[16]) );
  INV2 U315 ( .A(data_address[30]), .Q(n302) );
  MUX22 U316 ( .A(mem_data_alures[12]), .B(wb_data_memout[12]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[12]) );
  INV2 U317 ( .A(data_address[20]), .Q(n276) );
  INV2 U318 ( .A(data_address[28]), .Q(n296) );
  INV1 U319 ( .A(data_address[14]), .Q(n261) );
  INV2 U320 ( .A(data_address[24]), .Q(n286) );
  ADD22 U321 ( .A(add_x_4_n18), .B(instruction_address[14]), .CO(add_x_4_n17), 
        .S(u_fetch_jmux_i_addr_pc4_14_) );
  ADD22 U322 ( .A(add_x_4_n19), .B(instruction_address[13]), .CO(add_x_4_n18), 
        .S(u_fetch_jmux_i_addr_pc4_13_) );
  ADD22 U323 ( .A(instruction_address[2]), .B(instruction_address[3]), .CO(
        add_x_4_n28), .S(u_fetch_jmux_i_addr_pc4_3_) );
  ADD22 U324 ( .A(add_x_4_n9), .B(instruction_address[23]), .CO(add_x_4_n8), 
        .S(u_fetch_jmux_i_addr_pc4_23_) );
  ADD22 U325 ( .A(add_x_4_n10), .B(instruction_address[22]), .CO(add_x_4_n9), 
        .S(u_fetch_jmux_i_addr_pc4_22_) );
  NOR21 U326 ( .A(n282), .B(mem_data_pc4[23]), .Q(n284) );
  NOR21 U327 ( .A(n277), .B(mem_data_pc4[21]), .Q(n279) );
  NOR21 U328 ( .A(n272), .B(mem_data_pc4[19]), .Q(n274) );
  NOR21 U329 ( .A(n267), .B(mem_data_pc4[17]), .Q(n269) );
  NOR21 U330 ( .A(n262), .B(mem_data_pc4[15]), .Q(n264) );
  NOR21 U331 ( .A(n257), .B(mem_data_pc4[13]), .Q(n259) );
  NOR21 U332 ( .A(n252), .B(mem_data_pc4[11]), .Q(n254) );
  NOR21 U333 ( .A(n321), .B(mem_data_pc4[9]), .Q(n320) );
  NOR21 U334 ( .A(n315), .B(mem_data_pc4[7]), .Q(n317) );
  INV3 U335 ( .A(if_con_ifstall), .Q(n242) );
  AOI210 U336 ( .A(n292), .B(mem_data_pc4[27]), .C(n294), .Q(n293) );
  NOR21 U337 ( .A(n292), .B(mem_data_pc4[27]), .Q(n294) );
  NOR21 U338 ( .A(n287), .B(mem_data_pc4[25]), .Q(n289) );
  AOI210 U339 ( .A(n287), .B(mem_data_pc4[25]), .C(n289), .Q(n288) );
  AOI220 U340 ( .A(n245), .B(id_data_jr[0]), .C(n243), .D(if_addr_b[0]), .Q(
        n151) );
  AOI220 U341 ( .A(n245), .B(id_data_jr[1]), .C(n243), .D(if_addr_b[1]), .Q(
        n152) );
  NOR41 U342 ( .A(if_con_b), .B(if_con_j[0]), .C(n242), .D(n149), .Q(n245) );
  AOI210 U343 ( .A(n310), .B(mem_data_pc4[5]), .C(n312), .Q(n311) );
  AOI210 U344 ( .A(n315), .B(mem_data_pc4[7]), .C(n317), .Q(n316) );
  AOI210 U345 ( .A(n321), .B(mem_data_pc4[9]), .C(n320), .Q(n322) );
  AOI210 U346 ( .A(n252), .B(mem_data_pc4[11]), .C(n254), .Q(n253) );
  AOI210 U347 ( .A(n257), .B(mem_data_pc4[13]), .C(n259), .Q(n258) );
  AOI210 U348 ( .A(n262), .B(mem_data_pc4[15]), .C(n264), .Q(n263) );
  AOI210 U349 ( .A(n267), .B(mem_data_pc4[17]), .C(n269), .Q(n268) );
  AOI210 U350 ( .A(n272), .B(mem_data_pc4[19]), .C(n274), .Q(n273) );
  AOI210 U351 ( .A(n277), .B(mem_data_pc4[21]), .C(n279), .Q(n278) );
  AOI210 U352 ( .A(n282), .B(mem_data_pc4[23]), .C(n284), .Q(n283) );
  OAI210 U353 ( .A(n294), .B(mem_data_pc4[28]), .C(n297), .Q(n295) );
  IMUX20 U354 ( .A(n309), .B(n308), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[4]) );
  INV3 U355 ( .A(n304), .Q(n307) );
  IMUX20 U356 ( .A(n299), .B(mem_data_pc4[2]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[2]) );
  IMUX20 U357 ( .A(n314), .B(n313), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[6]) );
  MUX21 U358 ( .A(data_address[1]), .B(u_mem_pc8[1]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[1]) );
  MUX21 U359 ( .A(data_address[5]), .B(n311), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[5]) );
  MUX21 U360 ( .A(data_address[0]), .B(u_mem_pc8[0]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[0]) );
  MUX21 U361 ( .A(data_address[7]), .B(n316), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[7]) );
  IMUX20 U362 ( .A(n319), .B(n318), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[8]) );
  MUX21 U363 ( .A(data_address[9]), .B(n322), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[9]) );
  IMUX20 U364 ( .A(n251), .B(n250), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[10]) );
  MUX21 U365 ( .A(data_address[11]), .B(n253), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[11]) );
  IMUX20 U366 ( .A(n256), .B(n255), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[12]) );
  MUX21 U367 ( .A(data_address[13]), .B(n258), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[13]) );
  IMUX20 U368 ( .A(n261), .B(n260), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[14]) );
  MUX21 U369 ( .A(data_address[15]), .B(n263), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[15]) );
  IMUX20 U370 ( .A(n266), .B(n265), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[16]) );
  MUX21 U371 ( .A(data_address[17]), .B(n268), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[17]) );
  IMUX20 U372 ( .A(n271), .B(n270), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[18]) );
  MUX21 U373 ( .A(data_address[19]), .B(n273), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[19]) );
  IMUX20 U374 ( .A(n276), .B(n275), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[20]) );
  MUX21 U375 ( .A(data_address[21]), .B(n278), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[21]) );
  MUX21 U376 ( .A(data_address[23]), .B(n283), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[23]) );
  OAI2111 U377 ( .A(n249), .B(n163), .C(n162), .D(n161), .Q(n134) );
  OAI2111 U378 ( .A(n249), .B(n172), .C(n171), .D(n170), .Q(n131) );
  OAI2111 U379 ( .A(n249), .B(n166), .C(n165), .D(n164), .Q(n133) );
  OAI2111 U380 ( .A(n249), .B(n169), .C(n168), .D(n167), .Q(n132) );
  OAI2111 U381 ( .A(n249), .B(n238), .C(n237), .D(n236), .Q(n109) );
  OAI2111 U382 ( .A(n249), .B(n178), .C(n177), .D(n176), .Q(n129) );
  OAI2111 U383 ( .A(n249), .B(n175), .C(n174), .D(n173), .Q(n130) );
  AOI211 U384 ( .A(n297), .B(mem_data_pc4[29]), .C(n300), .Q(n298) );
  NAND22 U385 ( .A(n300), .B(mem_data_pc4[30]), .Q(n303) );
  NOR21 U386 ( .A(n297), .B(mem_data_pc4[29]), .Q(n300) );
  NAND22 U387 ( .A(n294), .B(mem_data_pc4[28]), .Q(n297) );
  NAND22 U388 ( .A(n289), .B(mem_data_pc4[26]), .Q(n292) );
  NAND22 U389 ( .A(n284), .B(mem_data_pc4[24]), .Q(n287) );
  NAND22 U390 ( .A(n279), .B(mem_data_pc4[22]), .Q(n282) );
  NAND22 U391 ( .A(n274), .B(mem_data_pc4[20]), .Q(n277) );
  NAND22 U392 ( .A(n269), .B(mem_data_pc4[18]), .Q(n272) );
  NAND22 U393 ( .A(n264), .B(mem_data_pc4[16]), .Q(n267) );
  NAND22 U394 ( .A(n259), .B(mem_data_pc4[14]), .Q(n262) );
  NAND22 U395 ( .A(n254), .B(mem_data_pc4[12]), .Q(n257) );
  NAND22 U396 ( .A(n320), .B(mem_data_pc4[10]), .Q(n252) );
  NAND22 U397 ( .A(n317), .B(mem_data_pc4[8]), .Q(n321) );
  NAND22 U398 ( .A(n312), .B(mem_data_pc4[6]), .Q(n315) );
  NOR21 U399 ( .A(n310), .B(mem_data_pc4[5]), .Q(n312) );
  NAND31 U400 ( .A(mem_data_pc4[2]), .B(mem_data_pc4[3]), .C(mem_data_pc4[4]), 
        .Q(n310) );
  OAI2111 U401 ( .A(n249), .B(n184), .C(n183), .D(n182), .Q(n127) );
  OAI2111 U402 ( .A(n249), .B(n211), .C(n210), .D(n209), .Q(n118) );
  OAI2111 U403 ( .A(n249), .B(n196), .C(n195), .D(n194), .Q(n123) );
  OAI2111 U404 ( .A(n249), .B(n205), .C(n204), .D(n203), .Q(n120) );
  OAI2111 U405 ( .A(n249), .B(n199), .C(n198), .D(n197), .Q(n122) );
  OAI2111 U406 ( .A(n249), .B(n202), .C(n201), .D(n200), .Q(n121) );
  OAI2111 U407 ( .A(n249), .B(n193), .C(n192), .D(n191), .Q(n124) );
  OAI2111 U408 ( .A(n249), .B(n208), .C(n207), .D(n206), .Q(n119) );
  OAI2111 U409 ( .A(n249), .B(n190), .C(n189), .D(n188), .Q(n125) );
  OAI2111 U410 ( .A(n249), .B(n187), .C(n186), .D(n185), .Q(n126) );
  OAI2111 U411 ( .A(n249), .B(n241), .C(n240), .D(n239), .Q(n108) );
  OAI2111 U412 ( .A(n249), .B(n248), .C(n247), .D(n246), .Q(n107) );
  OAI2111 U413 ( .A(n249), .B(n181), .C(n180), .D(n179), .Q(n128) );
  OAI2111 U414 ( .A(n249), .B(n220), .C(n219), .D(n218), .Q(n115) );
  OAI2111 U415 ( .A(n249), .B(n232), .C(n231), .D(n230), .Q(n111) );
  OAI2111 U416 ( .A(n249), .B(n235), .C(n234), .D(n233), .Q(n110) );
  OAI2111 U417 ( .A(n249), .B(n217), .C(n216), .D(n215), .Q(n116) );
  OAI2111 U418 ( .A(n249), .B(n229), .C(n228), .D(n227), .Q(n112) );
  OAI2111 U419 ( .A(n249), .B(n223), .C(n222), .D(n221), .Q(n114) );
  OAI2111 U420 ( .A(n249), .B(n214), .C(n213), .D(n212), .Q(n117) );
  OAI2111 U421 ( .A(n249), .B(n226), .C(n225), .D(n224), .Q(n113) );
  NAND22 U422 ( .A(if_con_b), .B(if_con_ifstall), .Q(n150) );
  INV3 U423 ( .A(if_con_j[0]), .Q(n155) );
  INV3 U424 ( .A(if_con_j[1]), .Q(n149) );
  LOGIC0 U425 ( .Q(n146) );
  AOI220 U426 ( .A(if_addr_b[31]), .B(n243), .C(instruction_address[31]), .D(
        n242), .Q(n157) );
  NOR40 U427 ( .A(if_con_b), .B(if_con_j[1]), .C(n242), .D(n155), .Q(n244) );
  AOI220 U428 ( .A(if_addr_b[2]), .B(n243), .C(instruction_address[2]), .D(
        n242), .Q(n160) );
  AOI220 U429 ( .A(n245), .B(id_data_jr[2]), .C(n147), .D(if_addr_j[2]), .Q(
        n159) );
  AOI220 U430 ( .A(if_addr_b[3]), .B(n243), .C(instruction_address[3]), .D(
        n242), .Q(n162) );
  AOI220 U431 ( .A(n245), .B(id_data_jr[3]), .C(n147), .D(if_addr_j[3]), .Q(
        n161) );
  AOI220 U432 ( .A(if_addr_b[4]), .B(n243), .C(instruction_address[4]), .D(
        n242), .Q(n165) );
  AOI220 U433 ( .A(n245), .B(id_data_jr[4]), .C(n147), .D(if_addr_j[4]), .Q(
        n164) );
  AOI220 U434 ( .A(if_addr_b[5]), .B(n243), .C(instruction_address[5]), .D(
        n242), .Q(n168) );
  AOI220 U435 ( .A(n245), .B(id_data_jr[5]), .C(n147), .D(if_addr_j[5]), .Q(
        n167) );
  AOI220 U436 ( .A(if_addr_b[6]), .B(n243), .C(instruction_address[6]), .D(
        n242), .Q(n171) );
  AOI220 U437 ( .A(n245), .B(id_data_jr[6]), .C(n147), .D(if_addr_j[6]), .Q(
        n170) );
  AOI220 U438 ( .A(if_addr_b[7]), .B(n243), .C(instruction_address[7]), .D(
        n242), .Q(n174) );
  AOI220 U439 ( .A(n245), .B(id_data_jr[7]), .C(n147), .D(if_addr_j[7]), .Q(
        n173) );
  AOI220 U440 ( .A(if_addr_b[8]), .B(n243), .C(instruction_address[8]), .D(
        n242), .Q(n177) );
  AOI220 U441 ( .A(n245), .B(id_data_jr[8]), .C(n147), .D(if_addr_j[8]), .Q(
        n176) );
  AOI220 U442 ( .A(if_addr_b[9]), .B(n243), .C(instruction_address[9]), .D(
        n242), .Q(n180) );
  AOI220 U443 ( .A(if_addr_b[10]), .B(n243), .C(instruction_address[10]), .D(
        n242), .Q(n183) );
  AOI220 U444 ( .A(if_addr_b[11]), .B(n243), .C(instruction_address[11]), .D(
        n242), .Q(n186) );
  AOI220 U445 ( .A(if_addr_b[12]), .B(n243), .C(instruction_address[12]), .D(
        n242), .Q(n189) );
  AOI220 U446 ( .A(if_addr_b[13]), .B(n243), .C(instruction_address[13]), .D(
        n242), .Q(n192) );
  AOI220 U447 ( .A(if_addr_b[14]), .B(n243), .C(instruction_address[14]), .D(
        n242), .Q(n195) );
  AOI220 U448 ( .A(if_addr_b[15]), .B(n243), .C(instruction_address[15]), .D(
        n242), .Q(n198) );
  AOI220 U449 ( .A(if_addr_b[16]), .B(n243), .C(instruction_address[16]), .D(
        n242), .Q(n201) );
  AOI220 U450 ( .A(n148), .B(id_data_jr[16]), .C(n147), .D(if_addr_j[16]), .Q(
        n200) );
  AOI220 U451 ( .A(if_addr_b[17]), .B(n243), .C(instruction_address[17]), .D(
        n242), .Q(n204) );
  AOI220 U452 ( .A(if_addr_b[18]), .B(n243), .C(instruction_address[18]), .D(
        n242), .Q(n207) );
  AOI220 U453 ( .A(if_addr_b[19]), .B(n243), .C(instruction_address[19]), .D(
        n242), .Q(n210) );
  AOI220 U454 ( .A(if_addr_b[20]), .B(n243), .C(instruction_address[20]), .D(
        n242), .Q(n213) );
  AOI220 U455 ( .A(n148), .B(id_data_jr[20]), .C(n147), .D(if_addr_j[20]), .Q(
        n212) );
  AOI220 U456 ( .A(if_addr_b[21]), .B(n243), .C(instruction_address[21]), .D(
        n242), .Q(n216) );
  AOI220 U457 ( .A(if_addr_b[22]), .B(n243), .C(instruction_address[22]), .D(
        n242), .Q(n219) );
  AOI220 U458 ( .A(n148), .B(id_data_jr[22]), .C(n147), .D(if_addr_j[22]), .Q(
        n218) );
  AOI220 U459 ( .A(if_addr_b[23]), .B(n243), .C(instruction_address[23]), .D(
        n242), .Q(n222) );
  AOI220 U460 ( .A(n148), .B(id_data_jr[23]), .C(n147), .D(if_addr_j[23]), .Q(
        n221) );
  AOI220 U461 ( .A(if_addr_b[24]), .B(n243), .C(instruction_address[24]), .D(
        n242), .Q(n225) );
  AOI220 U462 ( .A(n148), .B(id_data_jr[24]), .C(n147), .D(if_addr_j[24]), .Q(
        n224) );
  AOI220 U463 ( .A(if_addr_b[25]), .B(n243), .C(instruction_address[25]), .D(
        n242), .Q(n228) );
  AOI220 U464 ( .A(n148), .B(id_data_jr[25]), .C(n147), .D(if_addr_j[25]), .Q(
        n227) );
  AOI220 U465 ( .A(if_addr_b[26]), .B(n243), .C(instruction_address[26]), .D(
        n242), .Q(n231) );
  AOI220 U466 ( .A(n148), .B(id_data_jr[26]), .C(n147), .D(if_addr_j[26]), .Q(
        n230) );
  AOI220 U467 ( .A(if_addr_b[27]), .B(n243), .C(instruction_address[27]), .D(
        n242), .Q(n234) );
  AOI220 U468 ( .A(if_addr_b[28]), .B(n243), .C(instruction_address[28]), .D(
        n242), .Q(n237) );
  AOI220 U469 ( .A(n245), .B(id_data_jr[28]), .C(n147), .D(if_addr_j[28]), .Q(
        n236) );
  AOI220 U470 ( .A(if_addr_b[29]), .B(n243), .C(instruction_address[29]), .D(
        n242), .Q(n240) );
  AOI220 U471 ( .A(if_addr_b[30]), .B(n243), .C(instruction_address[30]), .D(
        n242), .Q(n247) );
  OAI210 U472 ( .A(n320), .B(mem_data_pc4[10]), .C(n252), .Q(n250) );
  OAI210 U473 ( .A(n254), .B(mem_data_pc4[12]), .C(n257), .Q(n255) );
  OAI210 U474 ( .A(n259), .B(mem_data_pc4[14]), .C(n262), .Q(n260) );
  OAI210 U475 ( .A(n264), .B(mem_data_pc4[16]), .C(n267), .Q(n265) );
  OAI210 U476 ( .A(n269), .B(mem_data_pc4[18]), .C(n272), .Q(n270) );
  OAI210 U477 ( .A(n274), .B(mem_data_pc4[20]), .C(n277), .Q(n275) );
  OAI210 U478 ( .A(n279), .B(mem_data_pc4[22]), .C(n282), .Q(n280) );
  OAI210 U479 ( .A(n284), .B(mem_data_pc4[24]), .C(n287), .Q(n285) );
  OAI210 U480 ( .A(n289), .B(mem_data_pc4[26]), .C(n292), .Q(n290) );
  OAI210 U481 ( .A(mem_data_pc4[2]), .B(mem_data_pc4[3]), .C(mem_con_Malupc8), 
        .Q(n306) );
  OAI220 U482 ( .A(n307), .B(n306), .C(mem_con_Malupc8), .D(n305), .Q(
        u_mem_resmux_o_data_alu[3]) );
  OAI210 U483 ( .A(n312), .B(mem_data_pc4[6]), .C(n315), .Q(n313) );
  OAI210 U484 ( .A(n317), .B(mem_data_pc4[8]), .C(n321), .Q(n318) );
endmodule

