
module F_jumpmux ( i_addr_j, i_addr_jr, i_addr_pc4, i_con_jump, o_addr_jumpmux
 );
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [31:0] i_addr_pc4;
  input [1:0] i_con_jump;
  output [31:0] o_addr_jumpmux;
  wire   n3, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n23,
         n24, n45, n46, n63, n64, n65, n66, n67, n68, n1, n2, n5, n6, n19, n20,
         n21, n22, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  AOI221 U1 ( .A(i_addr_pc4[0]), .B(n6), .C(i_addr_jr[0]), .D(n1), .Q(n67) );
  AOI221 U2 ( .A(i_addr_pc4[1]), .B(n6), .C(i_addr_jr[1]), .D(n1), .Q(n45) );
  AOI221 U3 ( .A(i_addr_pc4[2]), .B(n6), .C(i_addr_jr[2]), .D(n1), .Q(n23) );
  AOI221 U4 ( .A(i_addr_pc4[4]), .B(n5), .C(i_addr_jr[4]), .D(n1), .Q(n15) );
  AOI221 U5 ( .A(i_addr_pc4[6]), .B(n5), .C(i_addr_jr[6]), .D(n1), .Q(n11) );
  AOI221 U6 ( .A(i_addr_pc4[8]), .B(n5), .C(i_addr_jr[8]), .D(n1), .Q(n7) );
  AOI221 U7 ( .A(i_addr_pc4[9]), .B(n5), .C(i_addr_jr[9]), .D(n1), .Q(n3) );
  AOI221 U8 ( .A(i_addr_pc4[10]), .B(n6), .C(i_addr_jr[10]), .D(n2), .Q(n65)
         );
  AOI221 U9 ( .A(i_addr_pc4[11]), .B(n6), .C(i_addr_jr[11]), .D(n1), .Q(n63)
         );
  AOI221 U10 ( .A(i_addr_j[12]), .B(n20), .C(i_addr_pc4[12]), .D(n76), .Q(n28)
         );
  AOI221 U11 ( .A(i_addr_j[16]), .B(n19), .C(i_addr_pc4[16]), .D(n6), .Q(n36)
         );
  AOI221 U12 ( .A(i_addr_j[17]), .B(n19), .C(i_addr_pc4[17]), .D(n6), .Q(n38)
         );
  AOI221 U13 ( .A(i_addr_j[18]), .B(n19), .C(i_addr_pc4[18]), .D(n6), .Q(n40)
         );
  AOI221 U14 ( .A(i_addr_j[19]), .B(n19), .C(i_addr_pc4[19]), .D(n6), .Q(n42)
         );
  AOI221 U15 ( .A(i_addr_j[20]), .B(n19), .C(i_addr_pc4[20]), .D(n6), .Q(n44)
         );
  AOI221 U16 ( .A(i_addr_j[21]), .B(n19), .C(i_addr_pc4[21]), .D(n6), .Q(n48)
         );
  AOI221 U17 ( .A(i_addr_j[23]), .B(n19), .C(i_addr_pc4[23]), .D(n6), .Q(n52)
         );
  AOI221 U18 ( .A(i_addr_j[24]), .B(n19), .C(i_addr_pc4[24]), .D(n6), .Q(n54)
         );
  AOI221 U19 ( .A(i_addr_j[25]), .B(n19), .C(i_addr_pc4[25]), .D(n5), .Q(n56)
         );
  AOI221 U20 ( .A(i_addr_j[26]), .B(n19), .C(i_addr_pc4[26]), .D(n5), .Q(n58)
         );
  AOI221 U21 ( .A(i_addr_j[27]), .B(n19), .C(i_addr_pc4[27]), .D(n5), .Q(n60)
         );
  AOI221 U22 ( .A(i_addr_j[28]), .B(n19), .C(i_addr_pc4[28]), .D(n5), .Q(n62)
         );
  BUF2 U23 ( .A(n77), .Q(n19) );
  BUF2 U24 ( .A(n76), .Q(n5) );
  BUF2 U25 ( .A(n75), .Q(n1) );
  BUF2 U26 ( .A(n75), .Q(n2) );
  BUF2 U27 ( .A(n76), .Q(n6) );
  BUF2 U28 ( .A(n77), .Q(n20) );
  INV3 U29 ( .A(n26), .Q(n75) );
  NAND22 U30 ( .A(n67), .B(n68), .Q(o_addr_jumpmux[0]) );
  NAND22 U31 ( .A(i_addr_j[0]), .B(n20), .Q(n68) );
  NAND22 U32 ( .A(n45), .B(n46), .Q(o_addr_jumpmux[1]) );
  NAND22 U33 ( .A(i_addr_j[1]), .B(n77), .Q(n46) );
  NAND22 U34 ( .A(n23), .B(n24), .Q(o_addr_jumpmux[2]) );
  NAND22 U35 ( .A(i_addr_j[2]), .B(n20), .Q(n24) );
  NAND22 U36 ( .A(n15), .B(n16), .Q(o_addr_jumpmux[4]) );
  NAND22 U37 ( .A(i_addr_j[4]), .B(n20), .Q(n16) );
  NAND22 U38 ( .A(n11), .B(n12), .Q(o_addr_jumpmux[6]) );
  NAND22 U39 ( .A(i_addr_j[6]), .B(n20), .Q(n12) );
  NAND22 U40 ( .A(n7), .B(n8), .Q(o_addr_jumpmux[8]) );
  NAND22 U41 ( .A(i_addr_j[8]), .B(n20), .Q(n8) );
  NAND22 U42 ( .A(n3), .B(n4), .Q(o_addr_jumpmux[9]) );
  NAND22 U43 ( .A(i_addr_j[9]), .B(n20), .Q(n4) );
  NAND22 U44 ( .A(n65), .B(n66), .Q(o_addr_jumpmux[10]) );
  NAND22 U45 ( .A(i_addr_j[10]), .B(n20), .Q(n66) );
  NAND22 U46 ( .A(n63), .B(n64), .Q(o_addr_jumpmux[11]) );
  NAND22 U47 ( .A(i_addr_j[11]), .B(n20), .Q(n64) );
  NAND22 U48 ( .A(n17), .B(n18), .Q(o_addr_jumpmux[3]) );
  NAND22 U49 ( .A(i_addr_j[3]), .B(n20), .Q(n18) );
  AOI221 U50 ( .A(i_addr_pc4[3]), .B(n6), .C(i_addr_jr[3]), .D(n1), .Q(n17) );
  NAND22 U51 ( .A(n13), .B(n14), .Q(o_addr_jumpmux[5]) );
  NAND22 U52 ( .A(i_addr_j[5]), .B(n20), .Q(n14) );
  AOI221 U53 ( .A(i_addr_pc4[5]), .B(n5), .C(i_addr_jr[5]), .D(n1), .Q(n13) );
  NAND22 U54 ( .A(n9), .B(n10), .Q(o_addr_jumpmux[7]) );
  NAND22 U55 ( .A(i_addr_j[7]), .B(n20), .Q(n10) );
  AOI221 U56 ( .A(i_addr_pc4[7]), .B(n5), .C(i_addr_jr[7]), .D(n1), .Q(n9) );
  AOI221 U57 ( .A(i_addr_j[13]), .B(n20), .C(i_addr_pc4[13]), .D(n76), .Q(n30)
         );
  AOI221 U58 ( .A(i_addr_j[14]), .B(n19), .C(i_addr_pc4[14]), .D(n6), .Q(n32)
         );
  AOI221 U59 ( .A(i_addr_j[15]), .B(n19), .C(i_addr_pc4[15]), .D(n5), .Q(n34)
         );
  AOI221 U60 ( .A(i_addr_j[22]), .B(n19), .C(i_addr_pc4[22]), .D(n6), .Q(n50)
         );
  AOI221 U61 ( .A(i_addr_j[29]), .B(n19), .C(i_addr_pc4[29]), .D(n5), .Q(n70)
         );
  AOI221 U62 ( .A(i_addr_j[30]), .B(n19), .C(i_addr_pc4[30]), .D(n5), .Q(n72)
         );
  AOI221 U63 ( .A(i_addr_j[31]), .B(n20), .C(i_addr_pc4[31]), .D(n5), .Q(n74)
         );
  CLKIN3 U64 ( .A(i_con_jump[1]), .Q(n21) );
  NAND22 U65 ( .A(i_con_jump[0]), .B(n21), .Q(n22) );
  CLKIN3 U66 ( .A(n22), .Q(n77) );
  XNR21 U67 ( .A(i_con_jump[0]), .B(i_con_jump[1]), .Q(n76) );
  CLKIN3 U68 ( .A(i_con_jump[0]), .Q(n25) );
  NAND22 U69 ( .A(i_con_jump[1]), .B(n25), .Q(n26) );
  NAND22 U70 ( .A(i_addr_jr[12]), .B(n2), .Q(n27) );
  NAND22 U71 ( .A(n28), .B(n27), .Q(o_addr_jumpmux[12]) );
  NAND22 U72 ( .A(i_addr_jr[13]), .B(n75), .Q(n29) );
  NAND22 U73 ( .A(n30), .B(n29), .Q(o_addr_jumpmux[13]) );
  NAND22 U74 ( .A(i_addr_jr[14]), .B(n2), .Q(n31) );
  NAND22 U75 ( .A(n32), .B(n31), .Q(o_addr_jumpmux[14]) );
  NAND22 U76 ( .A(i_addr_jr[15]), .B(n75), .Q(n33) );
  NAND22 U77 ( .A(n34), .B(n33), .Q(o_addr_jumpmux[15]) );
  NAND22 U78 ( .A(i_addr_jr[16]), .B(n2), .Q(n35) );
  NAND22 U79 ( .A(n36), .B(n35), .Q(o_addr_jumpmux[16]) );
  NAND22 U80 ( .A(i_addr_jr[17]), .B(n75), .Q(n37) );
  NAND22 U81 ( .A(n38), .B(n37), .Q(o_addr_jumpmux[17]) );
  NAND22 U82 ( .A(i_addr_jr[18]), .B(n2), .Q(n39) );
  NAND22 U83 ( .A(n40), .B(n39), .Q(o_addr_jumpmux[18]) );
  NAND22 U84 ( .A(i_addr_jr[19]), .B(n75), .Q(n41) );
  NAND22 U85 ( .A(n42), .B(n41), .Q(o_addr_jumpmux[19]) );
  NAND22 U86 ( .A(i_addr_jr[20]), .B(n2), .Q(n43) );
  NAND22 U87 ( .A(n44), .B(n43), .Q(o_addr_jumpmux[20]) );
  NAND22 U88 ( .A(i_addr_jr[21]), .B(n75), .Q(n47) );
  NAND22 U89 ( .A(n48), .B(n47), .Q(o_addr_jumpmux[21]) );
  NAND22 U90 ( .A(i_addr_jr[22]), .B(n2), .Q(n49) );
  NAND22 U91 ( .A(n50), .B(n49), .Q(o_addr_jumpmux[22]) );
  NAND22 U92 ( .A(i_addr_jr[23]), .B(n75), .Q(n51) );
  NAND22 U93 ( .A(n52), .B(n51), .Q(o_addr_jumpmux[23]) );
  NAND22 U94 ( .A(i_addr_jr[24]), .B(n2), .Q(n53) );
  NAND22 U95 ( .A(n54), .B(n53), .Q(o_addr_jumpmux[24]) );
  NAND22 U96 ( .A(i_addr_jr[25]), .B(n75), .Q(n55) );
  NAND22 U97 ( .A(n56), .B(n55), .Q(o_addr_jumpmux[25]) );
  NAND22 U98 ( .A(i_addr_jr[26]), .B(n2), .Q(n57) );
  NAND22 U99 ( .A(n58), .B(n57), .Q(o_addr_jumpmux[26]) );
  NAND22 U100 ( .A(i_addr_jr[27]), .B(n1), .Q(n59) );
  NAND22 U101 ( .A(n60), .B(n59), .Q(o_addr_jumpmux[27]) );
  NAND22 U102 ( .A(i_addr_jr[28]), .B(n2), .Q(n61) );
  NAND22 U103 ( .A(n62), .B(n61), .Q(o_addr_jumpmux[28]) );
  NAND22 U104 ( .A(i_addr_jr[29]), .B(n1), .Q(n69) );
  NAND22 U105 ( .A(n70), .B(n69), .Q(o_addr_jumpmux[29]) );
  NAND22 U106 ( .A(i_addr_jr[30]), .B(n2), .Q(n71) );
  NAND22 U107 ( .A(n72), .B(n71), .Q(o_addr_jumpmux[30]) );
  NAND22 U108 ( .A(i_addr_jr[31]), .B(n75), .Q(n73) );
  NAND22 U109 ( .A(n74), .B(n73), .Q(o_addr_jumpmux[31]) );
endmodule


module F_branchmux ( i_addr_jumpmux, i_addr_b, i_con_ifbranch, o_addr_nextpc
 );
  input [31:0] i_addr_jumpmux;
  input [31:0] i_addr_b;
  output [31:0] o_addr_nextpc;
  input i_con_ifbranch;
  wire   n1, n2;

  MUX22 U1 ( .A(i_addr_jumpmux[31]), .B(i_addr_b[31]), .S(n2), .Q(
        o_addr_nextpc[31]) );
  BUF15 U2 ( .A(i_con_ifbranch), .Q(n1) );
  MUX22 U3 ( .A(i_addr_jumpmux[2]), .B(i_addr_b[2]), .S(n1), .Q(
        o_addr_nextpc[2]) );
  MUX22 U4 ( .A(i_addr_jumpmux[4]), .B(i_addr_b[4]), .S(n2), .Q(
        o_addr_nextpc[4]) );
  MUX22 U5 ( .A(i_addr_jumpmux[6]), .B(i_addr_b[6]), .S(n1), .Q(
        o_addr_nextpc[6]) );
  MUX22 U6 ( .A(i_addr_jumpmux[8]), .B(i_addr_b[8]), .S(n2), .Q(
        o_addr_nextpc[8]) );
  MUX22 U7 ( .A(i_addr_jumpmux[9]), .B(i_addr_b[9]), .S(n1), .Q(
        o_addr_nextpc[9]) );
  MUX22 U8 ( .A(i_addr_jumpmux[10]), .B(i_addr_b[10]), .S(n2), .Q(
        o_addr_nextpc[10]) );
  MUX22 U9 ( .A(i_addr_jumpmux[11]), .B(i_addr_b[11]), .S(n1), .Q(
        o_addr_nextpc[11]) );
  MUX22 U10 ( .A(i_addr_jumpmux[12]), .B(i_addr_b[12]), .S(n2), .Q(
        o_addr_nextpc[12]) );
  MUX22 U11 ( .A(i_addr_jumpmux[16]), .B(i_addr_b[16]), .S(n1), .Q(
        o_addr_nextpc[16]) );
  MUX22 U12 ( .A(i_addr_jumpmux[17]), .B(i_addr_b[17]), .S(n2), .Q(
        o_addr_nextpc[17]) );
  MUX22 U13 ( .A(i_addr_jumpmux[18]), .B(i_addr_b[18]), .S(n1), .Q(
        o_addr_nextpc[18]) );
  MUX22 U14 ( .A(i_addr_jumpmux[19]), .B(i_addr_b[19]), .S(n2), .Q(
        o_addr_nextpc[19]) );
  MUX22 U15 ( .A(i_addr_jumpmux[20]), .B(i_addr_b[20]), .S(n1), .Q(
        o_addr_nextpc[20]) );
  MUX22 U16 ( .A(i_addr_jumpmux[21]), .B(i_addr_b[21]), .S(n2), .Q(
        o_addr_nextpc[21]) );
  MUX22 U17 ( .A(i_addr_jumpmux[23]), .B(i_addr_b[23]), .S(n1), .Q(
        o_addr_nextpc[23]) );
  MUX22 U18 ( .A(i_addr_jumpmux[24]), .B(i_addr_b[24]), .S(n2), .Q(
        o_addr_nextpc[24]) );
  MUX22 U19 ( .A(i_addr_jumpmux[25]), .B(i_addr_b[25]), .S(n1), .Q(
        o_addr_nextpc[25]) );
  MUX22 U20 ( .A(i_addr_jumpmux[26]), .B(i_addr_b[26]), .S(n2), .Q(
        o_addr_nextpc[26]) );
  MUX22 U21 ( .A(i_addr_jumpmux[27]), .B(i_addr_b[27]), .S(n1), .Q(
        o_addr_nextpc[27]) );
  MUX22 U22 ( .A(i_addr_jumpmux[28]), .B(i_addr_b[28]), .S(n2), .Q(
        o_addr_nextpc[28]) );
  MUX22 U23 ( .A(i_addr_jumpmux[5]), .B(i_addr_b[5]), .S(n1), .Q(
        o_addr_nextpc[5]) );
  MUX22 U24 ( .A(i_addr_jumpmux[7]), .B(i_addr_b[7]), .S(n2), .Q(
        o_addr_nextpc[7]) );
  MUX22 U25 ( .A(i_addr_jumpmux[13]), .B(i_addr_b[13]), .S(n1), .Q(
        o_addr_nextpc[13]) );
  MUX22 U26 ( .A(i_addr_jumpmux[14]), .B(i_addr_b[14]), .S(n2), .Q(
        o_addr_nextpc[14]) );
  MUX22 U27 ( .A(i_addr_jumpmux[15]), .B(i_addr_b[15]), .S(n1), .Q(
        o_addr_nextpc[15]) );
  MUX22 U28 ( .A(i_addr_jumpmux[22]), .B(i_addr_b[22]), .S(n2), .Q(
        o_addr_nextpc[22]) );
  MUX22 U29 ( .A(i_addr_jumpmux[29]), .B(i_addr_b[29]), .S(n1), .Q(
        o_addr_nextpc[29]) );
  MUX22 U30 ( .A(i_addr_jumpmux[30]), .B(i_addr_b[30]), .S(n2), .Q(
        o_addr_nextpc[30]) );
  BUF15 U31 ( .A(i_con_ifbranch), .Q(n2) );
  MUX22 U32 ( .A(i_addr_jumpmux[0]), .B(i_addr_b[0]), .S(n1), .Q(
        o_addr_nextpc[0]) );
  MUX22 U33 ( .A(i_addr_jumpmux[1]), .B(i_addr_b[1]), .S(n1), .Q(
        o_addr_nextpc[1]) );
  MUX22 U34 ( .A(i_addr_jumpmux[3]), .B(i_addr_b[3]), .S(n2), .Q(
        o_addr_nextpc[3]) );
endmodule


module F_pc ( i_clk, i_rst_n, i_con_stall, i_addr_next_pc, o_addr_pc );
  input [31:0] i_addr_next_pc;
  output [31:0] o_addr_pc;
  input i_clk, i_rst_n, i_con_stall;


  DFEC3 program_counter_reg_25_ ( .D(i_addr_next_pc[25]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[25]) );
  DFEC3 program_counter_reg_24_ ( .D(i_addr_next_pc[24]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[24]) );
  DFEC3 program_counter_reg_23_ ( .D(i_addr_next_pc[23]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[23]) );
  DFEC3 program_counter_reg_31_ ( .D(i_addr_next_pc[31]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[31]) );
  DFEC3 program_counter_reg_30_ ( .D(i_addr_next_pc[30]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[30]) );
  DFEC3 program_counter_reg_27_ ( .D(i_addr_next_pc[27]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[27]) );
  DFEC3 program_counter_reg_29_ ( .D(i_addr_next_pc[29]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[29]) );
  DFEC3 program_counter_reg_28_ ( .D(i_addr_next_pc[28]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[28]) );
  DFEC3 program_counter_reg_22_ ( .D(i_addr_next_pc[22]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[22]) );
  DFEC3 program_counter_reg_21_ ( .D(i_addr_next_pc[21]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[21]) );
  DFEC3 program_counter_reg_18_ ( .D(i_addr_next_pc[18]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[18]) );
  DFEC3 program_counter_reg_17_ ( .D(i_addr_next_pc[17]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[17]) );
  DFEC3 program_counter_reg_2_ ( .D(i_addr_next_pc[2]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[2]) );
  DFEC3 program_counter_reg_15_ ( .D(i_addr_next_pc[15]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[15]) );
  DFEC3 program_counter_reg_19_ ( .D(i_addr_next_pc[19]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[19]) );
  DFEC3 program_counter_reg_9_ ( .D(i_addr_next_pc[9]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[9]) );
  DFEC3 program_counter_reg_7_ ( .D(i_addr_next_pc[7]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[7]) );
  DFEC3 program_counter_reg_5_ ( .D(i_addr_next_pc[5]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[5]) );
  DFEC3 program_counter_reg_10_ ( .D(i_addr_next_pc[10]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[10]) );
  DFEC3 program_counter_reg_14_ ( .D(i_addr_next_pc[14]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[14]) );
  DFEC3 program_counter_reg_6_ ( .D(i_addr_next_pc[6]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[6]) );
  DFEC3 program_counter_reg_11_ ( .D(i_addr_next_pc[11]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[11]) );
  DFEC3 program_counter_reg_8_ ( .D(i_addr_next_pc[8]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[8]) );
  DFEC3 program_counter_reg_12_ ( .D(i_addr_next_pc[12]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[12]) );
  DFEC3 program_counter_reg_16_ ( .D(i_addr_next_pc[16]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[16]) );
  DFEC3 program_counter_reg_4_ ( .D(i_addr_next_pc[4]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[4]) );
  DFEC3 program_counter_reg_20_ ( .D(i_addr_next_pc[20]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[20]) );
  DFEC3 program_counter_reg_3_ ( .D(i_addr_next_pc[3]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[3]) );
  DFEC3 program_counter_reg_1_ ( .D(i_addr_next_pc[1]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[1]) );
  DFEC3 program_counter_reg_0_ ( .D(i_addr_next_pc[0]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[0]) );
  DFEC3 program_counter_reg_26_ ( .D(i_addr_next_pc[26]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[26]) );
  DFEC3 program_counter_reg_13_ ( .D(i_addr_next_pc[13]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[13]) );
endmodule


module F_add4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  NAND22 U2 ( .A(n61), .B(n3), .Q(n70) );
  NAND22 U3 ( .A(n67), .B(A[14]), .Q(n66) );
  NAND22 U4 ( .A(n39), .B(n36), .Q(n49) );
  NAND22 U5 ( .A(n46), .B(A[21]), .Q(n47) );
  NAND22 U6 ( .A(n27), .B(n36), .Q(n37) );
  NAND22 U7 ( .A(n33), .B(A[25]), .Q(n34) );
  INV3 U8 ( .A(n58), .Q(n36) );
  NAND41 U9 ( .A(n59), .B(n60), .C(n61), .D(n62), .Q(n58) );
  NOR21 U10 ( .A(n64), .B(n65), .Q(n59) );
  NOR21 U11 ( .A(n63), .B(SUM[2]), .Q(n62) );
  XNR21 U12 ( .A(n68), .B(n64), .Q(SUM[13]) );
  XNR21 U13 ( .A(n56), .B(n51), .Q(SUM[17]) );
  XNR21 U14 ( .A(A[22]), .B(n47), .Q(SUM[22]) );
  XNR21 U15 ( .A(A[26]), .B(n34), .Q(SUM[26]) );
  XOR21 U16 ( .A(A[14]), .B(n67), .Q(SUM[14]) );
  XOR21 U17 ( .A(A[25]), .B(n33), .Q(SUM[25]) );
  XNR21 U18 ( .A(n55), .B(n52), .Q(SUM[18]) );
  XNR21 U19 ( .A(n74), .B(n75), .Q(SUM[10]) );
  NOR21 U20 ( .A(n64), .B(n69), .Q(n67) );
  NOR21 U21 ( .A(n51), .B(n57), .Q(n55) );
  NOR21 U22 ( .A(n8), .B(n10), .Q(n6) );
  NOR21 U23 ( .A(n76), .B(n2), .Q(n74) );
  INV3 U24 ( .A(n21), .Q(n24) );
  XNR21 U25 ( .A(n46), .B(n42), .Q(SUM[21]) );
  XNR21 U26 ( .A(n6), .B(n7), .Q(SUM[6]) );
  XNR21 U27 ( .A(n9), .B(n8), .Q(SUM[5]) );
  XNR21 U28 ( .A(n1), .B(n2), .Q(SUM[9]) );
  NOR31 U29 ( .A(n52), .B(n50), .C(n51), .Q(n39) );
  NAND22 U30 ( .A(A[19]), .B(A[16]), .Q(n50) );
  NAND31 U31 ( .A(A[15]), .B(A[12]), .C(A[3]), .Q(n63) );
  XNR21 U32 ( .A(A[20]), .B(n49), .Q(SUM[20]) );
  XNR21 U33 ( .A(A[24]), .B(n37), .Q(SUM[24]) );
  XNR21 U34 ( .A(A[16]), .B(n58), .Q(SUM[16]) );
  XNR21 U35 ( .A(A[28]), .B(n24), .Q(SUM[28]) );
  XOR21 U36 ( .A(A[29]), .B(n23), .Q(SUM[29]) );
  NOR21 U37 ( .A(n24), .B(n15), .Q(n23) );
  XNR21 U38 ( .A(A[15]), .B(n66), .Q(SUM[15]) );
  XOR21 U39 ( .A(n53), .B(n54), .Q(SUM[19]) );
  INV3 U40 ( .A(A[19]), .Q(n53) );
  NAND22 U41 ( .A(n55), .B(A[18]), .Q(n54) );
  XOR21 U42 ( .A(n44), .B(n45), .Q(SUM[23]) );
  INV3 U43 ( .A(A[23]), .Q(n44) );
  NAND31 U44 ( .A(A[21]), .B(n46), .C(A[22]), .Q(n45) );
  XOR21 U45 ( .A(n31), .B(n32), .Q(SUM[27]) );
  INV3 U46 ( .A(A[27]), .Q(n31) );
  NAND31 U47 ( .A(A[25]), .B(n33), .C(A[26]), .Q(n32) );
  XOR21 U48 ( .A(n18), .B(n19), .Q(SUM[30]) );
  INV3 U49 ( .A(A[30]), .Q(n18) );
  NAND22 U50 ( .A(n20), .B(n21), .Q(n19) );
  NOR21 U51 ( .A(n15), .B(n17), .Q(n20) );
  XOR21 U52 ( .A(n72), .B(n73), .Q(SUM[11]) );
  INV3 U53 ( .A(A[11]), .Q(n72) );
  NAND22 U54 ( .A(n74), .B(A[10]), .Q(n73) );
  XNR21 U55 ( .A(A[31]), .B(n13), .Q(SUM[31]) );
  INV3 U56 ( .A(n14), .Q(n13) );
  NOR31 U57 ( .A(n16), .B(n24), .C(n15), .Q(n14) );
  NAND22 U58 ( .A(A[30]), .B(A[29]), .Q(n16) );
  INV3 U59 ( .A(n77), .Q(n3) );
  NAND22 U60 ( .A(n78), .B(n60), .Q(n77) );
  NOR21 U61 ( .A(n81), .B(SUM[2]), .Q(n78) );
  INV3 U62 ( .A(A[3]), .Q(n81) );
  NOR21 U63 ( .A(n58), .B(n25), .Q(n21) );
  NAND22 U64 ( .A(n26), .B(n27), .Q(n25) );
  NOR31 U65 ( .A(n30), .B(n28), .C(n29), .Q(n26) );
  NAND22 U66 ( .A(A[27]), .B(A[24]), .Q(n28) );
  INV3 U67 ( .A(A[17]), .Q(n51) );
  NOR21 U68 ( .A(n79), .B(n80), .Q(n60) );
  NAND22 U69 ( .A(A[5]), .B(A[6]), .Q(n79) );
  NAND22 U70 ( .A(A[7]), .B(A[4]), .Q(n80) );
  INV3 U71 ( .A(A[18]), .Q(n52) );
  INV3 U72 ( .A(A[21]), .Q(n42) );
  INV3 U73 ( .A(A[22]), .Q(n43) );
  INV3 U74 ( .A(A[2]), .Q(SUM[2]) );
  INV3 U75 ( .A(n35), .Q(n33) );
  NAND31 U76 ( .A(n27), .B(n36), .C(A[24]), .Q(n35) );
  INV3 U77 ( .A(n48), .Q(n46) );
  NAND31 U78 ( .A(n39), .B(A[20]), .C(n36), .Q(n48) );
  INV3 U79 ( .A(n38), .Q(n27) );
  NAND22 U80 ( .A(n39), .B(n40), .Q(n38) );
  NOR31 U81 ( .A(n41), .B(n42), .C(n43), .Q(n40) );
  NAND22 U82 ( .A(A[23]), .B(A[20]), .Q(n41) );
  XOR21 U83 ( .A(n4), .B(n5), .Q(SUM[7]) );
  INV3 U84 ( .A(A[7]), .Q(n4) );
  NAND22 U85 ( .A(n6), .B(A[6]), .Q(n5) );
  INV3 U86 ( .A(n71), .Q(n61) );
  NAND41 U87 ( .A(A[11]), .B(A[8]), .C(A[10]), .D(A[9]), .Q(n71) );
  INV3 U88 ( .A(n12), .Q(n11) );
  NAND22 U89 ( .A(A[3]), .B(A[2]), .Q(n12) );
  INV3 U90 ( .A(n10), .Q(n9) );
  NAND22 U91 ( .A(A[4]), .B(n11), .Q(n10) );
  INV3 U92 ( .A(n57), .Q(n56) );
  NAND22 U93 ( .A(A[16]), .B(n36), .Q(n57) );
  INV3 U94 ( .A(n76), .Q(n1) );
  NAND22 U95 ( .A(A[8]), .B(n3), .Q(n76) );
  INV3 U96 ( .A(n69), .Q(n68) );
  NAND31 U97 ( .A(n61), .B(A[12]), .C(n3), .Q(n69) );
  INV3 U98 ( .A(A[13]), .Q(n64) );
  INV3 U99 ( .A(A[14]), .Q(n65) );
  XNR21 U100 ( .A(A[12]), .B(n70), .Q(SUM[12]) );
  XOR21 U101 ( .A(n3), .B(A[8]), .Q(SUM[8]) );
  XOR21 U102 ( .A(n11), .B(A[4]), .Q(SUM[4]) );
  XOR21 U103 ( .A(A[3]), .B(A[2]), .Q(SUM[3]) );
  INV3 U104 ( .A(A[28]), .Q(n15) );
  INV3 U105 ( .A(A[26]), .Q(n30) );
  INV3 U106 ( .A(A[5]), .Q(n8) );
  INV3 U107 ( .A(A[29]), .Q(n17) );
  INV3 U108 ( .A(A[9]), .Q(n2) );
  INV3 U109 ( .A(A[6]), .Q(n7) );
  INV3 U110 ( .A(A[10]), .Q(n75) );
  INV3 U111 ( .A(A[25]), .Q(n29) );
endmodule


module F_add4 ( i_addr_pc, o_addr_pcadd4 );
  input [31:0] i_addr_pc;
  output [31:0] o_addr_pcadd4;
  wire   n2, n1;

  F_add4_DW01_add_1 add_5 ( .A(i_addr_pc), .B({n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n2, n1, n1}), .CI(n1), .SUM(o_addr_pcadd4) );
  LOGIC0 U3 ( .Q(n1) );
  LOGIC1 U4 ( .Q(n2) );
endmodule


module fetch ( i_clk, i_nrst, i_addr_b, i_addr_j, i_addr_jr, i_con_b, i_con_j, 
        i_data_instr, i_con_ifstall, o_addr_pc, o_addr_pc4, o_data_instr );
  input [31:0] i_addr_b;
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [1:0] i_con_j;
  input [31:0] i_data_instr;
  output [31:0] o_addr_pc;
  output [31:0] o_addr_pc4;
  output [31:0] o_data_instr;
  input i_clk, i_nrst, i_con_b, i_con_ifstall;

  wire   [31:0] jmux_i_addr_pc4;
  wire   [31:0] bmux_i_addr_jumpmux;
  wire   [31:0] pc_i_addr_next_pc;

  DFC3 pipe_instr_reg_31_ ( .D(i_data_instr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[31]) );
  DFC3 pipe_instr_reg_30_ ( .D(i_data_instr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[30]) );
  DFC3 pipe_instr_reg_29_ ( .D(i_data_instr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[29]) );
  DFC3 pipe_instr_reg_28_ ( .D(i_data_instr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[28]) );
  DFC3 pipe_instr_reg_27_ ( .D(i_data_instr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[27]) );
  DFC3 pipe_instr_reg_26_ ( .D(i_data_instr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[26]) );
  DFC3 pipe_instr_reg_25_ ( .D(i_data_instr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[25]) );
  DFC3 pipe_instr_reg_24_ ( .D(i_data_instr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[24]) );
  DFC3 pipe_instr_reg_23_ ( .D(i_data_instr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[23]) );
  DFC3 pipe_instr_reg_22_ ( .D(i_data_instr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[22]) );
  DFC3 pipe_instr_reg_21_ ( .D(i_data_instr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[21]) );
  DFC3 pipe_instr_reg_20_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[20]) );
  DFC3 pipe_instr_reg_19_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[19]) );
  DFC3 pipe_instr_reg_18_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[18]) );
  DFC3 pipe_instr_reg_17_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[17]) );
  DFC3 pipe_instr_reg_16_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[16]) );
  DFC3 pipe_instr_reg_15_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[15]) );
  DFC3 pipe_instr_reg_14_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[14]) );
  DFC3 pipe_instr_reg_13_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[13]) );
  DFC3 pipe_instr_reg_12_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[12]) );
  DFC3 pipe_instr_reg_11_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[11]) );
  DFC3 pipe_instr_reg_10_ ( .D(i_data_instr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[10]) );
  DFC3 pipe_instr_reg_9_ ( .D(i_data_instr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[9]) );
  DFC3 pipe_instr_reg_8_ ( .D(i_data_instr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[8]) );
  DFC3 pipe_instr_reg_7_ ( .D(i_data_instr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[7]) );
  DFC3 pipe_instr_reg_6_ ( .D(i_data_instr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[6]) );
  DFC3 pipe_instr_reg_5_ ( .D(i_data_instr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[5]) );
  DFC3 pipe_instr_reg_4_ ( .D(i_data_instr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[4]) );
  DFC3 pipe_instr_reg_3_ ( .D(i_data_instr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[3]) );
  DFC3 pipe_instr_reg_2_ ( .D(i_data_instr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[2]) );
  DFC3 pipe_instr_reg_1_ ( .D(i_data_instr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[1]) );
  DFC3 pipe_instr_reg_0_ ( .D(i_data_instr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(jmux_i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(jmux_i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(jmux_i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(jmux_i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(jmux_i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(jmux_i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(jmux_i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(jmux_i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(jmux_i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(jmux_i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(jmux_i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(jmux_i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(jmux_i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(jmux_i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(jmux_i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(jmux_i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(jmux_i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(jmux_i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(jmux_i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(jmux_i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(jmux_i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(jmux_i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(jmux_i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(jmux_i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(jmux_i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(jmux_i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(jmux_i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(jmux_i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(jmux_i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(jmux_i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(jmux_i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(jmux_i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  F_jumpmux u_jumpmux ( .i_addr_j(i_addr_j), .i_addr_jr(i_addr_jr), 
        .i_addr_pc4(jmux_i_addr_pc4), .i_con_jump(i_con_j), .o_addr_jumpmux(
        bmux_i_addr_jumpmux) );
  F_branchmux u_branchmux ( .i_addr_jumpmux(bmux_i_addr_jumpmux), .i_addr_b(
        i_addr_b), .i_con_ifbranch(i_con_b), .o_addr_nextpc(pc_i_addr_next_pc)
         );
  F_pc u_pc ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_con_stall(i_con_ifstall), 
        .i_addr_next_pc(pc_i_addr_next_pc), .o_addr_pc(o_addr_pc) );
  F_add4 u_add4 ( .i_addr_pc(o_addr_pc), .o_addr_pcadd4(jmux_i_addr_pc4) );
endmodule


module D_control ( o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite, 
        o_con_alusrc, o_con_regwrite, o_con_ifsign, o_con_aluop, i_con_instru
 );
  output [5:0] o_con_aluop;
  input [5:0] i_con_instru;
  output o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite,
         o_con_alusrc, o_con_regwrite, o_con_ifsign;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n1, n2, n3, n5, n6, n7, n8, n9, n10;

  OAI212 U2 ( .A(i_con_instru[3]), .B(n11), .C(n12), .Q(o_con_regwrite) );
  OAI212 U3 ( .A(n5), .B(n13), .C(n3), .Q(n12) );
  OAI222 U6 ( .A(i_con_instru[3]), .B(n15), .C(i_con_instru[4]), .D(n17), .Q(
        o_con_memread) );
  OAI212 U23 ( .A(i_con_instru[5]), .B(n20), .C(n14), .Q(o_con_aluop[1]) );
  NAND22 U4 ( .A(n9), .B(n13), .Q(n11) );
  NAND31 U5 ( .A(n24), .B(n3), .C(n13), .Q(n14) );
  AOI211 U7 ( .A(n5), .B(n8), .C(o_con_memwrite), .Q(n18) );
  INV3 U8 ( .A(n20), .Q(n5) );
  INV3 U9 ( .A(n24), .Q(n9) );
  INV3 U10 ( .A(n21), .Q(n2) );
  NAND22 U11 ( .A(n20), .B(n15), .Q(o_con_alusrc) );
  NAND22 U12 ( .A(n15), .B(n16), .Q(o_con_memtoreg) );
  NOR21 U13 ( .A(n11), .B(n21), .Q(o_con_aluop[5]) );
  INV3 U14 ( .A(n16), .Q(o_con_memwrite) );
  NOR31 U15 ( .A(i_con_instru[2]), .B(i_con_instru[4]), .C(n27), .Q(n13) );
  XNR21 U16 ( .A(i_con_instru[1]), .B(n10), .Q(n27) );
  OAI2111 U17 ( .A(n9), .B(n18), .C(n19), .D(n15), .Q(o_con_ifsign) );
  NAND31 U18 ( .A(n9), .B(n5), .C(i_con_instru[2]), .Q(n19) );
  NAND22 U19 ( .A(i_con_instru[5]), .B(n7), .Q(n15) );
  INV3 U20 ( .A(n11), .Q(n7) );
  INV3 U21 ( .A(i_con_instru[0]), .Q(n10) );
  NAND22 U22 ( .A(i_con_instru[3]), .B(n3), .Q(n21) );
  NAND31 U24 ( .A(n2), .B(n9), .C(i_con_instru[2]), .Q(n17) );
  NAND31 U25 ( .A(i_con_instru[1]), .B(n10), .C(n2), .Q(n23) );
  NAND22 U26 ( .A(i_con_instru[0]), .B(i_con_instru[1]), .Q(n24) );
  NAND22 U27 ( .A(i_con_instru[3]), .B(n6), .Q(n20) );
  INV3 U28 ( .A(i_con_instru[4]), .Q(n6) );
  INV3 U29 ( .A(i_con_instru[2]), .Q(n8) );
  NAND22 U30 ( .A(i_con_instru[5]), .B(n5), .Q(n16) );
  AOI211 U31 ( .A(n23), .B(n25), .C(i_con_instru[4]), .Q(o_con_aluop[3]) );
  NAND31 U32 ( .A(n2), .B(i_con_instru[0]), .C(i_con_instru[2]), .Q(n25) );
  INV3 U33 ( .A(i_con_instru[5]), .Q(n3) );
  NOR21 U34 ( .A(i_con_instru[3]), .B(n14), .Q(o_con_regdst) );
  AOI211 U35 ( .A(n17), .B(n22), .C(i_con_instru[4]), .Q(o_con_aluop[4]) );
  NAND22 U36 ( .A(n1), .B(n8), .Q(n22) );
  INV3 U37 ( .A(n23), .Q(n1) );
  AOI2111 U38 ( .A(n24), .B(n26), .C(n21), .D(i_con_instru[4]), .Q(
        o_con_aluop[2]) );
  NAND22 U39 ( .A(i_con_instru[2]), .B(n10), .Q(n26) );
  NOR21 U40 ( .A(i_con_instru[4]), .B(n21), .Q(o_con_aluop[0]) );
endmodule


module D_jb_control ( o_con_jump, o_con_bop, o_con_aluPC4, o_con_ifstall, 
        i_con_instru, i_con_func, i_con_rt );
  output [1:0] o_con_jump;
  output [2:0] o_con_bop;
  input [5:0] i_con_instru;
  input [5:0] i_con_func;
  input i_con_rt;
  output o_con_aluPC4, o_con_ifstall;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n2, n3, n4,
         n5, n6;

  OAI222 U13 ( .A(n5), .B(n16), .C(n14), .D(n17), .Q(o_con_bop[1]) );
  NAND31 U3 ( .A(n5), .B(n3), .C(n6), .Q(n8) );
  NAND22 U4 ( .A(n7), .B(n8), .Q(o_con_jump[1]) );
  INV3 U5 ( .A(n7), .Q(n2) );
  NAND22 U6 ( .A(n7), .B(n4), .Q(n17) );
  OAI311 U7 ( .A(n4), .B(n2), .C(n14), .D(n16), .Q(o_con_bop[0]) );
  INV3 U8 ( .A(n13), .Q(o_con_ifstall) );
  AOI211 U9 ( .A(n3), .B(n14), .C(n2), .Q(n13) );
  OAI2111 U10 ( .A(n9), .B(n8), .C(n10), .D(n7), .Q(o_con_jump[0]) );
  NOR40 U11 ( .A(n11), .B(i_con_func[2]), .C(i_con_func[5]), .D(i_con_func[4]), 
        .Q(n9) );
  NAND22 U12 ( .A(i_con_instru[1]), .B(n3), .Q(n10) );
  NAND22 U14 ( .A(n12), .B(i_con_func[3]), .Q(n11) );
  NOR31 U15 ( .A(i_con_instru[3]), .B(i_con_instru[5]), .C(i_con_instru[4]), 
        .Q(n7) );
  INV3 U16 ( .A(i_con_instru[2]), .Q(n3) );
  INV3 U17 ( .A(i_con_instru[1]), .Q(n5) );
  INV3 U18 ( .A(i_con_instru[0]), .Q(n6) );
  NOR21 U19 ( .A(i_con_func[1]), .B(i_con_func[0]), .Q(n12) );
  NOR40 U20 ( .A(i_con_instru[2]), .B(n2), .C(n5), .D(n6), .Q(o_con_aluPC4) );
  NAND31 U21 ( .A(n7), .B(n6), .C(i_con_instru[2]), .Q(n16) );
  NAND22 U22 ( .A(i_con_instru[0]), .B(n5), .Q(n14) );
  NOR31 U23 ( .A(n15), .B(n2), .C(n6), .Q(o_con_bop[2]) );
  XNR21 U24 ( .A(n5), .B(i_con_instru[2]), .Q(n15) );
  INV3 U25 ( .A(n18), .Q(n4) );
  NOR21 U26 ( .A(i_con_instru[2]), .B(i_con_rt), .Q(n18) );
endmodule


module D_pcadd_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279;

  NAND22 U2 ( .A(n23), .B(n25), .Q(n26) );
  NAND22 U3 ( .A(n236), .B(n231), .Q(n246) );
  NAND22 U4 ( .A(n190), .B(n188), .Q(n220) );
  NAND22 U5 ( .A(n181), .B(n189), .Q(n215) );
  NAND22 U6 ( .A(n152), .B(n147), .Q(n170) );
  NAND22 U7 ( .A(n175), .B(n176), .Q(n106) );
  NOR21 U8 ( .A(n177), .B(n178), .Q(n176) );
  NOR21 U9 ( .A(n195), .B(n196), .Q(n175) );
  INV3 U10 ( .A(n179), .Q(n178) );
  INV3 U11 ( .A(B[30]), .Q(n9) );
  NAND22 U12 ( .A(n103), .B(n104), .Q(n67) );
  AOI211 U13 ( .A(n109), .B(n110), .C(n111), .Q(n103) );
  NAND22 U14 ( .A(n105), .B(n106), .Q(n104) );
  NOR21 U15 ( .A(n202), .B(n33), .Q(n195) );
  NAND31 U16 ( .A(n200), .B(n201), .C(n204), .Q(n202) );
  AOI211 U17 ( .A(n204), .B(n203), .C(n251), .Q(n16) );
  NAND22 U18 ( .A(n198), .B(n199), .Q(n251) );
  AOI211 U19 ( .A(n143), .B(n106), .C(n110), .Q(n139) );
  INV3 U20 ( .A(n107), .Q(n143) );
  OAI2111 U21 ( .A(n16), .B(n208), .C(n192), .D(n193), .Q(n228) );
  AOI311 U22 ( .A(n180), .B(n181), .C(n182), .D(n183), .Q(n179) );
  NOR21 U23 ( .A(n184), .B(n185), .Q(n183) );
  INV3 U24 ( .A(n191), .Q(n180) );
  OAI2111 U25 ( .A(n186), .B(n187), .C(n188), .D(n189), .Q(n182) );
  AOI211 U26 ( .A(n192), .B(n193), .C(n194), .Q(n177) );
  NAND22 U27 ( .A(n120), .B(n134), .Q(n129) );
  NAND22 U28 ( .A(n135), .B(n121), .Q(n134) );
  NAND22 U29 ( .A(n229), .B(n230), .Q(n193) );
  AOI211 U30 ( .A(n234), .B(n231), .C(n235), .Q(n229) );
  AOI311 U31 ( .A(n231), .B(n13), .C(n232), .D(n233), .Q(n230) );
  NAND22 U32 ( .A(n152), .B(n168), .Q(n163) );
  NAND22 U33 ( .A(n169), .B(n147), .Q(n168) );
  NAND22 U34 ( .A(n83), .B(n95), .Q(n90) );
  NAND22 U35 ( .A(n96), .B(n84), .Q(n95) );
  NAND22 U36 ( .A(n200), .B(n201), .Q(n197) );
  XOR21 U37 ( .A(n135), .B(n136), .Q(SUM[21]) );
  NOR21 U38 ( .A(n137), .B(n118), .Q(n136) );
  XOR21 U39 ( .A(n96), .B(n97), .Q(SUM[25]) );
  NOR21 U40 ( .A(n98), .B(n81), .Q(n97) );
  XOR21 U41 ( .A(n129), .B(n130), .Q(SUM[22]) );
  NOR21 U42 ( .A(n117), .B(n131), .Q(n130) );
  XOR21 U43 ( .A(n163), .B(n164), .Q(SUM[18]) );
  NOR21 U44 ( .A(n150), .B(n165), .Q(n164) );
  XOR21 U45 ( .A(n90), .B(n91), .Q(SUM[26]) );
  NOR21 U46 ( .A(n80), .B(n92), .Q(n91) );
  XNR21 U47 ( .A(n26), .B(n22), .Q(SUM[6]) );
  XNR21 U48 ( .A(n246), .B(n244), .Q(SUM[10]) );
  XNR21 U49 ( .A(n220), .B(n217), .Q(SUM[13]) );
  XNR21 U50 ( .A(n215), .B(n213), .Q(SUM[14]) );
  XOR21 U51 ( .A(n10), .B(n11), .Q(SUM[9]) );
  NAND22 U52 ( .A(n12), .B(n13), .Q(n10) );
  NAND22 U53 ( .A(n188), .B(n216), .Q(n213) );
  NAND22 U54 ( .A(n217), .B(n190), .Q(n216) );
  NOR21 U55 ( .A(n107), .B(n108), .Q(n105) );
  NAND22 U56 ( .A(n151), .B(n152), .Q(n149) );
  NOR21 U57 ( .A(n68), .B(n69), .Q(n66) );
  XNR21 U58 ( .A(n169), .B(n170), .Q(SUM[17]) );
  XOR21 U59 ( .A(n30), .B(n31), .Q(SUM[5]) );
  NOR21 U60 ( .A(n27), .B(n32), .Q(n31) );
  INV3 U61 ( .A(n29), .Q(n32) );
  XOR21 U62 ( .A(n44), .B(n57), .Q(SUM[2]) );
  NOR21 U63 ( .A(n58), .B(n46), .Q(n57) );
  INV3 U64 ( .A(n82), .Q(n126) );
  XOR21 U65 ( .A(n61), .B(n158), .Q(SUM[1]) );
  NOR21 U66 ( .A(n159), .B(n63), .Q(n158) );
  INV3 U67 ( .A(n151), .Q(n210) );
  NAND22 U68 ( .A(n59), .B(n60), .Q(n44) );
  NAND22 U69 ( .A(n61), .B(n62), .Q(n60) );
  INV3 U70 ( .A(n63), .Q(n62) );
  INV3 U71 ( .A(n46), .Q(n45) );
  NAND31 U72 ( .A(n181), .B(n190), .C(n205), .Q(n194) );
  NOR21 U73 ( .A(n206), .B(n207), .Q(n205) );
  NOR21 U74 ( .A(B[15]), .B(A[15]), .Q(n207) );
  NOR21 U75 ( .A(B[12]), .B(A[12]), .Q(n206) );
  NAND22 U76 ( .A(n54), .B(n55), .Q(n50) );
  NAND22 U77 ( .A(B[29]), .B(A[29]), .Q(n54) );
  NAND22 U78 ( .A(n64), .B(n65), .Q(n56) );
  AOI221 U79 ( .A(B[28]), .B(A[28]), .C(n70), .D(n71), .Q(n64) );
  NAND22 U80 ( .A(n66), .B(n67), .Q(n65) );
  INV3 U81 ( .A(n69), .Q(n71) );
  XOR21 U82 ( .A(n47), .B(n48), .Q(SUM[31]) );
  XNR21 U83 ( .A(B[31]), .B(A[31]), .Q(n47) );
  AOI211 U84 ( .A(n49), .B(n50), .C(n51), .Q(n48) );
  NOR21 U85 ( .A(n52), .B(n9), .Q(n51) );
  NOR21 U86 ( .A(A[20]), .B(B[20]), .Q(n140) );
  NAND22 U87 ( .A(n273), .B(n274), .Q(n23) );
  INV3 U88 ( .A(A[6]), .Q(n274) );
  INV3 U89 ( .A(B[6]), .Q(n273) );
  NOR21 U90 ( .A(A[4]), .B(B[4]), .Q(n34) );
  NOR21 U91 ( .A(A[5]), .B(B[5]), .Q(n27) );
  NAND22 U92 ( .A(B[19]), .B(A[19]), .Q(n146) );
  NOR21 U93 ( .A(A[19]), .B(B[19]), .Q(n145) );
  AOI311 U94 ( .A(n147), .B(n148), .C(n149), .D(n150), .Q(n144) );
  NAND22 U95 ( .A(n3), .B(n171), .Q(n147) );
  INV3 U96 ( .A(A[17]), .Q(n171) );
  INV3 U97 ( .A(B[17]), .Q(n3) );
  NAND22 U98 ( .A(B[27]), .B(A[27]), .Q(n77) );
  NOR21 U99 ( .A(A[27]), .B(B[27]), .Q(n76) );
  AOI211 U100 ( .A(n78), .B(n79), .C(n80), .Q(n75) );
  NAND31 U101 ( .A(n79), .B(n84), .C(n85), .Q(n68) );
  NOR21 U102 ( .A(n86), .B(n87), .Q(n85) );
  NOR21 U103 ( .A(B[27]), .B(A[27]), .Q(n87) );
  NOR21 U104 ( .A(B[24]), .B(A[24]), .Q(n86) );
  NOR21 U105 ( .A(A[12]), .B(B[12]), .Q(n222) );
  NAND22 U106 ( .A(B[10]), .B(A[10]), .Q(n231) );
  NAND22 U107 ( .A(n224), .B(n225), .Q(n190) );
  INV3 U108 ( .A(A[13]), .Q(n225) );
  INV3 U109 ( .A(B[13]), .Q(n224) );
  NAND22 U110 ( .A(B[24]), .B(A[24]), .Q(n82) );
  NAND22 U111 ( .A(B[16]), .B(A[16]), .Q(n151) );
  NAND31 U112 ( .A(n236), .B(n12), .C(n237), .Q(n208) );
  NOR21 U113 ( .A(n238), .B(n239), .Q(n237) );
  NOR21 U114 ( .A(B[11]), .B(A[11]), .Q(n238) );
  NOR21 U115 ( .A(B[8]), .B(A[8]), .Q(n239) );
  NAND22 U116 ( .A(n218), .B(n219), .Q(n181) );
  INV3 U117 ( .A(A[14]), .Q(n219) );
  INV3 U118 ( .A(B[14]), .Q(n218) );
  NAND22 U119 ( .A(n4), .B(n166), .Q(n148) );
  INV3 U120 ( .A(A[18]), .Q(n166) );
  INV3 U121 ( .A(B[18]), .Q(n4) );
  NAND22 U122 ( .A(B[22]), .B(A[22]), .Q(n133) );
  XOR21 U123 ( .A(n72), .B(n73), .Q(SUM[28]) );
  XNR21 U124 ( .A(B[28]), .B(A[28]), .Q(n72) );
  AOI211 U125 ( .A(n74), .B(n67), .C(n70), .Q(n73) );
  NAND22 U126 ( .A(B[18]), .B(A[18]), .Q(n167) );
  NAND22 U127 ( .A(B[17]), .B(A[17]), .Q(n152) );
  NAND22 U128 ( .A(B[6]), .B(A[6]), .Q(n25) );
  NAND22 U129 ( .A(B[14]), .B(A[14]), .Q(n189) );
  NAND22 U130 ( .A(B[13]), .B(A[13]), .Q(n188) );
  NAND22 U131 ( .A(B[9]), .B(A[9]), .Q(n13) );
  NAND22 U132 ( .A(B[20]), .B(A[20]), .Q(n119) );
  NOR21 U133 ( .A(A[3]), .B(B[3]), .Q(n267) );
  NOR21 U134 ( .A(A[8]), .B(B[8]), .Q(n250) );
  NAND22 U135 ( .A(B[23]), .B(A[23]), .Q(n114) );
  NOR21 U136 ( .A(A[23]), .B(B[23]), .Q(n113) );
  AOI211 U137 ( .A(n115), .B(n116), .C(n117), .Q(n112) );
  NAND22 U138 ( .A(B[7]), .B(A[7]), .Q(n199) );
  NOR21 U139 ( .A(A[28]), .B(B[28]), .Q(n69) );
  NAND22 U140 ( .A(B[21]), .B(A[21]), .Q(n120) );
  NAND22 U141 ( .A(B[25]), .B(A[25]), .Q(n83) );
  NAND22 U142 ( .A(n100), .B(n82), .Q(n96) );
  NAND22 U143 ( .A(n172), .B(n151), .Q(n169) );
  NOR21 U144 ( .A(n270), .B(n271), .Q(n204) );
  NAND22 U145 ( .A(n23), .B(n272), .Q(n270) );
  INV3 U146 ( .A(n27), .Q(n272) );
  NOR21 U147 ( .A(n267), .B(n268), .Q(n266) );
  NAND22 U148 ( .A(A[2]), .B(B[2]), .Q(n268) );
  NAND22 U149 ( .A(B[11]), .B(A[11]), .Q(n192) );
  NAND31 U150 ( .A(n116), .B(n121), .C(n122), .Q(n108) );
  NOR21 U151 ( .A(n123), .B(n124), .Q(n122) );
  NOR21 U152 ( .A(B[23]), .B(A[23]), .Q(n124) );
  NOR21 U153 ( .A(B[20]), .B(A[20]), .Q(n123) );
  XOR21 U154 ( .A(n20), .B(n21), .Q(SUM[7]) );
  XNR21 U155 ( .A(B[7]), .B(A[7]), .Q(n20) );
  AOI211 U156 ( .A(n22), .B(n23), .C(n24), .Q(n21) );
  XOR21 U157 ( .A(n242), .B(n243), .Q(SUM[11]) );
  XNR21 U158 ( .A(B[11]), .B(A[11]), .Q(n242) );
  AOI211 U159 ( .A(n244), .B(n236), .C(n245), .Q(n243) );
  XOR21 U160 ( .A(n211), .B(n212), .Q(SUM[15]) );
  XNR21 U161 ( .A(B[15]), .B(A[15]), .Q(n211) );
  AOI211 U162 ( .A(n213), .B(n181), .C(n214), .Q(n212) );
  XOR21 U163 ( .A(n161), .B(n162), .Q(SUM[19]) );
  XNR21 U164 ( .A(B[19]), .B(A[19]), .Q(n161) );
  AOI211 U165 ( .A(n163), .B(n148), .C(n150), .Q(n162) );
  XOR21 U166 ( .A(n127), .B(n128), .Q(SUM[23]) );
  XNR21 U167 ( .A(B[23]), .B(A[23]), .Q(n127) );
  AOI211 U168 ( .A(n129), .B(n116), .C(n117), .Q(n128) );
  XOR21 U169 ( .A(n88), .B(n89), .Q(SUM[27]) );
  XNR21 U170 ( .A(B[27]), .B(A[27]), .Q(n88) );
  AOI211 U171 ( .A(n90), .B(n79), .C(n80), .Q(n89) );
  XNR21 U172 ( .A(n50), .B(n1), .Q(SUM[30]) );
  XNR21 U173 ( .A(B[30]), .B(A[30]), .Q(n1) );
  XNR21 U174 ( .A(n56), .B(n2), .Q(SUM[29]) );
  XNR21 U175 ( .A(B[29]), .B(A[29]), .Q(n2) );
  NAND22 U176 ( .A(A[12]), .B(B[12]), .Q(n187) );
  NOR21 U177 ( .A(A[15]), .B(B[15]), .Q(n191) );
  NAND22 U178 ( .A(B[8]), .B(A[8]), .Q(n232) );
  NAND31 U179 ( .A(n148), .B(n147), .C(n153), .Q(n107) );
  NOR21 U180 ( .A(n154), .B(n155), .Q(n153) );
  NOR21 U181 ( .A(B[16]), .B(A[16]), .Q(n154) );
  NOR21 U182 ( .A(B[19]), .B(A[19]), .Q(n155) );
  NOR21 U183 ( .A(A[11]), .B(B[11]), .Q(n233) );
  IMUX21 U184 ( .A(n101), .B(n102), .S(n67), .Q(SUM[24]) );
  XNR21 U185 ( .A(B[24]), .B(A[24]), .Q(n101) );
  NOR21 U186 ( .A(n125), .B(n126), .Q(n102) );
  NOR21 U187 ( .A(B[24]), .B(A[24]), .Q(n125) );
  IMUX21 U188 ( .A(n141), .B(n142), .S(n139), .Q(SUM[20]) );
  XNR21 U189 ( .A(B[20]), .B(A[20]), .Q(n142) );
  NOR21 U190 ( .A(n156), .B(n157), .Q(n141) );
  NOR21 U191 ( .A(B[20]), .B(A[20]), .Q(n156) );
  IMUX21 U192 ( .A(n226), .B(n227), .S(n221), .Q(SUM[12]) );
  NOR21 U193 ( .A(n240), .B(n241), .Q(n226) );
  XNR21 U194 ( .A(B[12]), .B(A[12]), .Q(n227) );
  NOR21 U195 ( .A(B[12]), .B(A[12]), .Q(n240) );
  INV3 U196 ( .A(B[15]), .Q(n185) );
  INV3 U197 ( .A(A[15]), .Q(n184) );
  NAND22 U198 ( .A(B[26]), .B(A[26]), .Q(n94) );
  INV3 U199 ( .A(n252), .Q(n198) );
  AOI311 U200 ( .A(n25), .B(n253), .C(n254), .D(n255), .Q(n252) );
  NOR21 U201 ( .A(A[7]), .B(B[7]), .Q(n255) );
  NAND31 U202 ( .A(A[5]), .B(B[5]), .C(n23), .Q(n253) );
  NAND31 U203 ( .A(n256), .B(n257), .C(n258), .Q(n203) );
  NAND22 U204 ( .A(n260), .B(n261), .Q(n257) );
  NAND22 U205 ( .A(B[3]), .B(A[3]), .Q(n258) );
  NOR21 U206 ( .A(n265), .B(n266), .Q(n256) );
  NAND41 U207 ( .A(B[4]), .B(A[4]), .C(n272), .D(n23), .Q(n254) );
  NAND22 U208 ( .A(n247), .B(n248), .Q(n12) );
  INV3 U209 ( .A(A[9]), .Q(n248) );
  INV3 U210 ( .A(B[9]), .Q(n247) );
  NAND22 U211 ( .A(n275), .B(n276), .Q(n236) );
  INV3 U212 ( .A(A[10]), .Q(n276) );
  INV3 U213 ( .A(B[10]), .Q(n275) );
  NAND22 U214 ( .A(n6), .B(n132), .Q(n116) );
  INV3 U215 ( .A(A[22]), .Q(n132) );
  INV3 U216 ( .A(B[22]), .Q(n6) );
  NAND22 U217 ( .A(n8), .B(n93), .Q(n79) );
  INV3 U218 ( .A(A[26]), .Q(n93) );
  INV3 U219 ( .A(B[26]), .Q(n8) );
  NAND22 U220 ( .A(n5), .B(n138), .Q(n121) );
  INV3 U221 ( .A(A[21]), .Q(n138) );
  INV3 U222 ( .A(B[21]), .Q(n5) );
  NAND22 U223 ( .A(n7), .B(n99), .Q(n84) );
  INV3 U224 ( .A(A[25]), .Q(n99) );
  INV3 U225 ( .A(B[25]), .Q(n7) );
  NOR21 U226 ( .A(A[2]), .B(B[2]), .Q(n46) );
  NAND22 U227 ( .A(B[4]), .B(A[4]), .Q(n35) );
  NAND22 U228 ( .A(B[5]), .B(A[5]), .Q(n29) );
  NAND22 U229 ( .A(B[12]), .B(A[12]), .Q(n223) );
  NAND22 U230 ( .A(B[8]), .B(A[8]), .Q(n19) );
  NAND22 U231 ( .A(B[2]), .B(A[2]), .Q(n42) );
  XOR21 U232 ( .A(n40), .B(n41), .Q(SUM[3]) );
  NAND22 U233 ( .A(n42), .B(n43), .Q(n40) );
  XOR21 U234 ( .A(B[3]), .B(A[3]), .Q(n41) );
  NAND22 U235 ( .A(n44), .B(n45), .Q(n43) );
  IMUX21 U236 ( .A(n173), .B(n174), .S(n106), .Q(SUM[16]) );
  XNR21 U237 ( .A(B[16]), .B(A[16]), .Q(n173) );
  NOR21 U238 ( .A(n209), .B(n210), .Q(n174) );
  NOR21 U239 ( .A(B[16]), .B(A[16]), .Q(n209) );
  IMUX21 U240 ( .A(n14), .B(n15), .S(n16), .Q(SUM[8]) );
  NOR21 U241 ( .A(n17), .B(n18), .Q(n14) );
  XNR21 U242 ( .A(B[8]), .B(A[8]), .Q(n15) );
  NOR21 U243 ( .A(B[8]), .B(A[8]), .Q(n17) );
  IMUX21 U244 ( .A(n36), .B(n37), .S(n33), .Q(SUM[4]) );
  NOR21 U245 ( .A(n38), .B(n39), .Q(n36) );
  XNR21 U246 ( .A(B[4]), .B(A[4]), .Q(n37) );
  NOR21 U247 ( .A(B[4]), .B(A[4]), .Q(n38) );
  INV3 U248 ( .A(n53), .Q(n49) );
  NOR21 U249 ( .A(A[30]), .B(B[30]), .Q(n53) );
  NOR21 U250 ( .A(A[1]), .B(B[1]), .Q(n63) );
  INV3 U251 ( .A(B[0]), .Q(n277) );
  INV3 U252 ( .A(n279), .Q(n278) );
  NOR21 U253 ( .A(B[0]), .B(n259), .Q(n279) );
  INV3 U254 ( .A(A[30]), .Q(n52) );
  INV3 U255 ( .A(A[0]), .Q(n259) );
  NOR31 U256 ( .A(n269), .B(n46), .C(n267), .Q(n265) );
  NAND22 U257 ( .A(B[1]), .B(A[1]), .Q(n269) );
  AOI211 U258 ( .A(n263), .B(n264), .C(n63), .Q(n260) );
  INV3 U259 ( .A(A[3]), .Q(n264) );
  INV3 U260 ( .A(B[3]), .Q(n263) );
  NAND22 U261 ( .A(B[1]), .B(A[1]), .Q(n59) );
  NOR21 U262 ( .A(n46), .B(n262), .Q(n261) );
  NAND22 U263 ( .A(B[0]), .B(A[0]), .Q(n262) );
  INV3 U264 ( .A(n160), .Q(n61) );
  NAND22 U265 ( .A(B[0]), .B(A[0]), .Q(n160) );
  CLKIN3 U266 ( .A(n19), .Q(n18) );
  CLKIN3 U267 ( .A(n25), .Q(n24) );
  OAI212 U268 ( .A(n27), .B(n28), .C(n29), .Q(n22) );
  CLKIN3 U269 ( .A(n30), .Q(n28) );
  OAI212 U270 ( .A(n33), .B(n34), .C(n35), .Q(n30) );
  CLKIN3 U271 ( .A(n35), .Q(n39) );
  OAI212 U272 ( .A(A[29]), .B(B[29]), .C(n56), .Q(n55) );
  CLKIN3 U273 ( .A(n42), .Q(n58) );
  OAI212 U274 ( .A(n75), .B(n76), .C(n77), .Q(n70) );
  OAI212 U275 ( .A(n81), .B(n82), .C(n83), .Q(n78) );
  CLKIN3 U276 ( .A(n68), .Q(n74) );
  CLKIN3 U277 ( .A(n79), .Q(n92) );
  CLKIN3 U278 ( .A(n94), .Q(n80) );
  CLKIN3 U279 ( .A(n84), .Q(n81) );
  CLKIN3 U280 ( .A(n83), .Q(n98) );
  OAI212 U281 ( .A(A[24]), .B(B[24]), .C(n67), .Q(n100) );
  OAI212 U282 ( .A(n112), .B(n113), .C(n114), .Q(n111) );
  OAI212 U283 ( .A(n118), .B(n119), .C(n120), .Q(n115) );
  CLKIN3 U284 ( .A(n108), .Q(n109) );
  CLKIN3 U285 ( .A(n116), .Q(n131) );
  CLKIN3 U286 ( .A(n133), .Q(n117) );
  CLKIN3 U287 ( .A(n121), .Q(n118) );
  CLKIN3 U288 ( .A(n120), .Q(n137) );
  OAI212 U289 ( .A(n139), .B(n140), .C(n119), .Q(n135) );
  OAI212 U290 ( .A(n144), .B(n145), .C(n146), .Q(n110) );
  CLKIN3 U291 ( .A(n119), .Q(n157) );
  CLKIN3 U292 ( .A(n59), .Q(n159) );
  CLKIN3 U293 ( .A(n148), .Q(n165) );
  CLKIN3 U294 ( .A(n167), .Q(n150) );
  OAI212 U295 ( .A(A[16]), .B(B[16]), .C(n106), .Q(n172) );
  CLKIN3 U296 ( .A(n190), .Q(n186) );
  OAI222 U297 ( .A(n197), .B(n198), .C(n197), .D(n199), .Q(n196) );
  CLKIN3 U298 ( .A(n203), .Q(n33) );
  CLKIN3 U299 ( .A(n194), .Q(n201) );
  CLKIN3 U300 ( .A(n208), .Q(n200) );
  CLKIN3 U301 ( .A(n189), .Q(n214) );
  OAI212 U302 ( .A(n221), .B(n222), .C(n223), .Q(n217) );
  CLKIN3 U303 ( .A(n228), .Q(n221) );
  CLKIN3 U304 ( .A(n236), .Q(n235) );
  CLKIN3 U305 ( .A(n223), .Q(n241) );
  CLKIN3 U306 ( .A(n231), .Q(n245) );
  OAI212 U307 ( .A(n11), .B(n234), .C(n13), .Q(n244) );
  CLKIN3 U308 ( .A(n12), .Q(n234) );
  CLKIN3 U309 ( .A(n249), .Q(n11) );
  OAI212 U310 ( .A(n16), .B(n250), .C(n19), .Q(n249) );
  OAI222 U311 ( .A(B[7]), .B(A[7]), .C(B[4]), .D(A[4]), .Q(n271) );
  OAI212 U312 ( .A(A[0]), .B(n277), .C(n278), .Q(SUM[0]) );
endmodule


module D_pcadd ( i_addr_pcadd4E, i_data_immshiftl, o_addr_pcbranchE );
  input [31:0] i_addr_pcadd4E;
  input [31:0] i_data_immshiftl;
  output [31:0] o_addr_pcbranchE;
  wire   n1;

  D_pcadd_DW01_add_1 add_5 ( .A(i_addr_pcadd4E), .B(i_data_immshiftl), .CI(n1), 
        .SUM(o_addr_pcbranchE) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_addr_Rt, i_con_RegWr, 
        i_addr_Rd, i_data_Rd, o_data_Rs, o_data_Rt );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rt;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr;
  wire   n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856;
  wire   [1023:0] regs;

  DFEC1 regs_reg_30__31_ ( .D(i_data_Rd[31]), .E(n832), .C(i_clk), .RN(n810), 
        .Q(regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(i_data_Rd[30]), .E(n832), .C(i_clk), .RN(n810), 
        .Q(regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(i_data_Rd[29]), .E(n832), .C(i_clk), .RN(n810), 
        .Q(regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(i_data_Rd[28]), .E(n832), .C(i_clk), .RN(n810), 
        .Q(regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(i_data_Rd[27]), .E(n832), .C(i_clk), .RN(n811), 
        .Q(regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(i_data_Rd[26]), .E(n832), .C(i_clk), .RN(n811), 
        .Q(regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(i_data_Rd[25]), .E(n832), .C(i_clk), .RN(n811), 
        .Q(regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(i_data_Rd[24]), .E(n832), .C(i_clk), .RN(n811), 
        .Q(regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(i_data_Rd[23]), .E(n832), .C(i_clk), .RN(n811), 
        .Q(regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(i_data_Rd[22]), .E(n832), .C(i_clk), .RN(n811), 
        .Q(regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(i_data_Rd[21]), .E(n832), .C(i_clk), .RN(n811), 
        .Q(regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(i_data_Rd[20]), .E(n832), .C(i_clk), .RN(n811), 
        .Q(regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n832), .C(i_clk), .RN(n811), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(i_data_Rd[18]), .E(n832), .C(i_clk), .RN(n812), 
        .Q(regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(i_data_Rd[17]), .E(n832), .C(i_clk), .RN(n812), 
        .Q(regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(i_data_Rd[16]), .E(n832), .C(i_clk), .RN(n812), 
        .Q(regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(i_data_Rd[15]), .E(n832), .C(i_clk), .RN(n812), 
        .Q(regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(i_data_Rd[14]), .E(n832), .C(i_clk), .RN(n812), 
        .Q(regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(i_data_Rd[13]), .E(n832), .C(i_clk), .RN(n812), 
        .Q(regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(i_data_Rd[12]), .E(n832), .C(i_clk), .RN(n812), 
        .Q(regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(i_data_Rd[11]), .E(n832), .C(i_clk), .RN(n812), 
        .Q(regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(i_data_Rd[10]), .E(n832), .C(i_clk), .RN(n812), 
        .Q(regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(i_data_Rd[9]), .E(n832), .C(i_clk), .RN(n813), 
        .Q(regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(i_data_Rd[8]), .E(n832), .C(i_clk), .RN(n813), 
        .Q(regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(i_data_Rd[7]), .E(n832), .C(i_clk), .RN(n813), 
        .Q(regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n832), .C(i_clk), .RN(n813), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(i_data_Rd[5]), .E(n832), .C(i_clk), .RN(n813), 
        .Q(regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(i_data_Rd[4]), .E(n832), .C(i_clk), .RN(n813), 
        .Q(regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(i_data_Rd[3]), .E(n832), .C(i_clk), .RN(n813), 
        .Q(regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(i_data_Rd[2]), .E(n832), .C(i_clk), .RN(n813), 
        .Q(regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n832), .C(i_clk), .RN(n813), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(i_data_Rd[0]), .E(n832), .C(i_clk), .RN(n814), 
        .Q(regs[960]) );
  DFEC1 regs_reg_26__31_ ( .D(i_data_Rd[31]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(i_data_Rd[30]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(i_data_Rd[29]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(i_data_Rd[28]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(i_data_Rd[27]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(i_data_Rd[26]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(i_data_Rd[25]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(i_data_Rd[24]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(i_data_Rd[23]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(i_data_Rd[22]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(i_data_Rd[21]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(i_data_Rd[20]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(i_data_Rd[18]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(i_data_Rd[17]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(i_data_Rd[16]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(i_data_Rd[15]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(i_data_Rd[14]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(i_data_Rd[13]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(i_data_Rd[12]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(i_data_Rd[11]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(i_data_Rd[10]), .E(n828), .C(i_clk), .RN(i_rst_n), .Q(regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(i_data_Rd[9]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(i_data_Rd[8]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(i_data_Rd[7]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(i_data_Rd[5]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(i_data_Rd[4]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(i_data_Rd[3]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(i_data_Rd[2]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(i_data_Rd[0]), .E(n828), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[832]) );
  DFEC1 regs_reg_22__31_ ( .D(i_data_Rd[31]), .E(n820), .C(i_clk), .RN(n809), 
        .Q(regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(i_data_Rd[30]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(i_data_Rd[29]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(i_data_Rd[28]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(i_data_Rd[27]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(i_data_Rd[26]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(i_data_Rd[25]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(i_data_Rd[24]), .E(n820), .C(i_clk), .RN(n818), 
        .Q(regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(i_data_Rd[23]), .E(n820), .C(i_clk), .RN(n812), 
        .Q(regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(i_data_Rd[22]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(i_data_Rd[21]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(i_data_Rd[20]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(i_data_Rd[19]), .E(n820), .C(i_clk), .RN(n815), 
        .Q(regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(i_data_Rd[18]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(i_data_Rd[17]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(i_data_Rd[16]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(i_data_Rd[15]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(i_data_Rd[14]), .E(n820), .C(i_clk), .RN(n814), 
        .Q(regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(i_data_Rd[13]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(i_data_Rd[12]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(i_data_Rd[11]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(i_data_Rd[10]), .E(n820), .C(i_clk), .RN(i_rst_n), .Q(regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(i_data_Rd[9]), .E(n820), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(i_data_Rd[8]), .E(n820), .C(i_clk), .RN(n810), 
        .Q(regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(i_data_Rd[7]), .E(n820), .C(i_clk), .RN(n809), 
        .Q(regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(i_data_Rd[6]), .E(n820), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(i_data_Rd[5]), .E(n820), .C(i_clk), .RN(n818), 
        .Q(regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(i_data_Rd[4]), .E(n820), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(i_data_Rd[3]), .E(n820), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(i_data_Rd[2]), .E(n820), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(i_data_Rd[1]), .E(n820), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(i_data_Rd[0]), .E(n820), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[704]) );
  DFEC1 regs_reg_18__31_ ( .D(i_data_Rd[31]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(i_data_Rd[30]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(i_data_Rd[29]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(i_data_Rd[28]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(i_data_Rd[27]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(i_data_Rd[26]), .E(n824), .C(i_clk), .RN(n811), 
        .Q(regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(i_data_Rd[25]), .E(n824), .C(i_clk), .RN(n817), 
        .Q(regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(i_data_Rd[24]), .E(n824), .C(i_clk), .RN(n811), 
        .Q(regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(i_data_Rd[23]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(i_data_Rd[22]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(i_data_Rd[21]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(i_data_Rd[20]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(i_data_Rd[19]), .E(n824), .C(i_clk), .RN(n816), 
        .Q(regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(i_data_Rd[18]), .E(n824), .C(i_clk), .RN(n813), 
        .Q(regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(i_data_Rd[17]), .E(n824), .C(i_clk), .RN(n814), 
        .Q(regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(i_data_Rd[16]), .E(n824), .C(i_clk), .RN(n810), 
        .Q(regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(i_data_Rd[15]), .E(n824), .C(i_clk), .RN(n818), 
        .Q(regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(i_data_Rd[14]), .E(n824), .C(i_clk), .RN(n813), 
        .Q(regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(i_data_Rd[13]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(i_data_Rd[12]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(i_data_Rd[11]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(i_data_Rd[10]), .E(n824), .C(i_clk), .RN(i_rst_n), .Q(regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(i_data_Rd[9]), .E(n824), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(i_data_Rd[8]), .E(n824), .C(i_clk), .RN(n813), 
        .Q(regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(i_data_Rd[7]), .E(n824), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(i_data_Rd[6]), .E(n824), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(i_data_Rd[5]), .E(n824), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(i_data_Rd[4]), .E(n824), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(i_data_Rd[3]), .E(n824), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(i_data_Rd[2]), .E(n824), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(i_data_Rd[1]), .E(n824), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(i_data_Rd[0]), .E(n824), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[576]) );
  DFEC1 regs_reg_14__31_ ( .D(i_data_Rd[31]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(i_data_Rd[30]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(i_data_Rd[29]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(i_data_Rd[28]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(i_data_Rd[27]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(i_data_Rd[26]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(i_data_Rd[25]), .E(n837), .C(i_clk), .RN(n815), 
        .Q(regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(i_data_Rd[24]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(i_data_Rd[23]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(i_data_Rd[22]), .E(n837), .C(i_clk), .RN(n811), 
        .Q(regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(i_data_Rd[21]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(i_data_Rd[20]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(i_data_Rd[19]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(i_data_Rd[18]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(i_data_Rd[17]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(i_data_Rd[16]), .E(n837), .C(i_clk), .RN(n817), 
        .Q(regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(i_data_Rd[15]), .E(n837), .C(i_clk), .RN(n811), 
        .Q(regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n837), .C(i_clk), .RN(n812), 
        .Q(regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(i_data_Rd[13]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(i_data_Rd[12]), .E(n837), .C(i_clk), .RN(n812), 
        .Q(regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(i_data_Rd[11]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n837), .C(i_clk), .RN(i_rst_n), .Q(regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(i_data_Rd[9]), .E(n837), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(i_data_Rd[8]), .E(n837), .C(i_clk), .RN(n816), 
        .Q(regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(i_data_Rd[7]), .E(n837), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(i_data_Rd[6]), .E(n837), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(i_data_Rd[5]), .E(n837), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(i_data_Rd[4]), .E(n837), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(i_data_Rd[3]), .E(n837), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(i_data_Rd[2]), .E(n837), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(i_data_Rd[1]), .E(n837), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(i_data_Rd[0]), .E(n837), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[448]) );
  DFEC1 regs_reg_10__31_ ( .D(i_data_Rd[31]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(i_data_Rd[30]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(i_data_Rd[29]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(i_data_Rd[28]), .E(n841), .C(i_clk), .RN(n811), 
        .Q(regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(i_data_Rd[27]), .E(n841), .C(i_clk), .RN(n812), 
        .Q(regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(i_data_Rd[26]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(i_data_Rd[25]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(i_data_Rd[24]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(i_data_Rd[23]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(i_data_Rd[22]), .E(n841), .C(i_clk), .RN(n816), 
        .Q(regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(i_data_Rd[21]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(i_data_Rd[20]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(i_data_Rd[19]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(i_data_Rd[18]), .E(n841), .C(i_clk), .RN(n816), 
        .Q(regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(i_data_Rd[17]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(i_data_Rd[16]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(i_data_Rd[15]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(i_data_Rd[13]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(i_data_Rd[12]), .E(n841), .C(i_clk), .RN(n813), 
        .Q(regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(i_data_Rd[11]), .E(n841), .C(i_clk), .RN(i_rst_n), .Q(regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n841), .C(i_clk), .RN(n809), 
        .Q(regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(i_data_Rd[9]), .E(n841), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(i_data_Rd[8]), .E(n841), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(i_data_Rd[7]), .E(n841), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(i_data_Rd[6]), .E(n841), .C(i_clk), .RN(n818), 
        .Q(regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(i_data_Rd[5]), .E(n841), .C(i_clk), .RN(n817), 
        .Q(regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(i_data_Rd[4]), .E(n841), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(i_data_Rd[3]), .E(n841), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(i_data_Rd[2]), .E(n841), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(i_data_Rd[1]), .E(n841), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(i_data_Rd[0]), .E(n841), .C(i_clk), .RN(n815), 
        .Q(regs[320]) );
  DFEC1 regs_reg_6__31_ ( .D(i_data_Rd[31]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(i_data_Rd[30]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(i_data_Rd[29]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(i_data_Rd[28]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(i_data_Rd[27]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(i_data_Rd[26]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(i_data_Rd[25]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(i_data_Rd[24]), .E(n845), .C(i_clk), .RN(n809), 
        .Q(regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(i_data_Rd[23]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(i_data_Rd[22]), .E(n845), .C(i_clk), .RN(n811), 
        .Q(regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(i_data_Rd[21]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(i_data_Rd[20]), .E(n845), .C(i_clk), .RN(n817), 
        .Q(regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(i_data_Rd[19]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(i_data_Rd[18]), .E(n845), .C(i_clk), .RN(n811), 
        .Q(regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(i_data_Rd[17]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(i_data_Rd[16]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(i_data_Rd[15]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(i_data_Rd[14]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(i_data_Rd[13]), .E(n845), .C(i_clk), .RN(n818), 
        .Q(regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(i_data_Rd[12]), .E(n845), .C(i_clk), .RN(n809), 
        .Q(regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(i_data_Rd[11]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(i_data_Rd[10]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(i_data_Rd[9]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(i_data_Rd[8]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(i_data_Rd[7]), .E(n845), .C(i_clk), .RN(n815), .Q(
        regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(i_data_Rd[6]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(i_data_Rd[5]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(i_data_Rd[4]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(i_data_Rd[3]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(i_data_Rd[2]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(i_data_Rd[1]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(i_data_Rd[0]), .E(n845), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[192]) );
  DFEC1 regs_reg_2__31_ ( .D(i_data_Rd[31]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(i_data_Rd[30]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(i_data_Rd[29]), .E(n849), .C(i_clk), .RN(n809), 
        .Q(regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(i_data_Rd[28]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(i_data_Rd[27]), .E(n849), .C(i_clk), .RN(n815), 
        .Q(regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(i_data_Rd[26]), .E(n849), .C(i_clk), .RN(n809), 
        .Q(regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(i_data_Rd[25]), .E(n849), .C(i_clk), .RN(n813), 
        .Q(regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(i_data_Rd[24]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(i_data_Rd[23]), .E(n849), .C(i_clk), .RN(n814), 
        .Q(regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(i_data_Rd[22]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(i_data_Rd[21]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(i_data_Rd[20]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(i_data_Rd[19]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(i_data_Rd[18]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(i_data_Rd[17]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(i_data_Rd[16]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(i_data_Rd[15]), .E(n849), .C(i_clk), .RN(n818), 
        .Q(regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(i_data_Rd[14]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(i_data_Rd[13]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(i_data_Rd[12]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(i_data_Rd[11]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(i_data_Rd[10]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(i_data_Rd[9]), .E(n849), .C(i_clk), .RN(n810), .Q(
        regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(i_data_Rd[8]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(i_data_Rd[7]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(i_data_Rd[6]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(i_data_Rd[5]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(i_data_Rd[4]), .E(n849), .C(i_clk), .RN(n815), .Q(
        regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(i_data_Rd[3]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(i_data_Rd[2]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(i_data_Rd[1]), .E(n849), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(i_data_Rd[0]), .E(n849), .C(i_clk), .RN(n818), .Q(
        regs[64]) );
  DFEC1 regs_reg_31__31_ ( .D(i_data_Rd[31]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1023]) );
  DFEC1 regs_reg_31__30_ ( .D(i_data_Rd[30]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(i_data_Rd[29]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(i_data_Rd[28]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(i_data_Rd[27]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(i_data_Rd[26]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(i_data_Rd[25]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(i_data_Rd[24]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(i_data_Rd[23]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(i_data_Rd[22]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(i_data_Rd[21]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(i_data_Rd[20]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(i_data_Rd[18]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(i_data_Rd[17]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(i_data_Rd[16]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(i_data_Rd[15]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(i_data_Rd[14]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(i_data_Rd[13]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(i_data_Rd[12]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(i_data_Rd[11]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(i_data_Rd[10]), .E(n831), .C(i_clk), .RN(i_rst_n), .Q(regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(i_data_Rd[9]), .E(n831), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(i_data_Rd[8]), .E(n831), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(i_data_Rd[7]), .E(n831), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n831), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(i_data_Rd[5]), .E(n831), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(i_data_Rd[4]), .E(n831), .C(i_clk), .RN(n810), 
        .Q(regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(i_data_Rd[3]), .E(n831), .C(i_clk), .RN(n810), 
        .Q(regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(i_data_Rd[2]), .E(n831), .C(i_clk), .RN(n810), 
        .Q(regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n831), .C(i_clk), .RN(n810), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(i_data_Rd[0]), .E(n831), .C(i_clk), .RN(n810), 
        .Q(regs[992]) );
  DFEC1 regs_reg_29__31_ ( .D(i_data_Rd[31]), .E(n833), .C(i_clk), .RN(n814), 
        .Q(regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(i_data_Rd[30]), .E(n833), .C(i_clk), .RN(n814), 
        .Q(regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(i_data_Rd[29]), .E(n833), .C(i_clk), .RN(n814), 
        .Q(regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(i_data_Rd[28]), .E(n833), .C(i_clk), .RN(n814), 
        .Q(regs[956]) );
  DFEC1 regs_reg_29__27_ ( .D(i_data_Rd[27]), .E(n833), .C(i_clk), .RN(n814), 
        .Q(regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(i_data_Rd[26]), .E(n833), .C(i_clk), .RN(n814), 
        .Q(regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(i_data_Rd[25]), .E(n833), .C(i_clk), .RN(n814), 
        .Q(regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(i_data_Rd[24]), .E(n833), .C(i_clk), .RN(n814), 
        .Q(regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(i_data_Rd[23]), .E(n833), .C(i_clk), .RN(n815), 
        .Q(regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(i_data_Rd[22]), .E(n833), .C(i_clk), .RN(n815), 
        .Q(regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(i_data_Rd[21]), .E(n833), .C(i_clk), .RN(n815), 
        .Q(regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(i_data_Rd[20]), .E(n833), .C(i_clk), .RN(n815), 
        .Q(regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n833), .C(i_clk), .RN(n815), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(i_data_Rd[18]), .E(n833), .C(i_clk), .RN(n815), 
        .Q(regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(i_data_Rd[17]), .E(n833), .C(i_clk), .RN(n815), 
        .Q(regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(i_data_Rd[16]), .E(n833), .C(i_clk), .RN(n815), 
        .Q(regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(i_data_Rd[15]), .E(n833), .C(i_clk), .RN(n815), 
        .Q(regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(i_data_Rd[14]), .E(n833), .C(i_clk), .RN(n816), 
        .Q(regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(i_data_Rd[13]), .E(n833), .C(i_clk), .RN(n816), 
        .Q(regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(i_data_Rd[12]), .E(n833), .C(i_clk), .RN(n816), 
        .Q(regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(i_data_Rd[11]), .E(n833), .C(i_clk), .RN(n816), 
        .Q(regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(i_data_Rd[10]), .E(n833), .C(i_clk), .RN(n816), 
        .Q(regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(i_data_Rd[9]), .E(n833), .C(i_clk), .RN(n816), 
        .Q(regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(i_data_Rd[8]), .E(n833), .C(i_clk), .RN(n816), 
        .Q(regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(i_data_Rd[7]), .E(n833), .C(i_clk), .RN(n816), 
        .Q(regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n833), .C(i_clk), .RN(n816), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(i_data_Rd[5]), .E(n833), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(i_data_Rd[4]), .E(n833), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(i_data_Rd[3]), .E(n833), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(i_data_Rd[2]), .E(n833), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n833), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(i_data_Rd[0]), .E(n833), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[928]) );
  DFEC1 regs_reg_28__31_ ( .D(i_data_Rd[31]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(i_data_Rd[30]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(i_data_Rd[29]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(i_data_Rd[28]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(i_data_Rd[27]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(i_data_Rd[26]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(i_data_Rd[25]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(i_data_Rd[24]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(i_data_Rd[23]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(i_data_Rd[22]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(i_data_Rd[21]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(i_data_Rd[20]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(i_data_Rd[18]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(i_data_Rd[17]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(i_data_Rd[16]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(i_data_Rd[15]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(i_data_Rd[14]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(i_data_Rd[13]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(i_data_Rd[12]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(i_data_Rd[11]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(i_data_Rd[10]), .E(n834), .C(i_clk), .RN(i_rst_n), .Q(regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(i_data_Rd[9]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(i_data_Rd[8]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(i_data_Rd[7]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(i_data_Rd[5]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(i_data_Rd[4]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(i_data_Rd[3]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(i_data_Rd[2]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(i_data_Rd[0]), .E(n834), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(i_data_Rd[31]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(i_data_Rd[30]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(i_data_Rd[29]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(i_data_Rd[28]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(i_data_Rd[27]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(i_data_Rd[26]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(i_data_Rd[25]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(i_data_Rd[24]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(i_data_Rd[23]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(i_data_Rd[22]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(i_data_Rd[21]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(i_data_Rd[20]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(i_data_Rd[18]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(i_data_Rd[17]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(i_data_Rd[16]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(i_data_Rd[15]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(i_data_Rd[14]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(i_data_Rd[13]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(i_data_Rd[12]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(i_data_Rd[11]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(i_data_Rd[10]), .E(n827), .C(i_clk), .RN(i_rst_n), .Q(regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(i_data_Rd[9]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(i_data_Rd[8]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(i_data_Rd[7]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(i_data_Rd[5]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(i_data_Rd[4]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(i_data_Rd[3]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(i_data_Rd[2]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(i_data_Rd[1]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(i_data_Rd[0]), .E(n827), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[864]) );
  DFEC1 regs_reg_25__31_ ( .D(i_data_Rd[31]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(i_data_Rd[30]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(i_data_Rd[29]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(i_data_Rd[28]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(i_data_Rd[27]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(i_data_Rd[26]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(i_data_Rd[25]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(i_data_Rd[24]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(i_data_Rd[23]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(i_data_Rd[22]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(i_data_Rd[21]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(i_data_Rd[20]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(i_data_Rd[19]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(i_data_Rd[18]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(i_data_Rd[17]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(i_data_Rd[16]), .E(n829), .C(i_clk), .RN(n811), 
        .Q(regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(i_data_Rd[15]), .E(n829), .C(i_clk), .RN(n812), 
        .Q(regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(i_data_Rd[14]), .E(n829), .C(i_clk), .RN(n816), 
        .Q(regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(i_data_Rd[13]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(i_data_Rd[12]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(i_data_Rd[11]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(i_data_Rd[10]), .E(n829), .C(i_clk), .RN(i_rst_n), .Q(regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(i_data_Rd[9]), .E(n829), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(i_data_Rd[8]), .E(n829), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(i_data_Rd[7]), .E(n829), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(i_data_Rd[6]), .E(n829), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(i_data_Rd[5]), .E(n829), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(i_data_Rd[4]), .E(n829), .C(i_clk), .RN(n817), 
        .Q(regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(i_data_Rd[3]), .E(n829), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(i_data_Rd[2]), .E(n829), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(i_data_Rd[1]), .E(n829), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(i_data_Rd[0]), .E(n829), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[800]) );
  DFEC1 regs_reg_24__31_ ( .D(i_data_Rd[31]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(i_data_Rd[30]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(i_data_Rd[29]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(i_data_Rd[28]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(i_data_Rd[27]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(i_data_Rd[26]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(i_data_Rd[25]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(i_data_Rd[24]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(i_data_Rd[23]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(i_data_Rd[22]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(i_data_Rd[21]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(i_data_Rd[20]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(i_data_Rd[19]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(i_data_Rd[18]), .E(n830), .C(i_clk), .RN(n818), 
        .Q(regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(i_data_Rd[17]), .E(n830), .C(i_clk), .RN(n815), 
        .Q(regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(i_data_Rd[16]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(i_data_Rd[15]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(i_data_Rd[14]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(i_data_Rd[13]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(i_data_Rd[12]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(i_data_Rd[11]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(i_data_Rd[10]), .E(n830), .C(i_clk), .RN(i_rst_n), .Q(regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(i_data_Rd[9]), .E(n830), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(i_data_Rd[8]), .E(n830), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(i_data_Rd[7]), .E(n830), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(i_data_Rd[6]), .E(n830), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(i_data_Rd[5]), .E(n830), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(i_data_Rd[4]), .E(n830), .C(i_clk), .RN(n818), 
        .Q(regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(i_data_Rd[3]), .E(n830), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(i_data_Rd[2]), .E(n830), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(i_data_Rd[1]), .E(n830), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(i_data_Rd[0]), .E(n830), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(i_data_Rd[31]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(i_data_Rd[30]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(i_data_Rd[29]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(i_data_Rd[28]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(i_data_Rd[27]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(i_data_Rd[26]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(i_data_Rd[25]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(i_data_Rd[24]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(i_data_Rd[23]), .E(n819), .C(i_clk), .RN(n809), 
        .Q(regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(i_data_Rd[22]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(i_data_Rd[21]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(i_data_Rd[20]), .E(n819), .C(i_clk), .RN(n816), 
        .Q(regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(i_data_Rd[19]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(i_data_Rd[18]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(i_data_Rd[17]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(i_data_Rd[16]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(i_data_Rd[15]), .E(n819), .C(i_clk), .RN(n818), 
        .Q(regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(i_data_Rd[14]), .E(n819), .C(i_clk), .RN(n817), 
        .Q(regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(i_data_Rd[13]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(i_data_Rd[12]), .E(n819), .C(i_clk), .RN(n817), 
        .Q(regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(i_data_Rd[11]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(i_data_Rd[10]), .E(n819), .C(i_clk), .RN(i_rst_n), .Q(regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(i_data_Rd[9]), .E(n819), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(i_data_Rd[8]), .E(n819), .C(i_clk), .RN(n815), 
        .Q(regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(i_data_Rd[7]), .E(n819), .C(i_clk), .RN(n814), 
        .Q(regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(i_data_Rd[6]), .E(n819), .C(i_clk), .RN(n813), 
        .Q(regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(i_data_Rd[5]), .E(n819), .C(i_clk), .RN(n812), 
        .Q(regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(i_data_Rd[4]), .E(n819), .C(i_clk), .RN(n811), 
        .Q(regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(i_data_Rd[3]), .E(n819), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(i_data_Rd[2]), .E(n819), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(i_data_Rd[1]), .E(n819), .C(i_clk), .RN(n810), 
        .Q(regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(i_data_Rd[0]), .E(n819), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[736]) );
  DFEC1 regs_reg_21__31_ ( .D(i_data_Rd[31]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(i_data_Rd[30]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(i_data_Rd[29]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(i_data_Rd[28]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(i_data_Rd[27]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(i_data_Rd[26]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(i_data_Rd[25]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(i_data_Rd[24]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(i_data_Rd[23]), .E(n821), .C(i_clk), .RN(n809), 
        .Q(regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(i_data_Rd[22]), .E(n821), .C(i_clk), .RN(n810), 
        .Q(regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(i_data_Rd[21]), .E(n821), .C(i_clk), .RN(n809), 
        .Q(regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(i_data_Rd[20]), .E(n821), .C(i_clk), .RN(n818), 
        .Q(regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(i_data_Rd[19]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(i_data_Rd[18]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(i_data_Rd[17]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(i_data_Rd[16]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(i_data_Rd[15]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(i_data_Rd[14]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(i_data_Rd[13]), .E(n821), .C(i_clk), .RN(n814), 
        .Q(regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(i_data_Rd[12]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(i_data_Rd[11]), .E(n821), .C(i_clk), .RN(n817), 
        .Q(regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(i_data_Rd[10]), .E(n821), .C(i_clk), .RN(i_rst_n), .Q(regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(i_data_Rd[9]), .E(n821), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(i_data_Rd[8]), .E(n821), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(i_data_Rd[7]), .E(n821), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(i_data_Rd[6]), .E(n821), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(i_data_Rd[5]), .E(n821), .C(i_clk), .RN(n812), 
        .Q(regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(i_data_Rd[4]), .E(n821), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(i_data_Rd[3]), .E(n821), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(i_data_Rd[2]), .E(n821), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(i_data_Rd[1]), .E(n821), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(i_data_Rd[0]), .E(n821), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[672]) );
  DFEC1 regs_reg_20__31_ ( .D(i_data_Rd[31]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(i_data_Rd[30]), .E(n822), .C(i_clk), .RN(n810), 
        .Q(regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(i_data_Rd[29]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(i_data_Rd[28]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(i_data_Rd[27]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(i_data_Rd[26]), .E(n822), .C(i_clk), .RN(n817), 
        .Q(regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(i_data_Rd[25]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(i_data_Rd[24]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(i_data_Rd[23]), .E(n822), .C(i_clk), .RN(n809), 
        .Q(regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(i_data_Rd[22]), .E(n822), .C(i_clk), .RN(n817), 
        .Q(regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(i_data_Rd[21]), .E(n822), .C(i_clk), .RN(n818), 
        .Q(regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(i_data_Rd[20]), .E(n822), .C(i_clk), .RN(n815), 
        .Q(regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(i_data_Rd[19]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(i_data_Rd[18]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(i_data_Rd[17]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(i_data_Rd[16]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(i_data_Rd[15]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(i_data_Rd[14]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(i_data_Rd[13]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(i_data_Rd[12]), .E(n822), .C(i_clk), .RN(n811), 
        .Q(regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(i_data_Rd[11]), .E(n822), .C(i_clk), .RN(n809), 
        .Q(regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(i_data_Rd[10]), .E(n822), .C(i_clk), .RN(i_rst_n), .Q(regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(i_data_Rd[9]), .E(n822), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(i_data_Rd[8]), .E(n822), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(i_data_Rd[7]), .E(n822), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(i_data_Rd[6]), .E(n822), .C(i_clk), .RN(n817), 
        .Q(regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(i_data_Rd[5]), .E(n822), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(i_data_Rd[4]), .E(n822), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(i_data_Rd[3]), .E(n822), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(i_data_Rd[2]), .E(n822), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(i_data_Rd[1]), .E(n822), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(i_data_Rd[0]), .E(n822), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(i_data_Rd[31]), .E(n823), .C(i_clk), .RN(n812), 
        .Q(regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(i_data_Rd[30]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(i_data_Rd[29]), .E(n823), .C(i_clk), .RN(n815), 
        .Q(regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(i_data_Rd[28]), .E(n823), .C(i_clk), .RN(n810), 
        .Q(regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(i_data_Rd[27]), .E(n823), .C(i_clk), .RN(n809), 
        .Q(regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(i_data_Rd[26]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(i_data_Rd[25]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(i_data_Rd[24]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(i_data_Rd[23]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(i_data_Rd[22]), .E(n823), .C(i_clk), .RN(n809), 
        .Q(regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(i_data_Rd[21]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(i_data_Rd[20]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(i_data_Rd[19]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(i_data_Rd[18]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(i_data_Rd[17]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(i_data_Rd[16]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(i_data_Rd[15]), .E(n823), .C(i_clk), .RN(n818), 
        .Q(regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(i_data_Rd[14]), .E(n823), .C(i_clk), .RN(n817), 
        .Q(regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(i_data_Rd[13]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(i_data_Rd[12]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(i_data_Rd[11]), .E(n823), .C(i_clk), .RN(i_rst_n), .Q(regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(i_data_Rd[10]), .E(n823), .C(i_clk), .RN(n812), 
        .Q(regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(i_data_Rd[9]), .E(n823), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(i_data_Rd[8]), .E(n823), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(i_data_Rd[7]), .E(n823), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(i_data_Rd[6]), .E(n823), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(i_data_Rd[5]), .E(n823), .C(i_clk), .RN(n813), 
        .Q(regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(i_data_Rd[4]), .E(n823), .C(i_clk), .RN(n814), 
        .Q(regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(i_data_Rd[3]), .E(n823), .C(i_clk), .RN(n815), 
        .Q(regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(i_data_Rd[2]), .E(n823), .C(i_clk), .RN(n816), 
        .Q(regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(i_data_Rd[1]), .E(n823), .C(i_clk), .RN(n809), 
        .Q(regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(i_data_Rd[0]), .E(n823), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[608]) );
  DFEC1 regs_reg_17__31_ ( .D(i_data_Rd[31]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(i_data_Rd[30]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(i_data_Rd[29]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(i_data_Rd[28]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(i_data_Rd[27]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(i_data_Rd[26]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(i_data_Rd[25]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(i_data_Rd[24]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(i_data_Rd[23]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(i_data_Rd[22]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(i_data_Rd[21]), .E(n825), .C(i_clk), .RN(n818), 
        .Q(regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(i_data_Rd[20]), .E(n825), .C(i_clk), .RN(n809), 
        .Q(regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(i_data_Rd[19]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(i_data_Rd[18]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(i_data_Rd[17]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(i_data_Rd[16]), .E(n825), .C(i_clk), .RN(n814), 
        .Q(regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(i_data_Rd[15]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(i_data_Rd[14]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(i_data_Rd[13]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(i_data_Rd[12]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(i_data_Rd[11]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(i_data_Rd[10]), .E(n825), .C(i_clk), .RN(i_rst_n), .Q(regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(i_data_Rd[9]), .E(n825), .C(i_clk), .RN(n814), 
        .Q(regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(i_data_Rd[8]), .E(n825), .C(i_clk), .RN(n813), 
        .Q(regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(i_data_Rd[7]), .E(n825), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(i_data_Rd[6]), .E(n825), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(i_data_Rd[5]), .E(n825), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(i_data_Rd[4]), .E(n825), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(i_data_Rd[3]), .E(n825), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(i_data_Rd[2]), .E(n825), .C(i_clk), .RN(n816), 
        .Q(regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(i_data_Rd[1]), .E(n825), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(i_data_Rd[0]), .E(n825), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(i_data_Rd[31]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(i_data_Rd[30]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(i_data_Rd[29]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(i_data_Rd[28]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(i_data_Rd[27]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(i_data_Rd[26]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(i_data_Rd[25]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(i_data_Rd[24]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(i_data_Rd[23]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(i_data_Rd[22]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(i_data_Rd[21]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(i_data_Rd[20]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(i_data_Rd[19]), .E(n826), .C(i_clk), .RN(n818), 
        .Q(regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(i_data_Rd[18]), .E(n826), .C(i_clk), .RN(n817), 
        .Q(regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(i_data_Rd[17]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(i_data_Rd[16]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(i_data_Rd[15]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(i_data_Rd[14]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(i_data_Rd[13]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(i_data_Rd[12]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(i_data_Rd[11]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(i_data_Rd[10]), .E(n826), .C(i_clk), .RN(i_rst_n), .Q(regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(i_data_Rd[9]), .E(n826), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(i_data_Rd[8]), .E(n826), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(i_data_Rd[7]), .E(n826), .C(i_clk), .RN(n813), 
        .Q(regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(i_data_Rd[6]), .E(n826), .C(i_clk), .RN(n814), 
        .Q(regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(i_data_Rd[5]), .E(n826), .C(i_clk), .RN(n815), 
        .Q(regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(i_data_Rd[4]), .E(n826), .C(i_clk), .RN(n816), 
        .Q(regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(i_data_Rd[3]), .E(n826), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(i_data_Rd[2]), .E(n826), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(i_data_Rd[1]), .E(n826), .C(i_clk), .RN(n817), 
        .Q(regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(i_data_Rd[0]), .E(n826), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[512]) );
  DFEC1 regs_reg_15__31_ ( .D(i_data_Rd[31]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(i_data_Rd[30]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(i_data_Rd[29]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(i_data_Rd[28]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(i_data_Rd[27]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(i_data_Rd[26]), .E(n836), .C(i_clk), .RN(n810), 
        .Q(regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(i_data_Rd[25]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(i_data_Rd[24]), .E(n836), .C(i_clk), .RN(n815), 
        .Q(regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(i_data_Rd[23]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(i_data_Rd[22]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(i_data_Rd[21]), .E(n836), .C(i_clk), .RN(n814), 
        .Q(regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(i_data_Rd[20]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(i_data_Rd[19]), .E(n836), .C(i_clk), .RN(n812), 
        .Q(regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(i_data_Rd[18]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(i_data_Rd[17]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(i_data_Rd[16]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(i_data_Rd[15]), .E(n836), .C(i_clk), .RN(n814), 
        .Q(regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(i_data_Rd[13]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(i_data_Rd[12]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(i_data_Rd[11]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n836), .C(i_clk), .RN(i_rst_n), .Q(regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(i_data_Rd[9]), .E(n836), .C(i_clk), .RN(n812), 
        .Q(regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(i_data_Rd[8]), .E(n836), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(i_data_Rd[7]), .E(n836), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(i_data_Rd[6]), .E(n836), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(i_data_Rd[5]), .E(n836), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(i_data_Rd[4]), .E(n836), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(i_data_Rd[3]), .E(n836), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(i_data_Rd[2]), .E(n836), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(i_data_Rd[1]), .E(n836), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(i_data_Rd[0]), .E(n836), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[480]) );
  DFEC1 regs_reg_13__31_ ( .D(i_data_Rd[31]), .E(n838), .C(i_clk), .RN(n815), 
        .Q(regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(i_data_Rd[30]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(i_data_Rd[29]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(i_data_Rd[28]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[444]) );
  DFEC1 regs_reg_13__27_ ( .D(i_data_Rd[27]), .E(n838), .C(i_clk), .RN(n810), 
        .Q(regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(i_data_Rd[26]), .E(n838), .C(i_clk), .RN(n811), 
        .Q(regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(i_data_Rd[25]), .E(n838), .C(i_clk), .RN(n812), 
        .Q(regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(i_data_Rd[24]), .E(n838), .C(i_clk), .RN(n813), 
        .Q(regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(i_data_Rd[23]), .E(n838), .C(i_clk), .RN(n814), 
        .Q(regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(i_data_Rd[22]), .E(n838), .C(i_clk), .RN(n813), 
        .Q(regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(i_data_Rd[21]), .E(n838), .C(i_clk), .RN(n811), 
        .Q(regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(i_data_Rd[20]), .E(n838), .C(i_clk), .RN(n816), 
        .Q(regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(i_data_Rd[19]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(i_data_Rd[18]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(i_data_Rd[17]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(i_data_Rd[16]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(i_data_Rd[15]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(i_data_Rd[13]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(i_data_Rd[12]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(i_data_Rd[11]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n838), .C(i_clk), .RN(i_rst_n), .Q(regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(i_data_Rd[9]), .E(n838), .C(i_clk), .RN(n818), 
        .Q(regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(i_data_Rd[8]), .E(n838), .C(i_clk), .RN(n817), 
        .Q(regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(i_data_Rd[7]), .E(n838), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(i_data_Rd[6]), .E(n838), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(i_data_Rd[5]), .E(n838), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(i_data_Rd[4]), .E(n838), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(i_data_Rd[3]), .E(n838), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(i_data_Rd[2]), .E(n838), .C(i_clk), .RN(n816), 
        .Q(regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(i_data_Rd[1]), .E(n838), .C(i_clk), .RN(n816), 
        .Q(regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(i_data_Rd[0]), .E(n838), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[416]) );
  DFEC1 regs_reg_12__31_ ( .D(i_data_Rd[31]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(i_data_Rd[30]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(i_data_Rd[29]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(i_data_Rd[28]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(i_data_Rd[27]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(i_data_Rd[26]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(i_data_Rd[25]), .E(n839), .C(i_clk), .RN(n816), 
        .Q(regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(i_data_Rd[24]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(i_data_Rd[23]), .E(n839), .C(i_clk), .RN(n815), 
        .Q(regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(i_data_Rd[22]), .E(n839), .C(i_clk), .RN(n813), 
        .Q(regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(i_data_Rd[21]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(i_data_Rd[20]), .E(n839), .C(i_clk), .RN(n812), 
        .Q(regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(i_data_Rd[19]), .E(n839), .C(i_clk), .RN(n813), 
        .Q(regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(i_data_Rd[18]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(i_data_Rd[17]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(i_data_Rd[16]), .E(n839), .C(i_clk), .RN(n816), 
        .Q(regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(i_data_Rd[15]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(i_data_Rd[13]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(i_data_Rd[12]), .E(n839), .C(i_clk), .RN(n817), 
        .Q(regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(i_data_Rd[11]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n839), .C(i_clk), .RN(i_rst_n), .Q(regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(i_data_Rd[9]), .E(n839), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(i_data_Rd[8]), .E(n839), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(i_data_Rd[7]), .E(n839), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(i_data_Rd[6]), .E(n839), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(i_data_Rd[5]), .E(n839), .C(i_clk), .RN(n818), 
        .Q(regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(i_data_Rd[4]), .E(n839), .C(i_clk), .RN(n813), 
        .Q(regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(i_data_Rd[3]), .E(n839), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(i_data_Rd[2]), .E(n839), .C(i_clk), .RN(n817), 
        .Q(regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(i_data_Rd[1]), .E(n839), .C(i_clk), .RN(n810), 
        .Q(regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(i_data_Rd[0]), .E(n839), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[384]) );
  DFEC1 regs_reg_11__31_ ( .D(i_data_Rd[31]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(i_data_Rd[30]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(i_data_Rd[29]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(i_data_Rd[28]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(i_data_Rd[27]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(i_data_Rd[26]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(i_data_Rd[25]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(i_data_Rd[24]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(i_data_Rd[23]), .E(n840), .C(i_clk), .RN(n815), 
        .Q(regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(i_data_Rd[22]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(i_data_Rd[21]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(i_data_Rd[20]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(i_data_Rd[19]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(i_data_Rd[18]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(i_data_Rd[17]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(i_data_Rd[16]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(i_data_Rd[15]), .E(n840), .C(i_clk), .RN(n809), 
        .Q(regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(i_data_Rd[13]), .E(n840), .C(i_clk), .RN(n810), 
        .Q(regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(i_data_Rd[12]), .E(n840), .C(i_clk), .RN(n818), 
        .Q(regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(i_data_Rd[11]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(i_data_Rd[10]), .E(n840), .C(i_clk), .RN(i_rst_n), .Q(regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(i_data_Rd[9]), .E(n840), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(i_data_Rd[8]), .E(n840), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(i_data_Rd[7]), .E(n840), .C(i_clk), .RN(n811), 
        .Q(regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(i_data_Rd[6]), .E(n840), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(i_data_Rd[5]), .E(n840), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(i_data_Rd[4]), .E(n840), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(i_data_Rd[3]), .E(n840), .C(i_clk), .RN(n814), 
        .Q(regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(i_data_Rd[2]), .E(n840), .C(i_clk), .RN(n812), 
        .Q(regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(i_data_Rd[1]), .E(n840), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(i_data_Rd[0]), .E(n840), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[352]) );
  DFEC1 regs_reg_9__31_ ( .D(i_data_Rd[31]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(i_data_Rd[30]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(i_data_Rd[29]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(i_data_Rd[28]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(i_data_Rd[27]), .E(n842), .C(i_clk), .RN(n809), 
        .Q(regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(i_data_Rd[26]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(i_data_Rd[25]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(i_data_Rd[24]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(i_data_Rd[23]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(i_data_Rd[22]), .E(n842), .C(i_clk), .RN(n812), 
        .Q(regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(i_data_Rd[21]), .E(n842), .C(i_clk), .RN(n810), 
        .Q(regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(i_data_Rd[20]), .E(n842), .C(i_clk), .RN(n811), 
        .Q(regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(i_data_Rd[19]), .E(n842), .C(i_clk), .RN(n809), 
        .Q(regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(i_data_Rd[18]), .E(n842), .C(i_clk), .RN(n810), 
        .Q(regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(i_data_Rd[17]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(i_data_Rd[16]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(i_data_Rd[15]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(i_data_Rd[14]), .E(n842), .C(i_clk), .RN(n816), 
        .Q(regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(i_data_Rd[13]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(i_data_Rd[12]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(i_data_Rd[11]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(i_data_Rd[10]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(i_data_Rd[9]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(i_data_Rd[8]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(i_data_Rd[7]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(i_data_Rd[6]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(i_data_Rd[5]), .E(n842), .C(i_clk), .RN(n816), .Q(
        regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(i_data_Rd[4]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(i_data_Rd[3]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(i_data_Rd[2]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(i_data_Rd[1]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(i_data_Rd[0]), .E(n842), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[288]) );
  DFEC1 regs_reg_8__31_ ( .D(i_data_Rd[31]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(i_data_Rd[30]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(i_data_Rd[29]), .E(n843), .C(i_clk), .RN(n810), 
        .Q(regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(i_data_Rd[28]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(i_data_Rd[27]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(i_data_Rd[26]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(i_data_Rd[25]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(i_data_Rd[24]), .E(n843), .C(i_clk), .RN(n814), 
        .Q(regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(i_data_Rd[23]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(i_data_Rd[22]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(i_data_Rd[21]), .E(n843), .C(i_clk), .RN(n809), 
        .Q(regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(i_data_Rd[20]), .E(n843), .C(i_clk), .RN(n809), 
        .Q(regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(i_data_Rd[19]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(i_data_Rd[18]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(i_data_Rd[17]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(i_data_Rd[16]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(i_data_Rd[15]), .E(n843), .C(i_clk), .RN(n809), 
        .Q(regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(i_data_Rd[14]), .E(n843), .C(i_clk), .RN(n811), 
        .Q(regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(i_data_Rd[13]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(i_data_Rd[12]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(i_data_Rd[11]), .E(n843), .C(i_clk), .RN(n818), 
        .Q(regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(i_data_Rd[10]), .E(n843), .C(i_clk), .RN(n814), 
        .Q(regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(i_data_Rd[9]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(i_data_Rd[8]), .E(n843), .C(i_clk), .RN(n810), .Q(
        regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(i_data_Rd[7]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(i_data_Rd[6]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(i_data_Rd[5]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(i_data_Rd[4]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(i_data_Rd[3]), .E(n843), .C(i_clk), .RN(n809), .Q(
        regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(i_data_Rd[2]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(i_data_Rd[1]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(i_data_Rd[0]), .E(n843), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[256]) );
  DFEC1 regs_reg_7__31_ ( .D(i_data_Rd[31]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(i_data_Rd[30]), .E(n844), .C(i_clk), .RN(n812), 
        .Q(regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(i_data_Rd[29]), .E(n844), .C(i_clk), .RN(n817), 
        .Q(regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(i_data_Rd[28]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(i_data_Rd[27]), .E(n844), .C(i_clk), .RN(n817), 
        .Q(regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(i_data_Rd[26]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(i_data_Rd[25]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(i_data_Rd[24]), .E(n844), .C(i_clk), .RN(n818), 
        .Q(regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(i_data_Rd[23]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(i_data_Rd[22]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(i_data_Rd[21]), .E(n844), .C(i_clk), .RN(n815), 
        .Q(regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(i_data_Rd[20]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(i_data_Rd[19]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(i_data_Rd[18]), .E(n844), .C(i_clk), .RN(n818), 
        .Q(regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(i_data_Rd[17]), .E(n844), .C(i_clk), .RN(n817), 
        .Q(regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(i_data_Rd[16]), .E(n844), .C(i_clk), .RN(n810), 
        .Q(regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(i_data_Rd[15]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(i_data_Rd[14]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(i_data_Rd[13]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(i_data_Rd[12]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(i_data_Rd[11]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(i_data_Rd[10]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(i_data_Rd[9]), .E(n844), .C(i_clk), .RN(n813), .Q(
        regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(i_data_Rd[8]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(i_data_Rd[7]), .E(n844), .C(i_clk), .RN(n816), .Q(
        regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(i_data_Rd[6]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(i_data_Rd[5]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(i_data_Rd[4]), .E(n844), .C(i_clk), .RN(n813), .Q(
        regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(i_data_Rd[3]), .E(n844), .C(i_clk), .RN(n818), .Q(
        regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(i_data_Rd[2]), .E(n844), .C(i_clk), .RN(n817), .Q(
        regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(i_data_Rd[1]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(i_data_Rd[0]), .E(n844), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[224]) );
  DFEC1 regs_reg_5__31_ ( .D(i_data_Rd[31]), .E(n846), .C(i_clk), .RN(n813), 
        .Q(regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(i_data_Rd[30]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(i_data_Rd[29]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(i_data_Rd[28]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[188]) );
  DFEC1 regs_reg_5__27_ ( .D(i_data_Rd[27]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(i_data_Rd[26]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(i_data_Rd[25]), .E(n846), .C(i_clk), .RN(n818), 
        .Q(regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(i_data_Rd[24]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(i_data_Rd[23]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(i_data_Rd[22]), .E(n846), .C(i_clk), .RN(n811), 
        .Q(regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(i_data_Rd[21]), .E(n846), .C(i_clk), .RN(n818), 
        .Q(regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(i_data_Rd[20]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(i_data_Rd[19]), .E(n846), .C(i_clk), .RN(n818), 
        .Q(regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(i_data_Rd[18]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(i_data_Rd[17]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(i_data_Rd[16]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(i_data_Rd[15]), .E(n846), .C(i_clk), .RN(n816), 
        .Q(regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(i_data_Rd[14]), .E(n846), .C(i_clk), .RN(n811), 
        .Q(regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(i_data_Rd[13]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(i_data_Rd[12]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(i_data_Rd[11]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(i_data_Rd[10]), .E(n846), .C(i_clk), .RN(n812), 
        .Q(regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(i_data_Rd[9]), .E(n846), .C(i_clk), .RN(n809), .Q(
        regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(i_data_Rd[8]), .E(n846), .C(i_clk), .RN(n817), .Q(
        regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(i_data_Rd[7]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(i_data_Rd[6]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(i_data_Rd[5]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(i_data_Rd[4]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(i_data_Rd[3]), .E(n846), .C(i_clk), .RN(n815), .Q(
        regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(i_data_Rd[2]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(i_data_Rd[1]), .E(n846), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(i_data_Rd[0]), .E(n846), .C(i_clk), .RN(n813), .Q(
        regs[160]) );
  DFEC1 regs_reg_4__31_ ( .D(i_data_Rd[31]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(i_data_Rd[30]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(i_data_Rd[29]), .E(n847), .C(i_clk), .RN(n815), 
        .Q(regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(i_data_Rd[28]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(i_data_Rd[27]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(i_data_Rd[26]), .E(n847), .C(i_clk), .RN(n813), 
        .Q(regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(i_data_Rd[25]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(i_data_Rd[24]), .E(n847), .C(i_clk), .RN(n809), 
        .Q(regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(i_data_Rd[23]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(i_data_Rd[22]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(i_data_Rd[21]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(i_data_Rd[20]), .E(n847), .C(i_clk), .RN(n814), 
        .Q(regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(i_data_Rd[19]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(i_data_Rd[18]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(i_data_Rd[17]), .E(n847), .C(i_clk), .RN(n811), 
        .Q(regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(i_data_Rd[16]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(i_data_Rd[15]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(i_data_Rd[14]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(i_data_Rd[13]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(i_data_Rd[12]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(i_data_Rd[11]), .E(n847), .C(i_clk), .RN(n818), 
        .Q(regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(i_data_Rd[10]), .E(n847), .C(i_clk), .RN(n817), 
        .Q(regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(i_data_Rd[9]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(i_data_Rd[8]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(i_data_Rd[7]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(i_data_Rd[6]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(i_data_Rd[5]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(i_data_Rd[4]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(i_data_Rd[3]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(i_data_Rd[2]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(i_data_Rd[1]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(i_data_Rd[0]), .E(n847), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[128]) );
  DFEC1 regs_reg_3__31_ ( .D(i_data_Rd[31]), .E(n848), .C(i_clk), .RN(n810), 
        .Q(regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(i_data_Rd[30]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(i_data_Rd[29]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(i_data_Rd[28]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(i_data_Rd[27]), .E(n848), .C(i_clk), .RN(n816), 
        .Q(regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(i_data_Rd[26]), .E(n848), .C(i_clk), .RN(n811), 
        .Q(regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(i_data_Rd[25]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(i_data_Rd[24]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(i_data_Rd[23]), .E(n848), .C(i_clk), .RN(n812), 
        .Q(regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(i_data_Rd[22]), .E(n848), .C(i_clk), .RN(n810), 
        .Q(regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(i_data_Rd[21]), .E(n848), .C(i_clk), .RN(n814), 
        .Q(regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(i_data_Rd[20]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(i_data_Rd[19]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(i_data_Rd[18]), .E(n848), .C(i_clk), .RN(n817), 
        .Q(regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(i_data_Rd[17]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(i_data_Rd[16]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(i_data_Rd[15]), .E(n848), .C(i_clk), .RN(n809), 
        .Q(regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(i_data_Rd[14]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(i_data_Rd[13]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(i_data_Rd[12]), .E(n848), .C(i_clk), .RN(n817), 
        .Q(regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(i_data_Rd[11]), .E(n848), .C(i_clk), .RN(n814), 
        .Q(regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(i_data_Rd[10]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(i_data_Rd[9]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(i_data_Rd[8]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(i_data_Rd[7]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(i_data_Rd[6]), .E(n848), .C(i_clk), .RN(n810), .Q(
        regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(i_data_Rd[5]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(i_data_Rd[4]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(i_data_Rd[3]), .E(n848), .C(i_clk), .RN(n812), .Q(
        regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(i_data_Rd[2]), .E(n848), .C(i_clk), .RN(n818), .Q(
        regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(i_data_Rd[1]), .E(n848), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(i_data_Rd[0]), .E(n848), .C(i_clk), .RN(n809), .Q(
        regs[96]) );
  DFEC1 regs_reg_1__31_ ( .D(i_data_Rd[31]), .E(n850), .C(i_clk), .RN(n817), 
        .Q(regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(i_data_Rd[30]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(i_data_Rd[29]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(i_data_Rd[28]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(i_data_Rd[27]), .E(n850), .C(i_clk), .RN(n814), 
        .Q(regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(i_data_Rd[26]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(i_data_Rd[25]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(i_data_Rd[24]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(i_data_Rd[23]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(i_data_Rd[22]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(i_data_Rd[21]), .E(n850), .C(i_clk), .RN(n817), 
        .Q(regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(i_data_Rd[20]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(i_data_Rd[19]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(i_data_Rd[18]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(i_data_Rd[17]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(i_data_Rd[16]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(i_data_Rd[15]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(i_data_Rd[14]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(i_data_Rd[13]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(i_data_Rd[12]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(i_data_Rd[11]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(i_data_Rd[10]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(i_data_Rd[9]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(i_data_Rd[8]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(i_data_Rd[7]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(i_data_Rd[6]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(i_data_Rd[5]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(i_data_Rd[4]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(i_data_Rd[3]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(i_data_Rd[2]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(i_data_Rd[1]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(i_data_Rd[0]), .E(n850), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[32]) );
  DFEC1 regs_reg_0__31_ ( .D(i_data_Rd[31]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(i_data_Rd[30]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(i_data_Rd[29]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(i_data_Rd[28]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(i_data_Rd[27]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(i_data_Rd[26]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(i_data_Rd[25]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(i_data_Rd[24]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(i_data_Rd[23]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(i_data_Rd[22]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(i_data_Rd[21]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(i_data_Rd[20]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(i_data_Rd[19]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(i_data_Rd[18]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(i_data_Rd[17]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(i_data_Rd[16]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(i_data_Rd[15]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(i_data_Rd[14]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(i_data_Rd[13]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(i_data_Rd[12]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(i_data_Rd[11]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(i_data_Rd[10]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(i_data_Rd[9]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(i_data_Rd[8]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(i_data_Rd[7]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(i_data_Rd[6]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(i_data_Rd[5]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(i_data_Rd[4]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(i_data_Rd[3]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(i_data_Rd[2]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(i_data_Rd[1]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(i_data_Rd[0]), .E(n851), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[0]) );
  BUF2 U2 ( .A(i_addr_Rs[4]), .Q(n749) );
  BUF2 U3 ( .A(n809), .Q(n816) );
  BUF2 U4 ( .A(n817), .Q(n815) );
  BUF2 U5 ( .A(n817), .Q(n814) );
  BUF2 U6 ( .A(n817), .Q(n813) );
  BUF2 U7 ( .A(n818), .Q(n812) );
  BUF2 U8 ( .A(n818), .Q(n811) );
  BUF2 U9 ( .A(n818), .Q(n810) );
  BUF2 U10 ( .A(n809), .Q(n817) );
  BUF2 U11 ( .A(n816), .Q(n818) );
  BUF2 U12 ( .A(n806), .Q(n786) );
  BUF2 U13 ( .A(i_addr_Rs[0]), .Q(n787) );
  BUF2 U14 ( .A(n805), .Q(n788) );
  BUF2 U15 ( .A(n806), .Q(n789) );
  BUF2 U16 ( .A(n805), .Q(n790) );
  BUF2 U17 ( .A(n805), .Q(n791) );
  BUF2 U18 ( .A(n804), .Q(n792) );
  BUF2 U19 ( .A(n804), .Q(n793) );
  BUF2 U20 ( .A(n804), .Q(n794) );
  BUF2 U21 ( .A(n805), .Q(n795) );
  BUF2 U22 ( .A(n805), .Q(n796) );
  BUF2 U23 ( .A(n805), .Q(n797) );
  BUF2 U24 ( .A(n806), .Q(n798) );
  BUF2 U25 ( .A(n806), .Q(n799) );
  BUF2 U26 ( .A(n806), .Q(n800) );
  BUF2 U27 ( .A(n807), .Q(n801) );
  BUF2 U28 ( .A(n807), .Q(n802) );
  BUF2 U29 ( .A(n807), .Q(n803) );
  BUF2 U30 ( .A(n783), .Q(n766) );
  BUF2 U31 ( .A(n785), .Q(n767) );
  BUF2 U32 ( .A(n765), .Q(n768) );
  BUF2 U33 ( .A(n765), .Q(n769) );
  BUF2 U34 ( .A(n764), .Q(n770) );
  BUF2 U35 ( .A(n764), .Q(n771) );
  BUF2 U36 ( .A(n764), .Q(n772) );
  BUF2 U37 ( .A(n763), .Q(n773) );
  BUF2 U38 ( .A(n763), .Q(n774) );
  BUF2 U39 ( .A(n762), .Q(n775) );
  BUF2 U40 ( .A(n762), .Q(n776) );
  BUF2 U41 ( .A(n762), .Q(n777) );
  BUF2 U42 ( .A(n761), .Q(n778) );
  BUF2 U43 ( .A(n761), .Q(n779) );
  BUF2 U44 ( .A(n761), .Q(n780) );
  BUF2 U45 ( .A(n421), .Q(n408) );
  BUF2 U46 ( .A(n421), .Q(n409) );
  BUF2 U47 ( .A(n423), .Q(n410) );
  BUF2 U48 ( .A(n423), .Q(n411) );
  BUF2 U49 ( .A(n423), .Q(n412) );
  BUF2 U50 ( .A(n424), .Q(n413) );
  BUF2 U51 ( .A(n424), .Q(n414) );
  BUF2 U52 ( .A(n424), .Q(n415) );
  BUF2 U53 ( .A(n425), .Q(n416) );
  BUF2 U54 ( .A(n425), .Q(n417) );
  BUF2 U55 ( .A(n426), .Q(n418) );
  BUF2 U56 ( .A(n426), .Q(n419) );
  INV3 U57 ( .A(n47), .Q(n831) );
  NAND22 U58 ( .A(n48), .B(n42), .Q(n47) );
  BUF2 U59 ( .A(n406), .Q(n385) );
  BUF2 U60 ( .A(n382), .Q(n386) );
  BUF2 U61 ( .A(n405), .Q(n387) );
  BUF2 U62 ( .A(n384), .Q(n388) );
  BUF2 U63 ( .A(n384), .Q(n389) );
  BUF2 U64 ( .A(n384), .Q(n390) );
  BUF2 U65 ( .A(n383), .Q(n391) );
  BUF2 U66 ( .A(n383), .Q(n392) );
  BUF2 U67 ( .A(n382), .Q(n393) );
  BUF2 U68 ( .A(n382), .Q(n394) );
  BUF2 U69 ( .A(n382), .Q(n395) );
  BUF2 U70 ( .A(n381), .Q(n396) );
  BUF2 U71 ( .A(n381), .Q(n397) );
  BUF2 U72 ( .A(n381), .Q(n398) );
  BUF2 U73 ( .A(n380), .Q(n399) );
  BUF2 U74 ( .A(n380), .Q(n400) );
  BUF2 U75 ( .A(n380), .Q(n401) );
  BUF2 U76 ( .A(n379), .Q(n402) );
  BUF2 U77 ( .A(n379), .Q(n403) );
  BUF2 U78 ( .A(n379), .Q(n404) );
  BUF2 U79 ( .A(i_rst_n), .Q(n809) );
  BUF2 U80 ( .A(n760), .Q(n781) );
  BUF2 U81 ( .A(n760), .Q(n782) );
  BUF2 U82 ( .A(i_addr_Rs[0]), .Q(n804) );
  BUF2 U83 ( .A(i_addr_Rs[0]), .Q(n805) );
  BUF2 U84 ( .A(i_addr_Rs[0]), .Q(n806) );
  BUF2 U85 ( .A(i_addr_Rs[0]), .Q(n807) );
  BUF2 U86 ( .A(i_addr_Rs[0]), .Q(n808) );
  BUF2 U87 ( .A(n785), .Q(n765) );
  BUF2 U88 ( .A(n785), .Q(n764) );
  BUF2 U89 ( .A(n784), .Q(n763) );
  BUF2 U90 ( .A(n784), .Q(n762) );
  BUF2 U91 ( .A(n784), .Q(n761) );
  NOR31 U92 ( .A(n835), .B(n852), .C(n856), .Q(n42) );
  NOR31 U93 ( .A(n854), .B(n855), .C(n853), .Q(n48) );
  INV3 U94 ( .A(n39), .Q(n827) );
  NAND22 U95 ( .A(n42), .B(n57), .Q(n39) );
  INV3 U96 ( .A(n80), .Q(n830) );
  NAND22 U97 ( .A(n51), .B(n42), .Q(n80) );
  INV3 U98 ( .A(n81), .Q(n829) );
  NAND22 U99 ( .A(n53), .B(n42), .Q(n81) );
  INV3 U100 ( .A(n82), .Q(n828) );
  NAND22 U101 ( .A(n55), .B(n42), .Q(n82) );
  INV3 U102 ( .A(n40), .Q(n834) );
  NAND22 U103 ( .A(n41), .B(n42), .Q(n40) );
  INV3 U104 ( .A(n43), .Q(n833) );
  NAND22 U105 ( .A(n44), .B(n42), .Q(n43) );
  INV3 U106 ( .A(n45), .Q(n832) );
  NAND22 U107 ( .A(n46), .B(n42), .Q(n45) );
  INV3 U108 ( .A(n49), .Q(n851) );
  NAND22 U109 ( .A(n50), .B(n51), .Q(n49) );
  INV3 U110 ( .A(n56), .Q(n848) );
  NAND22 U111 ( .A(n50), .B(n57), .Q(n56) );
  INV3 U112 ( .A(n58), .Q(n847) );
  NAND22 U113 ( .A(n50), .B(n41), .Q(n58) );
  INV3 U114 ( .A(n59), .Q(n846) );
  NAND22 U115 ( .A(n50), .B(n44), .Q(n59) );
  INV3 U116 ( .A(n60), .Q(n845) );
  NAND22 U117 ( .A(n50), .B(n46), .Q(n60) );
  INV3 U118 ( .A(n61), .Q(n844) );
  NAND22 U119 ( .A(n50), .B(n48), .Q(n61) );
  INV3 U120 ( .A(n52), .Q(n850) );
  NAND22 U121 ( .A(n53), .B(n50), .Q(n52) );
  INV3 U122 ( .A(n54), .Q(n849) );
  NAND22 U123 ( .A(n55), .B(n50), .Q(n54) );
  INV3 U124 ( .A(n62), .Q(n843) );
  NAND22 U125 ( .A(n63), .B(n51), .Q(n62) );
  INV3 U126 ( .A(n64), .Q(n842) );
  NAND22 U127 ( .A(n63), .B(n53), .Q(n64) );
  INV3 U128 ( .A(n65), .Q(n841) );
  NAND22 U129 ( .A(n63), .B(n55), .Q(n65) );
  INV3 U130 ( .A(n66), .Q(n840) );
  NAND22 U131 ( .A(n63), .B(n57), .Q(n66) );
  INV3 U132 ( .A(n67), .Q(n839) );
  NAND22 U133 ( .A(n63), .B(n41), .Q(n67) );
  INV3 U134 ( .A(n68), .Q(n838) );
  NAND22 U135 ( .A(n63), .B(n44), .Q(n68) );
  INV3 U136 ( .A(n69), .Q(n837) );
  NAND22 U137 ( .A(n63), .B(n46), .Q(n69) );
  INV3 U138 ( .A(n70), .Q(n836) );
  NAND22 U139 ( .A(n63), .B(n48), .Q(n70) );
  INV3 U140 ( .A(n71), .Q(n826) );
  NAND22 U141 ( .A(n72), .B(n51), .Q(n71) );
  INV3 U142 ( .A(n73), .Q(n825) );
  NAND22 U143 ( .A(n72), .B(n53), .Q(n73) );
  INV3 U144 ( .A(n74), .Q(n824) );
  NAND22 U145 ( .A(n72), .B(n55), .Q(n74) );
  INV3 U146 ( .A(n75), .Q(n823) );
  NAND22 U147 ( .A(n72), .B(n57), .Q(n75) );
  INV3 U148 ( .A(n76), .Q(n822) );
  NAND22 U149 ( .A(n72), .B(n41), .Q(n76) );
  INV3 U150 ( .A(n77), .Q(n821) );
  NAND22 U151 ( .A(n72), .B(n44), .Q(n77) );
  INV3 U152 ( .A(n78), .Q(n820) );
  NAND22 U153 ( .A(n72), .B(n46), .Q(n78) );
  INV3 U154 ( .A(n79), .Q(n819) );
  NAND22 U155 ( .A(n72), .B(n48), .Q(n79) );
  BUF2 U156 ( .A(i_addr_Rt[0]), .Q(n420) );
  BUF2 U157 ( .A(i_addr_Rt[0]), .Q(n421) );
  BUF2 U158 ( .A(i_addr_Rt[0]), .Q(n422) );
  BUF2 U159 ( .A(i_addr_Rt[0]), .Q(n423) );
  BUF2 U160 ( .A(i_addr_Rt[0]), .Q(n424) );
  BUF2 U161 ( .A(i_addr_Rt[0]), .Q(n425) );
  BUF2 U162 ( .A(i_addr_Rt[0]), .Q(n426) );
  BUF2 U163 ( .A(i_addr_Rt[0]), .Q(n427) );
  BUF2 U164 ( .A(n407), .Q(n384) );
  BUF2 U165 ( .A(n407), .Q(n383) );
  BUF2 U166 ( .A(n407), .Q(n382) );
  BUF2 U167 ( .A(n406), .Q(n381) );
  BUF2 U168 ( .A(n406), .Q(n380) );
  BUF2 U169 ( .A(n406), .Q(n379) );
  IMUX40 U170 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n786), .S1(n784), .Q(n437) );
  IMUX40 U171 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n786), .S1(n783), .Q(n435) );
  IMUX40 U172 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n786), .S1(i_addr_Rs[1]), .Q(n434) );
  IMUX40 U173 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(n795), .S1(n767), .Q(n432) );
  IMUX40 U174 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(n796), .S1(n761), .Q(n430) );
  IMUX40 U175 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(n798), .S1(n763), .Q(n429) );
  IMUX40 U176 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n786), .S1(n764), .Q(n442) );
  IMUX40 U177 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n786), .S1(n763), .Q(n440) );
  IMUX40 U178 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n786), .S1(i_addr_Rs[1]), .Q(n439) );
  IMUX40 U179 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n786), .S1(n767), .Q(n447) );
  IMUX40 U180 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n786), .S1(n765), .Q(n445) );
  IMUX40 U181 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n786), .S1(n764), .Q(n444) );
  IMUX40 U182 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n787), .S1(n762), .Q(n452) );
  IMUX40 U183 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n787), .S1(n766), .Q(n450) );
  IMUX40 U184 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n787), .S1(n764), .Q(n449) );
  IMUX40 U185 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n787), .S1(n766), .Q(n457) );
  IMUX40 U186 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n787), .S1(n768), .Q(n455) );
  IMUX40 U187 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n787), .S1(n782), .Q(n454) );
  IMUX40 U188 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n787), .S1(n767), .Q(n462) );
  IMUX40 U189 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n787), .S1(n768), .Q(n460) );
  IMUX40 U190 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n787), .S1(n771), .Q(n459) );
  IMUX40 U191 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n788), .S1(n765), .Q(n467) );
  IMUX40 U192 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n788), .S1(n766), .Q(n465) );
  IMUX40 U193 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n788), .S1(n763), .Q(n472) );
  IMUX40 U194 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n788), .S1(i_addr_Rs[1]), .Q(n470) );
  IMUX40 U195 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n788), .S1(n764), .Q(n469) );
  IMUX40 U196 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n788), .S1(n761), .Q(n477) );
  IMUX40 U197 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n788), .S1(n762), .Q(n475) );
  IMUX40 U198 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n789), .S1(n762), .Q(n482) );
  IMUX40 U199 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n789), .S1(n766), .Q(n480) );
  IMUX40 U200 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n789), .S1(i_addr_Rs[1]), .Q(n479) );
  IMUX40 U201 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n789), .S1(n761), .Q(n487) );
  IMUX40 U202 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n789), .S1(n783), .Q(n485) );
  IMUX40 U203 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n789), .S1(n760), .Q(n492) );
  IMUX40 U204 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n789), .S1(n766), .Q(n490) );
  IMUX40 U205 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n789), .S1(n766), .Q(n489) );
  IMUX40 U206 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n790), .S1(n766), .Q(n497) );
  IMUX40 U207 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n790), .S1(n766), .Q(n495) );
  IMUX40 U208 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n790), .S1(n766), .Q(n502) );
  IMUX40 U209 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n790), .S1(n766), .Q(n500) );
  IMUX40 U210 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n790), .S1(n767), .Q(n499) );
  IMUX40 U211 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n790), .S1(n767), .Q(n507) );
  IMUX40 U212 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n790), .S1(n767), .Q(n505) );
  IMUX40 U213 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n791), .S1(n767), .Q(n512) );
  IMUX40 U214 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n791), .S1(n767), .Q(n510) );
  IMUX40 U215 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n791), .S1(n784), .Q(n509) );
  IMUX40 U216 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n791), .S1(n763), .Q(n517) );
  IMUX40 U217 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n791), .S1(n761), .Q(n515) );
  IMUX40 U218 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n791), .S1(n766), .Q(n522) );
  IMUX40 U219 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n791), .S1(n764), .Q(n520) );
  IMUX40 U220 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n791), .S1(n767), .Q(n519) );
  IMUX40 U221 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n792), .S1(i_addr_Rs[1]), .Q(n527) );
  IMUX40 U222 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n792), .S1(i_addr_Rs[1]), .Q(n525) );
  IMUX40 U223 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n792), .S1(n783), .Q(n532) );
  IMUX40 U224 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n792), .S1(n764), .Q(n530) );
  IMUX40 U225 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n792), .S1(n785), .Q(n529) );
  IMUX40 U226 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n792), .S1(n765), .Q(n537) );
  IMUX40 U227 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n792), .S1(n765), .Q(n535) );
  IMUX40 U228 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n793), .S1(n782), .Q(n542) );
  IMUX40 U229 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n793), .S1(n769), .Q(n540) );
  IMUX40 U230 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n793), .S1(n784), .Q(n539) );
  IMUX40 U231 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n793), .S1(n762), .Q(n547) );
  IMUX40 U232 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n793), .S1(n763), .Q(n545) );
  IMUX40 U233 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n793), .S1(i_addr_Rs[1]), .Q(n552) );
  IMUX40 U234 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n793), .S1(n765), .Q(n550) );
  IMUX40 U235 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n793), .S1(n763), .Q(n549) );
  IMUX40 U236 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n794), .S1(n767), .Q(n557) );
  IMUX40 U237 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n794), .S1(n762), .Q(n555) );
  IMUX40 U238 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n794), .S1(n769), .Q(n562) );
  IMUX40 U239 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n794), .S1(i_addr_Rs[1]), .Q(n560) );
  IMUX40 U240 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n794), .S1(n770), .Q(n559) );
  IMUX40 U241 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n794), .S1(i_addr_Rs[1]), .Q(n567) );
  IMUX40 U242 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n794), .S1(n772), .Q(n565) );
  IMUX40 U243 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n795), .S1(n768), .Q(n572) );
  IMUX40 U244 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n795), .S1(n768), .Q(n570) );
  IMUX40 U245 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n795), .S1(n768), .Q(n569) );
  IMUX40 U246 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n795), .S1(n768), .Q(n577) );
  IMUX40 U247 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n795), .S1(n768), .Q(n575) );
  IMUX40 U248 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n795), .S1(n768), .Q(n582) );
  IMUX40 U249 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n795), .S1(n769), .Q(n580) );
  IMUX40 U250 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n795), .S1(n769), .Q(n579) );
  IMUX40 U251 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n796), .S1(n769), .Q(n587) );
  IMUX40 U252 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n796), .S1(n769), .Q(n585) );
  IMUX40 U253 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n796), .S1(n769), .Q(n592) );
  IMUX40 U254 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n796), .S1(n769), .Q(n590) );
  IMUX40 U255 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n796), .S1(n770), .Q(n589) );
  IMUX40 U256 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n796), .S1(n770), .Q(n597) );
  IMUX40 U257 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n796), .S1(n770), .Q(n595) );
  IMUX40 U258 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n797), .S1(n770), .Q(n602) );
  IMUX40 U259 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n797), .S1(n770), .Q(n600) );
  IMUX40 U260 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n797), .S1(n771), .Q(n599) );
  IMUX40 U261 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n797), .S1(n771), .Q(n607) );
  IMUX40 U262 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n797), .S1(n771), .Q(n605) );
  IMUX40 U263 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n797), .S1(n771), .Q(n612) );
  IMUX40 U264 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n797), .S1(n771), .Q(n610) );
  IMUX40 U265 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n797), .S1(n771), .Q(n609) );
  IMUX40 U266 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n798), .S1(n772), .Q(n617) );
  IMUX40 U267 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n798), .S1(n772), .Q(n615) );
  IMUX40 U268 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n798), .S1(n772), .Q(n622) );
  IMUX40 U269 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n798), .S1(n772), .Q(n620) );
  IMUX40 U270 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n798), .S1(n772), .Q(n619) );
  IMUX40 U271 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n798), .S1(n772), .Q(n627) );
  IMUX40 U272 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n798), .S1(n773), .Q(n625) );
  IMUX40 U273 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n799), .S1(n773), .Q(n632) );
  IMUX40 U274 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n799), .S1(n773), .Q(n630) );
  IMUX40 U275 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n799), .S1(n773), .Q(n629) );
  IMUX40 U276 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n799), .S1(n773), .Q(n637) );
  IMUX40 U277 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n799), .S1(n773), .Q(n635) );
  IMUX40 U278 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n799), .S1(n772), .Q(n642) );
  IMUX40 U279 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n799), .S1(n776), .Q(n640) );
  IMUX40 U280 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n799), .S1(n770), .Q(n639) );
  IMUX40 U281 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n800), .S1(n779), .Q(n647) );
  IMUX40 U282 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n800), .S1(n762), .Q(n645) );
  IMUX40 U283 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n800), .S1(n774), .Q(n652) );
  IMUX40 U284 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n800), .S1(n774), .Q(n650) );
  IMUX40 U285 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n800), .S1(n774), .Q(n649) );
  IMUX40 U286 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n800), .S1(n774), .Q(n657) );
  IMUX40 U287 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n800), .S1(n774), .Q(n655) );
  IMUX40 U288 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n801), .S1(n775), .Q(n662) );
  IMUX40 U289 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n801), .S1(n775), .Q(n660) );
  IMUX40 U290 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n801), .S1(n775), .Q(n659) );
  IMUX40 U291 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n801), .S1(n775), .Q(n667) );
  IMUX40 U292 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n801), .S1(n775), .Q(n665) );
  IMUX40 U293 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n801), .S1(n775), .Q(n672) );
  IMUX40 U294 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n801), .S1(n776), .Q(n670) );
  IMUX40 U295 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n801), .S1(n776), .Q(n669) );
  IMUX40 U296 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n802), .S1(n776), .Q(n677) );
  IMUX40 U297 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n802), .S1(n776), .Q(n675) );
  IMUX40 U298 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n802), .S1(n776), .Q(n682) );
  IMUX40 U299 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n802), .S1(n776), .Q(n680) );
  IMUX40 U300 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n802), .S1(n777), .Q(n679) );
  IMUX40 U301 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n802), .S1(n777), .Q(n687) );
  IMUX40 U302 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n802), .S1(n777), .Q(n685) );
  IMUX40 U303 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n803), .S1(n777), .Q(n692) );
  IMUX40 U304 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n803), .S1(n777), .Q(n690) );
  IMUX40 U305 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n803), .S1(n778), .Q(n689) );
  IMUX40 U306 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n803), .S1(n778), .Q(n697) );
  IMUX40 U307 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n803), .S1(n778), .Q(n695) );
  IMUX40 U308 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n803), .S1(n778), .Q(n702) );
  IMUX40 U309 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n803), .S1(n778), .Q(n700) );
  IMUX40 U310 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n803), .S1(n778), .Q(n699) );
  IMUX40 U311 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n808), .S1(n779), .Q(n707) );
  IMUX40 U312 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n808), .S1(n779), .Q(n705) );
  IMUX40 U313 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n808), .S1(n779), .Q(n712) );
  IMUX40 U314 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n808), .S1(n779), .Q(n710) );
  IMUX40 U315 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n808), .S1(n779), .Q(n709) );
  IMUX40 U316 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n808), .S1(n779), .Q(n717) );
  IMUX40 U317 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n808), .S1(n780), .Q(n715) );
  IMUX40 U318 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n792), .S1(n780), .Q(n722) );
  IMUX40 U319 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n801), .S1(n780), .Q(n720) );
  IMUX40 U320 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n793), .S1(n780), .Q(n719) );
  IMUX40 U321 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n787), .S1(n780), .Q(n727) );
  IMUX40 U322 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n792), .S1(n780), .Q(n725) );
  IMUX40 U323 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n799), .S1(n781), .Q(n724) );
  IMUX40 U324 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n802), .S1(n781), .Q(n732) );
  IMUX40 U325 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n807), .S1(n781), .Q(n730) );
  IMUX40 U326 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n800), .S1(n781), .Q(n729) );
  IMUX40 U327 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n786), .S1(n782), .Q(n734) );
  IMUX40 U328 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n808), .S1(n781), .Q(n737) );
  IMUX40 U329 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n788), .S1(n781), .Q(n735) );
  IMUX40 U330 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n807), .S1(n782), .Q(n742) );
  IMUX40 U331 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n808), .S1(n782), .Q(n740) );
  IMUX40 U332 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n790), .S1(n782), .Q(n739) );
  IMUX40 U333 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n789), .S1(n782), .Q(n744) );
  IMUX40 U334 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n800), .S1(n782), .Q(n745) );
  IMUX40 U335 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n799), .S1(n782), .Q(n747) );
  IMUX40 U336 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n786), .S1(n761), .Q(n436) );
  IMUX40 U337 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(n794), .S1(n767), .Q(n431) );
  IMUX40 U338 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n786), .S1(n782), .Q(n441) );
  IMUX40 U339 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n787), .S1(n767), .Q(n451) );
  IMUX40 U340 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n787), .S1(n767), .Q(n461) );
  IMUX40 U341 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n788), .S1(n766), .Q(n466) );
  IMUX40 U342 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n788), .S1(n764), .Q(n471) );
  IMUX40 U343 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n788), .S1(n761), .Q(n476) );
  IMUX40 U344 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n789), .S1(n783), .Q(n481) );
  IMUX40 U345 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n789), .S1(n783), .Q(n486) );
  IMUX40 U346 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n789), .S1(n766), .Q(n491) );
  IMUX40 U347 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n790), .S1(n766), .Q(n496) );
  IMUX40 U348 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n790), .S1(n767), .Q(n501) );
  IMUX40 U349 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n790), .S1(n767), .Q(n506) );
  IMUX40 U350 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n791), .S1(n767), .Q(n511) );
  IMUX40 U351 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n791), .S1(n762), .Q(n516) );
  IMUX40 U352 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n791), .S1(n767), .Q(n521) );
  IMUX40 U353 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n792), .S1(i_addr_Rs[1]), .Q(n526) );
  IMUX40 U354 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n792), .S1(n760), .Q(n531) );
  IMUX40 U355 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n792), .S1(n768), .Q(n536) );
  IMUX40 U356 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n793), .S1(n761), .Q(n541) );
  IMUX40 U357 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n793), .S1(n769), .Q(n546) );
  IMUX40 U358 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n793), .S1(n768), .Q(n551) );
  IMUX40 U359 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n794), .S1(n781), .Q(n556) );
  IMUX40 U360 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n794), .S1(n781), .Q(n561) );
  IMUX40 U361 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n794), .S1(n781), .Q(n566) );
  IMUX40 U362 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n795), .S1(n768), .Q(n571) );
  IMUX40 U363 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n795), .S1(n768), .Q(n576) );
  IMUX40 U364 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n795), .S1(n769), .Q(n581) );
  IMUX40 U365 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n796), .S1(n769), .Q(n586) );
  IMUX40 U366 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n796), .S1(n770), .Q(n591) );
  IMUX40 U367 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n796), .S1(n770), .Q(n596) );
  IMUX40 U368 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n797), .S1(n770), .Q(n601) );
  IMUX40 U369 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n797), .S1(n771), .Q(n606) );
  IMUX40 U370 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n797), .S1(n771), .Q(n611) );
  IMUX40 U371 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n798), .S1(n772), .Q(n616) );
  IMUX40 U372 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n798), .S1(n772), .Q(n621) );
  IMUX40 U373 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n798), .S1(n773), .Q(n626) );
  IMUX40 U374 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n799), .S1(n773), .Q(n631) );
  IMUX40 U375 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n799), .S1(n774), .Q(n636) );
  IMUX40 U376 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n799), .S1(n775), .Q(n641) );
  IMUX40 U377 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n800), .S1(n777), .Q(n646) );
  IMUX40 U378 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n800), .S1(n774), .Q(n651) );
  IMUX40 U379 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n800), .S1(n774), .Q(n656) );
  IMUX40 U380 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n801), .S1(n775), .Q(n661) );
  IMUX40 U381 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n801), .S1(n775), .Q(n666) );
  IMUX40 U382 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n801), .S1(n776), .Q(n671) );
  IMUX40 U383 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n802), .S1(n776), .Q(n676) );
  IMUX40 U384 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n802), .S1(n777), .Q(n681) );
  IMUX40 U385 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n802), .S1(n777), .Q(n686) );
  IMUX40 U386 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n803), .S1(n777), .Q(n691) );
  IMUX40 U387 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n803), .S1(n778), .Q(n696) );
  IMUX40 U388 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n803), .S1(n778), .Q(n701) );
  IMUX40 U389 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n808), .S1(n779), .Q(n706) );
  IMUX40 U390 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n808), .S1(n779), .Q(n711) );
  IMUX40 U391 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n808), .S1(n780), .Q(n716) );
  IMUX40 U392 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n787), .S1(n780), .Q(n721) );
  IMUX40 U393 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n793), .S1(n781), .Q(n731) );
  IMUX40 U394 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n808), .S1(n782), .Q(n741) );
  BUF2 U395 ( .A(i_addr_Rs[3]), .Q(n751) );
  BUF2 U396 ( .A(i_addr_Rs[3]), .Q(n752) );
  BUF2 U397 ( .A(i_addr_Rs[3]), .Q(n753) );
  BUF2 U398 ( .A(i_addr_Rs[3]), .Q(n754) );
  MUX22 U399 ( .A(n433), .B(n428), .S(n748), .Q(o_data_Rs[0]) );
  IMUX40 U400 ( .A(n429), .B(n430), .C(n431), .D(n432), .S0(n750), .S1(n756), 
        .Q(n428) );
  IMUX40 U401 ( .A(n434), .B(n435), .C(n436), .D(n437), .S0(n750), .S1(n755), 
        .Q(n433) );
  MUX22 U402 ( .A(n443), .B(n438), .S(n748), .Q(o_data_Rs[1]) );
  IMUX40 U403 ( .A(n444), .B(n445), .C(n446), .D(n447), .S0(n750), .S1(n755), 
        .Q(n443) );
  IMUX40 U404 ( .A(n439), .B(n440), .C(n441), .D(n442), .S0(n750), .S1(n755), 
        .Q(n438) );
  IMUX40 U405 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n786), .S1(n767), .Q(n446) );
  MUX22 U406 ( .A(n453), .B(n448), .S(n748), .Q(o_data_Rs[2]) );
  IMUX40 U407 ( .A(n454), .B(n455), .C(n456), .D(n457), .S0(n751), .S1(n755), 
        .Q(n453) );
  IMUX40 U408 ( .A(n449), .B(n450), .C(n451), .D(n452), .S0(n751), .S1(n755), 
        .Q(n448) );
  IMUX40 U409 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n787), .S1(n767), .Q(n456) );
  MUX22 U410 ( .A(n463), .B(n458), .S(n748), .Q(o_data_Rs[3]) );
  IMUX40 U411 ( .A(n464), .B(n465), .C(n466), .D(n467), .S0(n751), .S1(n755), 
        .Q(n463) );
  IMUX40 U412 ( .A(n459), .B(n460), .C(n461), .D(n462), .S0(n751), .S1(n755), 
        .Q(n458) );
  IMUX40 U413 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n788), .S1(n766), .Q(n464) );
  MUX22 U414 ( .A(n473), .B(n468), .S(n748), .Q(o_data_Rs[4]) );
  IMUX40 U415 ( .A(n474), .B(n475), .C(n476), .D(n477), .S0(n751), .S1(n755), 
        .Q(n473) );
  IMUX40 U416 ( .A(n469), .B(n470), .C(n471), .D(n472), .S0(n751), .S1(n755), 
        .Q(n468) );
  IMUX40 U417 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n788), .S1(n763), .Q(n474) );
  MUX22 U418 ( .A(n483), .B(n478), .S(n748), .Q(o_data_Rs[5]) );
  IMUX40 U419 ( .A(n484), .B(n485), .C(n486), .D(n487), .S0(n751), .S1(
        i_addr_Rs[2]), .Q(n483) );
  IMUX40 U420 ( .A(n479), .B(n480), .C(n481), .D(n482), .S0(n751), .S1(
        i_addr_Rs[2]), .Q(n478) );
  IMUX40 U421 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n789), .S1(n762), .Q(n484) );
  MUX22 U422 ( .A(n493), .B(n488), .S(n749), .Q(o_data_Rs[6]) );
  IMUX40 U423 ( .A(n494), .B(n495), .C(n496), .D(n497), .S0(n751), .S1(
        i_addr_Rs[2]), .Q(n493) );
  IMUX40 U424 ( .A(n489), .B(n490), .C(n491), .D(n492), .S0(n751), .S1(n756), 
        .Q(n488) );
  IMUX40 U425 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n790), .S1(n766), .Q(n494) );
  MUX22 U426 ( .A(n503), .B(n498), .S(n749), .Q(o_data_Rs[7]) );
  IMUX40 U427 ( .A(n504), .B(n505), .C(n506), .D(n507), .S0(n751), .S1(
        i_addr_Rs[2]), .Q(n503) );
  IMUX40 U428 ( .A(n499), .B(n500), .C(n501), .D(n502), .S0(n751), .S1(
        i_addr_Rs[2]), .Q(n498) );
  IMUX40 U429 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n790), .S1(n767), .Q(n504) );
  MUX22 U430 ( .A(n513), .B(n508), .S(n749), .Q(o_data_Rs[8]) );
  IMUX40 U431 ( .A(n514), .B(n515), .C(n516), .D(n517), .S0(n752), .S1(
        i_addr_Rs[2]), .Q(n513) );
  IMUX40 U432 ( .A(n509), .B(n510), .C(n511), .D(n512), .S0(n752), .S1(
        i_addr_Rs[2]), .Q(n508) );
  IMUX40 U433 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n791), .S1(n766), .Q(n514) );
  MUX22 U434 ( .A(n523), .B(n518), .S(n749), .Q(o_data_Rs[9]) );
  IMUX40 U435 ( .A(n524), .B(n525), .C(n526), .D(n527), .S0(n752), .S1(n759), 
        .Q(n523) );
  IMUX40 U436 ( .A(n519), .B(n520), .C(n521), .D(n522), .S0(n752), .S1(
        i_addr_Rs[2]), .Q(n518) );
  IMUX40 U437 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n792), .S1(i_addr_Rs[1]), .Q(n524) );
  MUX22 U438 ( .A(n533), .B(n528), .S(n749), .Q(o_data_Rs[10]) );
  IMUX40 U439 ( .A(n534), .B(n535), .C(n536), .D(n537), .S0(n752), .S1(n757), 
        .Q(n533) );
  IMUX40 U440 ( .A(n529), .B(n530), .C(n531), .D(n532), .S0(n752), .S1(n755), 
        .Q(n528) );
  IMUX40 U441 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n792), .S1(n767), .Q(n534) );
  MUX22 U442 ( .A(n543), .B(n538), .S(n749), .Q(o_data_Rs[11]) );
  IMUX40 U443 ( .A(n544), .B(n545), .C(n546), .D(n547), .S0(n752), .S1(n758), 
        .Q(n543) );
  IMUX40 U444 ( .A(n539), .B(n540), .C(n541), .D(n542), .S0(n752), .S1(n756), 
        .Q(n538) );
  IMUX40 U445 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n793), .S1(n769), .Q(n544) );
  BUF2 U446 ( .A(i_addr_Rs[1]), .Q(n785) );
  BUF2 U447 ( .A(i_addr_Rs[1]), .Q(n784) );
  MUX22 U448 ( .A(n553), .B(n548), .S(n749), .Q(o_data_Rs[12]) );
  IMUX40 U449 ( .A(n554), .B(n555), .C(n556), .D(n557), .S0(n752), .S1(n758), 
        .Q(n553) );
  IMUX40 U450 ( .A(n549), .B(n550), .C(n551), .D(n552), .S0(n752), .S1(n759), 
        .Q(n548) );
  IMUX40 U451 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n794), .S1(n781), .Q(n554) );
  MUX22 U452 ( .A(n563), .B(n558), .S(n749), .Q(o_data_Rs[13]) );
  IMUX40 U453 ( .A(n564), .B(n565), .C(n566), .D(n567), .S0(n752), .S1(n755), 
        .Q(n563) );
  IMUX40 U454 ( .A(n559), .B(n560), .C(n561), .D(n562), .S0(n752), .S1(n757), 
        .Q(n558) );
  IMUX40 U455 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n794), .S1(n764), .Q(n564) );
  MUX22 U456 ( .A(n573), .B(n568), .S(n749), .Q(o_data_Rs[14]) );
  IMUX40 U457 ( .A(n574), .B(n575), .C(n576), .D(n577), .S0(n753), .S1(n756), 
        .Q(n573) );
  IMUX40 U458 ( .A(n569), .B(n570), .C(n571), .D(n572), .S0(n753), .S1(n756), 
        .Q(n568) );
  IMUX40 U459 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n795), .S1(n768), .Q(n574) );
  MUX22 U460 ( .A(n583), .B(n578), .S(n749), .Q(o_data_Rs[15]) );
  IMUX40 U461 ( .A(n584), .B(n585), .C(n586), .D(n587), .S0(n753), .S1(n756), 
        .Q(n583) );
  IMUX40 U462 ( .A(n579), .B(n580), .C(n581), .D(n582), .S0(n753), .S1(n756), 
        .Q(n578) );
  IMUX40 U463 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n796), .S1(n769), .Q(n584) );
  MUX22 U464 ( .A(n593), .B(n588), .S(n749), .Q(o_data_Rs[16]) );
  IMUX40 U465 ( .A(n594), .B(n595), .C(n596), .D(n597), .S0(n753), .S1(n756), 
        .Q(n593) );
  IMUX40 U466 ( .A(n589), .B(n590), .C(n591), .D(n592), .S0(n753), .S1(n756), 
        .Q(n588) );
  IMUX40 U467 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n796), .S1(n770), .Q(n594) );
  MUX22 U468 ( .A(n603), .B(n598), .S(n749), .Q(o_data_Rs[17]) );
  IMUX40 U469 ( .A(n604), .B(n605), .C(n606), .D(n607), .S0(n753), .S1(n756), 
        .Q(n603) );
  IMUX40 U470 ( .A(n599), .B(n600), .C(n601), .D(n602), .S0(n753), .S1(n756), 
        .Q(n598) );
  IMUX40 U471 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n797), .S1(n771), .Q(n604) );
  MUX22 U472 ( .A(n613), .B(n608), .S(n749), .Q(o_data_Rs[18]) );
  IMUX40 U473 ( .A(n614), .B(n615), .C(n616), .D(n617), .S0(n753), .S1(n757), 
        .Q(n613) );
  IMUX40 U474 ( .A(n609), .B(n610), .C(n611), .D(n612), .S0(n753), .S1(n756), 
        .Q(n608) );
  IMUX40 U475 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n798), .S1(n772), .Q(n614) );
  MUX22 U476 ( .A(n623), .B(n618), .S(n748), .Q(o_data_Rs[19]) );
  IMUX40 U477 ( .A(n624), .B(n625), .C(n626), .D(n627), .S0(n753), .S1(n757), 
        .Q(n623) );
  IMUX40 U478 ( .A(n619), .B(n620), .C(n621), .D(n622), .S0(n753), .S1(n757), 
        .Q(n618) );
  IMUX40 U479 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n798), .S1(n773), .Q(n624) );
  MUX22 U480 ( .A(n633), .B(n628), .S(n748), .Q(o_data_Rs[20]) );
  IMUX40 U481 ( .A(n634), .B(n635), .C(n636), .D(n637), .S0(n754), .S1(n757), 
        .Q(n633) );
  IMUX40 U482 ( .A(n629), .B(n630), .C(n631), .D(n632), .S0(n754), .S1(n757), 
        .Q(n628) );
  IMUX40 U483 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n799), .S1(n763), .Q(n634) );
  MUX22 U484 ( .A(n643), .B(n638), .S(n748), .Q(o_data_Rs[21]) );
  IMUX40 U485 ( .A(n644), .B(n645), .C(n646), .D(n647), .S0(n754), .S1(n757), 
        .Q(n643) );
  IMUX40 U486 ( .A(n639), .B(n640), .C(n641), .D(n642), .S0(n754), .S1(n757), 
        .Q(n638) );
  IMUX40 U487 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n800), .S1(n774), .Q(n644) );
  MUX22 U488 ( .A(n653), .B(n648), .S(n748), .Q(o_data_Rs[22]) );
  IMUX40 U489 ( .A(n654), .B(n655), .C(n656), .D(n657), .S0(n754), .S1(n757), 
        .Q(n653) );
  IMUX40 U490 ( .A(n649), .B(n650), .C(n651), .D(n652), .S0(n754), .S1(n757), 
        .Q(n648) );
  IMUX40 U491 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n800), .S1(n774), .Q(n654) );
  MUX22 U492 ( .A(n663), .B(n658), .S(n748), .Q(o_data_Rs[23]) );
  IMUX40 U493 ( .A(n664), .B(n665), .C(n666), .D(n667), .S0(n754), .S1(n758), 
        .Q(n663) );
  IMUX40 U494 ( .A(n659), .B(n660), .C(n661), .D(n662), .S0(n754), .S1(n758), 
        .Q(n658) );
  IMUX40 U495 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n801), .S1(n775), .Q(n664) );
  MUX22 U496 ( .A(n673), .B(n668), .S(i_addr_Rs[4]), .Q(o_data_Rs[24]) );
  IMUX40 U497 ( .A(n674), .B(n675), .C(n676), .D(n677), .S0(n754), .S1(n758), 
        .Q(n673) );
  IMUX40 U498 ( .A(n669), .B(n670), .C(n671), .D(n672), .S0(n754), .S1(n758), 
        .Q(n668) );
  IMUX40 U499 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n802), .S1(n776), .Q(n674) );
  MUX22 U500 ( .A(n683), .B(n678), .S(i_addr_Rs[4]), .Q(o_data_Rs[25]) );
  IMUX40 U501 ( .A(n684), .B(n685), .C(n686), .D(n687), .S0(n754), .S1(n758), 
        .Q(n683) );
  IMUX40 U502 ( .A(n679), .B(n680), .C(n681), .D(n682), .S0(n754), .S1(n758), 
        .Q(n678) );
  IMUX40 U503 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n802), .S1(n777), .Q(n684) );
  MUX22 U504 ( .A(n693), .B(n688), .S(i_addr_Rs[4]), .Q(o_data_Rs[26]) );
  IMUX40 U505 ( .A(n694), .B(n695), .C(n696), .D(n697), .S0(n754), .S1(n758), 
        .Q(n693) );
  IMUX40 U506 ( .A(n689), .B(n690), .C(n691), .D(n692), .S0(n750), .S1(n758), 
        .Q(n688) );
  IMUX40 U507 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n803), .S1(n778), .Q(n694) );
  MUX22 U508 ( .A(n703), .B(n698), .S(n748), .Q(o_data_Rs[27]) );
  IMUX40 U509 ( .A(n704), .B(n705), .C(n706), .D(n707), .S0(n750), .S1(n759), 
        .Q(n703) );
  IMUX40 U510 ( .A(n699), .B(n700), .C(n701), .D(n702), .S0(n750), .S1(n758), 
        .Q(n698) );
  IMUX40 U511 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n808), .S1(n779), .Q(n704) );
  MUX22 U512 ( .A(n713), .B(n708), .S(i_addr_Rs[4]), .Q(o_data_Rs[28]) );
  IMUX40 U513 ( .A(n714), .B(n715), .C(n716), .D(n717), .S0(i_addr_Rs[3]), 
        .S1(n759), .Q(n713) );
  IMUX40 U514 ( .A(n709), .B(n710), .C(n711), .D(n712), .S0(n750), .S1(n759), 
        .Q(n708) );
  IMUX40 U515 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n808), .S1(n780), .Q(n714) );
  MUX22 U516 ( .A(n723), .B(n718), .S(n748), .Q(o_data_Rs[29]) );
  IMUX40 U517 ( .A(n724), .B(n725), .C(n726), .D(n727), .S0(n753), .S1(n759), 
        .Q(n723) );
  IMUX40 U518 ( .A(n719), .B(n720), .C(n721), .D(n722), .S0(n750), .S1(n759), 
        .Q(n718) );
  IMUX40 U519 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n808), .S1(n781), .Q(n726) );
  MUX22 U520 ( .A(n733), .B(n728), .S(i_addr_Rs[4]), .Q(o_data_Rs[30]) );
  IMUX40 U521 ( .A(n734), .B(n735), .C(n736), .D(n737), .S0(i_addr_Rs[3]), 
        .S1(n759), .Q(n733) );
  IMUX40 U522 ( .A(n729), .B(n730), .C(n731), .D(n732), .S0(n750), .S1(n759), 
        .Q(n728) );
  IMUX40 U523 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n791), .S1(n781), .Q(n736) );
  MUX22 U524 ( .A(n743), .B(n738), .S(n748), .Q(o_data_Rs[31]) );
  IMUX40 U525 ( .A(n744), .B(n745), .C(n746), .D(n747), .S0(n750), .S1(n759), 
        .Q(n743) );
  IMUX40 U526 ( .A(n739), .B(n740), .C(n741), .D(n742), .S0(n750), .S1(n759), 
        .Q(n738) );
  IMUX40 U527 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n797), .S1(n782), .Q(n746) );
  BUF2 U528 ( .A(n783), .Q(n760) );
  BUF2 U529 ( .A(i_addr_Rs[1]), .Q(n783) );
  NOR31 U530 ( .A(i_addr_Rd[3]), .B(i_addr_Rd[4]), .C(n856), .Q(n50) );
  NOR31 U531 ( .A(n835), .B(i_addr_Rd[3]), .C(n856), .Q(n72) );
  NOR31 U532 ( .A(n852), .B(i_addr_Rd[4]), .C(n856), .Q(n63) );
  MUX22 U533 ( .A(n16), .B(n11), .S(n365), .Q(o_data_Rt[1]) );
  IMUX40 U534 ( .A(n17), .B(n18), .C(n19), .D(n20), .S0(n366), .S1(n371), .Q(
        n16) );
  IMUX40 U535 ( .A(n12), .B(n13), .C(n14), .D(n15), .S0(n366), .S1(n371), .Q(
        n11) );
  IMUX40 U536 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n408), .S1(n391), .Q(n17) );
  MUX22 U537 ( .A(n26), .B(n21), .S(n365), .Q(o_data_Rt[2]) );
  IMUX40 U538 ( .A(n27), .B(n28), .C(n29), .D(n30), .S0(n367), .S1(n371), .Q(
        n26) );
  IMUX40 U539 ( .A(n22), .B(n23), .C(n24), .D(n25), .S0(n367), .S1(n371), .Q(
        n21) );
  IMUX40 U540 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n409), .S1(n384), .Q(n27) );
  MUX22 U541 ( .A(n36), .B(n31), .S(n365), .Q(o_data_Rt[3]) );
  IMUX40 U542 ( .A(n37), .B(n38), .C(n83), .D(n84), .S0(n367), .S1(n371), .Q(
        n36) );
  IMUX40 U543 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(n367), .S1(n371), .Q(
        n31) );
  IMUX40 U544 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n423), .S1(n389), .Q(n37) );
  MUX22 U545 ( .A(n90), .B(n85), .S(n365), .Q(o_data_Rt[4]) );
  IMUX40 U546 ( .A(n91), .B(n92), .C(n93), .D(n94), .S0(n367), .S1(n371), .Q(
        n90) );
  IMUX40 U547 ( .A(n86), .B(n87), .C(n88), .D(n89), .S0(n367), .S1(n371), .Q(
        n85) );
  IMUX40 U548 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n424), .S1(n390), .Q(n91) );
  MUX22 U549 ( .A(n100), .B(n95), .S(n365), .Q(o_data_Rt[5]) );
  IMUX40 U550 ( .A(n101), .B(n102), .C(n103), .D(n104), .S0(n367), .S1(n372), 
        .Q(n100) );
  IMUX40 U551 ( .A(n96), .B(n97), .C(n98), .D(n99), .S0(n367), .S1(n372), .Q(
        n95) );
  IMUX40 U552 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n422), .S1(n405), .Q(n101) );
  MUX22 U553 ( .A(n110), .B(n105), .S(i_addr_Rt[4]), .Q(o_data_Rt[6]) );
  IMUX40 U554 ( .A(n111), .B(n112), .C(n113), .D(n114), .S0(n367), .S1(n372), 
        .Q(n110) );
  IMUX40 U555 ( .A(n106), .B(n107), .C(n108), .D(n109), .S0(n367), .S1(n372), 
        .Q(n105) );
  IMUX40 U556 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        i_addr_Rt[0]), .S1(n385), .Q(n111) );
  MUX22 U557 ( .A(n120), .B(n115), .S(i_addr_Rt[4]), .Q(o_data_Rt[7]) );
  IMUX40 U558 ( .A(n121), .B(n122), .C(n123), .D(n124), .S0(n367), .S1(n372), 
        .Q(n120) );
  IMUX40 U559 ( .A(n116), .B(n117), .C(n118), .D(n119), .S0(n367), .S1(n372), 
        .Q(n115) );
  IMUX40 U560 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        i_addr_Rt[0]), .S1(n386), .Q(n121) );
  MUX22 U561 ( .A(n130), .B(n125), .S(i_addr_Rt[4]), .Q(o_data_Rt[8]) );
  IMUX40 U562 ( .A(n131), .B(n132), .C(n133), .D(n134), .S0(n368), .S1(n372), 
        .Q(n130) );
  IMUX40 U563 ( .A(n126), .B(n127), .C(n128), .D(n129), .S0(n368), .S1(n372), 
        .Q(n125) );
  IMUX40 U564 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n425), .S1(n387), .Q(n131) );
  MUX22 U565 ( .A(n140), .B(n135), .S(i_addr_Rt[4]), .Q(o_data_Rt[9]) );
  IMUX40 U566 ( .A(n141), .B(n142), .C(n143), .D(n144), .S0(n368), .S1(n373), 
        .Q(n140) );
  IMUX40 U567 ( .A(n136), .B(n137), .C(n138), .D(n139), .S0(n368), .S1(n372), 
        .Q(n135) );
  IMUX40 U568 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n410), .S1(n388), .Q(n141) );
  MUX22 U569 ( .A(n150), .B(n145), .S(i_addr_Rt[4]), .Q(o_data_Rt[10]) );
  IMUX40 U570 ( .A(n151), .B(n152), .C(n153), .D(n154), .S0(n368), .S1(n373), 
        .Q(n150) );
  IMUX40 U571 ( .A(n146), .B(n147), .C(n148), .D(n149), .S0(n368), .S1(n373), 
        .Q(n145) );
  IMUX40 U572 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n410), .S1(n389), .Q(n151) );
  MUX22 U573 ( .A(n160), .B(n155), .S(i_addr_Rt[4]), .Q(o_data_Rt[11]) );
  IMUX40 U574 ( .A(n161), .B(n162), .C(n163), .D(n164), .S0(n368), .S1(n373), 
        .Q(n160) );
  IMUX40 U575 ( .A(n156), .B(n157), .C(n158), .D(n159), .S0(n368), .S1(n373), 
        .Q(n155) );
  IMUX40 U576 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n411), .S1(n390), .Q(n161) );
  MUX22 U577 ( .A(n170), .B(n165), .S(i_addr_Rt[4]), .Q(o_data_Rt[12]) );
  IMUX40 U578 ( .A(n171), .B(n172), .C(n173), .D(n174), .S0(n368), .S1(n373), 
        .Q(n170) );
  IMUX40 U579 ( .A(n166), .B(n167), .C(n168), .D(n169), .S0(n368), .S1(n373), 
        .Q(n165) );
  IMUX40 U580 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n412), .S1(n384), .Q(n171) );
  MUX22 U581 ( .A(n180), .B(n175), .S(i_addr_Rt[4]), .Q(o_data_Rt[13]) );
  IMUX40 U582 ( .A(n181), .B(n182), .C(n183), .D(n184), .S0(n368), .S1(n373), 
        .Q(n180) );
  IMUX40 U583 ( .A(n176), .B(n177), .C(n178), .D(n179), .S0(n368), .S1(n373), 
        .Q(n175) );
  IMUX40 U584 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n412), .S1(n407), .Q(n181) );
  MUX22 U585 ( .A(n190), .B(n185), .S(i_addr_Rt[4]), .Q(o_data_Rt[14]) );
  IMUX40 U586 ( .A(n191), .B(n192), .C(n193), .D(n194), .S0(n369), .S1(n374), 
        .Q(n190) );
  IMUX40 U587 ( .A(n186), .B(n187), .C(n188), .D(n189), .S0(n369), .S1(n374), 
        .Q(n185) );
  IMUX40 U588 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n413), .S1(n391), .Q(n191) );
  MUX22 U589 ( .A(n200), .B(n195), .S(i_addr_Rt[4]), .Q(o_data_Rt[15]) );
  IMUX40 U590 ( .A(n201), .B(n202), .C(n203), .D(n204), .S0(n369), .S1(n374), 
        .Q(n200) );
  IMUX40 U591 ( .A(n196), .B(n197), .C(n198), .D(n199), .S0(n369), .S1(n374), 
        .Q(n195) );
  IMUX40 U592 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n414), .S1(n392), .Q(n201) );
  MUX22 U593 ( .A(n210), .B(n205), .S(i_addr_Rt[4]), .Q(o_data_Rt[16]) );
  IMUX40 U594 ( .A(n211), .B(n212), .C(n213), .D(n214), .S0(n369), .S1(n374), 
        .Q(n210) );
  IMUX40 U595 ( .A(n206), .B(n207), .C(n208), .D(n209), .S0(n369), .S1(n374), 
        .Q(n205) );
  IMUX40 U596 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n414), .S1(n393), .Q(n211) );
  MUX22 U597 ( .A(n220), .B(n215), .S(i_addr_Rt[4]), .Q(o_data_Rt[17]) );
  IMUX40 U598 ( .A(n221), .B(n222), .C(n223), .D(n224), .S0(n369), .S1(n374), 
        .Q(n220) );
  IMUX40 U599 ( .A(n216), .B(n217), .C(n218), .D(n219), .S0(n369), .S1(n374), 
        .Q(n215) );
  IMUX40 U600 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n415), .S1(n394), .Q(n221) );
  MUX22 U601 ( .A(n230), .B(n225), .S(i_addr_Rt[4]), .Q(o_data_Rt[18]) );
  IMUX40 U602 ( .A(n231), .B(n232), .C(n233), .D(n234), .S0(n369), .S1(n375), 
        .Q(n230) );
  IMUX40 U603 ( .A(n226), .B(n227), .C(n228), .D(n229), .S0(n369), .S1(n374), 
        .Q(n225) );
  IMUX40 U604 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n416), .S1(n395), .Q(n231) );
  MUX22 U605 ( .A(n240), .B(n235), .S(n365), .Q(o_data_Rt[19]) );
  IMUX40 U606 ( .A(n241), .B(n242), .C(n243), .D(n244), .S0(n369), .S1(n375), 
        .Q(n240) );
  IMUX40 U607 ( .A(n236), .B(n237), .C(n238), .D(n239), .S0(n369), .S1(n375), 
        .Q(n235) );
  IMUX40 U608 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n416), .S1(n396), .Q(n241) );
  MUX22 U609 ( .A(n250), .B(n245), .S(n365), .Q(o_data_Rt[20]) );
  IMUX40 U610 ( .A(n251), .B(n252), .C(n253), .D(n254), .S0(n370), .S1(n375), 
        .Q(n250) );
  IMUX40 U611 ( .A(n246), .B(n247), .C(n248), .D(n249), .S0(n370), .S1(n375), 
        .Q(n245) );
  IMUX40 U612 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n417), .S1(n397), .Q(n251) );
  MUX22 U613 ( .A(n260), .B(n255), .S(n365), .Q(o_data_Rt[21]) );
  IMUX40 U614 ( .A(n261), .B(n262), .C(n263), .D(n264), .S0(n370), .S1(n375), 
        .Q(n260) );
  IMUX40 U615 ( .A(n256), .B(n257), .C(n258), .D(n259), .S0(n370), .S1(n375), 
        .Q(n255) );
  IMUX40 U616 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n421), .S1(n398), .Q(n261) );
  MUX22 U617 ( .A(n270), .B(n265), .S(n365), .Q(o_data_Rt[22]) );
  IMUX40 U618 ( .A(n271), .B(n272), .C(n273), .D(n274), .S0(n370), .S1(n375), 
        .Q(n270) );
  IMUX40 U619 ( .A(n266), .B(n267), .C(n268), .D(n269), .S0(n370), .S1(n375), 
        .Q(n265) );
  IMUX40 U620 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n422), .S1(n398), .Q(n271) );
  MUX22 U621 ( .A(n280), .B(n275), .S(n365), .Q(o_data_Rt[23]) );
  IMUX40 U622 ( .A(n281), .B(n282), .C(n283), .D(n284), .S0(n370), .S1(n376), 
        .Q(n280) );
  IMUX40 U623 ( .A(n276), .B(n277), .C(n278), .D(n279), .S0(n370), .S1(n376), 
        .Q(n275) );
  IMUX40 U624 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n418), .S1(n399), .Q(n281) );
  MUX22 U625 ( .A(n290), .B(n285), .S(n365), .Q(o_data_Rt[24]) );
  IMUX40 U626 ( .A(n291), .B(n292), .C(n293), .D(n294), .S0(n370), .S1(n376), 
        .Q(n290) );
  IMUX40 U627 ( .A(n286), .B(n287), .C(n288), .D(n289), .S0(n370), .S1(n376), 
        .Q(n285) );
  IMUX40 U628 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n419), .S1(n400), .Q(n291) );
  MUX22 U629 ( .A(n300), .B(n295), .S(n365), .Q(o_data_Rt[25]) );
  IMUX40 U630 ( .A(n301), .B(n302), .C(n303), .D(n304), .S0(n370), .S1(n376), 
        .Q(n300) );
  IMUX40 U631 ( .A(n296), .B(n297), .C(n298), .D(n299), .S0(n370), .S1(n376), 
        .Q(n295) );
  IMUX40 U632 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n419), .S1(n401), .Q(n301) );
  MUX22 U633 ( .A(n310), .B(n305), .S(i_addr_Rt[4]), .Q(o_data_Rt[26]) );
  IMUX40 U634 ( .A(n311), .B(n312), .C(n313), .D(n314), .S0(n366), .S1(n376), 
        .Q(n310) );
  IMUX40 U635 ( .A(n306), .B(n307), .C(n308), .D(n309), .S0(n366), .S1(n376), 
        .Q(n305) );
  IMUX40 U636 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n415), .S1(n402), .Q(n311) );
  MUX22 U637 ( .A(n320), .B(n315), .S(i_addr_Rt[4]), .Q(o_data_Rt[27]) );
  IMUX40 U638 ( .A(n321), .B(n322), .C(n323), .D(n324), .S0(n366), .S1(n377), 
        .Q(n320) );
  IMUX40 U639 ( .A(n316), .B(n317), .C(n318), .D(n319), .S0(n366), .S1(n376), 
        .Q(n315) );
  IMUX40 U640 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n427), .S1(n403), .Q(n321) );
  MUX22 U641 ( .A(n330), .B(n325), .S(i_addr_Rt[4]), .Q(o_data_Rt[28]) );
  IMUX40 U642 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(i_addr_Rt[3]), 
        .S1(n377), .Q(n330) );
  IMUX40 U643 ( .A(n326), .B(n327), .C(n328), .D(n329), .S0(n366), .S1(n377), 
        .Q(n325) );
  IMUX40 U644 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n427), .S1(n404), .Q(n331) );
  MUX22 U645 ( .A(n340), .B(n335), .S(i_addr_Rt[4]), .Q(o_data_Rt[29]) );
  IMUX40 U646 ( .A(n341), .B(n342), .C(n343), .D(n344), .S0(i_addr_Rt[3]), 
        .S1(n377), .Q(n340) );
  IMUX40 U647 ( .A(n336), .B(n337), .C(n338), .D(n339), .S0(n366), .S1(n377), 
        .Q(n335) );
  IMUX40 U648 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n413), .S1(n378), .Q(n341) );
  MUX22 U649 ( .A(n350), .B(n345), .S(i_addr_Rt[4]), .Q(o_data_Rt[30]) );
  IMUX40 U650 ( .A(n351), .B(n352), .C(n353), .D(n354), .S0(i_addr_Rt[3]), 
        .S1(n377), .Q(n350) );
  IMUX40 U651 ( .A(n346), .B(n347), .C(n348), .D(n349), .S0(n366), .S1(n377), 
        .Q(n345) );
  IMUX40 U652 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n420), .S1(i_addr_Rt[1]), .Q(n351) );
  MUX22 U653 ( .A(n360), .B(n355), .S(i_addr_Rt[4]), .Q(o_data_Rt[31]) );
  IMUX40 U654 ( .A(n361), .B(n362), .C(n363), .D(n364), .S0(i_addr_Rt[3]), 
        .S1(n377), .Q(n360) );
  IMUX40 U655 ( .A(n356), .B(n357), .C(n358), .D(n359), .S0(n366), .S1(n377), 
        .Q(n355) );
  IMUX40 U656 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n420), .S1(i_addr_Rt[1]), .Q(n361) );
  NOR31 U657 ( .A(n855), .B(i_addr_Rd[2]), .C(n854), .Q(n57) );
  NOR31 U658 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n853), .Q(n41) );
  NOR31 U659 ( .A(n855), .B(i_addr_Rd[1]), .C(n853), .Q(n44) );
  NOR31 U660 ( .A(n854), .B(i_addr_Rd[0]), .C(n853), .Q(n46) );
  NOR31 U661 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(i_addr_Rd[0]), .Q(n51)
         );
  NOR31 U662 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(n855), .Q(n53) );
  NOR31 U663 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[2]), .C(n854), .Q(n55) );
  IMUX40 U664 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n408), .S1(i_addr_Rt[1]), .Q(n10) );
  IMUX40 U665 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n408), .S1(i_addr_Rt[1]), .Q(n8) );
  IMUX40 U666 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n408), .S1(i_addr_Rt[1]), .Q(n7) );
  IMUX40 U667 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(n420), .S1(n380), .Q(n5) );
  IMUX40 U668 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(n417), .S1(n406), .Q(n3) );
  IMUX40 U669 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(n426), .S1(n393), .Q(n2) );
  IMUX40 U670 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n408), .S1(n382), .Q(n15) );
  IMUX40 U671 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n408), .S1(i_addr_Rt[1]), .Q(n13) );
  IMUX40 U672 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n408), .S1(i_addr_Rt[1]), .Q(n12) );
  IMUX40 U673 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n408), .S1(i_addr_Rt[1]), .Q(n20) );
  IMUX40 U674 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n408), .S1(n384), .Q(n18) );
  IMUX40 U675 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n409), .S1(n381), .Q(n25) );
  IMUX40 U676 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n409), .S1(n379), .Q(n23) );
  IMUX40 U677 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n409), .S1(i_addr_Rt[1]), .Q(n22) );
  IMUX40 U678 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n409), .S1(i_addr_Rt[1]), .Q(n30) );
  IMUX40 U679 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n409), .S1(n395), .Q(n28) );
  IMUX40 U680 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n409), .S1(n385), .Q(n35) );
  IMUX40 U681 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n409), .S1(n387), .Q(n33) );
  IMUX40 U682 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n409), .S1(n383), .Q(n32) );
  IMUX40 U683 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n420), .S1(n386), .Q(n84) );
  IMUX40 U684 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n409), .S1(n382), .Q(n38) );
  IMUX40 U685 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n422), .S1(n387), .Q(n89) );
  IMUX40 U686 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n423), .S1(n406), .Q(n87) );
  IMUX40 U687 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n427), .S1(n388), .Q(n86) );
  IMUX40 U688 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n426), .S1(n380), .Q(n94) );
  IMUX40 U689 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n425), .S1(i_addr_Rt[1]), .Q(n92) );
  IMUX40 U690 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n422), .S1(n385), .Q(n99) );
  IMUX40 U691 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n422), .S1(n405), .Q(n97) );
  IMUX40 U692 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n422), .S1(n392), .Q(n96) );
  IMUX40 U693 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n422), .S1(n405), .Q(n104) );
  IMUX40 U694 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n422), .S1(n391), .Q(n102) );
  IMUX40 U695 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n422), .S1(n378), .Q(n109) );
  IMUX40 U696 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n422), .S1(n385), .Q(n107) );
  IMUX40 U697 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n422), .S1(n385), .Q(n106) );
  IMUX40 U698 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n422), .S1(n385), .Q(n114) );
  IMUX40 U699 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n426), .S1(n385), .Q(n112) );
  IMUX40 U700 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n426), .S1(n385), .Q(n119) );
  IMUX40 U701 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n408), .S1(n385), .Q(n117) );
  IMUX40 U702 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n421), .S1(n386), .Q(n116) );
  IMUX40 U703 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n420), .S1(n386), .Q(n124) );
  IMUX40 U704 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n427), .S1(n386), .Q(n122) );
  IMUX40 U705 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n427), .S1(n386), .Q(n129) );
  IMUX40 U706 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n415), .S1(n386), .Q(n127) );
  IMUX40 U707 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n424), .S1(n387), .Q(n126) );
  IMUX40 U708 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n411), .S1(n387), .Q(n134) );
  IMUX40 U709 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n423), .S1(n387), .Q(n132) );
  IMUX40 U710 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n425), .S1(n387), .Q(n139) );
  IMUX40 U711 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n414), .S1(n387), .Q(n137) );
  IMUX40 U712 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n420), .S1(n387), .Q(n136) );
  IMUX40 U713 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n410), .S1(n388), .Q(n144) );
  IMUX40 U714 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n410), .S1(n388), .Q(n142) );
  IMUX40 U715 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n410), .S1(n388), .Q(n149) );
  IMUX40 U716 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n410), .S1(n388), .Q(n147) );
  IMUX40 U717 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n410), .S1(n388), .Q(n146) );
  IMUX40 U718 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n410), .S1(n388), .Q(n154) );
  IMUX40 U719 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n410), .S1(n389), .Q(n152) );
  IMUX40 U720 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n411), .S1(n389), .Q(n159) );
  IMUX40 U721 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n411), .S1(n389), .Q(n157) );
  IMUX40 U722 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n411), .S1(n389), .Q(n156) );
  IMUX40 U723 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n411), .S1(n389), .Q(n164) );
  IMUX40 U724 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n411), .S1(n389), .Q(n162) );
  IMUX40 U725 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n411), .S1(n390), .Q(n169) );
  IMUX40 U726 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n411), .S1(n390), .Q(n167) );
  IMUX40 U727 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n411), .S1(n390), .Q(n166) );
  IMUX40 U728 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n412), .S1(n390), .Q(n174) );
  IMUX40 U729 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n412), .S1(n390), .Q(n172) );
  IMUX40 U730 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n412), .S1(n378), .Q(n179) );
  IMUX40 U731 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n412), .S1(n378), .Q(n177) );
  IMUX40 U732 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n412), .S1(n405), .Q(n176) );
  IMUX40 U733 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n412), .S1(n379), .Q(n184) );
  IMUX40 U734 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n412), .S1(n382), .Q(n182) );
  IMUX40 U735 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n413), .S1(n391), .Q(n189) );
  IMUX40 U736 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n413), .S1(n391), .Q(n187) );
  IMUX40 U737 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n413), .S1(n391), .Q(n186) );
  IMUX40 U738 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n413), .S1(n391), .Q(n194) );
  IMUX40 U739 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n413), .S1(n391), .Q(n192) );
  IMUX40 U740 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n413), .S1(n391), .Q(n199) );
  IMUX40 U741 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n413), .S1(n392), .Q(n197) );
  IMUX40 U742 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n413), .S1(n392), .Q(n196) );
  IMUX40 U743 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n414), .S1(n392), .Q(n204) );
  IMUX40 U744 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n414), .S1(n392), .Q(n202) );
  IMUX40 U745 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n414), .S1(n392), .Q(n209) );
  IMUX40 U746 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n414), .S1(n392), .Q(n207) );
  IMUX40 U747 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n414), .S1(n393), .Q(n206) );
  IMUX40 U748 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n414), .S1(n393), .Q(n214) );
  IMUX40 U749 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n414), .S1(n393), .Q(n212) );
  IMUX40 U750 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n415), .S1(n393), .Q(n219) );
  IMUX40 U751 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n415), .S1(n393), .Q(n217) );
  IMUX40 U752 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n415), .S1(n394), .Q(n216) );
  IMUX40 U753 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n415), .S1(n394), .Q(n224) );
  IMUX40 U754 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n415), .S1(n394), .Q(n222) );
  IMUX40 U755 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n415), .S1(n394), .Q(n229) );
  IMUX40 U756 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n415), .S1(n394), .Q(n227) );
  IMUX40 U757 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n415), .S1(n394), .Q(n226) );
  IMUX40 U758 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n416), .S1(n395), .Q(n234) );
  IMUX40 U759 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n416), .S1(n395), .Q(n232) );
  IMUX40 U760 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n416), .S1(n395), .Q(n239) );
  IMUX40 U761 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n416), .S1(n395), .Q(n237) );
  IMUX40 U762 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n416), .S1(n395), .Q(n236) );
  IMUX40 U763 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n416), .S1(n395), .Q(n244) );
  IMUX40 U764 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n416), .S1(n396), .Q(n242) );
  IMUX40 U765 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n417), .S1(n396), .Q(n249) );
  IMUX40 U766 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n417), .S1(n396), .Q(n247) );
  IMUX40 U767 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n417), .S1(n396), .Q(n246) );
  IMUX40 U768 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n417), .S1(n396), .Q(n254) );
  IMUX40 U769 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n417), .S1(n396), .Q(n252) );
  IMUX40 U770 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n417), .S1(n397), .Q(n259) );
  IMUX40 U771 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n417), .S1(n397), .Q(n257) );
  IMUX40 U772 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n417), .S1(n397), .Q(n256) );
  IMUX40 U773 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n412), .S1(n397), .Q(n264) );
  IMUX40 U774 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n411), .S1(n397), .Q(n262) );
  IMUX40 U775 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n408), .S1(n398), .Q(n269) );
  IMUX40 U776 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n409), .S1(n398), .Q(n267) );
  IMUX40 U777 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n413), .S1(n398), .Q(n266) );
  IMUX40 U778 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n410), .S1(n398), .Q(n274) );
  IMUX40 U779 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n412), .S1(n398), .Q(n272) );
  IMUX40 U780 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n418), .S1(n399), .Q(n279) );
  IMUX40 U781 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n418), .S1(n399), .Q(n277) );
  IMUX40 U782 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n418), .S1(n399), .Q(n276) );
  IMUX40 U783 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n418), .S1(n399), .Q(n284) );
  IMUX40 U784 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n418), .S1(n399), .Q(n282) );
  IMUX40 U785 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n418), .S1(n399), .Q(n289) );
  IMUX40 U786 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n418), .S1(n400), .Q(n287) );
  IMUX40 U787 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n418), .S1(n400), .Q(n286) );
  IMUX40 U788 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n419), .S1(n400), .Q(n294) );
  IMUX40 U789 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n419), .S1(n400), .Q(n292) );
  IMUX40 U790 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n419), .S1(n400), .Q(n299) );
  IMUX40 U791 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n419), .S1(n400), .Q(n297) );
  IMUX40 U792 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n419), .S1(n401), .Q(n296) );
  IMUX40 U793 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n419), .S1(n401), .Q(n304) );
  IMUX40 U794 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n419), .S1(n401), .Q(n302) );
  IMUX40 U795 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n426), .S1(n401), .Q(n309) );
  IMUX40 U796 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n415), .S1(n401), .Q(n307) );
  IMUX40 U797 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n426), .S1(n402), .Q(n306) );
  IMUX40 U798 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n425), .S1(n402), .Q(n314) );
  IMUX40 U799 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n425), .S1(n402), .Q(n312) );
  IMUX40 U800 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n414), .S1(n402), .Q(n319) );
  IMUX40 U801 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n416), .S1(n402), .Q(n317) );
  IMUX40 U802 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n414), .S1(n402), .Q(n316) );
  IMUX40 U803 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n427), .S1(n403), .Q(n324) );
  IMUX40 U804 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n427), .S1(n403), .Q(n322) );
  IMUX40 U805 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n427), .S1(n403), .Q(n329) );
  IMUX40 U806 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n427), .S1(n403), .Q(n327) );
  IMUX40 U807 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n427), .S1(n403), .Q(n326) );
  IMUX40 U808 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n427), .S1(n403), .Q(n334) );
  IMUX40 U809 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n427), .S1(n404), .Q(n332) );
  IMUX40 U810 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n408), .S1(n404), .Q(n339) );
  IMUX40 U811 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n420), .S1(n404), .Q(n337) );
  IMUX40 U812 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n411), .S1(n404), .Q(n336) );
  IMUX40 U813 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n413), .S1(n404), .Q(n344) );
  IMUX40 U814 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n410), .S1(n404), .Q(n342) );
  IMUX40 U815 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n409), .S1(n378), .Q(n349) );
  IMUX40 U816 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n422), .S1(n378), .Q(n347) );
  IMUX40 U817 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n412), .S1(n378), .Q(n346) );
  IMUX40 U818 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n420), .S1(n378), .Q(n354) );
  IMUX40 U819 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n420), .S1(n378), .Q(n352) );
  IMUX40 U820 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n420), .S1(n384), .Q(n359) );
  IMUX40 U821 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n420), .S1(n383), .Q(n357) );
  IMUX40 U822 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n420), .S1(i_addr_Rt[1]), .Q(n356) );
  IMUX40 U823 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n420), .S1(i_addr_Rt[1]), .Q(n364) );
  IMUX40 U824 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n420), .S1(i_addr_Rt[1]), .Q(n362) );
  IMUX40 U825 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n408), .S1(i_addr_Rt[1]), .Q(n9) );
  IMUX40 U826 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(n420), .S1(n387), .Q(n4) );
  IMUX40 U827 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n408), .S1(n405), .Q(n14) );
  IMUX40 U828 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n408), .S1(n394), .Q(n19) );
  IMUX40 U829 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n409), .S1(n392), .Q(n24) );
  IMUX40 U830 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n409), .S1(n385), .Q(n29) );
  IMUX40 U831 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n409), .S1(n385), .Q(n34) );
  IMUX40 U832 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n413), .S1(n387), .Q(n83) );
  IMUX40 U833 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n422), .S1(n387), .Q(n88) );
  IMUX40 U834 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n424), .S1(n383), .Q(n93) );
  IMUX40 U835 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n422), .S1(n385), .Q(n98) );
  IMUX40 U836 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n422), .S1(n378), .Q(n103) );
  IMUX40 U837 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n422), .S1(n385), .Q(n108) );
  IMUX40 U838 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n427), .S1(n385), .Q(n113) );
  IMUX40 U839 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n422), .S1(n386), .Q(n118) );
  IMUX40 U840 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n421), .S1(n386), .Q(n123) );
  IMUX40 U841 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n420), .S1(n386), .Q(n128) );
  IMUX40 U842 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n410), .S1(n387), .Q(n133) );
  IMUX40 U843 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n427), .S1(n387), .Q(n138) );
  IMUX40 U844 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n410), .S1(n388), .Q(n143) );
  IMUX40 U845 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n410), .S1(n388), .Q(n148) );
  IMUX40 U846 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n410), .S1(n389), .Q(n153) );
  IMUX40 U847 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n411), .S1(n389), .Q(n158) );
  IMUX40 U848 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n411), .S1(n390), .Q(n163) );
  IMUX40 U849 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n411), .S1(n390), .Q(n168) );
  IMUX40 U850 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n412), .S1(n390), .Q(n173) );
  IMUX40 U851 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n412), .S1(n378), .Q(n178) );
  IMUX40 U852 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n412), .S1(n381), .Q(n183) );
  IMUX40 U853 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n413), .S1(n391), .Q(n188) );
  IMUX40 U854 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n413), .S1(n391), .Q(n193) );
  IMUX40 U855 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n413), .S1(n392), .Q(n198) );
  IMUX40 U856 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n414), .S1(n392), .Q(n203) );
  IMUX40 U857 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n414), .S1(n393), .Q(n208) );
  IMUX40 U858 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n414), .S1(n393), .Q(n213) );
  IMUX40 U859 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n415), .S1(n393), .Q(n218) );
  IMUX40 U860 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n415), .S1(n394), .Q(n223) );
  IMUX40 U861 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n415), .S1(n394), .Q(n228) );
  IMUX40 U862 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n416), .S1(n395), .Q(n233) );
  IMUX40 U863 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n416), .S1(n395), .Q(n238) );
  IMUX40 U864 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n416), .S1(n396), .Q(n243) );
  IMUX40 U865 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n417), .S1(n396), .Q(n248) );
  IMUX40 U866 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n417), .S1(n397), .Q(n253) );
  IMUX40 U867 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n417), .S1(n397), .Q(n258) );
  IMUX40 U868 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n422), .S1(n397), .Q(n263) );
  IMUX40 U869 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n420), .S1(n398), .Q(n268) );
  IMUX40 U870 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n422), .S1(n398), .Q(n273) );
  IMUX40 U871 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n418), .S1(n399), .Q(n278) );
  IMUX40 U872 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n418), .S1(n399), .Q(n283) );
  IMUX40 U873 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n418), .S1(n400), .Q(n288) );
  IMUX40 U874 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n419), .S1(n400), .Q(n293) );
  IMUX40 U875 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n419), .S1(n401), .Q(n298) );
  IMUX40 U876 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n419), .S1(n401), .Q(n303) );
  IMUX40 U877 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n418), .S1(n401), .Q(n308) );
  IMUX40 U878 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n417), .S1(n402), .Q(n313) );
  IMUX40 U879 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n419), .S1(n402), .Q(n318) );
  IMUX40 U880 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n427), .S1(n403), .Q(n323) );
  IMUX40 U881 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n427), .S1(n403), .Q(n328) );
  IMUX40 U882 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n427), .S1(n404), .Q(n333) );
  IMUX40 U883 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n427), .S1(n404), .Q(n338) );
  IMUX40 U884 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n415), .S1(n378), .Q(n343) );
  IMUX40 U885 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n427), .S1(n378), .Q(n348) );
  IMUX40 U886 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n420), .S1(n378), .Q(n353) );
  IMUX40 U887 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n420), .S1(n378), .Q(n358) );
  IMUX40 U888 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n420), .S1(n385), .Q(n363) );
  BUF2 U889 ( .A(i_addr_Rt[3]), .Q(n367) );
  BUF2 U890 ( .A(i_addr_Rt[3]), .Q(n368) );
  BUF2 U891 ( .A(i_addr_Rt[3]), .Q(n369) );
  BUF2 U892 ( .A(i_addr_Rt[3]), .Q(n370) );
  INV3 U893 ( .A(i_addr_Rd[0]), .Q(n855) );
  INV3 U894 ( .A(i_addr_Rd[1]), .Q(n854) );
  INV3 U895 ( .A(i_addr_Rd[2]), .Q(n853) );
  INV3 U896 ( .A(i_con_RegWr), .Q(n856) );
  BUF2 U897 ( .A(i_addr_Rs[4]), .Q(n748) );
  BUF2 U898 ( .A(i_addr_Rt[4]), .Q(n365) );
  BUF2 U899 ( .A(i_addr_Rt[2]), .Q(n371) );
  BUF2 U900 ( .A(i_addr_Rt[2]), .Q(n372) );
  BUF2 U901 ( .A(i_addr_Rt[2]), .Q(n373) );
  BUF2 U902 ( .A(i_addr_Rt[2]), .Q(n374) );
  BUF2 U903 ( .A(i_addr_Rt[2]), .Q(n375) );
  BUF2 U904 ( .A(i_addr_Rt[2]), .Q(n376) );
  BUF2 U905 ( .A(i_addr_Rt[2]), .Q(n377) );
  INV3 U906 ( .A(i_addr_Rd[4]), .Q(n835) );
  BUF2 U907 ( .A(i_addr_Rs[2]), .Q(n755) );
  BUF2 U908 ( .A(i_addr_Rs[2]), .Q(n756) );
  BUF2 U909 ( .A(i_addr_Rs[2]), .Q(n757) );
  BUF2 U910 ( .A(i_addr_Rs[2]), .Q(n758) );
  BUF2 U911 ( .A(i_addr_Rs[2]), .Q(n759) );
  INV3 U912 ( .A(i_addr_Rd[3]), .Q(n852) );
  BUF2 U913 ( .A(i_addr_Rt[3]), .Q(n366) );
  BUF2 U914 ( .A(i_addr_Rs[3]), .Q(n750) );
  BUF2 U915 ( .A(i_addr_Rt[1]), .Q(n407) );
  BUF2 U916 ( .A(i_addr_Rt[1]), .Q(n406) );
  BUF2 U917 ( .A(n405), .Q(n378) );
  BUF2 U918 ( .A(i_addr_Rt[1]), .Q(n405) );
  MUX22 U919 ( .A(n6), .B(n1), .S(n365), .Q(o_data_Rt[0]) );
  IMUX40 U920 ( .A(n2), .B(n3), .C(n4), .D(n5), .S0(n366), .S1(i_addr_Rt[2]), 
        .Q(n1) );
  IMUX40 U921 ( .A(n7), .B(n8), .C(n9), .D(n10), .S0(n366), .S1(n371), .Q(n6)
         );
endmodule


module D_shiftleft ( i_data_immE, o_data_immshiftl );
  input [15:0] i_data_immE;
  output [31:0] o_data_immshiftl;
  wire   n1;
  assign o_data_immshiftl[0] = o_data_immshiftl[1];
  assign o_data_immshiftl[24] = o_data_immshiftl[31];
  assign o_data_immshiftl[19] = o_data_immshiftl[31];
  assign o_data_immshiftl[25] = o_data_immshiftl[31];
  assign o_data_immshiftl[17] = o_data_immshiftl[31];
  assign o_data_immshiftl[21] = o_data_immshiftl[31];
  assign o_data_immshiftl[29] = o_data_immshiftl[31];
  assign o_data_immshiftl[20] = o_data_immshiftl[30];
  assign o_data_immshiftl[23] = o_data_immshiftl[30];
  assign o_data_immshiftl[27] = o_data_immshiftl[30];
  assign o_data_immshiftl[28] = o_data_immshiftl[30];
  assign o_data_immshiftl[26] = o_data_immshiftl[30];
  assign o_data_immshiftl[22] = o_data_immshiftl[30];
  assign o_data_immshiftl[18] = o_data_immshiftl[30];
  assign o_data_immshiftl[16] = i_data_immE[14];
  assign o_data_immshiftl[15] = i_data_immE[13];
  assign o_data_immshiftl[14] = i_data_immE[12];
  assign o_data_immshiftl[13] = i_data_immE[11];
  assign o_data_immshiftl[12] = i_data_immE[10];
  assign o_data_immshiftl[11] = i_data_immE[9];
  assign o_data_immshiftl[10] = i_data_immE[8];
  assign o_data_immshiftl[9] = i_data_immE[7];
  assign o_data_immshiftl[8] = i_data_immE[6];
  assign o_data_immshiftl[7] = i_data_immE[5];
  assign o_data_immshiftl[6] = i_data_immE[4];
  assign o_data_immshiftl[5] = i_data_immE[3];
  assign o_data_immshiftl[4] = i_data_immE[2];
  assign o_data_immshiftl[3] = i_data_immE[1];
  assign o_data_immshiftl[2] = i_data_immE[0];

  INV3 U2 ( .A(n1), .Q(o_data_immshiftl[30]) );
  INV3 U3 ( .A(n1), .Q(o_data_immshiftl[31]) );
  INV3 U4 ( .A(i_data_immE[15]), .Q(n1) );
  LOGIC0 U5 ( .Q(o_data_immshiftl[1]) );
endmodule


module D_sign_extend ( i_data_immD, i_con_signext, o_data_immD );
  input [15:0] i_data_immD;
  output [31:0] o_data_immD;
  input i_con_signext;
  wire   n2;
  assign o_data_immD[15] = i_data_immD[15];
  assign o_data_immD[14] = i_data_immD[14];
  assign o_data_immD[13] = i_data_immD[13];
  assign o_data_immD[12] = i_data_immD[12];
  assign o_data_immD[11] = i_data_immD[11];
  assign o_data_immD[10] = i_data_immD[10];
  assign o_data_immD[9] = i_data_immD[9];
  assign o_data_immD[8] = i_data_immD[8];
  assign o_data_immD[7] = i_data_immD[7];
  assign o_data_immD[6] = i_data_immD[6];
  assign o_data_immD[5] = i_data_immD[5];
  assign o_data_immD[4] = i_data_immD[4];
  assign o_data_immD[3] = i_data_immD[3];
  assign o_data_immD[2] = i_data_immD[2];
  assign o_data_immD[1] = i_data_immD[1];
  assign o_data_immD[0] = i_data_immD[0];
  assign o_data_immD[16] = o_data_immD[31];
  assign o_data_immD[17] = o_data_immD[31];
  assign o_data_immD[18] = o_data_immD[31];
  assign o_data_immD[19] = o_data_immD[31];
  assign o_data_immD[20] = o_data_immD[31];
  assign o_data_immD[21] = o_data_immD[31];
  assign o_data_immD[22] = o_data_immD[31];
  assign o_data_immD[23] = o_data_immD[31];
  assign o_data_immD[24] = o_data_immD[31];
  assign o_data_immD[25] = o_data_immD[31];
  assign o_data_immD[26] = o_data_immD[31];
  assign o_data_immD[27] = o_data_immD[31];
  assign o_data_immD[28] = o_data_immD[31];
  assign o_data_immD[29] = o_data_immD[31];
  assign o_data_immD[30] = o_data_immD[31];

  INV3 U2 ( .A(n2), .Q(o_data_immD[31]) );
  NAND22 U3 ( .A(i_con_signext), .B(i_data_immD[15]), .Q(n2) );
endmodule


module D_jump_ext ( i_addr_j, i_PC4_j, o_addr_j );
  input [25:0] i_addr_j;
  input [3:0] i_PC4_j;
  output [31:0] o_addr_j;

  assign o_addr_j[0] = o_addr_j[1];
  assign o_addr_j[31] = i_PC4_j[3];
  assign o_addr_j[30] = i_PC4_j[2];
  assign o_addr_j[29] = i_PC4_j[1];
  assign o_addr_j[28] = i_PC4_j[0];
  assign o_addr_j[27] = i_addr_j[25];
  assign o_addr_j[26] = i_addr_j[24];
  assign o_addr_j[25] = i_addr_j[23];
  assign o_addr_j[24] = i_addr_j[22];
  assign o_addr_j[23] = i_addr_j[21];
  assign o_addr_j[22] = i_addr_j[20];
  assign o_addr_j[21] = i_addr_j[19];
  assign o_addr_j[20] = i_addr_j[18];
  assign o_addr_j[19] = i_addr_j[17];
  assign o_addr_j[18] = i_addr_j[16];
  assign o_addr_j[17] = i_addr_j[15];
  assign o_addr_j[16] = i_addr_j[14];
  assign o_addr_j[15] = i_addr_j[13];
  assign o_addr_j[14] = i_addr_j[12];
  assign o_addr_j[13] = i_addr_j[11];
  assign o_addr_j[12] = i_addr_j[10];
  assign o_addr_j[11] = i_addr_j[9];
  assign o_addr_j[10] = i_addr_j[8];
  assign o_addr_j[9] = i_addr_j[7];
  assign o_addr_j[8] = i_addr_j[6];
  assign o_addr_j[7] = i_addr_j[5];
  assign o_addr_j[6] = i_addr_j[4];
  assign o_addr_j[5] = i_addr_j[3];
  assign o_addr_j[4] = i_addr_j[2];
  assign o_addr_j[3] = i_addr_j[1];
  assign o_addr_j[2] = i_addr_j[0];

  LOGIC0 U2 ( .Q(o_addr_j[1]) );
endmodule


module D_forward ( i_addr_rs, i_addr_rt, i_addr_rdE, i_addr_rdM, i_addr_rtM, 
        i_addr_rtW, i_con_regwriteE, i_con_regwriteM, i_con_memreadM, 
        i_con_memreadW, o_con_fa, o_con_fb );
  input [4:0] i_addr_rs;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rdE;
  input [4:0] i_addr_rdM;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  output [2:0] o_con_fa;
  output [2:0] o_con_fb;
  input i_con_regwriteE, i_con_regwriteM, i_con_memreadM, i_con_memreadW;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;

  XNR21 U1 ( .A(i_addr_rt[4]), .B(i_addr_rtM[4]), .Q(n39) );
  CLKIN1 U2 ( .A(i_addr_rdE[3]), .Q(n28) );
  NAND41 U3 ( .A(n55), .B(i_con_regwriteE), .C(n56), .D(n57), .Q(n46) );
  NOR31 U4 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  OAI310 U5 ( .A(n1), .B(n2), .C(n3), .D(n4), .Q(o_con_fb[2]) );
  NOR40 U6 ( .A(n5), .B(n6), .C(n7), .D(n8), .Q(o_con_fb[1]) );
  CLKIN0 U7 ( .A(n9), .Q(n6) );
  NAND20 U8 ( .A(n4), .B(n10), .Q(o_con_fb[0]) );
  NAND40 U9 ( .A(n11), .B(i_con_regwriteM), .C(n12), .D(n13), .Q(n10) );
  NOR40 U10 ( .A(n14), .B(n15), .C(n16), .D(n17), .Q(n13) );
  XOR20 U11 ( .A(i_addr_rdM[4]), .B(i_addr_rt[4]), .Q(n17) );
  XNR20 U12 ( .A(n18), .B(i_addr_rt[2]), .Q(n16) );
  XNR20 U13 ( .A(n19), .B(i_addr_rt[1]), .Q(n15) );
  XNR20 U14 ( .A(n20), .B(i_addr_rt[0]), .Q(n14) );
  CLKIN0 U15 ( .A(n21), .Q(n12) );
  OAI210 U16 ( .A(n8), .B(n7), .C(n9), .Q(n21) );
  NAND40 U17 ( .A(n22), .B(n23), .C(n24), .D(n25), .Q(n7) );
  XNR20 U18 ( .A(i_addr_rt[0]), .B(i_addr_rdE[0]), .Q(n25) );
  NOR20 U19 ( .A(n26), .B(n27), .Q(n24) );
  XNR20 U20 ( .A(n28), .B(i_addr_rt[3]), .Q(n27) );
  XOR20 U21 ( .A(i_addr_rdE[1]), .B(i_addr_rt[1]), .Q(n26) );
  XNR20 U22 ( .A(i_addr_rt[2]), .B(i_addr_rdE[2]), .Q(n23) );
  XNR20 U23 ( .A(i_addr_rt[4]), .B(i_addr_rdE[4]), .Q(n22) );
  CLKIN0 U24 ( .A(i_con_regwriteE), .Q(n8) );
  XNR20 U25 ( .A(i_addr_rt[3]), .B(i_addr_rdM[3]), .Q(n11) );
  NAND20 U26 ( .A(n9), .B(n5), .Q(n4) );
  CLKIN0 U27 ( .A(n29), .Q(n5) );
  NAND40 U28 ( .A(n30), .B(i_con_memreadW), .C(n31), .D(n32), .Q(n29) );
  NOR30 U29 ( .A(n33), .B(n34), .C(n35), .Q(n32) );
  XOR20 U30 ( .A(i_addr_rtW[2]), .B(i_addr_rt[2]), .Q(n35) );
  XOR20 U31 ( .A(i_addr_rtW[4]), .B(i_addr_rt[4]), .Q(n34) );
  XOR20 U32 ( .A(i_addr_rtW[3]), .B(i_addr_rt[3]), .Q(n33) );
  XNR20 U33 ( .A(i_addr_rt[0]), .B(i_addr_rtW[0]), .Q(n31) );
  XNR20 U34 ( .A(i_addr_rt[1]), .B(i_addr_rtW[1]), .Q(n30) );
  AOI210 U35 ( .A(n36), .B(i_con_memreadM), .C(n2), .Q(n9) );
  NOR30 U36 ( .A(i_addr_rt[0]), .B(i_addr_rt[1]), .C(n37), .Q(n2) );
  CLKIN0 U37 ( .A(n38), .Q(n37) );
  NOR30 U38 ( .A(i_addr_rt[2]), .B(i_addr_rt[4]), .C(i_addr_rt[3]), .Q(n38) );
  CLKIN0 U39 ( .A(n3), .Q(n36) );
  NAND40 U40 ( .A(n39), .B(n40), .C(n41), .D(n42), .Q(n3) );
  XNR20 U41 ( .A(i_addr_rt[0]), .B(i_addr_rtM[0]), .Q(n42) );
  NOR20 U42 ( .A(n43), .B(n44), .Q(n41) );
  XOR20 U43 ( .A(i_addr_rtM[3]), .B(i_addr_rt[3]), .Q(n44) );
  XNR20 U44 ( .A(n45), .B(i_addr_rt[1]), .Q(n43) );
  XNR20 U45 ( .A(i_addr_rt[2]), .B(i_addr_rtM[2]), .Q(n40) );
  NOR20 U46 ( .A(o_con_fa[2]), .B(n46), .Q(o_con_fa[1]) );
  OAI210 U47 ( .A(n47), .B(n48), .C(n49), .Q(o_con_fa[0]) );
  NAND20 U48 ( .A(n50), .B(n51), .Q(n49) );
  NOR40 U49 ( .A(o_con_fa[2]), .B(n52), .C(n53), .D(n54), .Q(n51) );
  XNR20 U50 ( .A(n20), .B(i_addr_rs[0]), .Q(n54) );
  CLKIN0 U51 ( .A(i_addr_rdM[0]), .Q(n20) );
  CLKIN0 U52 ( .A(i_con_regwriteM), .Q(n53) );
  CLKIN0 U53 ( .A(n46), .Q(n52) );
  XNR20 U54 ( .A(n28), .B(i_addr_rs[3]), .Q(n60) );
  XOR20 U55 ( .A(i_addr_rdE[2]), .B(i_addr_rs[2]), .Q(n59) );
  IMUX20 U56 ( .A(n61), .B(i_addr_rs[4]), .S(i_addr_rdE[4]), .Q(n58) );
  NOR20 U57 ( .A(n62), .B(i_addr_rs[4]), .Q(n61) );
  NOR40 U58 ( .A(i_addr_rdE[3]), .B(i_addr_rdE[2]), .C(i_addr_rdE[1]), .D(
        i_addr_rdE[0]), .Q(n62) );
  XNR20 U59 ( .A(i_addr_rs[0]), .B(i_addr_rdE[0]), .Q(n56) );
  XNR20 U60 ( .A(i_addr_rs[1]), .B(i_addr_rdE[1]), .Q(n55) );
  NAND20 U61 ( .A(n63), .B(n48), .Q(o_con_fa[2]) );
  NOR40 U62 ( .A(n64), .B(n65), .C(n66), .D(n67), .Q(n50) );
  IMUX20 U63 ( .A(n68), .B(i_addr_rs[4]), .S(i_addr_rdM[4]), .Q(n67) );
  NOR20 U64 ( .A(n69), .B(i_addr_rs[4]), .Q(n68) );
  NOR40 U65 ( .A(i_addr_rdM[3]), .B(i_addr_rdM[2]), .C(i_addr_rdM[1]), .D(
        i_addr_rdM[0]), .Q(n69) );
  XOR20 U66 ( .A(i_addr_rdM[3]), .B(i_addr_rs[3]), .Q(n66) );
  XNR20 U67 ( .A(n18), .B(i_addr_rs[2]), .Q(n65) );
  CLKIN0 U68 ( .A(i_addr_rdM[2]), .Q(n18) );
  XNR20 U69 ( .A(n19), .B(i_addr_rs[1]), .Q(n64) );
  CLKIN0 U70 ( .A(i_addr_rdM[1]), .Q(n19) );
  NAND40 U71 ( .A(n70), .B(n71), .C(n72), .D(n73), .Q(n48) );
  NOR40 U72 ( .A(n74), .B(n75), .C(n76), .D(n77), .Q(n73) );
  XOR20 U73 ( .A(i_addr_rtW[1]), .B(i_addr_rs[1]), .Q(n77) );
  XOR20 U74 ( .A(i_addr_rtW[0]), .B(i_addr_rs[0]), .Q(n76) );
  CLKIN0 U75 ( .A(i_con_memreadW), .Q(n75) );
  XNR20 U76 ( .A(i_addr_rtW[3]), .B(i_addr_rs[3]), .Q(n72) );
  XNR20 U77 ( .A(i_addr_rtW[4]), .B(i_addr_rs[4]), .Q(n71) );
  XNR20 U78 ( .A(i_addr_rtW[2]), .B(i_addr_rs[2]), .Q(n70) );
  CLKIN0 U79 ( .A(n63), .Q(n47) );
  NAND40 U80 ( .A(n78), .B(n79), .C(n80), .D(n81), .Q(n63) );
  NOR40 U81 ( .A(n74), .B(n1), .C(n82), .D(n83), .Q(n81) );
  XNR20 U82 ( .A(n45), .B(i_addr_rs[1]), .Q(n83) );
  CLKIN0 U83 ( .A(i_addr_rtM[1]), .Q(n45) );
  XOR20 U84 ( .A(i_addr_rtM[0]), .B(i_addr_rs[0]), .Q(n82) );
  CLKIN0 U85 ( .A(i_con_memreadM), .Q(n1) );
  NOR30 U86 ( .A(i_addr_rs[0]), .B(i_addr_rs[1]), .C(n84), .Q(n74) );
  CLKIN0 U87 ( .A(n85), .Q(n84) );
  NOR30 U88 ( .A(i_addr_rs[2]), .B(i_addr_rs[4]), .C(i_addr_rs[3]), .Q(n85) );
  XNR20 U89 ( .A(i_addr_rtM[3]), .B(i_addr_rs[3]), .Q(n80) );
  XNR20 U90 ( .A(i_addr_rtM[4]), .B(i_addr_rs[4]), .Q(n79) );
  XNR20 U91 ( .A(i_addr_rtM[2]), .B(i_addr_rs[2]), .Q(n78) );
endmodule


module decode ( i_clk, i_nrst, i_addr_pc4, i_data_instr, i_con_Wregwrite, 
        i_data_Wregwrite, i_addr_Wregwrite, i_addr_Erd, i_addr_Mrd, 
        i_con_Eregwrite, i_con_Mregwrite, i_addr_rtM, i_addr_rtW, 
        i_con_memreadM, i_con_memreadW, i_data_Wmemout, o_data_rs, o_data_rt, 
        o_addr_rd, o_addr_rt, o_data_jr, o_con_jump, o_addr_pc4, o_addr_branch, 
        o_addr_jump, o_con_Ealuop, o_con_Ealusrc, o_con_Eregdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_con_ifstall, o_con_Ebop, o_data_signext, 
        o_con_Efamux, o_con_Efbmux, o_data_Fmemout );
  input [31:0] i_addr_pc4;
  input [31:0] i_data_instr;
  input [31:0] i_data_Wregwrite;
  input [4:0] i_addr_Wregwrite;
  input [4:0] i_addr_Erd;
  input [4:0] i_addr_Mrd;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  input [31:0] i_data_Wmemout;
  output [31:0] o_data_rs;
  output [31:0] o_data_rt;
  output [4:0] o_addr_rd;
  output [4:0] o_addr_rt;
  output [31:0] o_data_jr;
  output [1:0] o_con_jump;
  output [31:0] o_addr_pc4;
  output [31:0] o_addr_branch;
  output [31:0] o_addr_jump;
  output [5:0] o_con_Ealuop;
  output [2:0] o_con_Ebop;
  output [31:0] o_data_signext;
  output [2:0] o_con_Efamux;
  output [2:0] o_con_Efbmux;
  output [31:0] o_data_Fmemout;
  input i_clk, i_nrst, i_con_Wregwrite, i_con_Eregwrite, i_con_Mregwrite,
         i_con_memreadM, i_con_memreadW;
  output o_con_Ealusrc, o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite,
         o_con_Malupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall;
  wire   control_o_con_alusrc, control_o_con_regdst, jbcon_o_con_aluPC4,
         control_o_con_memread, control_o_con_memwrite, control_o_con_memtoreg,
         control_o_con_regwrite, signext_i_con_signext, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;
  wire   [31:0] regbank_o_data_Rt;
  wire   [5:0] control_o_con_aluop;
  wire   [31:0] signext_o_data_immD;
  wire   [2:0] for_o_con_fa;
  wire   [2:0] for_o_con_fb;
  wire   [31:0] pcadd_o_addr_pcbranchE;
  wire   [2:0] jbcon_o_con_bop;
  wire   [31:2] pcadd_i_data_immshiftl;
  assign o_addr_jump[1] = o_addr_jump[0];

  DFC3 pipe_bop_reg_2_ ( .D(jbcon_o_con_bop[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[2]) );
  DFC3 pipe_bop_reg_1_ ( .D(jbcon_o_con_bop[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[1]) );
  DFC3 pipe_bop_reg_0_ ( .D(jbcon_o_con_bop[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[0]) );
  DFC3 pipe_data_rs_reg_29_ ( .D(o_data_jr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[29]) );
  DFC3 pipe_data_rs_reg_17_ ( .D(o_data_jr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[17]) );
  DFC3 pipe_data_rs_reg_11_ ( .D(o_data_jr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[11]) );
  DFC3 pipe_data_rs_reg_10_ ( .D(o_data_jr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[10]) );
  DFC3 pipe_data_rs_reg_9_ ( .D(o_data_jr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[9]) );
  DFC3 pipe_data_rs_reg_8_ ( .D(o_data_jr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[8]) );
  DFC3 pipe_data_rs_reg_6_ ( .D(o_data_jr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[6]) );
  DFC3 pipe_data_rs_reg_4_ ( .D(o_data_jr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[4]) );
  DFC3 pipe_data_rs_reg_3_ ( .D(o_data_jr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[3]) );
  DFC3 pipe_data_rs_reg_2_ ( .D(o_data_jr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[2]) );
  DFC3 pipe_data_rs_reg_1_ ( .D(o_data_jr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[1]) );
  DFC3 pipe_data_rs_reg_0_ ( .D(o_data_jr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[0]) );
  DFC3 pipe_data_rt_reg_31_ ( .D(regbank_o_data_Rt[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[31]) );
  DFC3 pipe_data_rt_reg_30_ ( .D(regbank_o_data_Rt[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC3 pipe_data_rt_reg_29_ ( .D(regbank_o_data_Rt[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[29]) );
  DFC3 pipe_data_rt_reg_28_ ( .D(regbank_o_data_Rt[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28]) );
  DFC3 pipe_data_rt_reg_27_ ( .D(regbank_o_data_Rt[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27]) );
  DFC3 pipe_data_rt_reg_26_ ( .D(regbank_o_data_Rt[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26]) );
  DFC3 pipe_data_rt_reg_25_ ( .D(regbank_o_data_Rt[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25]) );
  DFC3 pipe_data_rt_reg_24_ ( .D(regbank_o_data_Rt[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24]) );
  DFC3 pipe_data_rt_reg_23_ ( .D(regbank_o_data_Rt[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23]) );
  DFC3 pipe_data_rt_reg_22_ ( .D(regbank_o_data_Rt[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC3 pipe_data_rt_reg_21_ ( .D(regbank_o_data_Rt[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21]) );
  DFC3 pipe_data_rt_reg_20_ ( .D(regbank_o_data_Rt[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20]) );
  DFC3 pipe_data_rt_reg_19_ ( .D(regbank_o_data_Rt[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19]) );
  DFC3 pipe_data_rt_reg_18_ ( .D(regbank_o_data_Rt[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18]) );
  DFC3 pipe_data_rt_reg_17_ ( .D(regbank_o_data_Rt[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17]) );
  DFC3 pipe_data_rt_reg_16_ ( .D(regbank_o_data_Rt[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC3 pipe_data_rt_reg_15_ ( .D(regbank_o_data_Rt[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15]) );
  DFC3 pipe_data_rt_reg_14_ ( .D(regbank_o_data_Rt[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14]) );
  DFC3 pipe_data_rt_reg_13_ ( .D(regbank_o_data_Rt[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC3 pipe_data_rt_reg_12_ ( .D(regbank_o_data_Rt[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12]) );
  DFC3 pipe_data_rt_reg_11_ ( .D(regbank_o_data_Rt[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11]) );
  DFC3 pipe_data_rt_reg_10_ ( .D(regbank_o_data_Rt[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC3 pipe_data_rt_reg_9_ ( .D(regbank_o_data_Rt[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[9]) );
  DFC3 pipe_data_rt_reg_8_ ( .D(regbank_o_data_Rt[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[8]) );
  DFC3 pipe_data_rt_reg_7_ ( .D(regbank_o_data_Rt[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[7]) );
  DFC3 pipe_data_rt_reg_6_ ( .D(regbank_o_data_Rt[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[6]) );
  DFC3 pipe_data_rt_reg_5_ ( .D(regbank_o_data_Rt[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[5]) );
  DFC3 pipe_data_rt_reg_4_ ( .D(regbank_o_data_Rt[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[4]) );
  DFC3 pipe_data_rt_reg_3_ ( .D(regbank_o_data_Rt[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[3]) );
  DFC3 pipe_data_rt_reg_2_ ( .D(regbank_o_data_Rt[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[2]) );
  DFC3 pipe_data_rt_reg_0_ ( .D(regbank_o_data_Rt[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[0]) );
  DFC3 pipe_addr_rd_reg_4_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[4]) );
  DFC3 pipe_addr_rd_reg_3_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[3]) );
  DFC3 pipe_addr_rd_reg_2_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[2]) );
  DFC3 pipe_addr_rd_reg_1_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[1]) );
  DFC3 pipe_addr_rd_reg_0_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[0]) );
  DFC3 pipe_addr_rt_reg_4_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[0]) );
  DFC3 pipe_addr_pc4_reg_31_ ( .D(i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_addr_pc4_reg_30_ ( .D(i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_addr_pc4_reg_29_ ( .D(i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_addr_pc4_reg_28_ ( .D(i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_addr_pc4_reg_27_ ( .D(i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_addr_pc4_reg_26_ ( .D(i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_addr_pc4_reg_25_ ( .D(i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_addr_pc4_reg_24_ ( .D(i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_addr_pc4_reg_23_ ( .D(i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_addr_pc4_reg_22_ ( .D(i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_addr_pc4_reg_21_ ( .D(i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_addr_pc4_reg_20_ ( .D(i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_addr_pc4_reg_19_ ( .D(i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_addr_pc4_reg_18_ ( .D(i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_addr_pc4_reg_17_ ( .D(i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_addr_pc4_reg_16_ ( .D(i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_addr_pc4_reg_15_ ( .D(i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_addr_pc4_reg_14_ ( .D(i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_addr_pc4_reg_13_ ( .D(i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_addr_pc4_reg_12_ ( .D(i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_addr_pc4_reg_11_ ( .D(i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_addr_pc4_reg_10_ ( .D(i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_addr_pc4_reg_9_ ( .D(i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_addr_pc4_reg_8_ ( .D(i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_addr_pc4_reg_7_ ( .D(i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_addr_pc4_reg_6_ ( .D(i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_addr_pc4_reg_5_ ( .D(i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_addr_pc4_reg_4_ ( .D(i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_addr_pc4_reg_3_ ( .D(i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_addr_pc4_reg_2_ ( .D(i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_addr_pc4_reg_1_ ( .D(i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_addr_pc4_reg_0_ ( .D(i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  DFC3 pipe_con_Ealuop_reg_5_ ( .D(control_o_con_aluop[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[5]) );
  DFC3 pipe_con_Ealuop_reg_4_ ( .D(control_o_con_aluop[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[4]) );
  DFC3 pipe_con_Ealuop_reg_3_ ( .D(control_o_con_aluop[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[3]) );
  DFC3 pipe_con_Ealuop_reg_2_ ( .D(control_o_con_aluop[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[2]) );
  DFC3 pipe_con_Ealuop_reg_1_ ( .D(control_o_con_aluop[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[1]) );
  DFC3 pipe_con_Ealuop_reg_0_ ( .D(control_o_con_aluop[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[0]) );
  DFC3 pipe_con_Ealusrc_reg ( .D(control_o_con_alusrc), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Ealusrc) );
  DFC3 pipe_con_MaluPC4_reg ( .D(jbcon_o_con_aluPC4), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Malupc8) );
  DFC3 pipe_con_Mmemread_reg ( .D(control_o_con_memread), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(control_o_con_memwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(control_o_con_memtoreg), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(control_o_con_regwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wregwrite) );
  DFC3 pipe_signext_o_data_immD_reg_31_ ( .D(signext_o_data_immD[31]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[31]) );
  DFC3 pipe_signext_o_data_immD_reg_30_ ( .D(signext_o_data_immD[30]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[30]) );
  DFC3 pipe_signext_o_data_immD_reg_29_ ( .D(signext_o_data_immD[29]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[29]) );
  DFC3 pipe_signext_o_data_immD_reg_28_ ( .D(signext_o_data_immD[28]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[28]) );
  DFC3 pipe_signext_o_data_immD_reg_27_ ( .D(signext_o_data_immD[27]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[27]) );
  DFC3 pipe_signext_o_data_immD_reg_26_ ( .D(signext_o_data_immD[26]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[26]) );
  DFC3 pipe_signext_o_data_immD_reg_25_ ( .D(signext_o_data_immD[25]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[25]) );
  DFC3 pipe_signext_o_data_immD_reg_24_ ( .D(signext_o_data_immD[24]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[24]) );
  DFC3 pipe_signext_o_data_immD_reg_23_ ( .D(signext_o_data_immD[23]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[23]) );
  DFC3 pipe_signext_o_data_immD_reg_22_ ( .D(signext_o_data_immD[22]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[22]) );
  DFC3 pipe_signext_o_data_immD_reg_21_ ( .D(signext_o_data_immD[21]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[21]) );
  DFC3 pipe_signext_o_data_immD_reg_20_ ( .D(signext_o_data_immD[20]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[20]) );
  DFC3 pipe_signext_o_data_immD_reg_19_ ( .D(signext_o_data_immD[19]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[19]) );
  DFC3 pipe_signext_o_data_immD_reg_18_ ( .D(signext_o_data_immD[18]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[18]) );
  DFC3 pipe_signext_o_data_immD_reg_17_ ( .D(signext_o_data_immD[17]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[17]) );
  DFC3 pipe_signext_o_data_immD_reg_16_ ( .D(signext_o_data_immD[16]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[16]) );
  DFC3 pipe_signext_o_data_immD_reg_15_ ( .D(signext_o_data_immD[15]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[15]) );
  DFC3 pipe_signext_o_data_immD_reg_14_ ( .D(signext_o_data_immD[14]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[14]) );
  DFC3 pipe_signext_o_data_immD_reg_13_ ( .D(signext_o_data_immD[13]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[13]) );
  DFC3 pipe_signext_o_data_immD_reg_12_ ( .D(signext_o_data_immD[12]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[12]) );
  DFC3 pipe_signext_o_data_immD_reg_11_ ( .D(signext_o_data_immD[11]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[11]) );
  DFC3 pipe_signext_o_data_immD_reg_10_ ( .D(signext_o_data_immD[10]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[10]) );
  DFC3 pipe_signext_o_data_immD_reg_9_ ( .D(signext_o_data_immD[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[9]) );
  DFC3 pipe_signext_o_data_immD_reg_8_ ( .D(signext_o_data_immD[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[8]) );
  DFC3 pipe_signext_o_data_immD_reg_7_ ( .D(signext_o_data_immD[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[7]) );
  DFC3 pipe_signext_o_data_immD_reg_6_ ( .D(signext_o_data_immD[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[6]) );
  DFC3 pipe_signext_o_data_immD_reg_5_ ( .D(signext_o_data_immD[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[5]) );
  DFC3 pipe_signext_o_data_immD_reg_4_ ( .D(signext_o_data_immD[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[4]) );
  DFC3 pipe_signext_o_data_immD_reg_3_ ( .D(signext_o_data_immD[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[3]) );
  DFC3 pipe_signext_o_data_immD_reg_2_ ( .D(signext_o_data_immD[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[2]) );
  DFC3 pipe_signext_o_data_immD_reg_1_ ( .D(signext_o_data_immD[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[1]) );
  DFC3 pipe_signext_o_data_immD_reg_0_ ( .D(signext_o_data_immD[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[0]) );
  DFC3 pipe_con_Efamux_reg_2_ ( .D(for_o_con_fa[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[2]) );
  DFC3 pipe_con_Efamux_reg_1_ ( .D(for_o_con_fa[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[1]) );
  DFC3 pipe_con_Efamux_reg_0_ ( .D(for_o_con_fa[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[0]) );
  DFC3 pipe_con_Efbmux_reg_2_ ( .D(for_o_con_fb[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[2]) );
  DFC3 pipe_con_Efbmux_reg_1_ ( .D(for_o_con_fb[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[1]) );
  DFC3 pipe_con_Efbmux_reg_0_ ( .D(for_o_con_fb[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[0]) );
  DFC3 pipe_FWmemout_reg_31_ ( .D(i_data_Wmemout[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[31]) );
  DFC3 pipe_FWmemout_reg_30_ ( .D(i_data_Wmemout[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[30]) );
  DFC3 pipe_FWmemout_reg_28_ ( .D(i_data_Wmemout[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[28]) );
  DFC3 pipe_FWmemout_reg_25_ ( .D(i_data_Wmemout[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[25]) );
  DFC3 pipe_FWmemout_reg_24_ ( .D(i_data_Wmemout[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[24]) );
  DFC3 pipe_FWmemout_reg_23_ ( .D(i_data_Wmemout[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[23]) );
  DFC3 pipe_FWmemout_reg_22_ ( .D(i_data_Wmemout[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[22]) );
  DFC3 pipe_FWmemout_reg_21_ ( .D(i_data_Wmemout[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[21]) );
  DFC3 pipe_FWmemout_reg_15_ ( .D(i_data_Wmemout[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[15]) );
  DFC3 pipe_FWmemout_reg_12_ ( .D(i_data_Wmemout[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[12]) );
  DFC3 pipe_FWmemout_reg_10_ ( .D(i_data_Wmemout[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[10]) );
  DFC3 pipe_FWmemout_reg_9_ ( .D(i_data_Wmemout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[9]) );
  DFC3 pipe_FWmemout_reg_8_ ( .D(i_data_Wmemout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[8]) );
  DFC3 pipe_FWmemout_reg_7_ ( .D(i_data_Wmemout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[7]) );
  DFC3 pipe_FWmemout_reg_6_ ( .D(i_data_Wmemout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[6]) );
  DFC3 pipe_FWmemout_reg_5_ ( .D(i_data_Wmemout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[5]) );
  DFC3 pipe_FWmemout_reg_4_ ( .D(i_data_Wmemout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[4]) );
  DFC3 pipe_FWmemout_reg_2_ ( .D(i_data_Wmemout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[2]) );
  DFC3 pipe_FWmemout_reg_1_ ( .D(i_data_Wmemout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[1]) );
  DFC3 pipe_FWmemout_reg_0_ ( .D(i_data_Wmemout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[0]) );
  DFC3 pipe_addr_branch_reg_31_ ( .D(pcadd_o_addr_pcbranchE[31]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[31]) );
  DFC3 pipe_addr_branch_reg_30_ ( .D(pcadd_o_addr_pcbranchE[30]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[30]) );
  DFC3 pipe_addr_branch_reg_29_ ( .D(pcadd_o_addr_pcbranchE[29]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[29]) );
  DFC3 pipe_addr_branch_reg_28_ ( .D(pcadd_o_addr_pcbranchE[28]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[28]) );
  DFC3 pipe_addr_branch_reg_27_ ( .D(pcadd_o_addr_pcbranchE[27]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[27]) );
  DFC3 pipe_addr_branch_reg_26_ ( .D(pcadd_o_addr_pcbranchE[26]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[26]) );
  DFC3 pipe_addr_branch_reg_25_ ( .D(pcadd_o_addr_pcbranchE[25]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[25]) );
  DFC3 pipe_addr_branch_reg_24_ ( .D(pcadd_o_addr_pcbranchE[24]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[24]) );
  DFC3 pipe_addr_branch_reg_23_ ( .D(pcadd_o_addr_pcbranchE[23]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[23]) );
  DFC3 pipe_addr_branch_reg_22_ ( .D(pcadd_o_addr_pcbranchE[22]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[22]) );
  DFC3 pipe_addr_branch_reg_21_ ( .D(pcadd_o_addr_pcbranchE[21]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[21]) );
  DFC3 pipe_addr_branch_reg_20_ ( .D(pcadd_o_addr_pcbranchE[20]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[20]) );
  DFC3 pipe_addr_branch_reg_19_ ( .D(pcadd_o_addr_pcbranchE[19]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[19]) );
  DFC3 pipe_addr_branch_reg_18_ ( .D(pcadd_o_addr_pcbranchE[18]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[18]) );
  DFC3 pipe_addr_branch_reg_17_ ( .D(pcadd_o_addr_pcbranchE[17]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[17]) );
  DFC3 pipe_addr_branch_reg_16_ ( .D(pcadd_o_addr_pcbranchE[16]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[16]) );
  DFC3 pipe_addr_branch_reg_15_ ( .D(pcadd_o_addr_pcbranchE[15]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[15]) );
  DFC3 pipe_addr_branch_reg_14_ ( .D(pcadd_o_addr_pcbranchE[14]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[14]) );
  DFC3 pipe_addr_branch_reg_13_ ( .D(pcadd_o_addr_pcbranchE[13]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[13]) );
  DFC3 pipe_addr_branch_reg_12_ ( .D(pcadd_o_addr_pcbranchE[12]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[12]) );
  DFC3 pipe_addr_branch_reg_11_ ( .D(pcadd_o_addr_pcbranchE[11]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[11]) );
  DFC3 pipe_addr_branch_reg_10_ ( .D(pcadd_o_addr_pcbranchE[10]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[10]) );
  DFC3 pipe_addr_branch_reg_9_ ( .D(pcadd_o_addr_pcbranchE[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[9]) );
  DFC3 pipe_addr_branch_reg_8_ ( .D(pcadd_o_addr_pcbranchE[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[8]) );
  DFC3 pipe_addr_branch_reg_7_ ( .D(pcadd_o_addr_pcbranchE[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[7]) );
  DFC3 pipe_addr_branch_reg_6_ ( .D(pcadd_o_addr_pcbranchE[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[6]) );
  DFC3 pipe_addr_branch_reg_5_ ( .D(pcadd_o_addr_pcbranchE[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[5]) );
  DFC3 pipe_addr_branch_reg_4_ ( .D(pcadd_o_addr_pcbranchE[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[4]) );
  DFC3 pipe_addr_branch_reg_3_ ( .D(pcadd_o_addr_pcbranchE[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[3]) );
  DFC3 pipe_addr_branch_reg_2_ ( .D(pcadd_o_addr_pcbranchE[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[2]) );
  DFC3 pipe_addr_branch_reg_1_ ( .D(pcadd_o_addr_pcbranchE[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[1]) );
  DFC3 pipe_addr_branch_reg_0_ ( .D(pcadd_o_addr_pcbranchE[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[0]) );
  D_control u_control ( .o_con_regdst(control_o_con_regdst), .o_con_memread(
        control_o_con_memread), .o_con_memtoreg(control_o_con_memtoreg), 
        .o_con_memwrite(control_o_con_memwrite), .o_con_alusrc(
        control_o_con_alusrc), .o_con_regwrite(control_o_con_regwrite), 
        .o_con_ifsign(signext_i_con_signext), .o_con_aluop(control_o_con_aluop), .i_con_instru(i_data_instr[31:26]) );
  D_jb_control u_jb_control ( .o_con_jump(o_con_jump), .o_con_bop(
        jbcon_o_con_bop), .o_con_aluPC4(jbcon_o_con_aluPC4), .o_con_ifstall(
        o_con_ifstall), .i_con_instru(i_data_instr[31:26]), .i_con_func(
        i_data_instr[5:0]), .i_con_rt(i_data_instr[16]) );
  D_pcadd u_pcadd ( .i_addr_pcadd4E(i_addr_pc4), .i_data_immshiftl({
        pcadd_i_data_immshiftl, o_addr_jump[0], o_addr_jump[0]}), 
        .o_addr_pcbranchE(pcadd_o_addr_pcbranchE) );
  D_register_bank u_regbank ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_addr_Rs(
        i_data_instr[25:21]), .i_addr_Rt(i_data_instr[20:16]), .i_con_RegWr(
        i_con_Wregwrite), .i_addr_Rd(i_addr_Wregwrite), .i_data_Rd(
        i_data_Wregwrite), .o_data_Rs(o_data_jr), .o_data_Rt(regbank_o_data_Rt) );
  D_shiftleft u_sl ( .i_data_immE(i_data_instr[15:0]), .o_data_immshiftl({
        pcadd_i_data_immshiftl, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}) );
  D_sign_extend u_signext ( .i_data_immD(i_data_instr[15:0]), .i_con_signext(
        signext_i_con_signext), .o_data_immD(signext_o_data_immD) );
  D_jump_ext u_jump_ext ( .i_addr_j(i_data_instr[25:0]), .i_PC4_j(
        i_addr_pc4[31:28]), .o_addr_j({o_addr_jump[31:2], 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4}) );
  D_forward u_forward ( .i_addr_rs(i_data_instr[25:21]), .i_addr_rt(
        i_data_instr[20:16]), .i_addr_rdE(i_addr_Erd), .i_addr_rdM(i_addr_Mrd), 
        .i_addr_rtM(i_addr_rtM), .i_addr_rtW(i_addr_rtW), .i_con_regwriteE(
        i_con_Eregwrite), .i_con_regwriteM(i_con_Mregwrite), .i_con_memreadM(
        i_con_memreadM), .i_con_memreadW(i_con_memreadW), .o_con_fa(
        for_o_con_fa), .o_con_fb(for_o_con_fb) );
  DFC1 pipe_con_Eregdst_reg ( .D(control_o_con_regdst), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Eregdst) );
  DFC1 pipe_data_rs_reg_19_ ( .D(o_data_jr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[19]) );
  DFC1 pipe_FWmemout_reg_27_ ( .D(i_data_Wmemout[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[27]) );
  DFC1 pipe_FWmemout_reg_3_ ( .D(i_data_Wmemout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[3]) );
  DFC1 pipe_FWmemout_reg_17_ ( .D(i_data_Wmemout[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[17]) );
  DFC1 pipe_FWmemout_reg_13_ ( .D(i_data_Wmemout[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[13]) );
  DFC1 pipe_FWmemout_reg_14_ ( .D(i_data_Wmemout[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[14]) );
  DFC1 pipe_FWmemout_reg_29_ ( .D(i_data_Wmemout[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[29]) );
  DFC1 pipe_FWmemout_reg_19_ ( .D(i_data_Wmemout[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[19]) );
  DFC1 pipe_data_rs_reg_28_ ( .D(o_data_jr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[28]) );
  DFC1 pipe_data_rs_reg_25_ ( .D(o_data_jr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[25]) );
  DFC1 pipe_data_rs_reg_13_ ( .D(o_data_jr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[13]) );
  DFC1 pipe_data_rs_reg_31_ ( .D(o_data_jr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[31]) );
  DFC1 pipe_data_rs_reg_26_ ( .D(o_data_jr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[26]) );
  DFC1 pipe_data_rs_reg_15_ ( .D(o_data_jr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[15]) );
  DFC1 pipe_data_rs_reg_24_ ( .D(o_data_jr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[24]) );
  DFC1 pipe_data_rs_reg_23_ ( .D(o_data_jr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[23]) );
  DFC1 pipe_data_rs_reg_22_ ( .D(o_data_jr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[22]) );
  DFC1 pipe_data_rs_reg_21_ ( .D(o_data_jr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[21]) );
  DFC1 pipe_data_rs_reg_16_ ( .D(o_data_jr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[16]) );
  DFC1 pipe_data_rs_reg_14_ ( .D(o_data_jr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[14]) );
  DFC1 pipe_data_rs_reg_7_ ( .D(o_data_jr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[7]) );
  DFC1 pipe_data_rs_reg_5_ ( .D(o_data_jr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[5]) );
  DFC1 pipe_data_rs_reg_30_ ( .D(o_data_jr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[30]) );
  DFC1 pipe_data_rs_reg_12_ ( .D(o_data_jr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[12]) );
  DFC1 pipe_FWmemout_reg_26_ ( .D(i_data_Wmemout[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[26]) );
  DFC1 pipe_data_rt_reg_1_ ( .D(regbank_o_data_Rt[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[1]) );
  DFC3 pipe_data_rs_reg_20_ ( .D(o_data_jr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[20]) );
  DFC3 pipe_data_rs_reg_18_ ( .D(o_data_jr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[18]) );
  DFC3 pipe_data_rs_reg_27_ ( .D(o_data_jr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[27]) );
  DFC1 pipe_FWmemout_reg_16_ ( .D(i_data_Wmemout[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[16]) );
  DFC1 pipe_FWmemout_reg_18_ ( .D(i_data_Wmemout[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[18]) );
  DFC3 pipe_FWmemout_reg_20_ ( .D(i_data_Wmemout[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[20]) );
  DFC1 pipe_FWmemout_reg_11_ ( .D(i_data_Wmemout[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[11]) );
  LOGIC0 U3 ( .Q(o_addr_jump[0]) );
endmodule


module E_alu_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233;

  NAND22 U3 ( .A(n129), .B(n125), .Q(n143) );
  XOR22 U4 ( .A(n193), .B(n194), .Q(DIFF[10]) );
  NAND23 U5 ( .A(B[9]), .B(n231), .Q(n27) );
  AOI312 U6 ( .A(n35), .B(n223), .C(n224), .D(n225), .Q(n1) );
  NOR20 U7 ( .A(A[4]), .B(n50), .Q(n47) );
  NOR20 U8 ( .A(A[4]), .B(n50), .Q(n54) );
  CLKIN3 U9 ( .A(A[4]), .Q(n229) );
  NOR22 U10 ( .A(A[4]), .B(n50), .Q(n204) );
  INV3 U11 ( .A(n147), .Q(n109) );
  INV6 U12 ( .A(n96), .Q(n127) );
  XOR22 U13 ( .A(n140), .B(n141), .Q(DIFF[13]) );
  NOR24 U14 ( .A(n154), .B(n146), .Q(n153) );
  INV4 U15 ( .A(n149), .Q(n222) );
  INV3 U16 ( .A(n37), .Q(n225) );
  AOI2111 U17 ( .A(n142), .B(n44), .C(n143), .D(n144), .Q(n141) );
  NAND22 U18 ( .A(A[1]), .B(n216), .Q(n63) );
  NAND24 U19 ( .A(n203), .B(n4), .Q(n96) );
  NOR22 U20 ( .A(n134), .B(n135), .Q(n133) );
  INV3 U21 ( .A(n132), .Q(n190) );
  NAND23 U22 ( .A(n221), .B(n222), .Q(n78) );
  INV3 U23 ( .A(n59), .Q(n212) );
  NAND24 U24 ( .A(B[2]), .B(n219), .Q(n59) );
  NAND24 U25 ( .A(B[1]), .B(n220), .Q(n66) );
  INV3 U26 ( .A(n119), .Q(n2) );
  NOR24 U27 ( .A(n212), .B(n63), .Q(n214) );
  NAND22 U28 ( .A(A[9]), .B(n168), .Q(n28) );
  NAND24 U29 ( .A(n214), .B(n215), .Q(n137) );
  NAND23 U30 ( .A(n60), .B(n215), .Q(n136) );
  INV3 U31 ( .A(n3), .Q(n4) );
  NOR23 U32 ( .A(n204), .B(n205), .Q(n203) );
  NAND22 U33 ( .A(n42), .B(n35), .Q(n3) );
  INV3 U34 ( .A(n165), .Q(n152) );
  NAND22 U35 ( .A(n39), .B(n40), .Q(n34) );
  INV6 U36 ( .A(n217), .Q(n215) );
  NOR23 U37 ( .A(A[3]), .B(n208), .Q(n217) );
  NOR21 U38 ( .A(A[9]), .B(n168), .Q(n167) );
  INV3 U39 ( .A(B[15]), .Q(n89) );
  INV3 U40 ( .A(n79), .Q(n98) );
  INV3 U41 ( .A(n129), .Q(n121) );
  CLKIN6 U42 ( .A(B[9]), .Q(n168) );
  NAND23 U43 ( .A(n97), .B(n98), .Q(n76) );
  INV3 U44 ( .A(A[13]), .Q(n156) );
  NAND22 U45 ( .A(B[14]), .B(n139), .Q(n87) );
  NAND22 U46 ( .A(n78), .B(n199), .Q(n198) );
  INV3 U47 ( .A(A[10]), .Q(n20) );
  INV12 U48 ( .A(n187), .Q(n44) );
  NAND20 U49 ( .A(n72), .B(B[0]), .Q(n232) );
  INV3 U50 ( .A(n71), .Q(n233) );
  CLKIN3 U51 ( .A(A[0]), .Q(n72) );
  INV3 U52 ( .A(B[0]), .Q(n70) );
  NOR21 U53 ( .A(B[0]), .B(n72), .Q(n71) );
  INV3 U54 ( .A(n66), .Q(n211) );
  NAND33 U55 ( .A(n59), .B(n191), .C(n66), .Q(n132) );
  NAND22 U56 ( .A(n209), .B(n210), .Q(n131) );
  NOR22 U57 ( .A(n211), .B(n212), .Q(n210) );
  NAND21 U58 ( .A(n87), .B(n94), .Q(n111) );
  NAND33 U59 ( .A(n87), .B(n94), .C(n99), .Q(n79) );
  INV3 U60 ( .A(n117), .Q(n125) );
  NAND24 U61 ( .A(n136), .B(n137), .Q(n189) );
  NAND22 U62 ( .A(A[2]), .B(n218), .Q(n67) );
  INV2 U63 ( .A(B[2]), .Q(n218) );
  NOR24 U64 ( .A(n7), .B(n192), .Q(n191) );
  NOR22 U65 ( .A(n172), .B(n173), .Q(n171) );
  INV2 U66 ( .A(n28), .Q(n195) );
  AOI212 U67 ( .A(n183), .B(n24), .C(n186), .Q(n194) );
  INV2 U68 ( .A(B[10]), .Q(n17) );
  NAND21 U69 ( .A(A[13]), .B(n155), .Q(n90) );
  INV1 U70 ( .A(B[13]), .Q(n155) );
  NOR32 U71 ( .A(n147), .B(n148), .C(n1), .Q(n117) );
  INV3 U72 ( .A(B[11]), .Q(n18) );
  INV8 U73 ( .A(B[3]), .Q(n208) );
  CLKIN2 U74 ( .A(B[1]), .Q(n216) );
  IMUX23 U75 ( .A(n157), .B(n158), .S(n159), .Q(DIFF[12]) );
  XNR21 U76 ( .A(n38), .B(n34), .Q(DIFF[6]) );
  NOR24 U77 ( .A(n100), .B(n101), .Q(n99) );
  NOR24 U78 ( .A(A[15]), .B(n89), .Q(n101) );
  NOR24 U79 ( .A(n70), .B(A[0]), .Q(n7) );
  AOI311 U80 ( .A(n127), .B(n109), .C(n128), .D(n121), .Q(n126) );
  INV1 U81 ( .A(n148), .Q(n221) );
  XOR22 U82 ( .A(n176), .B(n177), .Q(DIFF[11]) );
  AOI212 U83 ( .A(n178), .B(n179), .C(n180), .Q(n176) );
  XNR22 U84 ( .A(n32), .B(n33), .Q(DIFF[7]) );
  NAND22 U85 ( .A(n120), .B(n93), .Q(n144) );
  NAND22 U86 ( .A(A[12]), .B(n19), .Q(n93) );
  INV1 U87 ( .A(A[5]), .Q(n207) );
  INV2 U88 ( .A(A[9]), .Q(n231) );
  OAI212 U89 ( .A(B[4]), .B(n229), .C(n46), .Q(n223) );
  INV6 U90 ( .A(B[8]), .Q(n16) );
  NAND43 U91 ( .A(n151), .B(n152), .C(n27), .D(n153), .Q(n147) );
  NOR22 U92 ( .A(n167), .B(n165), .Q(n162) );
  NOR23 U93 ( .A(n10), .B(n11), .Q(n12) );
  INV3 U94 ( .A(n24), .Q(n11) );
  NOR22 U95 ( .A(n192), .B(n233), .Q(n209) );
  NAND23 U96 ( .A(B[6]), .B(n230), .Q(n35) );
  NOR21 U97 ( .A(n169), .B(n96), .Q(n14) );
  INV6 U98 ( .A(n27), .Q(n172) );
  NAND21 U99 ( .A(n65), .B(n66), .Q(n64) );
  NAND22 U100 ( .A(n13), .B(n131), .Q(n201) );
  OAI2111 U101 ( .A(n84), .B(n85), .C(n86), .D(n87), .Q(n80) );
  NAND22 U102 ( .A(n63), .B(n64), .Q(n58) );
  AOI312 U103 ( .A(n42), .B(n43), .C(n44), .D(n45), .Q(n39) );
  NAND42 U104 ( .A(n2), .B(n93), .C(n125), .D(n126), .Q(n124) );
  NOR22 U105 ( .A(n12), .B(n95), .Q(n159) );
  INV0 U106 ( .A(n46), .Q(n45) );
  NAND22 U107 ( .A(A[5]), .B(n228), .Q(n46) );
  NAND22 U108 ( .A(A[10]), .B(n17), .Q(n166) );
  NAND41 U109 ( .A(n13), .B(n131), .C(n132), .D(n133), .Q(n128) );
  OAI2112 U110 ( .A(n211), .B(n213), .C(n136), .D(n137), .Q(n200) );
  NOR24 U111 ( .A(A[11]), .B(n18), .Q(n165) );
  NOR24 U112 ( .A(n189), .B(n190), .Q(n5) );
  NOR24 U113 ( .A(n6), .B(n188), .Q(n187) );
  INV6 U114 ( .A(n5), .Q(n6) );
  OAI2112 U115 ( .A(n200), .B(n201), .C(n202), .D(n127), .Q(n199) );
  INV0 U116 ( .A(n192), .Q(n202) );
  CLKIN3 U117 ( .A(n8), .Q(n9) );
  NAND22 U118 ( .A(n119), .B(n118), .Q(n115) );
  NAND22 U119 ( .A(n114), .B(n116), .Q(n8) );
  NAND22 U120 ( .A(n115), .B(n9), .Q(n104) );
  CLKIN3 U121 ( .A(n169), .Q(n97) );
  CLKIN3 U122 ( .A(n111), .Q(n118) );
  NOR32 U123 ( .A(n104), .B(n105), .C(n106), .Q(n103) );
  NOR23 U124 ( .A(A[3]), .B(n208), .Q(n192) );
  NAND21 U125 ( .A(n117), .B(n118), .Q(n116) );
  INV1 U126 ( .A(n97), .Q(n10) );
  INV6 U127 ( .A(n197), .Q(n24) );
  NAND22 U128 ( .A(n130), .B(n131), .Q(n188) );
  NAND21 U129 ( .A(n127), .B(n44), .Q(n184) );
  CLKIN3 U130 ( .A(n47), .Q(n43) );
  NAND20 U131 ( .A(A[3]), .B(n208), .Q(n130) );
  NAND20 U132 ( .A(A[3]), .B(n208), .Q(n13) );
  INV2 U133 ( .A(B[5]), .Q(n228) );
  NOR21 U134 ( .A(A[0]), .B(n70), .Q(n69) );
  CLKIN3 U135 ( .A(n227), .Q(n224) );
  NAND22 U136 ( .A(n121), .B(n118), .Q(n114) );
  INV0 U137 ( .A(n91), .Q(n113) );
  OAI2112 U138 ( .A(n160), .B(n79), .C(n80), .D(n81), .Q(n74) );
  NAND20 U139 ( .A(n94), .B(n90), .Q(n140) );
  NAND22 U140 ( .A(B[13]), .B(n156), .Q(n94) );
  NOR20 U141 ( .A(n26), .B(n172), .Q(n183) );
  NOR20 U142 ( .A(n150), .B(n186), .Q(n185) );
  INV3 U143 ( .A(n181), .Q(n186) );
  NOR20 U144 ( .A(n93), .B(n111), .Q(n105) );
  NAND20 U145 ( .A(n41), .B(n42), .Q(n40) );
  AOI210 U146 ( .A(n112), .B(n87), .C(n113), .Q(n107) );
  NOR21 U147 ( .A(n92), .B(n93), .Q(n84) );
  NOR20 U148 ( .A(A[8]), .B(n16), .Q(n26) );
  NAND20 U149 ( .A(n181), .B(n182), .Q(n179) );
  NAND20 U150 ( .A(n27), .B(n28), .Q(n21) );
  INV0 U151 ( .A(n26), .Q(n23) );
  NAND20 U152 ( .A(n42), .B(n46), .Q(n48) );
  AOI210 U153 ( .A(n43), .B(n44), .C(n41), .Q(n49) );
  NAND20 U154 ( .A(n151), .B(n166), .Q(n193) );
  XNR20 U155 ( .A(n68), .B(n65), .Q(DIFF[1]) );
  NAND20 U156 ( .A(A[8]), .B(n16), .Q(n196) );
  NAND20 U157 ( .A(n59), .B(n67), .Q(n61) );
  NAND20 U158 ( .A(n87), .B(n91), .Q(n122) );
  NOR20 U159 ( .A(B[15]), .B(n83), .Q(n82) );
  INV0 U160 ( .A(A[15]), .Q(n83) );
  NAND22 U161 ( .A(n14), .B(n98), .Q(n15) );
  AOI210 U162 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  INV6 U163 ( .A(B[7]), .Q(n206) );
  NAND20 U164 ( .A(A[4]), .B(n50), .Q(n55) );
  INV3 U165 ( .A(n183), .Q(n182) );
  NAND22 U166 ( .A(n109), .B(n150), .Q(n129) );
  INV3 U167 ( .A(B[12]), .Q(n19) );
  INV3 U168 ( .A(n120), .Q(n119) );
  INV3 U169 ( .A(n88), .Q(n86) );
  NAND22 U170 ( .A(n90), .B(n91), .Q(n85) );
  INV3 U171 ( .A(n15), .Q(n73) );
  NAND22 U172 ( .A(n95), .B(n145), .Q(n120) );
  INV3 U173 ( .A(n146), .Q(n145) );
  INV0 U174 ( .A(A[11]), .Q(n164) );
  XOR21 U175 ( .A(n122), .B(n123), .Q(DIFF[14]) );
  NAND22 U176 ( .A(n170), .B(n171), .Q(n169) );
  NOR21 U177 ( .A(n165), .B(n154), .Q(n170) );
  XOR21 U178 ( .A(n48), .B(n49), .Q(DIFF[5]) );
  XOR21 U179 ( .A(n21), .B(n22), .Q(DIFF[9]) );
  AOI211 U180 ( .A(n23), .B(n24), .C(n25), .Q(n22) );
  INV3 U181 ( .A(n166), .Q(n180) );
  AOI311 U182 ( .A(n78), .B(n184), .C(n185), .D(n173), .Q(n178) );
  IMUX21 U183 ( .A(n29), .B(n30), .S(n24), .Q(DIFF[8]) );
  XOR21 U184 ( .A(n102), .B(n103), .Q(DIFF[15]) );
  NOR22 U185 ( .A(A[8]), .B(n16), .Q(n154) );
  NAND22 U186 ( .A(n107), .B(n108), .Q(n106) );
  NAND31 U187 ( .A(n109), .B(n110), .C(n44), .Q(n108) );
  NOR23 U188 ( .A(n150), .B(n198), .Q(n197) );
  INV3 U189 ( .A(A[8]), .Q(n31) );
  NAND22 U190 ( .A(n232), .B(n233), .Q(DIFF[0]) );
  INV3 U191 ( .A(n82), .Q(n81) );
  NOR21 U192 ( .A(A[7]), .B(n206), .Q(n205) );
  INV3 U193 ( .A(A[14]), .Q(n139) );
  NAND22 U194 ( .A(A[14]), .B(n138), .Q(n91) );
  INV3 U195 ( .A(B[14]), .Q(n138) );
  IMUX21 U196 ( .A(n51), .B(n52), .S(n53), .Q(DIFF[4]) );
  NOR21 U197 ( .A(n54), .B(n41), .Q(n51) );
  NOR21 U198 ( .A(n174), .B(n175), .Q(n157) );
  XNR21 U199 ( .A(n56), .B(n57), .Q(DIFF[3]) );
  INV3 U200 ( .A(B[4]), .Q(n50) );
  XOR21 U201 ( .A(n61), .B(n62), .Q(DIFF[2]) );
  NAND22 U202 ( .A(n233), .B(n69), .Q(n65) );
  OAI212 U203 ( .A(B[8]), .B(n31), .C(n28), .Q(n161) );
  INV3 U204 ( .A(A[1]), .Q(n220) );
  INV1 U205 ( .A(A[2]), .Q(n219) );
  NAND22 U206 ( .A(A[6]), .B(n226), .Q(n37) );
  CLKIN0 U207 ( .A(n37), .Q(n36) );
  NAND20 U208 ( .A(n66), .B(n63), .Q(n68) );
  NAND20 U209 ( .A(n35), .B(n37), .Q(n38) );
  NOR20 U210 ( .A(n147), .B(n96), .Q(n142) );
  NOR20 U211 ( .A(n111), .B(n96), .Q(n110) );
  XNR20 U212 ( .A(B[3]), .B(A[3]), .Q(n56) );
  NAND23 U213 ( .A(B[10]), .B(n20), .Q(n151) );
  INV1 U214 ( .A(B[6]), .Q(n226) );
  NAND22 U215 ( .A(B[5]), .B(n207), .Q(n42) );
  CLKIN2 U216 ( .A(A[6]), .Q(n230) );
  NOR21 U217 ( .A(A[5]), .B(n228), .Q(n227) );
  NAND21 U218 ( .A(A[7]), .B(n206), .Q(n77) );
  NOR21 U219 ( .A(A[7]), .B(n206), .Q(n148) );
  XNR20 U220 ( .A(B[7]), .B(A[7]), .Q(n32) );
  AOI210 U221 ( .A(B[8]), .B(n31), .C(n25), .Q(n30) );
  XOR20 U222 ( .A(B[8]), .B(A[8]), .Q(n29) );
  XOR20 U223 ( .A(B[15]), .B(A[15]), .Q(n102) );
  NOR21 U224 ( .A(A[15]), .B(n89), .Q(n88) );
  XOR20 U225 ( .A(B[11]), .B(A[11]), .Q(n177) );
  OAI210 U226 ( .A(A[0]), .B(n70), .C(n59), .Q(n213) );
  NOR21 U227 ( .A(A[12]), .B(n19), .Q(n174) );
  XOR20 U228 ( .A(B[12]), .B(A[12]), .Q(n158) );
  NOR22 U229 ( .A(A[12]), .B(n19), .Q(n146) );
  NOR22 U230 ( .A(A[12]), .B(n19), .Q(n100) );
  XOR20 U231 ( .A(B[4]), .B(A[4]), .Q(n52) );
  AOI212 U232 ( .A(n34), .B(n35), .C(n36), .Q(n33) );
  CLKIN3 U233 ( .A(n44), .Q(n53) );
  CLKIN3 U234 ( .A(n55), .Q(n41) );
  CLKIN3 U235 ( .A(n58), .Q(n62) );
  AOI2112 U236 ( .A(n73), .B(n44), .C(n74), .D(n75), .Q(DIFF[16]) );
  OAI222 U237 ( .A(n76), .B(n77), .C(n76), .D(n78), .Q(n75) );
  CLKIN3 U238 ( .A(n94), .Q(n92) );
  AOI212 U239 ( .A(n124), .B(n94), .C(n112), .Q(n123) );
  CLKIN3 U240 ( .A(n90), .Q(n112) );
  CLKIN3 U241 ( .A(n136), .Q(n135) );
  CLKIN3 U242 ( .A(n137), .Q(n134) );
  CLKIN6 U243 ( .A(n160), .Q(n95) );
  AOI312 U244 ( .A(n151), .B(n161), .C(n162), .D(n163), .Q(n160) );
  OAI222 U245 ( .A(B[11]), .B(n164), .C(n165), .D(n166), .Q(n163) );
  CLKIN3 U246 ( .A(n151), .Q(n173) );
  CLKIN3 U247 ( .A(n93), .Q(n175) );
  CLKIN3 U248 ( .A(n77), .Q(n150) );
  OAI212 U249 ( .A(n195), .B(n25), .C(n27), .Q(n181) );
  CLKIN3 U250 ( .A(n196), .Q(n25) );
  CLKIN3 U251 ( .A(n67), .Q(n60) );
  AOI312 U252 ( .A(n35), .B(n223), .C(n224), .D(n225), .Q(n149) );
endmodule


module E_alu_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74;

  CLKIN2 U2 ( .A(A[4]), .Q(n13) );
  CLKIN3 U3 ( .A(n40), .Q(n38) );
  AOI222 U4 ( .A(B[7]), .B(A[7]), .C(n24), .D(n25), .Q(n3) );
  NOR23 U5 ( .A(n61), .B(n16), .Q(n6) );
  NAND20 U6 ( .A(B[4]), .B(A[4]), .Q(n46) );
  NAND24 U7 ( .A(n44), .B(n45), .Q(n31) );
  NAND22 U8 ( .A(A[1]), .B(B[1]), .Q(n56) );
  NAND33 U9 ( .A(n21), .B(n22), .C(n23), .Q(n5) );
  NAND22 U10 ( .A(n17), .B(n18), .Q(n16) );
  NOR21 U11 ( .A(n19), .B(n20), .Q(n17) );
  CLKIN0 U12 ( .A(A[7]), .Q(n9) );
  XOR21 U13 ( .A(n40), .B(n43), .Q(SUM[5]) );
  NAND31 U14 ( .A(B[4]), .B(A[4]), .C(n31), .Q(n27) );
  AOI211 U15 ( .A(n13), .B(n14), .C(n15), .Q(n7) );
  NAND26 U16 ( .A(n41), .B(n42), .Q(n12) );
  NAND20 U17 ( .A(B[0]), .B(A[0]), .Q(n60) );
  NAND20 U18 ( .A(B[0]), .B(A[0]), .Q(n74) );
  INV3 U19 ( .A(n39), .Q(n30) );
  INV3 U20 ( .A(n57), .Q(n18) );
  BUF6 U21 ( .A(A[2]), .Q(n2) );
  INV3 U22 ( .A(B[5]), .Q(n44) );
  NAND24 U23 ( .A(n46), .B(n47), .Q(n40) );
  AOI212 U24 ( .A(n9), .B(n10), .C(n11), .Q(n8) );
  NAND21 U25 ( .A(B[3]), .B(A[3]), .Q(n21) );
  XNR22 U26 ( .A(n64), .B(n65), .Q(SUM[3]) );
  INV2 U27 ( .A(n74), .Q(n72) );
  CLKIN6 U28 ( .A(B[6]), .Q(n41) );
  INV2 U29 ( .A(A[5]), .Q(n45) );
  NAND22 U30 ( .A(B[5]), .B(A[5]), .Q(n39) );
  CLKIN1 U31 ( .A(A[0]), .Q(n20) );
  OAI2112 U32 ( .A(n26), .B(n27), .C(n28), .D(n29), .Q(n25) );
  NAND21 U33 ( .A(n30), .B(n12), .Q(n28) );
  NOR24 U34 ( .A(A[3]), .B(B[3]), .Q(n57) );
  CLKIN1 U35 ( .A(B[7]), .Q(n10) );
  XNR21 U36 ( .A(n37), .B(n35), .Q(SUM[6]) );
  NAND21 U37 ( .A(n66), .B(n67), .Q(n64) );
  INV2 U38 ( .A(n59), .Q(n51) );
  NOR30 U39 ( .A(n60), .B(n57), .C(n61), .Q(n59) );
  NOR20 U40 ( .A(n30), .B(n15), .Q(n43) );
  IMUX20 U41 ( .A(n49), .B(n50), .S(n48), .Q(SUM[4]) );
  IMUX20 U42 ( .A(n19), .B(B[0]), .S(A[0]), .Q(SUM[0]) );
  NAND22 U43 ( .A(n51), .B(n52), .Q(n48) );
  NOR21 U44 ( .A(n53), .B(n54), .Q(n52) );
  XNR21 U45 ( .A(n68), .B(n69), .Q(SUM[2]) );
  XOR21 U46 ( .A(n33), .B(n34), .Q(SUM[7]) );
  NAND22 U47 ( .A(n70), .B(n71), .Q(n68) );
  NOR21 U48 ( .A(n62), .B(n63), .Q(n50) );
  INV3 U49 ( .A(n46), .Q(n63) );
  INV3 U50 ( .A(B[4]), .Q(n14) );
  INV3 U51 ( .A(A[6]), .Q(n42) );
  XNR21 U52 ( .A(n72), .B(n73), .Q(SUM[1]) );
  NOR22 U53 ( .A(B[2]), .B(n2), .Q(n58) );
  INV3 U54 ( .A(B[0]), .Q(n19) );
  NAND20 U55 ( .A(B[1]), .B(A[1]), .Q(n70) );
  OAI212 U56 ( .A(A[4]), .B(B[4]), .C(n48), .Q(n47) );
  NAND24 U57 ( .A(n3), .B(n4), .Q(SUM[8]) );
  CLKIN1 U58 ( .A(n23), .Q(n53) );
  CLKIN2 U59 ( .A(n12), .Q(n11) );
  CLKIN1 U60 ( .A(n29), .Q(n36) );
  NAND22 U61 ( .A(n22), .B(n21), .Q(n54) );
  OAI222 U62 ( .A(B[2]), .B(n2), .C(B[1]), .D(A[1]), .Q(n61) );
  NAND20 U63 ( .A(n12), .B(n29), .Q(n37) );
  INV2 U64 ( .A(n12), .Q(n26) );
  XNR20 U65 ( .A(B[3]), .B(A[3]), .Q(n65) );
  OAI210 U66 ( .A(B[1]), .B(A[1]), .C(n70), .Q(n73) );
  OAI210 U67 ( .A(B[1]), .B(A[1]), .C(n72), .Q(n71) );
  INV3 U68 ( .A(n32), .Q(n24) );
  NOR20 U69 ( .A(B[4]), .B(A[4]), .Q(n62) );
  NAND22 U70 ( .A(B[6]), .B(A[6]), .Q(n29) );
  XNR20 U71 ( .A(B[7]), .B(A[7]), .Q(n33) );
  NOR20 U72 ( .A(A[7]), .B(B[7]), .Q(n32) );
  OAI2111 U73 ( .A(B[3]), .B(A[3]), .C(n2), .D(B[2]), .Q(n22) );
  OAI210 U74 ( .A(B[2]), .B(n2), .C(n68), .Q(n67) );
  NAND20 U75 ( .A(B[2]), .B(n2), .Q(n66) );
  OAI210 U76 ( .A(B[2]), .B(n2), .C(n66), .Q(n69) );
  XNR20 U77 ( .A(B[4]), .B(A[4]), .Q(n49) );
  INV6 U78 ( .A(n55), .Q(n23) );
  OAI2112 U79 ( .A(n5), .B(n6), .C(n7), .D(n8), .Q(n4) );
  AOI212 U80 ( .A(n35), .B(n12), .C(n36), .Q(n34) );
  OAI212 U81 ( .A(n15), .B(n38), .C(n39), .Q(n35) );
  CLKIN3 U82 ( .A(n31), .Q(n15) );
  NOR33 U83 ( .A(n56), .B(n58), .C(n57), .Q(n55) );
endmodule


module E_alu_DW01_add_12 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79;

  NOR22 U2 ( .A(A[3]), .B(B[3]), .Q(n49) );
  NOR23 U3 ( .A(n45), .B(n46), .Q(n44) );
  AOI311 U4 ( .A(A[0]), .B(B[0]), .C(n71), .D(n73), .Q(n68) );
  INV2 U5 ( .A(n25), .Q(n71) );
  NOR22 U6 ( .A(A[1]), .B(B[1]), .Q(n25) );
  XOR21 U7 ( .A(n60), .B(n61), .Q(SUM[3]) );
  NAND22 U8 ( .A(n47), .B(n48), .Q(n17) );
  NOR21 U9 ( .A(n36), .B(n37), .Q(n15) );
  NAND22 U10 ( .A(n68), .B(n69), .Q(n63) );
  XNR21 U11 ( .A(n1), .B(n2), .Q(SUM[4]) );
  NOR21 U12 ( .A(B[0]), .B(A[0]), .Q(n28) );
  AOI311 U13 ( .A(n9), .B(n10), .C(n11), .D(n12), .Q(n8) );
  NAND41 U14 ( .A(n16), .B(n17), .C(n18), .D(n19), .Q(n11) );
  NOR21 U15 ( .A(n49), .B(n50), .Q(n48) );
  NOR22 U16 ( .A(B[2]), .B(A[2]), .Q(n50) );
  INV2 U17 ( .A(n76), .Q(n73) );
  AOI222 U18 ( .A(n53), .B(n54), .C(n55), .D(n56), .Q(n43) );
  NOR21 U19 ( .A(n58), .B(n49), .Q(n55) );
  NAND21 U20 ( .A(B[0]), .B(A[0]), .Q(n57) );
  OAI2111 U21 ( .A(A[3]), .B(B[3]), .C(A[2]), .D(B[2]), .Q(n16) );
  XOR22 U22 ( .A(n7), .B(n8), .Q(SUM[7]) );
  AOI212 U23 ( .A(n62), .B(n63), .C(n64), .Q(n61) );
  XOR22 U24 ( .A(n3), .B(n39), .Q(SUM[5]) );
  INV1 U25 ( .A(B[1]), .Q(n52) );
  NAND24 U26 ( .A(n43), .B(n44), .Q(n35) );
  NAND21 U27 ( .A(n72), .B(n77), .Q(n74) );
  XOR21 U28 ( .A(n74), .B(n75), .Q(SUM[1]) );
  INV2 U29 ( .A(n33), .Q(n10) );
  INV0 U30 ( .A(n38), .Q(n40) );
  XOR20 U31 ( .A(B[4]), .B(A[4]), .Q(n2) );
  INV2 U32 ( .A(n72), .Q(n70) );
  CLKIN2 U33 ( .A(n35), .Q(n1) );
  INV2 U34 ( .A(n28), .Q(n20) );
  CLKIN0 U35 ( .A(n27), .Q(n21) );
  XNR20 U36 ( .A(B[3]), .B(A[3]), .Q(n60) );
  NAND21 U37 ( .A(n29), .B(n30), .Q(n18) );
  NOR20 U38 ( .A(B[2]), .B(A[2]), .Q(n26) );
  NOR20 U39 ( .A(B[2]), .B(A[2]), .Q(n58) );
  NOR20 U40 ( .A(B[2]), .B(A[2]), .Q(n66) );
  NAND20 U41 ( .A(B[3]), .B(A[3]), .Q(n24) );
  NAND20 U42 ( .A(B[2]), .B(A[2]), .Q(n65) );
  OAI210 U43 ( .A(B[2]), .B(A[2]), .C(n65), .Q(n67) );
  NOR20 U44 ( .A(n32), .B(n49), .Q(n29) );
  NOR20 U45 ( .A(B[2]), .B(A[2]), .Q(n32) );
  NOR20 U46 ( .A(B[2]), .B(A[2]), .Q(n59) );
  INV0 U47 ( .A(A[0]), .Q(n5) );
  NAND20 U48 ( .A(B[0]), .B(A[0]), .Q(n31) );
  NOR20 U49 ( .A(A[0]), .B(B[0]), .Q(n72) );
  NAND20 U50 ( .A(B[0]), .B(A[0]), .Q(n77) );
  NOR20 U51 ( .A(n42), .B(n6), .Q(n41) );
  INV0 U52 ( .A(A[4]), .Q(n42) );
  NAND20 U53 ( .A(B[1]), .B(A[1]), .Q(n76) );
  INV0 U54 ( .A(B[0]), .Q(n79) );
  XNR20 U55 ( .A(B[5]), .B(A[5]), .Q(n3) );
  NAND22 U56 ( .A(n16), .B(n24), .Q(n46) );
  INV3 U57 ( .A(n66), .Q(n62) );
  NOR21 U58 ( .A(B[3]), .B(A[3]), .Q(n27) );
  NOR21 U59 ( .A(n25), .B(n59), .Q(n54) );
  AOI311 U60 ( .A(n20), .B(n21), .C(n22), .D(n23), .Q(n19) );
  NOR21 U61 ( .A(n27), .B(n28), .Q(n53) );
  XNR21 U62 ( .A(n63), .B(n67), .Q(SUM[2]) );
  NAND22 U63 ( .A(n78), .B(n77), .Q(SUM[0]) );
  NAND22 U64 ( .A(n5), .B(n79), .Q(n78) );
  NAND22 U65 ( .A(n13), .B(n14), .Q(n12) );
  NOR21 U66 ( .A(n38), .B(n36), .Q(n9) );
  NOR21 U67 ( .A(A[4]), .B(B[4]), .Q(n38) );
  NAND22 U68 ( .A(n70), .B(n71), .Q(n69) );
  NOR21 U69 ( .A(n25), .B(n57), .Q(n56) );
  NOR21 U70 ( .A(n51), .B(n52), .Q(n47) );
  INV3 U71 ( .A(A[1]), .Q(n51) );
  NAND22 U72 ( .A(n15), .B(n10), .Q(n13) );
  XNR21 U73 ( .A(n4), .B(n34), .Q(SUM[6]) );
  XOR20 U74 ( .A(B[6]), .B(A[6]), .Q(n4) );
  INV3 U75 ( .A(B[4]), .Q(n6) );
  NOR20 U76 ( .A(n73), .B(n25), .Q(n75) );
  NOR20 U77 ( .A(n25), .B(n26), .Q(n22) );
  NOR20 U78 ( .A(n25), .B(n31), .Q(n30) );
  XNR20 U79 ( .A(B[7]), .B(A[7]), .Q(n7) );
  NOR21 U80 ( .A(A[5]), .B(B[5]), .Q(n36) );
  AOI220 U81 ( .A(B[5]), .B(A[5]), .C(B[4]), .D(A[4]), .Q(n37) );
  NOR20 U82 ( .A(A[6]), .B(B[6]), .Q(n33) );
  NAND20 U83 ( .A(B[6]), .B(A[6]), .Q(n14) );
  CLKIN3 U84 ( .A(n24), .Q(n23) );
  AOI212 U85 ( .A(n9), .B(n35), .C(n15), .Q(n34) );
  AOI212 U86 ( .A(n40), .B(n35), .C(n41), .Q(n39) );
  CLKIN3 U87 ( .A(n17), .Q(n45) );
  CLKIN3 U88 ( .A(n65), .Q(n64) );
endmodule


module E_alu_DW01_add_13 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;

  NOR22 U2 ( .A(A[1]), .B(B[1]), .Q(n17) );
  NOR22 U3 ( .A(n41), .B(n42), .Q(n40) );
  NOR21 U4 ( .A(B[2]), .B(A[2]), .Q(n42) );
  NOR21 U5 ( .A(n59), .B(n17), .Q(n60) );
  NAND22 U6 ( .A(n35), .B(n36), .Q(n26) );
  NAND22 U7 ( .A(B[1]), .B(A[1]), .Q(n61) );
  AOI221 U8 ( .A(B[5]), .B(A[5]), .C(B[4]), .D(A[4]), .Q(n28) );
  INV1 U9 ( .A(B[1]), .Q(n44) );
  AOI212 U10 ( .A(n6), .B(n26), .C(n12), .Q(n25) );
  AOI212 U11 ( .A(n32), .B(n26), .C(n33), .Q(n31) );
  OAI210 U12 ( .A(B[2]), .B(A[2]), .C(n54), .Q(n56) );
  NAND20 U13 ( .A(B[2]), .B(A[2]), .Q(n54) );
  NOR20 U14 ( .A(B[2]), .B(A[2]), .Q(n55) );
  NOR20 U15 ( .A(B[2]), .B(A[2]), .Q(n21) );
  NOR20 U16 ( .A(B[2]), .B(A[2]), .Q(n48) );
  OAI2111 U17 ( .A(A[3]), .B(B[3]), .C(A[2]), .D(B[2]), .Q(n13) );
  NOR23 U18 ( .A(A[3]), .B(B[3]), .Q(n41) );
  NOR21 U19 ( .A(A[3]), .B(B[3]), .Q(n22) );
  NAND21 U20 ( .A(B[3]), .B(A[3]), .Q(n16) );
  NAND22 U21 ( .A(B[0]), .B(A[0]), .Q(n47) );
  INV1 U22 ( .A(n17), .Q(n58) );
  NOR20 U23 ( .A(n17), .B(n20), .Q(n19) );
  INV3 U24 ( .A(n57), .Q(n52) );
  INV2 U25 ( .A(n23), .Q(n7) );
  NOR21 U26 ( .A(n21), .B(n22), .Q(n18) );
  NAND41 U27 ( .A(n13), .B(n14), .C(n15), .D(n16), .Q(n8) );
  NOR21 U28 ( .A(n48), .B(n22), .Q(n45) );
  XNR20 U29 ( .A(n26), .B(n1), .Q(SUM[4]) );
  NAND20 U30 ( .A(B[0]), .B(A[0]), .Q(n20) );
  INV3 U31 ( .A(n54), .Q(n53) );
  NOR22 U32 ( .A(n37), .B(n38), .Q(n36) );
  INV0 U33 ( .A(n29), .Q(n32) );
  MUX21 U34 ( .A(B[0]), .B(n63), .S(A[0]), .Q(SUM[0]) );
  XNR20 U35 ( .A(B[4]), .B(A[4]), .Q(n1) );
  NOR20 U36 ( .A(n34), .B(n3), .Q(n33) );
  INV0 U37 ( .A(A[4]), .Q(n34) );
  NAND20 U38 ( .A(B[0]), .B(A[0]), .Q(n62) );
  INV0 U39 ( .A(B[0]), .Q(n63) );
  NAND22 U40 ( .A(n13), .B(n16), .Q(n38) );
  XNR21 U41 ( .A(n52), .B(n56), .Q(SUM[2]) );
  XNR21 U42 ( .A(B[3]), .B(A[3]), .Q(n49) );
  AOI211 U43 ( .A(n51), .B(n52), .C(n53), .Q(n50) );
  INV3 U44 ( .A(n55), .Q(n51) );
  NAND22 U45 ( .A(n45), .B(n46), .Q(n35) );
  NAND22 U46 ( .A(n18), .B(n19), .Q(n15) );
  XOR21 U47 ( .A(n4), .B(n5), .Q(SUM[7]) );
  AOI311 U48 ( .A(n6), .B(n7), .C(n8), .D(n9), .Q(n5) );
  NOR21 U49 ( .A(n17), .B(n47), .Q(n46) );
  NOR21 U50 ( .A(n29), .B(n27), .Q(n6) );
  NOR21 U51 ( .A(A[4]), .B(B[4]), .Q(n29) );
  NAND22 U52 ( .A(n39), .B(n40), .Q(n14) );
  NOR21 U53 ( .A(n43), .B(n44), .Q(n39) );
  INV3 U54 ( .A(A[1]), .Q(n43) );
  XNR21 U55 ( .A(n62), .B(n60), .Q(SUM[1]) );
  NOR21 U56 ( .A(n27), .B(n28), .Q(n12) );
  XOR21 U57 ( .A(n30), .B(n31), .Q(SUM[5]) );
  XOR21 U58 ( .A(n24), .B(n25), .Q(SUM[6]) );
  NAND22 U59 ( .A(n10), .B(n11), .Q(n9) );
  NAND22 U60 ( .A(n12), .B(n7), .Q(n10) );
  INV3 U61 ( .A(B[4]), .Q(n3) );
  XNR20 U62 ( .A(B[6]), .B(A[6]), .Q(n24) );
  XNR21 U63 ( .A(B[7]), .B(A[7]), .Q(n4) );
  AOI311 U64 ( .A(A[0]), .B(B[0]), .C(n58), .D(n59), .Q(n57) );
  NOR21 U65 ( .A(A[5]), .B(B[5]), .Q(n27) );
  XNR20 U66 ( .A(B[5]), .B(A[5]), .Q(n30) );
  XOR21 U67 ( .A(n49), .B(n50), .Q(SUM[3]) );
  NOR20 U68 ( .A(A[6]), .B(B[6]), .Q(n23) );
  NAND20 U69 ( .A(B[6]), .B(A[6]), .Q(n11) );
  CLKIN3 U70 ( .A(n14), .Q(n37) );
  CLKIN3 U71 ( .A(n61), .Q(n59) );
endmodule


module E_alu_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   ML_int_1__31_, ML_int_1__30_, ML_int_1__29_, ML_int_1__28_,
         ML_int_1__27_, ML_int_1__26_, ML_int_1__25_, ML_int_1__24_,
         ML_int_1__23_, ML_int_1__22_, ML_int_1__21_, ML_int_1__20_,
         ML_int_1__19_, ML_int_1__18_, ML_int_1__17_, ML_int_1__16_,
         ML_int_1__15_, ML_int_1__14_, ML_int_1__13_, ML_int_1__12_,
         ML_int_1__11_, ML_int_1__10_, ML_int_1__9_, ML_int_1__8_,
         ML_int_1__7_, ML_int_1__6_, ML_int_1__5_, ML_int_1__4_, ML_int_1__3_,
         ML_int_1__2_, ML_int_1__1_, ML_int_1__0_, ML_int_2__31_,
         ML_int_2__30_, ML_int_2__29_, ML_int_2__28_, ML_int_2__27_,
         ML_int_2__26_, ML_int_2__25_, ML_int_2__24_, ML_int_2__23_,
         ML_int_2__22_, ML_int_2__21_, ML_int_2__20_, ML_int_2__19_,
         ML_int_2__18_, ML_int_2__17_, ML_int_2__16_, ML_int_2__15_,
         ML_int_2__14_, ML_int_2__13_, ML_int_2__12_, ML_int_2__11_,
         ML_int_2__10_, ML_int_2__9_, ML_int_2__8_, ML_int_2__7_, ML_int_2__6_,
         ML_int_2__5_, ML_int_2__4_, ML_int_2__3_, ML_int_2__2_, ML_int_2__1_,
         ML_int_2__0_, ML_int_3__31_, ML_int_3__30_, ML_int_3__29_,
         ML_int_3__28_, ML_int_3__27_, ML_int_3__26_, ML_int_3__25_,
         ML_int_3__24_, ML_int_3__23_, ML_int_3__22_, ML_int_3__21_,
         ML_int_3__20_, ML_int_3__19_, ML_int_3__18_, ML_int_3__17_,
         ML_int_3__16_, ML_int_3__15_, ML_int_3__14_, ML_int_3__13_,
         ML_int_3__12_, ML_int_3__11_, ML_int_3__10_, ML_int_3__9_,
         ML_int_3__8_, ML_int_3__7_, ML_int_3__6_, ML_int_3__5_, ML_int_3__4_,
         ML_int_3__3_, ML_int_3__2_, ML_int_3__1_, ML_int_3__0_, ML_int_4__31_,
         ML_int_4__30_, ML_int_4__29_, ML_int_4__28_, ML_int_4__27_,
         ML_int_4__26_, ML_int_4__25_, ML_int_4__24_, ML_int_4__23_,
         ML_int_4__22_, ML_int_4__21_, ML_int_4__20_, ML_int_4__19_,
         ML_int_4__18_, ML_int_4__17_, ML_int_4__16_, ML_int_4__15_,
         ML_int_4__14_, ML_int_4__13_, ML_int_4__12_, ML_int_4__11_,
         ML_int_4__10_, ML_int_4__9_, ML_int_4__8_, ML_int_4__7_, ML_int_4__6_,
         ML_int_4__5_, ML_int_4__4_, ML_int_4__3_, ML_int_4__2_, ML_int_4__1_,
         ML_int_4__0_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53;

  MUX21 M1_0_2 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Q(ML_int_1__2_) );
  MUX21 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n34), .Q(ML_int_1__7_) );
  MUX21 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n32), .Q(ML_int_1__11_) );
  MUX21 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n32), .Q(ML_int_1__10_) );
  MUX21 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n35), .Q(ML_int_1__8_) );
  MUX21 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n32), .Q(ML_int_1__4_) );
  MUX21 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n35), .Q(ML_int_1__6_) );
  MUX21 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n32), .Q(ML_int_1__12_) );
  MUX21 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n33), .Q(ML_int_1__19_) );
  MUX21 M1_0_1 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Q(ML_int_1__1_) );
  MUX22 M1_1_13 ( .A(ML_int_1__13_), .B(ML_int_1__11_), .S(n38), .Q(
        ML_int_2__13_) );
  MUX21 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n33), .Q(ML_int_1__17_) );
  MUX21 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n33), .Q(ML_int_1__16_) );
  MUX22 M1_2_29 ( .A(ML_int_2__29_), .B(ML_int_2__25_), .S(n42), .Q(
        ML_int_3__29_) );
  MUX22 M1_3_29 ( .A(ML_int_3__29_), .B(ML_int_3__21_), .S(n49), .Q(
        ML_int_4__29_) );
  MUX22 M1_2_28 ( .A(ML_int_2__28_), .B(ML_int_2__24_), .S(n42), .Q(
        ML_int_3__28_) );
  MUX22 M1_4_28 ( .A(ML_int_4__28_), .B(ML_int_4__12_), .S(n51), .Q(B[28]) );
  MUX22 M1_1_31 ( .A(ML_int_1__31_), .B(ML_int_1__29_), .S(n37), .Q(
        ML_int_2__31_) );
  MUX22 M1_2_31 ( .A(ML_int_2__31_), .B(ML_int_2__27_), .S(n43), .Q(
        ML_int_3__31_) );
  MUX22 M1_3_27 ( .A(ML_int_3__27_), .B(ML_int_3__19_), .S(n49), .Q(
        ML_int_4__27_) );
  MUX22 M1_2_26 ( .A(ML_int_2__26_), .B(ML_int_2__22_), .S(n42), .Q(
        ML_int_3__26_) );
  MUX22 M1_3_26 ( .A(ML_int_3__26_), .B(ML_int_3__18_), .S(n49), .Q(
        ML_int_4__26_) );
  MUX22 M1_3_24 ( .A(ML_int_3__24_), .B(ML_int_3__16_), .S(n48), .Q(
        ML_int_4__24_) );
  MUX22 M1_3_20 ( .A(ML_int_3__20_), .B(ML_int_3__12_), .S(n48), .Q(
        ML_int_4__20_) );
  MUX22 M1_4_20 ( .A(ML_int_4__20_), .B(ML_int_4__4_), .S(n51), .Q(B[20]) );
  MUX22 M1_1_30 ( .A(ML_int_1__30_), .B(ML_int_1__28_), .S(n38), .Q(
        ML_int_2__30_) );
  MUX22 M1_2_30 ( .A(ML_int_2__30_), .B(ML_int_2__26_), .S(n43), .Q(
        ML_int_3__30_) );
  MUX22 M1_3_30 ( .A(ML_int_3__30_), .B(ML_int_3__22_), .S(n50), .Q(
        ML_int_4__30_) );
  MUX22 M1_4_30 ( .A(ML_int_4__30_), .B(ML_int_4__14_), .S(n51), .Q(B[30]) );
  MUX22 M1_2_25 ( .A(ML_int_2__25_), .B(ML_int_2__21_), .S(n42), .Q(
        ML_int_3__25_) );
  MUX22 M1_3_25 ( .A(ML_int_3__25_), .B(ML_int_3__17_), .S(n49), .Q(
        ML_int_4__25_) );
  MUX22 M1_4_25 ( .A(ML_int_4__25_), .B(ML_int_4__9_), .S(n51), .Q(B[25]) );
  MUX22 M1_4_17 ( .A(ML_int_4__17_), .B(ML_int_4__1_), .S(n52), .Q(B[17]) );
  MUX22 M1_3_16 ( .A(ML_int_3__16_), .B(ML_int_3__8_), .S(n47), .Q(
        ML_int_4__16_) );
  MUX22 M1_4_16 ( .A(ML_int_4__16_), .B(ML_int_4__0_), .S(n52), .Q(B[16]) );
  MUX22 M1_4_18 ( .A(ML_int_4__18_), .B(ML_int_4__2_), .S(n52), .Q(B[18]) );
  MUX21 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n32), .Q(ML_int_1__13_) );
  MUX22 M1_4_19 ( .A(ML_int_4__19_), .B(ML_int_4__3_), .S(n51), .Q(B[19]) );
  MUX22 M1_2_19 ( .A(ML_int_2__19_), .B(ML_int_2__15_), .S(n41), .Q(
        ML_int_3__19_) );
  MUX22 M1_1_10 ( .A(ML_int_1__10_), .B(ML_int_1__8_), .S(SH[1]), .Q(
        ML_int_2__10_) );
  MUX22 M1_3_12 ( .A(ML_int_3__12_), .B(ML_int_3__4_), .S(n46), .Q(
        ML_int_4__12_) );
  MUX22 M1_3_14 ( .A(ML_int_3__14_), .B(ML_int_3__6_), .S(n46), .Q(
        ML_int_4__14_) );
  MUX22 M1_3_13 ( .A(ML_int_3__13_), .B(ML_int_3__5_), .S(n46), .Q(
        ML_int_4__13_) );
  MUX22 M1_2_7 ( .A(ML_int_2__7_), .B(ML_int_2__3_), .S(n40), .Q(ML_int_3__7_)
         );
  MUX22 M1_3_11 ( .A(ML_int_3__11_), .B(ML_int_3__3_), .S(n46), .Q(
        ML_int_4__11_) );
  MUX22 M1_2_5 ( .A(ML_int_2__5_), .B(ML_int_2__1_), .S(n40), .Q(ML_int_3__5_)
         );
  MUX22 M1_3_8 ( .A(ML_int_3__8_), .B(ML_int_3__0_), .S(n45), .Q(ML_int_4__8_)
         );
  MUX22 M1_3_10 ( .A(ML_int_3__10_), .B(ML_int_3__2_), .S(n46), .Q(
        ML_int_4__10_) );
  MUX22 M1_2_11 ( .A(ML_int_2__11_), .B(ML_int_2__7_), .S(n43), .Q(
        ML_int_3__11_) );
  MUX22 M1_2_23 ( .A(ML_int_2__23_), .B(ML_int_2__19_), .S(n41), .Q(
        ML_int_3__23_) );
  MUX22 M1_1_24 ( .A(ML_int_1__24_), .B(ML_int_1__22_), .S(n38), .Q(
        ML_int_2__24_) );
  MUX22 M1_1_23 ( .A(ML_int_1__23_), .B(ML_int_1__21_), .S(n38), .Q(
        ML_int_2__23_) );
  MUX22 M1_1_27 ( .A(ML_int_1__27_), .B(ML_int_1__25_), .S(n38), .Q(
        ML_int_2__27_) );
  MUX22 M1_2_22 ( .A(ML_int_2__22_), .B(ML_int_2__18_), .S(n41), .Q(
        ML_int_3__22_) );
  MUX22 M1_1_26 ( .A(ML_int_1__26_), .B(ML_int_1__24_), .S(n37), .Q(
        ML_int_2__26_) );
  MUX22 M1_2_20 ( .A(ML_int_2__20_), .B(ML_int_2__16_), .S(n41), .Q(
        ML_int_3__20_) );
  MUX22 M1_2_21 ( .A(ML_int_2__21_), .B(ML_int_2__17_), .S(n41), .Q(
        ML_int_3__21_) );
  MUX22 M1_2_16 ( .A(ML_int_2__16_), .B(ML_int_2__12_), .S(SH[2]), .Q(
        ML_int_3__16_) );
  MUX22 M1_2_12 ( .A(ML_int_2__12_), .B(ML_int_2__8_), .S(n41), .Q(
        ML_int_3__12_) );
  MUX22 M1_1_22 ( .A(ML_int_1__22_), .B(ML_int_1__20_), .S(n38), .Q(
        ML_int_2__22_) );
  MUX22 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n35), .Q(ML_int_1__29_) );
  MUX22 M1_1_20 ( .A(ML_int_1__20_), .B(ML_int_1__18_), .S(n38), .Q(
        ML_int_2__20_) );
  MUX22 M1_2_13 ( .A(ML_int_2__13_), .B(ML_int_2__9_), .S(n42), .Q(
        ML_int_3__13_) );
  MUX22 M1_1_4 ( .A(ML_int_1__4_), .B(ML_int_1__2_), .S(n36), .Q(ML_int_2__4_)
         );
  MUX22 M1_1_3 ( .A(ML_int_1__3_), .B(ML_int_1__1_), .S(n36), .Q(ML_int_2__3_)
         );
  MUX22 M1_1_18 ( .A(ML_int_1__18_), .B(ML_int_1__16_), .S(n37), .Q(
        ML_int_2__18_) );
  MUX22 M1_1_16 ( .A(ML_int_1__16_), .B(ML_int_1__14_), .S(n37), .Q(
        ML_int_2__16_) );
  MUX22 M1_1_12 ( .A(ML_int_1__12_), .B(ML_int_1__10_), .S(SH[1]), .Q(
        ML_int_2__12_) );
  MUX22 M1_1_7 ( .A(ML_int_1__7_), .B(ML_int_1__5_), .S(n36), .Q(ML_int_2__7_)
         );
  MUX22 M1_2_8 ( .A(ML_int_2__8_), .B(ML_int_2__4_), .S(n40), .Q(ML_int_3__8_)
         );
  MUX22 M1_1_11 ( .A(ML_int_1__11_), .B(ML_int_1__9_), .S(n36), .Q(
        ML_int_2__11_) );
  MUX22 M1_2_10 ( .A(ML_int_2__10_), .B(ML_int_2__6_), .S(n42), .Q(
        ML_int_3__10_) );
  MUX22 M1_3_23 ( .A(ML_int_3__23_), .B(ML_int_3__15_), .S(n48), .Q(
        ML_int_4__23_) );
  MUX22 M1_4_23 ( .A(ML_int_4__23_), .B(ML_int_4__7_), .S(n51), .Q(B[23]) );
  MUX21 M1_3_19 ( .A(ML_int_3__19_), .B(ML_int_3__11_), .S(n47), .Q(
        ML_int_4__19_) );
  MUX21 M1_3_17 ( .A(ML_int_3__17_), .B(ML_int_3__9_), .S(n47), .Q(
        ML_int_4__17_) );
  MUX21 M1_3_31 ( .A(ML_int_3__31_), .B(ML_int_3__23_), .S(n50), .Q(
        ML_int_4__31_) );
  MUX21 M1_4_31 ( .A(ML_int_4__31_), .B(ML_int_4__15_), .S(n51), .Q(B[31]) );
  MUX21 M1_2_27 ( .A(ML_int_2__27_), .B(ML_int_2__23_), .S(n42), .Q(
        ML_int_3__27_) );
  MUX21 M1_4_27 ( .A(ML_int_4__27_), .B(ML_int_4__11_), .S(n51), .Q(B[27]) );
  MUX21 M1_4_26 ( .A(ML_int_4__26_), .B(ML_int_4__10_), .S(n51), .Q(B[26]) );
  MUX21 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n34), .Q(ML_int_1__30_) );
  MUX21 M1_3_18 ( .A(ML_int_3__18_), .B(ML_int_3__10_), .S(n47), .Q(
        ML_int_4__18_) );
  MUX21 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n33), .Q(ML_int_1__15_) );
  MUX21 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n34), .Q(ML_int_1__22_) );
  MUX21 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n35), .Q(ML_int_1__25_) );
  MUX21 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n33), .Q(ML_int_1__18_) );
  MUX21 M1_1_9 ( .A(ML_int_1__9_), .B(ML_int_1__7_), .S(SH[1]), .Q(
        ML_int_2__9_) );
  MUX21 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n35), .Q(ML_int_1__28_) );
  MUX21 M1_1_5 ( .A(ML_int_1__5_), .B(ML_int_1__3_), .S(SH[1]), .Q(
        ML_int_2__5_) );
  MUX21 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n35), .Q(ML_int_1__26_) );
  MUX21 M1_1_8 ( .A(ML_int_1__8_), .B(ML_int_1__6_), .S(n37), .Q(ML_int_2__8_)
         );
  MUX21 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n34), .Q(ML_int_1__24_) );
  MUX21 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n34), .Q(ML_int_1__23_) );
  MUX21 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n32), .Q(ML_int_1__14_) );
  MUX21 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n34), .Q(ML_int_1__21_) );
  MUX21 M1_1_2 ( .A(ML_int_1__2_), .B(ML_int_1__0_), .S(n36), .Q(ML_int_2__2_)
         );
  MUX22 M1_2_24 ( .A(ML_int_2__24_), .B(ML_int_2__20_), .S(n41), .Q(
        ML_int_3__24_) );
  MUX22 M1_3_22 ( .A(ML_int_3__22_), .B(ML_int_3__14_), .S(n48), .Q(
        ML_int_4__22_) );
  MUX22 M1_4_22 ( .A(ML_int_4__22_), .B(ML_int_4__6_), .S(n51), .Q(B[22]) );
  MUX22 M1_2_9 ( .A(ML_int_2__9_), .B(ML_int_2__5_), .S(n40), .Q(ML_int_3__9_)
         );
  MUX22 M1_2_17 ( .A(ML_int_2__17_), .B(ML_int_2__13_), .S(n39), .Q(
        ML_int_3__17_) );
  MUX22 M1_2_15 ( .A(ML_int_2__15_), .B(ML_int_2__11_), .S(n43), .Q(
        ML_int_3__15_) );
  MUX22 M1_1_25 ( .A(ML_int_1__25_), .B(ML_int_1__23_), .S(n38), .Q(
        ML_int_2__25_) );
  MUX22 M1_3_15 ( .A(ML_int_3__15_), .B(ML_int_3__7_), .S(n47), .Q(
        ML_int_4__15_) );
  MUX22 M1_1_21 ( .A(ML_int_1__21_), .B(ML_int_1__19_), .S(n38), .Q(
        ML_int_2__21_) );
  MUX22 M1_3_9 ( .A(ML_int_3__9_), .B(ML_int_3__1_), .S(n45), .Q(ML_int_4__9_)
         );
  MUX22 M1_2_4 ( .A(ML_int_2__4_), .B(ML_int_2__0_), .S(n39), .Q(ML_int_3__4_)
         );
  MUX22 M1_4_24 ( .A(ML_int_4__24_), .B(ML_int_4__8_), .S(n51), .Q(B[24]) );
  MUX22 M1_3_28 ( .A(ML_int_3__28_), .B(ML_int_3__20_), .S(n49), .Q(
        ML_int_4__28_) );
  MUX21 M1_1_17 ( .A(ML_int_1__17_), .B(ML_int_1__15_), .S(n37), .Q(
        ML_int_2__17_) );
  MUX21 M1_2_6 ( .A(ML_int_2__6_), .B(ML_int_2__2_), .S(n40), .Q(ML_int_3__6_)
         );
  MUX22 M1_1_14 ( .A(ML_int_1__14_), .B(ML_int_1__12_), .S(SH[1]), .Q(
        ML_int_2__14_) );
  MUX22 M1_2_18 ( .A(ML_int_2__18_), .B(ML_int_2__14_), .S(n43), .Q(
        ML_int_3__18_) );
  MUX22 M1_1_6 ( .A(ML_int_1__6_), .B(ML_int_1__4_), .S(SH[1]), .Q(
        ML_int_2__6_) );
  MUX22 M1_2_14 ( .A(ML_int_2__14_), .B(ML_int_2__10_), .S(n41), .Q(
        ML_int_3__14_) );
  MUX21 M1_4_29 ( .A(ML_int_4__29_), .B(ML_int_4__13_), .S(n51), .Q(B[29]) );
  MUX22 M1_1_28 ( .A(ML_int_1__28_), .B(ML_int_1__26_), .S(n38), .Q(
        ML_int_2__28_) );
  MUX21 M1_3_21 ( .A(ML_int_3__21_), .B(ML_int_3__13_), .S(n48), .Q(
        ML_int_4__21_) );
  MUX22 M1_4_21 ( .A(ML_int_4__21_), .B(ML_int_4__5_), .S(n51), .Q(B[21]) );
  MUX21 M1_1_19 ( .A(ML_int_1__19_), .B(ML_int_1__17_), .S(n37), .Q(
        ML_int_2__19_) );
  MUX21 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n33), .Q(ML_int_1__3_) );
  MUX22 M1_1_29 ( .A(ML_int_1__29_), .B(ML_int_1__27_), .S(n37), .Q(
        ML_int_2__29_) );
  MUX21 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n32), .Q(ML_int_1__9_) );
  MUX22 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n35), .Q(ML_int_1__31_) );
  MUX22 M1_1_15 ( .A(ML_int_1__15_), .B(ML_int_1__13_), .S(n37), .Q(
        ML_int_2__15_) );
  MUX22 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n35), .Q(ML_int_1__27_) );
  MUX21 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n34), .Q(ML_int_1__20_) );
  MUX22 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n33), .Q(ML_int_1__5_) );
  NOR22 U3 ( .A(n36), .B(n29), .Q(ML_int_2__0_) );
  INV3 U4 ( .A(ML_int_2__1_), .Q(n27) );
  CLKIN3 U5 ( .A(ML_int_3__1_), .Q(n23) );
  CLKIN3 U6 ( .A(ML_int_4__15_), .Q(n1) );
  INV1 U7 ( .A(ML_int_1__1_), .Q(n31) );
  INV1 U8 ( .A(ML_int_4__7_), .Q(n9) );
  INV3 U9 ( .A(ML_int_2__3_), .Q(n25) );
  INV3 U10 ( .A(ML_int_3__5_), .Q(n19) );
  INV2 U11 ( .A(ML_int_4__4_), .Q(n12) );
  INV2 U12 ( .A(ML_int_4__0_), .Q(n16) );
  INV2 U13 ( .A(ML_int_1__0_), .Q(n29) );
  INV2 U14 ( .A(ML_int_3__0_), .Q(n24) );
  INV2 U15 ( .A(ML_int_3__2_), .Q(n22) );
  INV2 U16 ( .A(ML_int_4__1_), .Q(n15) );
  INV2 U17 ( .A(ML_int_2__2_), .Q(n26) );
  INV2 U18 ( .A(ML_int_4__2_), .Q(n14) );
  NOR22 U19 ( .A(n39), .B(n25), .Q(ML_int_3__3_) );
  INV0 U20 ( .A(ML_int_3__3_), .Q(n21) );
  INV2 U21 ( .A(ML_int_4__5_), .Q(n11) );
  INV2 U22 ( .A(ML_int_4__3_), .Q(n13) );
  BUF2 U23 ( .A(SH[4]), .Q(n51) );
  NOR21 U24 ( .A(n52), .B(n6), .Q(B[10]) );
  INV3 U25 ( .A(ML_int_4__10_), .Q(n6) );
  NOR21 U26 ( .A(n36), .B(n31), .Q(ML_int_2__1_) );
  NOR21 U27 ( .A(n34), .B(n30), .Q(ML_int_1__0_) );
  INV3 U28 ( .A(A[0]), .Q(n30) );
  NOR21 U29 ( .A(n45), .B(n19), .Q(ML_int_4__5_) );
  NOR21 U30 ( .A(n45), .B(n18), .Q(ML_int_4__6_) );
  INV3 U31 ( .A(ML_int_3__6_), .Q(n18) );
  NOR21 U32 ( .A(n45), .B(n17), .Q(ML_int_4__7_) );
  INV3 U33 ( .A(ML_int_3__7_), .Q(n17) );
  NOR21 U34 ( .A(n39), .B(n28), .Q(ML_int_3__0_) );
  INV3 U35 ( .A(ML_int_2__0_), .Q(n28) );
  NOR21 U36 ( .A(n39), .B(n27), .Q(ML_int_3__1_) );
  NOR21 U37 ( .A(n39), .B(n26), .Q(ML_int_3__2_) );
  NOR21 U38 ( .A(n44), .B(n24), .Q(ML_int_4__0_) );
  NOR21 U39 ( .A(n44), .B(n23), .Q(ML_int_4__1_) );
  NOR21 U40 ( .A(n44), .B(n22), .Q(ML_int_4__2_) );
  NOR21 U41 ( .A(n44), .B(n20), .Q(ML_int_4__4_) );
  INV3 U42 ( .A(ML_int_3__4_), .Q(n20) );
  NOR21 U43 ( .A(n44), .B(n21), .Q(ML_int_4__3_) );
  NOR21 U44 ( .A(n52), .B(n1), .Q(B[15]) );
  NOR21 U45 ( .A(n53), .B(n16), .Q(B[0]) );
  NOR21 U46 ( .A(n52), .B(n5), .Q(B[11]) );
  INV3 U47 ( .A(ML_int_4__11_), .Q(n5) );
  NOR21 U48 ( .A(n52), .B(n9), .Q(B[7]) );
  NOR21 U49 ( .A(n52), .B(n3), .Q(B[13]) );
  INV3 U50 ( .A(ML_int_4__13_), .Q(n3) );
  NOR21 U51 ( .A(n52), .B(n10), .Q(B[6]) );
  INV3 U52 ( .A(ML_int_4__6_), .Q(n10) );
  NOR21 U53 ( .A(n52), .B(n8), .Q(B[8]) );
  INV3 U54 ( .A(ML_int_4__8_), .Q(n8) );
  NOR21 U55 ( .A(n52), .B(n7), .Q(B[9]) );
  INV3 U56 ( .A(ML_int_4__9_), .Q(n7) );
  NOR21 U57 ( .A(n52), .B(n4), .Q(B[12]) );
  INV3 U58 ( .A(ML_int_4__12_), .Q(n4) );
  NOR21 U59 ( .A(n52), .B(n2), .Q(B[14]) );
  INV3 U60 ( .A(ML_int_4__14_), .Q(n2) );
  NOR21 U61 ( .A(n53), .B(n15), .Q(B[1]) );
  NOR21 U62 ( .A(n53), .B(n13), .Q(B[3]) );
  NOR21 U63 ( .A(n53), .B(n12), .Q(B[4]) );
  NOR21 U64 ( .A(n53), .B(n11), .Q(B[5]) );
  NOR21 U65 ( .A(n53), .B(n14), .Q(B[2]) );
  BUF2 U66 ( .A(SH[0]), .Q(n35) );
  BUF2 U67 ( .A(SH[1]), .Q(n37) );
  BUF2 U68 ( .A(SH[1]), .Q(n38) );
  BUF2 U69 ( .A(SH[1]), .Q(n36) );
  BUF2 U70 ( .A(SH[0]), .Q(n34) );
  BUF2 U71 ( .A(SH[0]), .Q(n32) );
  BUF2 U72 ( .A(SH[0]), .Q(n33) );
  BUF2 U73 ( .A(SH[4]), .Q(n52) );
  BUF2 U74 ( .A(SH[4]), .Q(n53) );
  BUF2 U75 ( .A(SH[3]), .Q(n46) );
  BUF2 U76 ( .A(SH[3]), .Q(n48) );
  BUF2 U77 ( .A(SH[3]), .Q(n49) );
  BUF2 U78 ( .A(SH[2]), .Q(n41) );
  BUF2 U79 ( .A(SH[2]), .Q(n42) );
  BUF2 U80 ( .A(SH[3]), .Q(n47) );
  BUF2 U81 ( .A(SH[2]), .Q(n40) );
  BUF2 U82 ( .A(SH[3]), .Q(n45) );
  BUF2 U83 ( .A(SH[2]), .Q(n39) );
  BUF2 U84 ( .A(SH[3]), .Q(n44) );
  BUF2 U85 ( .A(SH[3]), .Q(n50) );
  BUF2 U86 ( .A(SH[2]), .Q(n43) );
endmodule


module E_alu_DW01_add_18 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89;

  CLKIN1 U2 ( .A(A[0]), .Q(n9) );
  NAND20 U3 ( .A(B[0]), .B(A[0]), .Q(n24) );
  NAND20 U4 ( .A(B[0]), .B(A[0]), .Q(n86) );
  NOR22 U5 ( .A(n2), .B(n19), .Q(n17) );
  AOI212 U6 ( .A(n49), .B(n58), .C(n55), .Q(n57) );
  NAND22 U7 ( .A(n78), .B(n7), .Q(n32) );
  AOI311 U8 ( .A(n21), .B(B[5]), .C(A[5]), .D(n38), .Q(n37) );
  NAND22 U9 ( .A(n29), .B(n30), .Q(n22) );
  NAND26 U10 ( .A(n13), .B(n12), .Q(SUM[8]) );
  NAND24 U11 ( .A(n62), .B(n63), .Q(n21) );
  INV3 U12 ( .A(n21), .Q(n36) );
  INV1 U13 ( .A(B[0]), .Q(n6) );
  XOR21 U14 ( .A(n40), .B(n41), .Q(SUM[7]) );
  CLKIN3 U15 ( .A(n32), .Q(n47) );
  INV2 U16 ( .A(A[2]), .Q(n11) );
  NOR21 U17 ( .A(n7), .B(n10), .Q(n23) );
  NOR21 U18 ( .A(B[7]), .B(A[7]), .Q(n19) );
  CLKIN3 U19 ( .A(n11), .Q(n10) );
  INV6 U20 ( .A(n8), .Q(n7) );
  AOI211 U21 ( .A(n65), .B(n58), .C(n66), .Q(n64) );
  NAND22 U22 ( .A(n88), .B(n89), .Q(n30) );
  INV2 U23 ( .A(n30), .Q(n5) );
  OAI212 U24 ( .A(n7), .B(n10), .C(n26), .Q(n25) );
  NOR21 U25 ( .A(n20), .B(n36), .Q(n16) );
  INV2 U26 ( .A(B[6]), .Q(n62) );
  NOR21 U27 ( .A(n28), .B(n11), .Q(n78) );
  NAND21 U28 ( .A(B[3]), .B(A[3]), .Q(n31) );
  INV1 U29 ( .A(B[1]), .Q(n88) );
  NOR21 U30 ( .A(A[5]), .B(B[5]), .Q(n18) );
  NAND22 U31 ( .A(B[1]), .B(A[1]), .Q(n27) );
  NOR24 U32 ( .A(A[3]), .B(B[3]), .Q(n28) );
  BUF6 U33 ( .A(n27), .Q(n1) );
  BUF6 U34 ( .A(n18), .Q(n2) );
  NAND22 U35 ( .A(B[4]), .B(A[4]), .Q(n35) );
  NOR21 U36 ( .A(n77), .B(n47), .Q(n71) );
  INV1 U37 ( .A(n60), .Q(n68) );
  INV3 U38 ( .A(n55), .Q(n44) );
  XOR22 U39 ( .A(n56), .B(n57), .Q(SUM[6]) );
  XOR20 U40 ( .A(n87), .B(n86), .Q(SUM[1]) );
  CLKIN3 U41 ( .A(n43), .Q(n38) );
  NAND20 U42 ( .A(B[0]), .B(A[0]), .Q(n52) );
  IMUX20 U43 ( .A(n6), .B(B[0]), .S(A[0]), .Q(SUM[0]) );
  NAND33 U44 ( .A(n73), .B(n74), .C(n75), .Q(n72) );
  NOR20 U45 ( .A(n9), .B(n6), .Q(n75) );
  CLKIN0 U46 ( .A(n61), .Q(n65) );
  OAI312 U47 ( .A(n22), .B(n23), .C(n24), .D(n25), .Q(n15) );
  IMUX20 U48 ( .A(n69), .B(n70), .S(n58), .Q(SUM[4]) );
  NOR20 U49 ( .A(B[4]), .B(A[4]), .Q(n79) );
  CLKIN3 U50 ( .A(n39), .Q(n33) );
  INV3 U51 ( .A(n76), .Q(n74) );
  XNR21 U52 ( .A(n85), .B(n4), .Q(SUM[2]) );
  XNR21 U53 ( .A(n67), .B(n64), .Q(SUM[5]) );
  NOR21 U54 ( .A(n2), .B(n61), .Q(n49) );
  NAND20 U55 ( .A(A[4]), .B(B[4]), .Q(n59) );
  OAI311 U56 ( .A(n46), .B(n47), .C(n48), .D(n49), .Q(n45) );
  INV3 U57 ( .A(n31), .Q(n48) );
  OAI311 U58 ( .A(n50), .B(n51), .C(n52), .D(n53), .Q(n46) );
  NAND20 U59 ( .A(B[4]), .B(A[4]), .Q(n80) );
  NAND20 U60 ( .A(B[5]), .B(A[5]), .Q(n60) );
  NOR20 U61 ( .A(A[4]), .B(B[4]), .Q(n61) );
  NOR21 U62 ( .A(n79), .B(n66), .Q(n70) );
  XNR20 U63 ( .A(B[4]), .B(A[4]), .Q(n69) );
  NAND22 U64 ( .A(n31), .B(n32), .Q(n14) );
  NAND22 U65 ( .A(n30), .B(n1), .Q(n87) );
  NAND22 U66 ( .A(n29), .B(n30), .Q(n50) );
  OAI212 U67 ( .A(n86), .B(n5), .C(n1), .Q(n4) );
  NOR20 U68 ( .A(B[4]), .B(A[4]), .Q(n20) );
  INV3 U69 ( .A(B[2]), .Q(n8) );
  XOR21 U70 ( .A(n81), .B(n82), .Q(SUM[3]) );
  AOI211 U71 ( .A(n74), .B(n4), .C(n83), .Q(n82) );
  INV3 U72 ( .A(A[6]), .Q(n63) );
  OAI210 U73 ( .A(n7), .B(n10), .C(n84), .Q(n85) );
  NAND22 U74 ( .A(n7), .B(n10), .Q(n84) );
  NOR21 U75 ( .A(n7), .B(n10), .Q(n76) );
  NOR21 U76 ( .A(n7), .B(n10), .Q(n51) );
  CLKIN2 U77 ( .A(n28), .Q(n29) );
  AOI2110 U78 ( .A(n11), .B(n8), .C(n1), .D(n28), .Q(n77) );
  NOR21 U79 ( .A(n5), .B(n28), .Q(n73) );
  NOR20 U80 ( .A(n1), .B(n28), .Q(n54) );
  NOR21 U81 ( .A(n1), .B(n28), .Q(n26) );
  NAND20 U82 ( .A(n21), .B(n43), .Q(n56) );
  NAND22 U83 ( .A(B[6]), .B(A[6]), .Q(n43) );
  AOI211 U84 ( .A(n42), .B(n21), .C(n38), .Q(n41) );
  NAND22 U85 ( .A(n44), .B(n45), .Q(n42) );
  NOR20 U86 ( .A(n68), .B(n2), .Q(n67) );
  AOI222 U87 ( .A(B[7]), .B(A[7]), .C(n33), .D(n34), .Q(n12) );
  XNR20 U88 ( .A(B[7]), .B(A[7]), .Q(n40) );
  NOR21 U89 ( .A(A[7]), .B(B[7]), .Q(n39) );
  INV3 U90 ( .A(A[1]), .Q(n89) );
  XNR20 U91 ( .A(B[3]), .B(A[3]), .Q(n81) );
  OAI2112 U92 ( .A(n14), .B(n15), .C(n16), .D(n17), .Q(n13) );
  OAI312 U93 ( .A(n35), .B(n2), .C(n36), .D(n37), .Q(n34) );
  OAI212 U94 ( .A(n7), .B(n10), .C(n54), .Q(n53) );
  OAI212 U95 ( .A(n2), .B(n59), .C(n60), .Q(n55) );
  NAND33 U96 ( .A(n71), .B(n72), .C(n31), .Q(n58) );
  CLKIN3 U97 ( .A(n80), .Q(n66) );
  CLKIN3 U98 ( .A(n84), .Q(n83) );
endmodule


module E_alu_DW01_add_17 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106;

  OAI312 U2 ( .A(n47), .B(n48), .C(n49), .D(n50), .Q(n46) );
  NOR21 U3 ( .A(n2), .B(n5), .Q(n56) );
  INV6 U4 ( .A(n3), .Q(n2) );
  NOR22 U5 ( .A(A[5]), .B(B[5]), .Q(n13) );
  NOR20 U6 ( .A(A[0]), .B(B[0]), .Q(n101) );
  CLKIN6 U7 ( .A(n25), .Q(n82) );
  IMUX21 U8 ( .A(n74), .B(n75), .S(n63), .Q(SUM[4]) );
  NOR21 U9 ( .A(n2), .B(n5), .Q(n87) );
  INV6 U10 ( .A(n6), .Q(n5) );
  NOR21 U11 ( .A(n4), .B(n1), .Q(n86) );
  INV1 U12 ( .A(A[0]), .Q(n4) );
  INV3 U13 ( .A(B[0]), .Q(n1) );
  NOR21 U14 ( .A(B[0]), .B(A[0]), .Q(n31) );
  XOR21 U15 ( .A(n41), .B(n42), .Q(SUM[7]) );
  AOI211 U16 ( .A(n43), .B(n16), .C(n39), .Q(n42) );
  NAND22 U17 ( .A(B[1]), .B(A[1]), .Q(n22) );
  NAND21 U18 ( .A(n24), .B(n25), .Q(n55) );
  NAND21 U19 ( .A(n54), .B(n25), .Q(n51) );
  NAND26 U20 ( .A(n7), .B(n8), .Q(SUM[8]) );
  INV3 U21 ( .A(A[2]), .Q(n6) );
  NAND24 U22 ( .A(n104), .B(n105), .Q(n25) );
  NAND33 U23 ( .A(n76), .B(n77), .C(n78), .Q(n63) );
  XOR21 U24 ( .A(n92), .B(n93), .Q(SUM[3]) );
  AOI211 U25 ( .A(n85), .B(n94), .C(n95), .Q(n93) );
  OAI311 U26 ( .A(n55), .B(n56), .C(n57), .D(n58), .Q(n47) );
  NOR31 U27 ( .A(n31), .B(n82), .C(n32), .Q(n80) );
  OAI311 U28 ( .A(n17), .B(n18), .C(n19), .D(n20), .Q(n10) );
  NOR22 U29 ( .A(n88), .B(n48), .Q(n76) );
  NOR23 U30 ( .A(A[3]), .B(B[3]), .Q(n23) );
  NAND22 U31 ( .A(n89), .B(n2), .Q(n29) );
  INV3 U32 ( .A(n29), .Q(n48) );
  NAND22 U33 ( .A(n67), .B(n68), .Q(n16) );
  AOI2111 U34 ( .A(n6), .B(n3), .C(n22), .D(n23), .Q(n88) );
  AOI221 U35 ( .A(B[7]), .B(A[7]), .C(n33), .D(n34), .Q(n7) );
  NOR22 U36 ( .A(n23), .B(n6), .Q(n89) );
  OAI2112 U37 ( .A(n9), .B(n10), .C(n11), .D(n12), .Q(n8) );
  OAI2112 U38 ( .A(n26), .B(n27), .C(n28), .D(n29), .Q(n9) );
  INV1 U39 ( .A(B[1]), .Q(n104) );
  NAND20 U40 ( .A(n101), .B(n19), .Q(n103) );
  NAND22 U41 ( .A(n19), .B(n101), .Q(n99) );
  CLKIN2 U42 ( .A(n83), .Q(n79) );
  AOI212 U43 ( .A(n50), .B(n63), .C(n60), .Q(n62) );
  INV3 U44 ( .A(n98), .Q(n94) );
  NAND20 U45 ( .A(n25), .B(n22), .Q(n102) );
  NOR20 U46 ( .A(n2), .B(n5), .Q(n53) );
  NOR20 U47 ( .A(B[0]), .B(A[0]), .Q(n52) );
  NAND20 U48 ( .A(n2), .B(n5), .Q(n96) );
  NAND20 U49 ( .A(B[0]), .B(A[0]), .Q(n57) );
  NOR20 U50 ( .A(n2), .B(n5), .Q(n83) );
  NAND33 U51 ( .A(n84), .B(n85), .C(n86), .Q(n77) );
  NOR20 U52 ( .A(n73), .B(n13), .Q(n72) );
  CLKIN0 U53 ( .A(n66), .Q(n70) );
  CLKIN2 U54 ( .A(n40), .Q(n33) );
  NAND20 U55 ( .A(n16), .B(n44), .Q(n61) );
  NOR20 U56 ( .A(B[4]), .B(A[4]), .Q(n90) );
  XOR21 U57 ( .A(n97), .B(n98), .Q(SUM[2]) );
  NAND22 U58 ( .A(n106), .B(n19), .Q(SUM[0]) );
  NAND22 U59 ( .A(n4), .B(n1), .Q(n106) );
  INV3 U60 ( .A(n87), .Q(n85) );
  XNR21 U61 ( .A(n72), .B(n69), .Q(SUM[5]) );
  NOR21 U62 ( .A(n13), .B(n66), .Q(n50) );
  INV3 U63 ( .A(n60), .Q(n45) );
  NAND20 U64 ( .A(A[4]), .B(B[4]), .Q(n64) );
  NAND22 U65 ( .A(n54), .B(n25), .Q(n26) );
  CLKIN3 U66 ( .A(n31), .Q(n30) );
  OAI311 U67 ( .A(n51), .B(n52), .C(n53), .D(n28), .Q(n49) );
  OAI311 U68 ( .A(n35), .B(n36), .C(n37), .D(n38), .Q(n34) );
  NOR21 U69 ( .A(A[5]), .B(B[5]), .Q(n36) );
  NAND20 U70 ( .A(B[4]), .B(A[4]), .Q(n35) );
  INV3 U71 ( .A(n16), .Q(n37) );
  NAND22 U72 ( .A(B[0]), .B(A[0]), .Q(n19) );
  NOR21 U73 ( .A(n2), .B(n5), .Q(n18) );
  NAND22 U74 ( .A(n24), .B(n25), .Q(n17) );
  AOI311 U75 ( .A(n16), .B(B[5]), .C(A[5]), .D(n39), .Q(n38) );
  NOR20 U76 ( .A(A[4]), .B(B[4]), .Q(n66) );
  NAND22 U77 ( .A(B[5]), .B(A[5]), .Q(n65) );
  NOR21 U78 ( .A(n90), .B(n71), .Q(n75) );
  XNR20 U79 ( .A(B[4]), .B(A[4]), .Q(n74) );
  XNR21 U80 ( .A(n102), .B(n103), .Q(SUM[1]) );
  NAND20 U81 ( .A(B[4]), .B(A[4]), .Q(n91) );
  NOR21 U82 ( .A(n13), .B(n14), .Q(n12) );
  NAND22 U83 ( .A(n45), .B(n46), .Q(n43) );
  INV3 U84 ( .A(n23), .Q(n24) );
  AOI211 U85 ( .A(n99), .B(n25), .C(n100), .Q(n98) );
  INV3 U86 ( .A(n22), .Q(n100) );
  NOR21 U87 ( .A(n15), .B(n37), .Q(n11) );
  NOR20 U88 ( .A(B[4]), .B(A[4]), .Q(n15) );
  INV3 U89 ( .A(B[2]), .Q(n3) );
  INV3 U90 ( .A(A[6]), .Q(n68) );
  INV3 U91 ( .A(B[6]), .Q(n67) );
  NAND22 U92 ( .A(B[6]), .B(A[6]), .Q(n44) );
  OAI222 U93 ( .A(n79), .B(n81), .C(n80), .D(n81), .Q(n78) );
  OAI212 U94 ( .A(n2), .B(n5), .C(n30), .Q(n27) );
  NOR21 U95 ( .A(B[3]), .B(A[3]), .Q(n32) );
  NAND21 U96 ( .A(B[3]), .B(A[3]), .Q(n28) );
  XNR20 U97 ( .A(B[7]), .B(A[7]), .Q(n41) );
  NOR21 U98 ( .A(B[7]), .B(A[7]), .Q(n14) );
  NOR21 U99 ( .A(A[7]), .B(B[7]), .Q(n40) );
  NOR21 U100 ( .A(n82), .B(n23), .Q(n84) );
  NOR21 U101 ( .A(n22), .B(n23), .Q(n59) );
  NOR21 U102 ( .A(n22), .B(n23), .Q(n21) );
  INV3 U103 ( .A(A[1]), .Q(n105) );
  INV2 U104 ( .A(n32), .Q(n54) );
  XNR20 U105 ( .A(B[3]), .B(A[3]), .Q(n92) );
  OAI212 U106 ( .A(n2), .B(n5), .C(n21), .Q(n20) );
  CLKIN3 U107 ( .A(n44), .Q(n39) );
  OAI212 U108 ( .A(n2), .B(n5), .C(n59), .Q(n58) );
  XOR22 U109 ( .A(n61), .B(n62), .Q(SUM[6]) );
  OAI212 U110 ( .A(n13), .B(n64), .C(n65), .Q(n60) );
  AOI212 U111 ( .A(n70), .B(n63), .C(n71), .Q(n69) );
  CLKIN3 U112 ( .A(n65), .Q(n73) );
  CLKIN3 U113 ( .A(n28), .Q(n81) );
  CLKIN3 U114 ( .A(n91), .Q(n71) );
  CLKIN3 U115 ( .A(n96), .Q(n95) );
  OAI212 U116 ( .A(n2), .B(n5), .C(n96), .Q(n97) );
endmodule


module E_alu_DW01_cmp2_2 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271;

  AOI312 U1 ( .A(n43), .B(n44), .C(n45), .D(n33), .Q(n42) );
  INV0 U2 ( .A(A[10]), .Q(n16) );
  INV2 U3 ( .A(n98), .Q(n94) );
  NAND22 U4 ( .A(n161), .B(n162), .Q(n110) );
  INV3 U5 ( .A(n104), .Q(n141) );
  INV3 U6 ( .A(n115), .Q(n109) );
  INV8 U7 ( .A(n266), .Q(n106) );
  NAND22 U8 ( .A(A[17]), .B(n228), .Q(n105) );
  NAND21 U9 ( .A(n252), .B(n229), .Q(n215) );
  NAND21 U10 ( .A(B[9]), .B(n252), .Q(n251) );
  CLKIN0 U11 ( .A(B[11]), .Q(n4) );
  NAND42 U12 ( .A(n104), .B(n105), .C(n119), .D(n120), .Q(n118) );
  NAND20 U13 ( .A(A[9]), .B(n163), .Q(n161) );
  INV3 U14 ( .A(B[5]), .Q(n73) );
  NAND42 U15 ( .A(n131), .B(n132), .C(n125), .D(n133), .Q(n39) );
  CLKIN4 U16 ( .A(n106), .Q(n125) );
  NAND20 U17 ( .A(n174), .B(n115), .Q(n171) );
  NAND41 U18 ( .A(n115), .B(n116), .C(n117), .D(B[7]), .Q(n113) );
  NAND20 U19 ( .A(n116), .B(n115), .Q(n134) );
  NAND24 U20 ( .A(A[25]), .B(n260), .Q(n115) );
  NAND24 U21 ( .A(n257), .B(n182), .Q(n119) );
  NAND22 U22 ( .A(A[15]), .B(n130), .Q(n138) );
  NAND22 U23 ( .A(B[23]), .B(n258), .Q(n182) );
  NAND22 U24 ( .A(n46), .B(n30), .Q(n33) );
  INV3 U25 ( .A(B[23]), .Q(n10) );
  NOR21 U26 ( .A(A[22]), .B(n103), .Q(n225) );
  INV2 U27 ( .A(B[27]), .Q(n13) );
  INV3 U28 ( .A(n119), .Q(n102) );
  INV3 U29 ( .A(n116), .Q(n103) );
  INV3 U30 ( .A(n1), .Q(n157) );
  NAND22 U31 ( .A(n153), .B(n138), .Q(n253) );
  INV3 U32 ( .A(B[25]), .Q(n260) );
  NOR22 U33 ( .A(n37), .B(n38), .Q(n21) );
  INV3 U34 ( .A(B[10]), .Q(n3) );
  NOR21 U35 ( .A(n250), .B(n251), .Q(n249) );
  NOR21 U36 ( .A(n109), .B(n103), .Q(n256) );
  NOR21 U37 ( .A(n220), .B(n221), .Q(n219) );
  NAND23 U38 ( .A(A[26]), .B(n12), .Q(n174) );
  NOR31 U39 ( .A(n109), .B(n103), .C(n3), .Q(n200) );
  NAND22 U40 ( .A(A[27]), .B(n13), .Q(n173) );
  NOR21 U41 ( .A(n106), .B(n107), .Q(n43) );
  NAND31 U42 ( .A(n124), .B(n125), .C(n126), .Q(n40) );
  NOR21 U43 ( .A(n146), .B(n147), .Q(n145) );
  NOR31 U44 ( .A(n155), .B(n106), .C(n156), .Q(n146) );
  NOR31 U45 ( .A(n148), .B(n106), .C(n149), .Q(n147) );
  NOR22 U46 ( .A(n212), .B(n213), .Q(n19) );
  INV1 U47 ( .A(B[20]), .Q(n8) );
  NAND41 U48 ( .A(n104), .B(n105), .C(n119), .D(n201), .Q(n195) );
  NAND41 U49 ( .A(n105), .B(n60), .C(n104), .D(n262), .Q(n261) );
  NOR21 U50 ( .A(n263), .B(n264), .Q(n262) );
  INV0 U51 ( .A(B[0]), .Q(n88) );
  INV3 U52 ( .A(A[12]), .Q(n233) );
  INV3 U53 ( .A(n252), .Q(n114) );
  NOR32 U54 ( .A(n253), .B(n254), .C(n255), .Q(n252) );
  NAND42 U55 ( .A(n54), .B(n55), .C(n56), .D(n57), .Q(n53) );
  NAND42 U56 ( .A(n39), .B(n40), .C(n41), .D(n42), .Q(n38) );
  AOI221 U57 ( .A(B[6]), .B(n76), .C(n96), .D(n97), .Q(n50) );
  NAND33 U58 ( .A(n234), .B(n235), .C(n236), .Q(n212) );
  NAND33 U59 ( .A(n237), .B(n125), .C(n238), .Q(n236) );
  CLKIN1 U60 ( .A(B[9]), .Q(n163) );
  NAND41 U61 ( .A(n115), .B(n116), .C(n117), .D(B[8]), .Q(n160) );
  NAND24 U62 ( .A(A[21]), .B(n9), .Q(n104) );
  NOR20 U63 ( .A(B[1]), .B(n91), .Q(n90) );
  AOI312 U64 ( .A(n19), .B(n20), .C(n21), .D(n22), .Q(LT_LE) );
  NOR21 U65 ( .A(n5), .B(n233), .Q(n254) );
  INV1 U66 ( .A(B[12]), .Q(n6) );
  NAND21 U67 ( .A(n119), .B(n104), .Q(n240) );
  NAND21 U68 ( .A(n60), .B(n61), .Q(n122) );
  INV1 U69 ( .A(B[16]), .Q(n7) );
  NOR21 U70 ( .A(n121), .B(n122), .Q(n120) );
  NAND22 U71 ( .A(A[14]), .B(n135), .Q(n153) );
  INV1 U72 ( .A(B[14]), .Q(n135) );
  NAND22 U73 ( .A(n62), .B(n63), .Q(n58) );
  OAI311 U74 ( .A(n195), .B(n106), .C(n196), .D(n197), .Q(n187) );
  NOR21 U75 ( .A(n141), .B(n247), .Q(n246) );
  CLKIN3 U76 ( .A(B[21]), .Q(n9) );
  NOR21 U77 ( .A(n106), .B(n118), .Q(n111) );
  INV3 U78 ( .A(B[17]), .Q(n228) );
  NAND21 U79 ( .A(A[10]), .B(n3), .Q(n62) );
  NAND21 U80 ( .A(n60), .B(n61), .Q(n167) );
  NAND22 U81 ( .A(n61), .B(n265), .Q(n264) );
  NAND22 U82 ( .A(A[11]), .B(n4), .Q(n61) );
  NAND21 U83 ( .A(n256), .B(n119), .Q(n250) );
  NAND22 U84 ( .A(A[20]), .B(n8), .Q(n210) );
  NAND42 U85 ( .A(n104), .B(n105), .C(n119), .D(n165), .Q(n164) );
  NOR21 U86 ( .A(n106), .B(n164), .Q(n158) );
  NAND31 U87 ( .A(n116), .B(n119), .C(n157), .Q(n155) );
  INV2 U88 ( .A(A[3]), .Q(n95) );
  NOR20 U89 ( .A(n136), .B(n137), .Q(n132) );
  NAND24 U90 ( .A(A[24]), .B(n11), .Q(n180) );
  NOR31 U91 ( .A(n134), .B(n102), .C(n135), .Q(n133) );
  NOR20 U92 ( .A(n136), .B(n232), .Q(n231) );
  NAND22 U93 ( .A(n62), .B(n123), .Q(n121) );
  NOR20 U94 ( .A(n141), .B(n102), .Q(n230) );
  NAND21 U95 ( .A(n252), .B(n200), .Q(n196) );
  NOR20 U96 ( .A(n141), .B(n209), .Q(n208) );
  NAND22 U97 ( .A(n252), .B(n108), .Q(n107) );
  NOR21 U98 ( .A(n109), .B(n110), .Q(n108) );
  AOI2111 U99 ( .A(n186), .B(n180), .C(n187), .D(n188), .Q(n20) );
  INV0 U100 ( .A(A[18]), .Q(n18) );
  NAND20 U101 ( .A(n174), .B(n180), .Q(n179) );
  NOR31 U102 ( .A(n178), .B(n109), .C(n179), .Q(n177) );
  NOR21 U103 ( .A(n106), .B(n261), .Q(n248) );
  NOR31 U104 ( .A(n101), .B(n102), .C(n103), .Q(n44) );
  CLKIN2 U105 ( .A(B[24]), .Q(n11) );
  NAND22 U106 ( .A(A[16]), .B(n7), .Q(n60) );
  NAND30 U107 ( .A(n105), .B(n241), .C(n60), .Q(n239) );
  NAND42 U108 ( .A(n142), .B(n143), .C(n144), .D(n145), .Q(n37) );
  NOR20 U109 ( .A(A[26]), .B(n12), .Q(n194) );
  NAND20 U110 ( .A(n181), .B(n173), .Q(n178) );
  NOR20 U111 ( .A(A[27]), .B(n13), .Q(n193) );
  NOR20 U112 ( .A(A[24]), .B(n199), .Q(n198) );
  NAND26 U113 ( .A(A[23]), .B(n10), .Q(n116) );
  NAND20 U114 ( .A(B[21]), .B(n173), .Q(n172) );
  NAND20 U115 ( .A(n246), .B(n119), .Q(n244) );
  CLKIN2 U116 ( .A(n271), .Q(n269) );
  INV0 U117 ( .A(A[11]), .Q(n241) );
  NOR20 U118 ( .A(A[20]), .B(n141), .Q(n207) );
  INV0 U119 ( .A(A[15]), .Q(n129) );
  INV0 U120 ( .A(A[16]), .Q(n17) );
  NAND20 U121 ( .A(B[18]), .B(n115), .Q(n156) );
  NAND20 U122 ( .A(n62), .B(n168), .Q(n166) );
  NAND20 U123 ( .A(n210), .B(n211), .Q(n209) );
  NAND20 U124 ( .A(A[28]), .B(n14), .Q(n34) );
  NOR20 U125 ( .A(A[28]), .B(n14), .Q(n192) );
  NOR24 U126 ( .A(n267), .B(n268), .Q(n266) );
  INV0 U127 ( .A(B[1]), .Q(n100) );
  NOR20 U128 ( .A(A[1]), .B(n94), .Q(n97) );
  INV0 U129 ( .A(A[0]), .Q(n92) );
  NOR20 U130 ( .A(B[3]), .B(n95), .Q(n81) );
  INV0 U131 ( .A(A[17]), .Q(n227) );
  NAND20 U132 ( .A(n104), .B(n227), .Q(n226) );
  NOR20 U133 ( .A(B[3]), .B(n95), .Q(n93) );
  NOR30 U134 ( .A(n94), .B(A[0]), .C(n93), .Q(n86) );
  NAND20 U135 ( .A(n138), .B(n139), .Q(n137) );
  NAND21 U136 ( .A(n60), .B(n61), .Q(n59) );
  NOR21 U137 ( .A(n58), .B(n59), .Q(n57) );
  CLKIN0 U138 ( .A(A[19]), .Q(n211) );
  INV0 U139 ( .A(B[3]), .Q(n80) );
  CLKIN0 U140 ( .A(B[7]), .Q(n64) );
  NOR21 U141 ( .A(n175), .B(n109), .Q(n224) );
  INV3 U142 ( .A(n6), .Q(n5) );
  NAND22 U143 ( .A(n23), .B(n24), .Q(n22) );
  NOR21 U144 ( .A(n192), .B(n193), .Q(n191) );
  INV3 U145 ( .A(n194), .Q(n190) );
  NAND22 U146 ( .A(n243), .B(n125), .Q(n235) );
  NAND22 U147 ( .A(n248), .B(n249), .Q(n234) );
  NOR21 U148 ( .A(n136), .B(n202), .Q(n201) );
  NAND22 U149 ( .A(n61), .B(n16), .Q(n202) );
  NOR21 U150 ( .A(n176), .B(n177), .Q(n142) );
  NAND22 U151 ( .A(A[26]), .B(n12), .Q(n270) );
  INV3 U152 ( .A(B[26]), .Q(n12) );
  NAND22 U153 ( .A(n111), .B(n112), .Q(n41) );
  NOR21 U154 ( .A(n140), .B(n141), .Q(n131) );
  INV3 U155 ( .A(n75), .Q(n54) );
  NAND22 U156 ( .A(n65), .B(n66), .Q(n56) );
  INV3 U157 ( .A(n71), .Q(n55) );
  NAND31 U158 ( .A(n105), .B(n129), .C(n60), .Q(n127) );
  NOR21 U159 ( .A(n239), .B(n240), .Q(n238) );
  NAND22 U160 ( .A(n230), .B(n231), .Q(n214) );
  NOR21 U161 ( .A(n127), .B(n128), .Q(n126) );
  NAND20 U162 ( .A(n119), .B(n104), .Q(n128) );
  INV3 U163 ( .A(A[23]), .Q(n258) );
  NOR21 U164 ( .A(n242), .B(n114), .Q(n237) );
  NAND41 U165 ( .A(n105), .B(n60), .C(n104), .D(n150), .Q(n149) );
  NOR21 U166 ( .A(n171), .B(n172), .Q(n170) );
  NOR21 U167 ( .A(n244), .B(n245), .Q(n243) );
  NOR31 U168 ( .A(n77), .B(n78), .C(n79), .Q(n52) );
  NAND22 U169 ( .A(n68), .B(n84), .Q(n77) );
  NOR21 U170 ( .A(n81), .B(n82), .Q(n78) );
  NOR21 U171 ( .A(n151), .B(n152), .Q(n150) );
  NAND22 U172 ( .A(n153), .B(n154), .Q(n152) );
  NAND22 U173 ( .A(n105), .B(n233), .Q(n232) );
  NOR21 U174 ( .A(n183), .B(n184), .Q(n176) );
  NAND22 U175 ( .A(B[25]), .B(n173), .Q(n184) );
  NAND22 U176 ( .A(n174), .B(n185), .Q(n183) );
  INV3 U177 ( .A(A[25]), .Q(n185) );
  NOR21 U178 ( .A(n166), .B(n167), .Q(n165) );
  INV3 U179 ( .A(A[8]), .Q(n168) );
  NAND22 U180 ( .A(n158), .B(n159), .Q(n144) );
  NAND22 U181 ( .A(n105), .B(n17), .Q(n247) );
  NOR21 U182 ( .A(B[13]), .B(n154), .Q(n255) );
  NOR21 U183 ( .A(n25), .B(n26), .Q(n24) );
  NOR21 U184 ( .A(n27), .B(n47), .Q(n26) );
  NOR21 U185 ( .A(n47), .B(n28), .Q(n25) );
  XNR21 U186 ( .A(B[31]), .B(A[31]), .Q(n27) );
  NOR21 U187 ( .A(n31), .B(n32), .Q(n23) );
  NOR21 U188 ( .A(n33), .B(n34), .Q(n32) );
  NOR21 U189 ( .A(n33), .B(n35), .Q(n31) );
  INV3 U190 ( .A(B[31]), .Q(n15) );
  INV3 U191 ( .A(n47), .Q(n30) );
  NOR21 U192 ( .A(A[31]), .B(n15), .Q(n47) );
  INV3 U193 ( .A(B[15]), .Q(n130) );
  NAND22 U194 ( .A(n222), .B(n174), .Q(n221) );
  NAND22 U195 ( .A(n224), .B(n225), .Q(n220) );
  NOR21 U196 ( .A(n223), .B(n189), .Q(n222) );
  INV3 U197 ( .A(B[22]), .Q(n223) );
  INV3 U198 ( .A(B[29]), .Q(n36) );
  INV3 U199 ( .A(n110), .Q(n117) );
  INV3 U200 ( .A(B[30]), .Q(n29) );
  NOR21 U201 ( .A(n81), .B(n100), .Q(n96) );
  NOR21 U202 ( .A(B[22]), .B(n259), .Q(n257) );
  INV3 U203 ( .A(A[22]), .Q(n259) );
  NOR21 U204 ( .A(n48), .B(n49), .Q(n46) );
  NAND22 U205 ( .A(A[8]), .B(n2), .Q(n162) );
  NAND22 U206 ( .A(B[4]), .B(n70), .Q(n84) );
  INV3 U207 ( .A(A[14]), .Q(n139) );
  NAND22 U208 ( .A(n86), .B(n87), .Q(n51) );
  NOR31 U209 ( .A(n88), .B(n89), .C(n90), .Q(n87) );
  INV3 U210 ( .A(A[4]), .Q(n70) );
  INV3 U211 ( .A(B[28]), .Q(n14) );
  NAND20 U212 ( .A(A[29]), .B(n36), .Q(n35) );
  CLKIN2 U213 ( .A(B[8]), .Q(n2) );
  NOR21 U214 ( .A(n113), .B(n114), .Q(n112) );
  INV0 U215 ( .A(A[9]), .Q(n265) );
  INV1 U216 ( .A(A[13]), .Q(n154) );
  INV2 U217 ( .A(A[1]), .Q(n91) );
  NAND20 U218 ( .A(A[5]), .B(n73), .Q(n72) );
  INV0 U219 ( .A(A[5]), .Q(n85) );
  INV0 U220 ( .A(A[2]), .Q(n83) );
  NAND20 U221 ( .A(A[2]), .B(n99), .Q(n98) );
  NOR20 U222 ( .A(A[30]), .B(n29), .Q(n49) );
  NAND22 U223 ( .A(n18), .B(n104), .Q(n1) );
  NOR21 U224 ( .A(n160), .B(n114), .Q(n159) );
  NOR21 U225 ( .A(n69), .B(n70), .Q(n65) );
  NOR21 U226 ( .A(n69), .B(n72), .Q(n71) );
  NAND41 U227 ( .A(n116), .B(n115), .C(B[13]), .D(n119), .Q(n148) );
  NOR20 U228 ( .A(B[0]), .B(n92), .Q(n89) );
  NOR20 U229 ( .A(B[6]), .B(n76), .Q(n75) );
  CLKIN0 U230 ( .A(B[6]), .Q(n74) );
  NOR20 U231 ( .A(B[19]), .B(n211), .Q(n271) );
  NOR21 U232 ( .A(A[3]), .B(n80), .Q(n79) );
  NAND21 U233 ( .A(B[5]), .B(n85), .Q(n68) );
  NOR31 U234 ( .A(n226), .B(n102), .C(n103), .Q(n218) );
  AOI311 U235 ( .A(n217), .B(n125), .C(n218), .D(n219), .Q(n216) );
  NAND21 U236 ( .A(n104), .B(n105), .Q(n101) );
  NOR21 U237 ( .A(B[4]), .B(n67), .Q(n66) );
  CLKIN0 U238 ( .A(A[6]), .Q(n76) );
  NOR21 U239 ( .A(A[6]), .B(n74), .Q(n69) );
  CLKIN0 U240 ( .A(A[7]), .Q(n123) );
  NAND20 U241 ( .A(A[7]), .B(n64), .Q(n63) );
  NAND20 U242 ( .A(B[2]), .B(n83), .Q(n82) );
  INV1 U243 ( .A(B[2]), .Q(n99) );
  NAND31 U244 ( .A(n116), .B(n119), .C(n208), .Q(n203) );
  NAND31 U245 ( .A(n116), .B(n119), .C(n207), .Q(n205) );
  NAND40 U246 ( .A(n169), .B(n116), .C(n119), .D(n170), .Q(n143) );
  NAND30 U247 ( .A(B[16]), .B(n116), .C(n115), .Q(n245) );
  NAND30 U248 ( .A(B[11]), .B(n116), .C(n115), .Q(n242) );
  NOR21 U249 ( .A(A[29]), .B(n36), .Q(n48) );
  NOR21 U250 ( .A(A[21]), .B(n175), .Q(n169) );
  NAND20 U251 ( .A(A[30]), .B(n29), .Q(n28) );
  NAND40 U252 ( .A(B[24]), .B(n173), .C(n115), .D(n198), .Q(n197) );
  NAND40 U253 ( .A(B[20]), .B(n173), .C(n174), .D(n115), .Q(n206) );
  NAND40 U254 ( .A(B[19]), .B(n173), .C(n174), .D(n115), .Q(n204) );
  NOR21 U255 ( .A(n109), .B(n228), .Q(n217) );
  NOR31 U256 ( .A(n109), .B(n103), .C(n130), .Q(n124) );
  NOR31 U257 ( .A(n109), .B(n103), .C(n6), .Q(n229) );
  AOI312 U258 ( .A(n50), .B(n51), .C(n52), .D(n53), .Q(n45) );
  CLKIN3 U259 ( .A(n68), .Q(n67) );
  CLKIN3 U260 ( .A(n105), .Q(n140) );
  CLKIN3 U261 ( .A(n138), .Q(n151) );
  CLKIN3 U262 ( .A(n182), .Q(n181) );
  OAI212 U263 ( .A(n189), .B(n190), .C(n191), .Q(n188) );
  CLKIN3 U264 ( .A(n174), .Q(n199) );
  OAI222 U265 ( .A(n203), .B(n204), .C(n205), .D(n206), .Q(n186) );
  OAI312 U266 ( .A(n214), .B(n106), .C(n215), .D(n216), .Q(n213) );
  CLKIN3 U267 ( .A(n173), .Q(n189) );
  CLKIN3 U268 ( .A(n180), .Q(n175) );
  CLKIN3 U269 ( .A(n60), .Q(n136) );
  CLKIN3 U270 ( .A(n62), .Q(n263) );
  NAND33 U271 ( .A(n269), .B(n270), .C(n173), .Q(n268) );
  OAI2112 U272 ( .A(B[18]), .B(n18), .C(n210), .D(n180), .Q(n267) );
endmodule


module E_alu_DW01_add_15 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91;

  NOR22 U2 ( .A(n68), .B(n66), .Q(n25) );
  OAI210 U3 ( .A(B[2]), .B(A[2]), .C(n78), .Q(n83) );
  NAND24 U4 ( .A(n23), .B(n24), .Q(n9) );
  NOR32 U5 ( .A(n67), .B(n68), .C(n69), .Q(n27) );
  INV3 U6 ( .A(n25), .Q(n24) );
  NOR22 U7 ( .A(n26), .B(n27), .Q(n23) );
  NAND22 U8 ( .A(n48), .B(n49), .Q(n33) );
  INV3 U9 ( .A(B[2]), .Q(n3) );
  INV1 U10 ( .A(n19), .Q(n87) );
  NOR22 U11 ( .A(A[1]), .B(B[1]), .Q(n19) );
  NAND28 U12 ( .A(n8), .B(n7), .Q(SUM[8]) );
  INV3 U13 ( .A(n5), .Q(n4) );
  NOR23 U14 ( .A(A[3]), .B(B[3]), .Q(n68) );
  AOI211 U15 ( .A(n37), .B(n33), .C(n38), .Q(n31) );
  INV3 U16 ( .A(A[2]), .Q(n6) );
  NOR21 U17 ( .A(n13), .B(n14), .Q(n12) );
  AOI211 U18 ( .A(n15), .B(n16), .C(n17), .Q(n11) );
  NAND22 U19 ( .A(n60), .B(n61), .Q(n34) );
  XOR21 U20 ( .A(n46), .B(n47), .Q(SUM[6]) );
  INV3 U21 ( .A(n44), .Q(n37) );
  NAND22 U22 ( .A(B[5]), .B(A[5]), .Q(n44) );
  NAND22 U23 ( .A(B[6]), .B(A[6]), .Q(n50) );
  INV3 U24 ( .A(n2), .Q(n69) );
  NOR21 U25 ( .A(n27), .B(n25), .Q(n65) );
  AOI211 U26 ( .A(n59), .B(n53), .C(n56), .Q(n58) );
  INV2 U27 ( .A(B[5]), .Q(n60) );
  NAND21 U28 ( .A(n56), .B(n34), .Q(n43) );
  INV2 U29 ( .A(n75), .Q(n56) );
  CLKIN3 U30 ( .A(B[4]), .Q(n5) );
  NAND22 U31 ( .A(B[0]), .B(A[0]), .Q(n22) );
  NAND23 U32 ( .A(n3), .B(n6), .Q(n2) );
  NAND22 U33 ( .A(A[1]), .B(B[1]), .Q(n67) );
  NOR20 U34 ( .A(n54), .B(n17), .Q(n52) );
  INV2 U35 ( .A(n34), .Q(n17) );
  NOR21 U36 ( .A(n68), .B(n22), .Q(n21) );
  NOR21 U37 ( .A(n68), .B(n73), .Q(n71) );
  CLKIN2 U38 ( .A(B[7]), .Q(n16) );
  INV3 U39 ( .A(n18), .Q(n10) );
  INV1 U40 ( .A(A[7]), .Q(n15) );
  NOR21 U41 ( .A(n4), .B(A[4]), .Q(n13) );
  NAND21 U42 ( .A(n86), .B(n87), .Q(n85) );
  INV3 U43 ( .A(n90), .Q(n86) );
  AOI211 U44 ( .A(n70), .B(n71), .C(n26), .Q(n64) );
  NOR20 U45 ( .A(n36), .B(n5), .Q(n35) );
  CLKIN2 U46 ( .A(n82), .Q(n80) );
  XNR20 U47 ( .A(n81), .B(n83), .Q(SUM[2]) );
  NAND20 U48 ( .A(n34), .B(n44), .Q(n57) );
  CLKIN0 U49 ( .A(n54), .Q(n59) );
  AOI212 U50 ( .A(n28), .B(n29), .C(n30), .Q(n7) );
  NOR20 U51 ( .A(n38), .B(n14), .Q(n47) );
  NAND21 U52 ( .A(n45), .B(n51), .Q(n46) );
  NAND22 U53 ( .A(n31), .B(n32), .Q(n29) );
  IMUX20 U54 ( .A(n91), .B(B[0]), .S(A[0]), .Q(SUM[0]) );
  INV2 U55 ( .A(B[0]), .Q(n91) );
  NOR20 U56 ( .A(n74), .B(n56), .Q(n63) );
  NAND20 U57 ( .A(n4), .B(A[4]), .Q(n75) );
  IMUX20 U58 ( .A(n62), .B(n63), .S(n53), .Q(SUM[4]) );
  NAND22 U59 ( .A(A[2]), .B(B[2]), .Q(n66) );
  XOR21 U60 ( .A(n86), .B(n88), .Q(SUM[1]) );
  NAND22 U61 ( .A(n64), .B(n65), .Q(n53) );
  NAND22 U62 ( .A(n84), .B(n85), .Q(n81) );
  NOR21 U63 ( .A(n15), .B(n16), .Q(n30) );
  NAND22 U64 ( .A(n52), .B(n53), .Q(n45) );
  XOR21 U65 ( .A(n40), .B(n41), .Q(SUM[7]) );
  AOI211 U66 ( .A(n42), .B(n33), .C(n38), .Q(n41) );
  NAND31 U67 ( .A(n43), .B(n44), .C(n45), .Q(n42) );
  XOR21 U68 ( .A(n76), .B(n77), .Q(SUM[3]) );
  NAND22 U69 ( .A(n78), .B(n79), .Q(n76) );
  NAND22 U70 ( .A(n80), .B(n81), .Q(n79) );
  XOR21 U71 ( .A(n57), .B(n58), .Q(SUM[5]) );
  NOR21 U72 ( .A(n37), .B(n55), .Q(n51) );
  NAND31 U73 ( .A(n33), .B(n34), .C(n35), .Q(n32) );
  INV3 U74 ( .A(n33), .Q(n14) );
  INV3 U75 ( .A(n39), .Q(n28) );
  NAND22 U76 ( .A(n20), .B(n21), .Q(n18) );
  AOI210 U77 ( .A(n6), .B(n3), .C(n19), .Q(n20) );
  INV3 U78 ( .A(A[6]), .Q(n49) );
  NAND21 U79 ( .A(B[0]), .B(A[0]), .Q(n73) );
  NAND21 U80 ( .A(B[0]), .B(A[0]), .Q(n90) );
  NAND20 U81 ( .A(B[1]), .B(A[1]), .Q(n84) );
  INV2 U82 ( .A(A[5]), .Q(n61) );
  NAND21 U83 ( .A(B[3]), .B(A[3]), .Q(n72) );
  CLKIN3 U84 ( .A(B[6]), .Q(n48) );
  INV2 U85 ( .A(A[4]), .Q(n36) );
  NOR20 U86 ( .A(B[2]), .B(A[2]), .Q(n82) );
  NAND20 U87 ( .A(B[2]), .B(A[2]), .Q(n78) );
  XNR20 U88 ( .A(B[7]), .B(A[7]), .Q(n40) );
  NOR21 U89 ( .A(A[7]), .B(B[7]), .Q(n39) );
  NOR21 U90 ( .A(n89), .B(n19), .Q(n88) );
  AOI210 U91 ( .A(n6), .B(n3), .C(n19), .Q(n70) );
  XOR20 U92 ( .A(B[3]), .B(A[3]), .Q(n77) );
  NOR21 U93 ( .A(n4), .B(A[4]), .Q(n74) );
  NOR21 U94 ( .A(A[4]), .B(n4), .Q(n54) );
  XNR20 U95 ( .A(n4), .B(A[4]), .Q(n62) );
  OAI2112 U96 ( .A(n9), .B(n10), .C(n11), .D(n12), .Q(n8) );
  CLKIN3 U97 ( .A(n50), .Q(n38) );
  CLKIN3 U98 ( .A(n43), .Q(n55) );
  CLKIN3 U99 ( .A(n72), .Q(n26) );
  CLKIN3 U100 ( .A(n84), .Q(n89) );
endmodule


module E_alu_DW01_add_16 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95;

  NAND21 U2 ( .A(n15), .B(n49), .Q(n50) );
  NAND23 U3 ( .A(n19), .B(n20), .Q(n10) );
  NAND26 U4 ( .A(n7), .B(n8), .Q(SUM[8]) );
  OAI210 U5 ( .A(B[2]), .B(A[2]), .C(n81), .Q(n85) );
  NAND21 U6 ( .A(A[2]), .B(B[2]), .Q(n71) );
  NOR21 U7 ( .A(n27), .B(n28), .Q(n26) );
  CLKIN3 U8 ( .A(B[4]), .Q(n5) );
  NOR21 U9 ( .A(n23), .B(n73), .Q(n22) );
  NAND22 U10 ( .A(n29), .B(n30), .Q(n9) );
  NOR24 U11 ( .A(B[2]), .B(A[2]), .Q(n73) );
  NAND22 U12 ( .A(A[1]), .B(B[1]), .Q(n72) );
  AOI211 U13 ( .A(n6), .B(n3), .C(n24), .Q(n74) );
  NOR23 U14 ( .A(B[0]), .B(A[0]), .Q(n23) );
  CLKIN3 U15 ( .A(n62), .Q(n51) );
  NOR22 U16 ( .A(n27), .B(n71), .Q(n31) );
  NAND22 U17 ( .A(n74), .B(n26), .Q(n19) );
  NAND22 U18 ( .A(n21), .B(n22), .Q(n20) );
  NOR21 U19 ( .A(n24), .B(n25), .Q(n21) );
  NAND22 U20 ( .A(n67), .B(n68), .Q(n62) );
  XOR21 U21 ( .A(n46), .B(n47), .Q(SUM[7]) );
  INV3 U22 ( .A(B[2]), .Q(n3) );
  INV3 U23 ( .A(A[2]), .Q(n6) );
  AOI210 U24 ( .A(n74), .B(n75), .C(n32), .Q(n67) );
  NAND31 U25 ( .A(n15), .B(n39), .C(n40), .Q(n38) );
  AOI211 U26 ( .A(n42), .B(n15), .C(n43), .Q(n37) );
  INV2 U27 ( .A(B[7]), .Q(n17) );
  NOR24 U28 ( .A(A[3]), .B(B[3]), .Q(n27) );
  NOR23 U29 ( .A(A[1]), .B(B[1]), .Q(n24) );
  NAND22 U30 ( .A(B[6]), .B(A[6]), .Q(n49) );
  AOI211 U31 ( .A(n16), .B(n17), .C(n18), .Q(n11) );
  INV1 U32 ( .A(B[5]), .Q(n63) );
  NOR22 U33 ( .A(n13), .B(n14), .Q(n12) );
  NAND22 U34 ( .A(B[5]), .B(A[5]), .Q(n44) );
  NOR21 U35 ( .A(n27), .B(n77), .Q(n75) );
  NOR31 U36 ( .A(n72), .B(n27), .C(n73), .Q(n2) );
  AOI211 U37 ( .A(n61), .B(n62), .C(n54), .Q(n60) );
  NOR21 U38 ( .A(B[3]), .B(A[3]), .Q(n25) );
  OAI2112 U39 ( .A(n51), .B(n52), .C(n53), .D(n44), .Q(n48) );
  NOR32 U40 ( .A(n72), .B(n27), .C(n73), .Q(n33) );
  AOI212 U41 ( .A(n48), .B(n15), .C(n43), .Q(n47) );
  NAND21 U42 ( .A(n54), .B(n39), .Q(n53) );
  INV2 U43 ( .A(n78), .Q(n54) );
  NOR20 U44 ( .A(n56), .B(n18), .Q(n55) );
  INV1 U45 ( .A(A[7]), .Q(n16) );
  XNR21 U46 ( .A(n50), .B(n48), .Q(SUM[6]) );
  INV0 U47 ( .A(n86), .Q(n91) );
  NAND22 U48 ( .A(n63), .B(n64), .Q(n39) );
  INV2 U49 ( .A(n45), .Q(n34) );
  NOR20 U50 ( .A(n41), .B(n5), .Q(n40) );
  NOR21 U51 ( .A(n4), .B(A[4]), .Q(n13) );
  NAND20 U52 ( .A(B[2]), .B(A[2]), .Q(n81) );
  XNR20 U53 ( .A(n84), .B(n85), .Q(SUM[2]) );
  AOI212 U54 ( .A(n34), .B(n35), .C(n36), .Q(n7) );
  XOR20 U55 ( .A(n88), .B(n90), .Q(SUM[1]) );
  CLKIN0 U56 ( .A(n56), .Q(n61) );
  NOR20 U57 ( .A(A[0]), .B(B[0]), .Q(n93) );
  AOI210 U58 ( .A(n41), .B(n5), .C(n54), .Q(n65) );
  IMUX20 U59 ( .A(n65), .B(n66), .S(n51), .Q(SUM[4]) );
  INV3 U60 ( .A(n5), .Q(n4) );
  NOR21 U61 ( .A(n23), .B(n73), .Q(n70) );
  INV3 U62 ( .A(n73), .Q(n83) );
  INV3 U63 ( .A(B[0]), .Q(n95) );
  XOR21 U64 ( .A(n59), .B(n60), .Q(SUM[5]) );
  NAND22 U65 ( .A(n39), .B(n44), .Q(n59) );
  NOR21 U66 ( .A(n91), .B(n24), .Q(n90) );
  INV3 U67 ( .A(n55), .Q(n52) );
  NAND22 U68 ( .A(n86), .B(n87), .Q(n84) );
  NAND22 U69 ( .A(n88), .B(n89), .Q(n87) );
  INV3 U70 ( .A(n24), .Q(n89) );
  NAND22 U71 ( .A(n92), .B(n93), .Q(n88) );
  NOR21 U72 ( .A(n16), .B(n17), .Q(n36) );
  NOR21 U73 ( .A(n24), .B(n25), .Q(n69) );
  AOI2111 U74 ( .A(n69), .B(n70), .C(n2), .D(n31), .Q(n68) );
  XOR21 U75 ( .A(n79), .B(n80), .Q(SUM[3]) );
  NAND22 U76 ( .A(n81), .B(n82), .Q(n79) );
  NAND22 U77 ( .A(n83), .B(n84), .Q(n82) );
  NAND22 U78 ( .A(n37), .B(n38), .Q(n35) );
  INV3 U79 ( .A(n31), .Q(n30) );
  NOR21 U80 ( .A(n32), .B(n33), .Q(n29) );
  NAND22 U81 ( .A(n94), .B(n92), .Q(SUM[0]) );
  NAND22 U82 ( .A(n1), .B(n95), .Q(n94) );
  INV3 U83 ( .A(A[0]), .Q(n1) );
  INV3 U84 ( .A(n39), .Q(n18) );
  NAND22 U85 ( .A(n57), .B(n58), .Q(n15) );
  INV3 U86 ( .A(A[6]), .Q(n58) );
  INV3 U87 ( .A(B[6]), .Q(n57) );
  NAND20 U88 ( .A(n4), .B(A[4]), .Q(n78) );
  NAND21 U89 ( .A(B[0]), .B(A[0]), .Q(n92) );
  NAND21 U90 ( .A(B[0]), .B(A[0]), .Q(n77) );
  NAND22 U91 ( .A(B[0]), .B(A[0]), .Q(n28) );
  NAND20 U92 ( .A(B[1]), .B(A[1]), .Q(n86) );
  INV2 U93 ( .A(A[5]), .Q(n64) );
  NAND21 U94 ( .A(B[3]), .B(A[3]), .Q(n76) );
  INV2 U95 ( .A(A[4]), .Q(n41) );
  XNR20 U96 ( .A(B[7]), .B(A[7]), .Q(n46) );
  NOR21 U97 ( .A(A[7]), .B(B[7]), .Q(n45) );
  XOR20 U98 ( .A(B[3]), .B(A[3]), .Q(n80) );
  XNR20 U99 ( .A(n4), .B(A[4]), .Q(n66) );
  NOR21 U100 ( .A(A[4]), .B(n4), .Q(n56) );
  OAI2112 U101 ( .A(n9), .B(n10), .C(n11), .D(n12), .Q(n8) );
  CLKIN3 U102 ( .A(n15), .Q(n14) );
  CLKIN3 U103 ( .A(n44), .Q(n42) );
  CLKIN3 U104 ( .A(n49), .Q(n43) );
  CLKIN3 U105 ( .A(n76), .Q(n32) );
endmodule


module E_alu_DW_rash_3 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n2, n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n147, n148,
         n149, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357;

  NAND23 U3 ( .A(n267), .B(n268), .Q(n162) );
  NAND22 U4 ( .A(n299), .B(n300), .Q(n144) );
  INV3 U5 ( .A(n314), .Q(n195) );
  NOR21 U6 ( .A(n173), .B(n192), .Q(B[22]) );
  NOR21 U7 ( .A(n173), .B(n225), .Q(B[18]) );
  NAND24 U8 ( .A(n295), .B(n296), .Q(n145) );
  AOI221 U9 ( .A(A[27]), .B(n15), .C(A[28]), .D(n21), .Q(n296) );
  AOI221 U10 ( .A(A[25]), .B(n18), .C(A[26]), .D(n21), .Q(n268) );
  AOI221 U11 ( .A(A[27]), .B(n260), .C(A[28]), .D(n261), .Q(n267) );
  INV3 U12 ( .A(n147), .Q(n84) );
  NAND22 U13 ( .A(n155), .B(n156), .Q(n227) );
  NAND23 U14 ( .A(n331), .B(n332), .Q(n152) );
  NAND22 U15 ( .A(n315), .B(n316), .Q(n149) );
  AOI221 U16 ( .A(A[26]), .B(n14), .C(A[27]), .D(n22), .Q(n316) );
  NAND23 U17 ( .A(n335), .B(n336), .Q(n166) );
  NAND22 U18 ( .A(n343), .B(n344), .Q(n71) );
  NAND22 U19 ( .A(n19), .B(n107), .Q(n156) );
  NAND22 U20 ( .A(n94), .B(n95), .Q(n86) );
  AOI221 U21 ( .A(A[20]), .B(n15), .C(A[21]), .D(n22), .Q(n344) );
  NAND23 U22 ( .A(n337), .B(n338), .Q(n168) );
  AOI222 U23 ( .A(A[30]), .B(n260), .C(A[31]), .D(n261), .Q(n337) );
  NAND31 U24 ( .A(n37), .B(n38), .C(n143), .Q(n36) );
  INV3 U25 ( .A(A[20]), .Q(n24) );
  INV2 U26 ( .A(A[19]), .Q(n23) );
  MUX22 U27 ( .A(n333), .B(n334), .S(n29), .Q(B[0]) );
  CLKIN3 U28 ( .A(n125), .Q(n124) );
  NAND22 U29 ( .A(n83), .B(n38), .Q(n116) );
  NAND22 U30 ( .A(n256), .B(n257), .Q(n52) );
  AOI221 U31 ( .A(A[23]), .B(n260), .C(A[24]), .D(n261), .Q(n256) );
  NAND22 U32 ( .A(n221), .B(n222), .Q(n304) );
  AOI221 U33 ( .A(n260), .B(A[18]), .C(n21), .D(A[17]), .Q(n340) );
  NAND24 U34 ( .A(n139), .B(n168), .Q(n239) );
  AOI221 U35 ( .A(A[24]), .B(n260), .C(A[25]), .D(n261), .Q(n331) );
  AOI222 U36 ( .A(A[29]), .B(n260), .C(A[30]), .D(n261), .Q(n295) );
  NAND22 U37 ( .A(n157), .B(n158), .Q(n226) );
  AOI222 U38 ( .A(A[30]), .B(n15), .C(A[31]), .D(n22), .Q(n314) );
  AOI222 U39 ( .A(A[28]), .B(n260), .C(A[29]), .D(n261), .Q(n315) );
  NAND21 U40 ( .A(n19), .B(n162), .Q(n44) );
  AOI221 U41 ( .A(A[23]), .B(n13), .C(A[24]), .D(n21), .Q(n300) );
  NAND21 U42 ( .A(n143), .B(n166), .Q(n127) );
  AOI220 U43 ( .A(A[17]), .B(n16), .C(A[18]), .D(n21), .Q(n273) );
  AOI221 U44 ( .A(A[22]), .B(n260), .C(A[23]), .D(n261), .Q(n343) );
  AOI221 U45 ( .A(A[22]), .B(n18), .C(A[23]), .D(n22), .Q(n332) );
  NAND22 U46 ( .A(n237), .B(n3), .Q(n334) );
  NAND33 U47 ( .A(n239), .B(n240), .C(n238), .Q(n2) );
  INV2 U48 ( .A(n2), .Q(n3) );
  CLKIN0 U49 ( .A(n178), .Q(n175) );
  NAND22 U50 ( .A(n143), .B(n144), .Q(n136) );
  CLKIN2 U51 ( .A(n167), .Q(n165) );
  CLKIN0 U52 ( .A(n177), .Q(n176) );
  NAND21 U53 ( .A(n219), .B(n220), .Q(n305) );
  NAND21 U54 ( .A(n62), .B(n63), .Q(n61) );
  AOI221 U55 ( .A(n139), .B(n56), .C(n83), .D(n54), .Q(n212) );
  CLKIN2 U56 ( .A(n50), .Q(n45) );
  AOI221 U57 ( .A(n67), .B(n57), .C(n58), .D(n59), .Q(B[8]) );
  CLKIN3 U58 ( .A(n105), .Q(n193) );
  NAND22 U59 ( .A(n104), .B(n103), .Q(n194) );
  CLKIN3 U60 ( .A(n114), .Q(n198) );
  CLKIN2 U61 ( .A(n65), .Q(n182) );
  AOI221 U62 ( .A(A[20]), .B(n260), .C(A[21]), .D(n261), .Q(n329) );
  NOR21 U63 ( .A(n226), .B(n227), .Q(n225) );
  NAND40 U64 ( .A(n135), .B(n136), .C(n137), .D(n138), .Q(n134) );
  NAND40 U65 ( .A(n155), .B(n156), .C(n157), .D(n158), .Q(n154) );
  AOI220 U66 ( .A(n53), .B(n54), .C(n55), .D(n56), .Q(n33) );
  NOR21 U67 ( .A(n29), .B(n85), .Q(n186) );
  NAND41 U68 ( .A(n309), .B(n310), .C(n311), .D(n312), .Q(B[10]) );
  NAND20 U69 ( .A(n284), .B(n168), .Q(n281) );
  CLKIN2 U70 ( .A(n291), .Q(n290) );
  AOI220 U71 ( .A(n260), .B(A[17]), .C(A[18]), .D(n261), .Q(n306) );
  NAND20 U72 ( .A(n126), .B(n127), .Q(n123) );
  INV2 U73 ( .A(n252), .Q(n251) );
  NAND20 U74 ( .A(n20), .B(n166), .Q(n65) );
  NOR30 U75 ( .A(n147), .B(n9), .C(n148), .Q(n244) );
  NAND21 U76 ( .A(n143), .B(n52), .Q(n210) );
  AOI210 U77 ( .A(n139), .B(n38), .C(n233), .Q(n204) );
  AOI220 U78 ( .A(n51), .B(n152), .C(n48), .D(n107), .Q(n309) );
  NAND20 U79 ( .A(n139), .B(n38), .Q(n229) );
  CLKIN0 U80 ( .A(n208), .Q(n207) );
  CLKIN0 U81 ( .A(n209), .Q(n206) );
  NAND20 U82 ( .A(n51), .B(n71), .Q(n62) );
  NAND20 U83 ( .A(n55), .B(n76), .Q(n67) );
  CLKIN3 U84 ( .A(n115), .Q(n197) );
  NAND21 U85 ( .A(n143), .B(n71), .Q(n237) );
  NAND21 U86 ( .A(n143), .B(n152), .Q(n155) );
  CLKIN3 U87 ( .A(n64), .Q(n183) );
  NAND20 U88 ( .A(n81), .B(n82), .Q(n80) );
  NAND20 U89 ( .A(n83), .B(n84), .Q(n81) );
  NAND30 U90 ( .A(n114), .B(n115), .C(n116), .Q(n113) );
  CLKIN3 U91 ( .A(n89), .Q(n88) );
  NAND20 U92 ( .A(n51), .B(n52), .Q(n50) );
  NAND20 U93 ( .A(n48), .B(n52), .Q(n255) );
  INV2 U94 ( .A(n186), .Q(n185) );
  MUX22 U95 ( .A(n153), .B(n154), .S(n29), .Q(B[2]) );
  NAND20 U96 ( .A(n55), .B(n107), .Q(n248) );
  AOI220 U97 ( .A(n48), .B(n152), .C(n53), .D(n106), .Q(n249) );
  AOI220 U98 ( .A(A[14]), .B(n260), .C(A[15]), .D(n261), .Q(n347) );
  AOI220 U99 ( .A(A[12]), .B(n18), .C(A[13]), .D(n22), .Q(n348) );
  AOI220 U100 ( .A(A[18]), .B(n13), .C(A[19]), .D(n22), .Q(n330) );
  AOI220 U101 ( .A(A[13]), .B(n13), .C(A[14]), .D(n21), .Q(n266) );
  AOI2110 U102 ( .A(n144), .B(n48), .C(n243), .D(n244), .Q(n242) );
  NOR20 U103 ( .A(n92), .B(n247), .Q(n246) );
  AOI220 U104 ( .A(n83), .B(n90), .C(n139), .D(n97), .Q(n141) );
  AOI220 U105 ( .A(A[13]), .B(n260), .C(A[14]), .D(n261), .Q(n301) );
  NAND20 U106 ( .A(n55), .B(n72), .Q(n122) );
  AOI220 U107 ( .A(n53), .B(n76), .C(n55), .D(n73), .Q(n282) );
  MUX22 U108 ( .A(n133), .B(n134), .S(n29), .Q(B[3]) );
  NOR20 U109 ( .A(n29), .B(n172), .Q(n170) );
  NOR20 U110 ( .A(n92), .B(n131), .Q(n303) );
  AOI220 U111 ( .A(n51), .B(n162), .C(n53), .D(n56), .Q(n254) );
  INV0 U112 ( .A(n76), .Q(n130) );
  NAND20 U113 ( .A(n53), .B(n72), .Q(n68) );
  NAND21 U114 ( .A(n143), .B(n162), .Q(n114) );
  AOI220 U115 ( .A(n48), .B(n106), .C(n51), .D(n107), .Q(n99) );
  NAND20 U116 ( .A(n143), .B(n38), .Q(n180) );
  MUX22 U117 ( .A(n202), .B(n203), .S(n29), .Q(B[1]) );
  NOR20 U118 ( .A(n30), .B(n151), .Q(B[30]) );
  NAND20 U119 ( .A(n294), .B(n84), .Q(n291) );
  INV2 U120 ( .A(n342), .Q(n339) );
  NAND33 U121 ( .A(n339), .B(n340), .C(n341), .Q(n73) );
  NAND33 U122 ( .A(n273), .B(n274), .C(n275), .Q(n49) );
  NAND20 U123 ( .A(A[1]), .B(n21), .Q(n353) );
  NAND20 U124 ( .A(A[15]), .B(n14), .Q(n307) );
  NAND20 U125 ( .A(A[1]), .B(n14), .Q(n264) );
  CLKIN3 U126 ( .A(n169), .Q(B[27]) );
  NAND20 U127 ( .A(n142), .B(n168), .Q(n167) );
  CLKIN3 U128 ( .A(n356), .Q(n260) );
  NAND20 U129 ( .A(SH[0]), .B(n26), .Q(n357) );
  CLKIN3 U130 ( .A(SH[0]), .Q(n25) );
  INV0 U131 ( .A(SH[2]), .Q(n27) );
  NAND22 U132 ( .A(A[19]), .B(n13), .Q(n222) );
  NAND22 U133 ( .A(n139), .B(n84), .Q(n135) );
  NAND22 U134 ( .A(n127), .B(n126), .Q(n200) );
  INV3 U135 ( .A(n210), .Q(n233) );
  NOR21 U136 ( .A(n9), .B(n151), .Q(n252) );
  NOR21 U137 ( .A(n9), .B(n148), .Q(n284) );
  INV3 U138 ( .A(n10), .Q(n37) );
  NAND22 U139 ( .A(n219), .B(n220), .Q(n218) );
  NAND22 U140 ( .A(n221), .B(n222), .Q(n217) );
  INV3 U141 ( .A(n272), .Q(n261) );
  NOR21 U142 ( .A(n304), .B(n305), .Q(n92) );
  NAND22 U143 ( .A(n142), .B(n71), .Q(n126) );
  INV3 U144 ( .A(n231), .Q(n230) );
  NOR21 U145 ( .A(n232), .B(n233), .Q(n228) );
  NAND22 U146 ( .A(n101), .B(n102), .Q(n100) );
  NAND31 U147 ( .A(n103), .B(n104), .C(n105), .Q(n102) );
  NAND22 U148 ( .A(n142), .B(n195), .Q(n151) );
  NAND22 U149 ( .A(n142), .B(n144), .Q(n82) );
  NAND22 U150 ( .A(n83), .B(n195), .Q(n105) );
  AOI211 U151 ( .A(n116), .B(n196), .C(n179), .Q(B[21]) );
  NAND22 U152 ( .A(n143), .B(n195), .Q(n177) );
  NAND22 U153 ( .A(n83), .B(n166), .Q(n240) );
  NAND22 U154 ( .A(n139), .B(n195), .Q(n157) );
  NAND22 U155 ( .A(n20), .B(n52), .Q(n115) );
  NAND22 U156 ( .A(n19), .B(n152), .Q(n103) );
  AOI221 U157 ( .A(n77), .B(n10), .C(n78), .D(n77), .Q(B[7]) );
  NOR21 U158 ( .A(n79), .B(n80), .Q(n78) );
  NOR31 U159 ( .A(n86), .B(n87), .C(n88), .Q(n77) );
  NAND22 U160 ( .A(A[20]), .B(n21), .Q(n221) );
  NOR21 U161 ( .A(n272), .B(n24), .Q(n276) );
  NOR21 U162 ( .A(n272), .B(n23), .Q(n342) );
  NAND22 U163 ( .A(n239), .B(n240), .Q(n235) );
  NAND22 U164 ( .A(n237), .B(n238), .Q(n236) );
  NOR21 U165 ( .A(n9), .B(n172), .Q(n289) );
  NOR21 U166 ( .A(n193), .B(n194), .Q(n192) );
  NOR21 U167 ( .A(n206), .B(n207), .Q(n205) );
  NOR21 U168 ( .A(n182), .B(n183), .Q(n181) );
  NAND22 U169 ( .A(n111), .B(n112), .Q(B[5]) );
  NAND22 U170 ( .A(n101), .B(n113), .Q(n112) );
  INV3 U171 ( .A(n117), .Q(n111) );
  NAND22 U172 ( .A(n208), .B(n209), .Q(n232) );
  NOR21 U173 ( .A(n60), .B(n61), .Q(n59) );
  NAND22 U174 ( .A(n64), .B(n65), .Q(n60) );
  NOR21 U175 ( .A(n69), .B(n70), .Q(n57) );
  NAND22 U176 ( .A(n63), .B(n10), .Q(n69) );
  NAND22 U177 ( .A(n68), .B(n62), .Q(n70) );
  NOR21 U178 ( .A(n197), .B(n198), .Q(n196) );
  NAND22 U179 ( .A(n55), .B(n90), .Q(n89) );
  INV3 U180 ( .A(n313), .Q(n312) );
  INV3 U181 ( .A(n43), .Q(n35) );
  NOR21 U182 ( .A(n44), .B(n10), .Q(n43) );
  INV3 U183 ( .A(n66), .Q(n58) );
  NAND22 U184 ( .A(n67), .B(n68), .Q(n66) );
  INV3 U185 ( .A(n142), .Q(n148) );
  INV3 U186 ( .A(n201), .Q(n139) );
  INV3 U187 ( .A(n8), .Q(n9) );
  INV3 U188 ( .A(n8), .Q(n10) );
  BUF2 U189 ( .A(n11), .Q(n13) );
  BUF2 U190 ( .A(n11), .Q(n14) );
  BUF2 U191 ( .A(n12), .Q(n16) );
  BUF2 U192 ( .A(n258), .Q(n18) );
  BUF2 U193 ( .A(n258), .Q(n17) );
  BUF2 U194 ( .A(n12), .Q(n15) );
  NOR21 U195 ( .A(n9), .B(n148), .Q(n269) );
  NAND22 U196 ( .A(n118), .B(n119), .Q(n117) );
  NAND31 U197 ( .A(n254), .B(n255), .C(n253), .Q(B[13]) );
  NAND22 U198 ( .A(SH[1]), .B(SH[0]), .Q(n272) );
  AOI221 U199 ( .A(A[21]), .B(n14), .C(A[22]), .D(n22), .Q(n257) );
  NAND41 U200 ( .A(n285), .B(n286), .C(n287), .D(n288), .Q(B[11]) );
  NAND22 U201 ( .A(n55), .B(n97), .Q(n285) );
  INV3 U202 ( .A(n303), .Q(n286) );
  NOR21 U203 ( .A(n289), .B(n290), .Q(n288) );
  NAND22 U204 ( .A(n329), .B(n330), .Q(n107) );
  NAND22 U205 ( .A(n347), .B(n348), .Q(n76) );
  NAND41 U206 ( .A(n33), .B(n34), .C(n35), .D(n36), .Q(B[9]) );
  NOR21 U207 ( .A(n45), .B(n46), .Q(n34) );
  AOI221 U208 ( .A(A[24]), .B(n17), .C(A[25]), .D(n22), .Q(n336) );
  AOI221 U209 ( .A(A[26]), .B(n260), .C(A[27]), .D(n261), .Q(n335) );
  NAND41 U210 ( .A(n248), .B(n249), .C(n250), .D(n251), .Q(B[14]) );
  NAND22 U211 ( .A(n51), .B(n149), .Q(n250) );
  AOI221 U212 ( .A(A[25]), .B(n260), .C(A[26]), .D(n261), .Q(n299) );
  NAND22 U213 ( .A(n83), .B(n162), .Q(n209) );
  NAND22 U214 ( .A(n265), .B(n266), .Q(n56) );
  AOI221 U215 ( .A(n83), .B(n72), .C(n139), .D(n76), .Q(n346) );
  AOI221 U216 ( .A(n83), .B(n110), .C(n139), .D(n106), .Q(n160) );
  NAND22 U217 ( .A(n270), .B(n271), .Q(n38) );
  NAND22 U218 ( .A(A[31]), .B(n260), .Q(n270) );
  AOI221 U219 ( .A(A[29]), .B(n17), .C(A[30]), .D(n21), .Q(n271) );
  NAND22 U220 ( .A(A[31]), .B(n16), .Q(n147) );
  NAND22 U221 ( .A(n301), .B(n302), .Q(n90) );
  NAND22 U222 ( .A(A[21]), .B(n260), .Q(n220) );
  NAND22 U223 ( .A(n20), .B(n49), .Q(n208) );
  NAND31 U224 ( .A(n99), .B(n100), .C(n98), .Q(B[6]) );
  NAND22 U225 ( .A(n184), .B(n185), .Q(B[23]) );
  NAND22 U226 ( .A(n83), .B(n168), .Q(n125) );
  NAND31 U227 ( .A(n120), .B(n121), .C(n122), .Q(B[4]) );
  BUF2 U228 ( .A(n259), .Q(n22) );
  BUF2 U229 ( .A(n259), .Q(n21) );
  NAND22 U230 ( .A(n20), .B(n73), .Q(n238) );
  NAND31 U231 ( .A(n282), .B(n283), .C(n281), .Q(B[12]) );
  NAND22 U232 ( .A(n48), .B(n73), .Q(n63) );
  NAND22 U233 ( .A(n83), .B(n149), .Q(n158) );
  NAND22 U234 ( .A(n143), .B(n168), .Q(n64) );
  AOI211 U235 ( .A(n180), .B(n44), .C(n179), .Q(B[25]) );
  NAND22 U236 ( .A(n345), .B(n346), .Q(n333) );
  NAND22 U237 ( .A(n142), .B(n149), .Q(n178) );
  NAND22 U238 ( .A(A[22]), .B(n261), .Q(n219) );
  NAND22 U239 ( .A(n143), .B(n149), .Q(n104) );
  NOR21 U240 ( .A(n170), .B(n171), .Q(n169) );
  NAND22 U241 ( .A(n48), .B(n97), .Q(n94) );
  NAND22 U242 ( .A(n53), .B(n96), .Q(n95) );
  NOR21 U243 ( .A(n29), .B(n136), .Q(n215) );
  NOR21 U244 ( .A(n92), .B(n93), .Q(n87) );
  NOR21 U245 ( .A(n29), .B(n137), .Q(n216) );
  NAND22 U246 ( .A(n55), .B(n106), .Q(n311) );
  NAND22 U247 ( .A(n53), .B(n110), .Q(n310) );
  NOR21 U248 ( .A(n181), .B(n30), .Q(B[24]) );
  NAND22 U249 ( .A(n241), .B(n242), .Q(B[15]) );
  AOI211 U250 ( .A(n53), .B(n97), .C(n246), .Q(n241) );
  NOR21 U251 ( .A(n245), .B(n93), .Q(n243) );
  NOR21 U252 ( .A(n29), .B(n138), .Q(n224) );
  NOR21 U253 ( .A(n187), .B(n188), .Q(n184) );
  INV3 U254 ( .A(n189), .Q(n187) );
  NOR21 U255 ( .A(n29), .B(n82), .Q(n188) );
  NAND22 U256 ( .A(n190), .B(n84), .Q(n189) );
  NAND22 U257 ( .A(n213), .B(n214), .Q(B[19]) );
  AOI211 U258 ( .A(n223), .B(n84), .C(n224), .Q(n213) );
  NOR21 U259 ( .A(n215), .B(n216), .Q(n214) );
  NOR21 U260 ( .A(n29), .B(n201), .Q(n223) );
  NOR21 U261 ( .A(n130), .B(n131), .Q(n129) );
  NOR21 U262 ( .A(n132), .B(n93), .Q(n128) );
  NOR21 U263 ( .A(n234), .B(n173), .Q(B[16]) );
  NOR21 U264 ( .A(n235), .B(n236), .Q(n234) );
  NOR21 U265 ( .A(n179), .B(n199), .Q(B[20]) );
  NOR21 U266 ( .A(n124), .B(n200), .Q(n199) );
  INV3 U267 ( .A(n47), .Q(n46) );
  NAND22 U268 ( .A(n48), .B(n49), .Q(n47) );
  NOR21 U269 ( .A(n9), .B(n42), .Q(n294) );
  NAND22 U270 ( .A(n140), .B(n141), .Q(n133) );
  NAND22 U271 ( .A(n211), .B(n212), .Q(n202) );
  NAND22 U272 ( .A(n204), .B(n205), .Q(n203) );
  NOR31 U273 ( .A(n163), .B(n30), .C(n148), .Q(B[29]) );
  NAND22 U274 ( .A(n159), .B(n160), .Q(n153) );
  NOR21 U275 ( .A(SH[3]), .B(SH[2]), .Q(n142) );
  NAND22 U276 ( .A(SH[3]), .B(SH[2]), .Q(n201) );
  NOR21 U277 ( .A(SH[3]), .B(SH[2]), .Q(n19) );
  NOR21 U278 ( .A(SH[3]), .B(SH[2]), .Q(n20) );
  INV3 U279 ( .A(n191), .Q(n83) );
  INV3 U280 ( .A(n42), .Q(n143) );
  INV3 U281 ( .A(n247), .Q(n55) );
  NOR21 U282 ( .A(SH[1]), .B(SH[0]), .Q(n12) );
  NOR21 U283 ( .A(SH[1]), .B(SH[0]), .Q(n258) );
  NOR21 U284 ( .A(SH[1]), .B(SH[0]), .Q(n11) );
  INV3 U285 ( .A(n131), .Q(n48) );
  INV3 U286 ( .A(n93), .Q(n51) );
  NOR21 U287 ( .A(n29), .B(n191), .Q(n190) );
  INV3 U288 ( .A(n41), .Q(n8) );
  INV3 U289 ( .A(n30), .Q(n41) );
  INV3 U290 ( .A(n30), .Q(n231) );
  INV3 U291 ( .A(n322), .Q(n321) );
  NOR21 U292 ( .A(n272), .B(n323), .Q(n322) );
  NAND31 U293 ( .A(n306), .B(n307), .C(n308), .Q(n97) );
  AOI221 U294 ( .A(A[28]), .B(n16), .C(A[29]), .D(n22), .Q(n338) );
  NAND31 U295 ( .A(n262), .B(n263), .C(n264), .Q(n40) );
  NAND31 U296 ( .A(n319), .B(n320), .C(n321), .Q(n108) );
  NAND22 U297 ( .A(A[4]), .B(n260), .Q(n320) );
  NAND22 U298 ( .A(A[19]), .B(n260), .Q(n274) );
  INV3 U299 ( .A(n276), .Q(n275) );
  NAND22 U300 ( .A(n324), .B(n325), .Q(n106) );
  AOI220 U301 ( .A(A[14]), .B(n17), .C(A[15]), .D(n22), .Q(n325) );
  NAND22 U302 ( .A(n326), .B(n327), .Q(n110) );
  AOI220 U303 ( .A(A[12]), .B(n260), .C(A[13]), .D(n261), .Q(n326) );
  NAND22 U304 ( .A(n349), .B(n350), .Q(n72) );
  NAND22 U305 ( .A(n277), .B(n278), .Q(n54) );
  INV3 U306 ( .A(n164), .Q(B[28]) );
  NAND31 U307 ( .A(n353), .B(n354), .C(n355), .Q(n75) );
  NAND22 U308 ( .A(n297), .B(n298), .Q(n96) );
  NAND22 U309 ( .A(n165), .B(n32), .Q(n164) );
  NOR21 U310 ( .A(n173), .B(n174), .Q(B[26]) );
  INV3 U311 ( .A(n31), .Q(n173) );
  NOR21 U312 ( .A(n175), .B(n176), .Q(n174) );
  NAND22 U313 ( .A(SH[2]), .B(n28), .Q(n42) );
  NAND22 U314 ( .A(n139), .B(n32), .Q(n93) );
  NAND22 U315 ( .A(n83), .B(n32), .Q(n131) );
  NAND22 U316 ( .A(SH[1]), .B(n25), .Q(n356) );
  INV3 U317 ( .A(n31), .Q(n29) );
  NAND22 U318 ( .A(n143), .B(n32), .Q(n247) );
  NAND22 U319 ( .A(SH[3]), .B(n27), .Q(n191) );
  INV3 U320 ( .A(n31), .Q(n30) );
  INV3 U321 ( .A(n328), .Q(n53) );
  NAND22 U322 ( .A(n19), .B(n32), .Q(n328) );
  INV3 U323 ( .A(n31), .Q(n179) );
  INV3 U324 ( .A(SH[1]), .Q(n26) );
  INV3 U325 ( .A(SH[4]), .Q(n31) );
  INV3 U326 ( .A(SH[4]), .Q(n32) );
  INV3 U327 ( .A(SH[3]), .Q(n28) );
  OAI222 U328 ( .A(n228), .B(n230), .C(n229), .D(n230), .Q(B[17]) );
  NAND22 U329 ( .A(n143), .B(n145), .Q(n85) );
  NAND22 U330 ( .A(n83), .B(n145), .Q(n138) );
  INV3 U331 ( .A(n145), .Q(n245) );
  NAND22 U332 ( .A(n20), .B(n145), .Q(n172) );
  AOI220 U333 ( .A(A[8]), .B(n17), .C(A[9]), .D(n22), .Q(n350) );
  AOI220 U334 ( .A(A[16]), .B(n260), .C(A[17]), .D(n261), .Q(n324) );
  AOI220 U335 ( .A(A[15]), .B(n260), .C(A[16]), .D(n261), .Q(n265) );
  NAND20 U336 ( .A(A[16]), .B(n21), .Q(n308) );
  NAND22 U337 ( .A(A[16]), .B(n13), .Q(n341) );
  AOI220 U338 ( .A(n48), .B(n71), .C(n51), .D(n166), .Q(n283) );
  NOR30 U339 ( .A(n147), .B(n30), .C(n42), .Q(n171) );
  NOR31 U340 ( .A(n147), .B(n30), .C(n148), .Q(B[31]) );
  AOI221 U341 ( .A(n53), .B(n109), .C(n55), .D(n110), .Q(n98) );
  AOI220 U342 ( .A(n53), .B(n90), .C(n51), .D(n144), .Q(n287) );
  AOI220 U343 ( .A(n51), .B(n49), .C(n48), .D(n56), .Q(n118) );
  AOI220 U344 ( .A(n55), .B(n49), .C(n269), .D(n38), .Q(n253) );
  NAND22 U345 ( .A(n292), .B(n293), .Q(n91) );
  NAND22 U346 ( .A(n279), .B(n280), .Q(n39) );
  NAND22 U347 ( .A(n317), .B(n318), .Q(n109) );
  NAND22 U348 ( .A(n351), .B(n352), .Q(n74) );
  AOI220 U349 ( .A(n20), .B(n91), .C(n143), .D(n96), .Q(n140) );
  AOI221 U350 ( .A(n53), .B(n39), .C(n55), .D(n54), .Q(n119) );
  AOI221 U351 ( .A(n143), .B(n39), .C(n19), .D(n40), .Q(n211) );
  AOI221 U352 ( .A(n19), .B(n108), .C(n143), .D(n109), .Q(n159) );
  AOI2111 U353 ( .A(n53), .B(n74), .C(n128), .D(n129), .Q(n120) );
  AOI221 U354 ( .A(n20), .B(n75), .C(n143), .D(n74), .Q(n345) );
  NAND20 U355 ( .A(n15), .B(A[0]), .Q(n355) );
  AOI220 U356 ( .A(A[11]), .B(n260), .C(A[12]), .D(n261), .Q(n277) );
  AOI220 U357 ( .A(A[11]), .B(n16), .C(A[12]), .D(n21), .Q(n302) );
  CLKIN0 U358 ( .A(A[5]), .Q(n323) );
  AOI220 U359 ( .A(A[3]), .B(n260), .C(A[4]), .D(n261), .Q(n263) );
  AOI220 U360 ( .A(A[3]), .B(n17), .C(A[4]), .D(n22), .Q(n293) );
  AOI220 U361 ( .A(A[4]), .B(n16), .C(A[5]), .D(n21), .Q(n352) );
  NAND20 U362 ( .A(A[2]), .B(n21), .Q(n262) );
  AOI220 U363 ( .A(A[7]), .B(n260), .C(A[8]), .D(n261), .Q(n279) );
  AOI220 U364 ( .A(A[8]), .B(n260), .C(A[9]), .D(n261), .Q(n317) );
  AOI220 U365 ( .A(A[7]), .B(n14), .C(A[8]), .D(n21), .Q(n298) );
  AOI220 U366 ( .A(A[10]), .B(n260), .C(A[11]), .D(n261), .Q(n349) );
  AOI220 U367 ( .A(A[10]), .B(n14), .C(A[11]), .D(n22), .Q(n327) );
  AOI220 U368 ( .A(A[9]), .B(n15), .C(A[10]), .D(n21), .Q(n278) );
  AOI220 U369 ( .A(A[9]), .B(n260), .C(A[10]), .D(n261), .Q(n297) );
  AOI220 U370 ( .A(A[5]), .B(n260), .C(A[6]), .D(n261), .Q(n292) );
  AOI220 U371 ( .A(A[5]), .B(n18), .C(A[6]), .D(n21), .Q(n280) );
  AOI220 U372 ( .A(A[6]), .B(n13), .C(A[7]), .D(n22), .Q(n318) );
  AOI220 U373 ( .A(A[6]), .B(n260), .C(A[7]), .D(n261), .Q(n351) );
  AOI220 U374 ( .A(A[2]), .B(n18), .C(A[3]), .D(n22), .Q(n319) );
  AOI220 U375 ( .A(A[2]), .B(n260), .C(A[3]), .D(n261), .Q(n354) );
  CLKIN3 U376 ( .A(n85), .Q(n79) );
  OAI212 U377 ( .A(n123), .B(n124), .C(n101), .Q(n121) );
  CLKIN3 U378 ( .A(n10), .Q(n101) );
  CLKIN3 U379 ( .A(n38), .Q(n163) );
  CLKIN3 U380 ( .A(n73), .Q(n132) );
  OAI212 U381 ( .A(n217), .B(n218), .C(n19), .Q(n137) );
  OAI222 U382 ( .A(n10), .B(n178), .C(n10), .D(n177), .Q(n313) );
  CLKIN3 U383 ( .A(n357), .Q(n259) );
endmodule


module E_alu_DW01_sub_10 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182;

  NOR22 U3 ( .A(A[9]), .B(n139), .Q(n138) );
  XOR22 U4 ( .A(n28), .B(n29), .Q(DIFF[9]) );
  CLKIN2 U5 ( .A(A[0]), .Q(n23) );
  AOI222 U6 ( .A(n127), .B(n134), .C(n118), .D(n128), .Q(n126) );
  AOI312 U7 ( .A(n48), .B(n50), .C(n49), .D(n8), .Q(n47) );
  NOR22 U8 ( .A(n110), .B(n121), .Q(n120) );
  NOR23 U9 ( .A(n109), .B(n110), .Q(n101) );
  NAND34 U10 ( .A(n134), .B(n135), .C(n136), .Q(n110) );
  NOR22 U11 ( .A(A[4]), .B(n17), .Q(n173) );
  XNR21 U12 ( .A(n147), .B(n12), .Q(DIFF[11]) );
  INV3 U13 ( .A(A[2]), .Q(n24) );
  AOI312 U14 ( .A(n135), .B(n141), .C(n142), .D(n143), .Q(n103) );
  NAND23 U15 ( .A(n97), .B(n98), .Q(n84) );
  NOR33 U16 ( .A(n7), .B(n8), .C(n181), .Q(n6) );
  AOI312 U17 ( .A(n79), .B(n163), .C(n168), .D(n169), .Q(n112) );
  INV3 U18 ( .A(A[10]), .Q(n27) );
  INV3 U19 ( .A(B[7]), .Q(n19) );
  INV3 U20 ( .A(B[9]), .Q(n139) );
  INV3 U21 ( .A(B[5]), .Q(n18) );
  NAND22 U22 ( .A(A[6]), .B(n182), .Q(n51) );
  INV6 U23 ( .A(B[6]), .Q(n182) );
  NAND22 U24 ( .A(A[2]), .B(n15), .Q(n75) );
  NOR22 U25 ( .A(n131), .B(n6), .Q(n130) );
  INV3 U26 ( .A(n162), .Q(n5) );
  NAND22 U27 ( .A(B[7]), .B(n179), .Q(n124) );
  NOR21 U28 ( .A(B[4]), .B(n25), .Q(n181) );
  NAND22 U29 ( .A(n71), .B(n163), .Q(n115) );
  NOR21 U30 ( .A(B[3]), .B(n167), .Q(n169) );
  NOR21 U31 ( .A(n173), .B(n174), .Q(n172) );
  NAND22 U32 ( .A(n70), .B(n75), .Q(n72) );
  NOR21 U33 ( .A(n42), .B(n36), .Q(n41) );
  INV3 U34 ( .A(A[4]), .Q(n25) );
  INV3 U35 ( .A(B[8]), .Q(n20) );
  INV3 U36 ( .A(n52), .Q(n7) );
  INV3 U37 ( .A(A[8]), .Q(n26) );
  IMUX20 U38 ( .A(n13), .B(n14), .S(A[0]), .Q(DIFF[0]) );
  INV3 U39 ( .A(n51), .Q(n8) );
  NAND22 U40 ( .A(n45), .B(n4), .Q(n154) );
  INV2 U41 ( .A(n4), .Q(n65) );
  NAND22 U42 ( .A(n58), .B(n4), .Q(n53) );
  NAND33 U43 ( .A(n163), .B(n70), .C(n164), .Q(n116) );
  INV3 U44 ( .A(n74), .Q(n164) );
  NOR22 U45 ( .A(A[3]), .B(n16), .Q(n166) );
  CLKIN6 U46 ( .A(B[3]), .Q(n16) );
  INV1 U47 ( .A(B[10]), .Q(n21) );
  INV3 U48 ( .A(n48), .Q(n131) );
  NOR22 U49 ( .A(n30), .B(n31), .Q(n29) );
  AOI212 U50 ( .A(n32), .B(n33), .C(n34), .Q(n31) );
  XNR22 U51 ( .A(n11), .B(n126), .Q(DIFF[12]) );
  INV2 U52 ( .A(B[1]), .Q(n165) );
  NAND21 U53 ( .A(n54), .B(n53), .Q(n57) );
  AOI212 U54 ( .A(n57), .B(n49), .C(n7), .Q(n56) );
  NAND22 U55 ( .A(B[2]), .B(n24), .Q(n70) );
  NAND22 U56 ( .A(B[10]), .B(n27), .Q(n135) );
  XOR22 U57 ( .A(n157), .B(n158), .Q(DIFF[10]) );
  INV2 U58 ( .A(B[0]), .Q(n14) );
  NOR32 U59 ( .A(n23), .B(n13), .C(n170), .Q(n168) );
  INV3 U60 ( .A(n100), .Q(n108) );
  XOR22 U61 ( .A(n81), .B(n80), .Q(DIFF[15]) );
  NAND23 U62 ( .A(B[12]), .B(n105), .Q(n100) );
  NAND24 U63 ( .A(n112), .B(n5), .Q(n4) );
  INV3 U64 ( .A(B[4]), .Q(n17) );
  NAND22 U65 ( .A(n111), .B(n112), .Q(n99) );
  NOR23 U66 ( .A(n137), .B(n138), .Q(n136) );
  NOR22 U67 ( .A(A[8]), .B(n20), .Q(n137) );
  NAND21 U68 ( .A(B[1]), .B(n171), .Q(n79) );
  NAND21 U69 ( .A(A[1]), .B(n165), .Q(n2) );
  NAND22 U70 ( .A(A[1]), .B(n165), .Q(n74) );
  NOR21 U71 ( .A(A[2]), .B(n15), .Q(n170) );
  NAND22 U72 ( .A(A[5]), .B(n18), .Q(n52) );
  NAND20 U73 ( .A(A[5]), .B(n18), .Q(n3) );
  NOR22 U74 ( .A(n152), .B(n159), .Q(n158) );
  INV2 U75 ( .A(n146), .Q(n141) );
  INV0 U76 ( .A(A[3]), .Q(n167) );
  CLKIN0 U77 ( .A(n103), .Q(n127) );
  NOR21 U78 ( .A(A[11]), .B(n22), .Q(n107) );
  NOR20 U79 ( .A(A[11]), .B(n22), .Q(n140) );
  AOI210 U80 ( .A(n58), .B(n4), .C(n61), .Q(n60) );
  INV0 U81 ( .A(A[1]), .Q(n171) );
  INV0 U82 ( .A(B[13]), .Q(n95) );
  NAND21 U83 ( .A(B[8]), .B(n26), .Q(n35) );
  XOR20 U84 ( .A(B[8]), .B(A[8]), .Q(n40) );
  AOI210 U85 ( .A(B[8]), .B(n26), .C(n30), .Q(n39) );
  INV2 U86 ( .A(n140), .Q(n134) );
  NAND20 U87 ( .A(n49), .B(n3), .Q(n59) );
  NAND21 U88 ( .A(A[4]), .B(n17), .Q(n54) );
  NAND20 U89 ( .A(n151), .B(n144), .Q(n150) );
  NAND20 U90 ( .A(A[11]), .B(n22), .Q(n145) );
  NAND20 U91 ( .A(n135), .B(n144), .Q(n157) );
  NAND20 U92 ( .A(A[8]), .B(n20), .Q(n46) );
  NAND20 U93 ( .A(n37), .B(n38), .Q(n28) );
  NAND21 U94 ( .A(n153), .B(n154), .Q(n149) );
  INV0 U95 ( .A(n135), .Q(n155) );
  CLKIN3 U96 ( .A(n62), .Q(n58) );
  NAND30 U97 ( .A(n133), .B(n124), .C(n48), .Q(n177) );
  NAND20 U98 ( .A(n79), .B(n2), .Q(n76) );
  XOR22 U99 ( .A(n55), .B(n56), .Q(DIFF[6]) );
  NAND20 U100 ( .A(n48), .B(n51), .Q(n55) );
  IMUX20 U101 ( .A(n63), .B(n64), .S(n65), .Q(DIFF[4]) );
  XOR20 U102 ( .A(B[4]), .B(A[4]), .Q(n64) );
  NOR20 U103 ( .A(n66), .B(n61), .Q(n63) );
  NOR20 U104 ( .A(A[4]), .B(n17), .Q(n66) );
  XNR20 U105 ( .A(B[7]), .B(A[7]), .Q(n9) );
  NAND20 U106 ( .A(n124), .B(n48), .Q(n123) );
  NAND21 U107 ( .A(n82), .B(n84), .Q(n91) );
  XOR20 U108 ( .A(n96), .B(n84), .Q(DIFF[13]) );
  AOI210 U109 ( .A(n69), .B(n70), .C(n71), .Q(n68) );
  NOR21 U110 ( .A(n107), .B(n108), .Q(n106) );
  CLKIN3 U111 ( .A(n106), .Q(n104) );
  XNR20 U112 ( .A(B[12]), .B(A[12]), .Q(n11) );
  NAND22 U113 ( .A(B[6]), .B(n178), .Q(n48) );
  INV3 U114 ( .A(n78), .Q(n77) );
  NOR21 U115 ( .A(n13), .B(n23), .Q(n78) );
  NAND22 U116 ( .A(n45), .B(n4), .Q(n33) );
  IMUX21 U117 ( .A(n39), .B(n40), .S(n41), .Q(DIFF[8]) );
  NAND22 U118 ( .A(n152), .B(n135), .Q(n151) );
  NAND22 U119 ( .A(n144), .B(n145), .Q(n143) );
  OAI2111 U120 ( .A(n65), .B(n109), .C(n44), .D(n43), .Q(n128) );
  NAND22 U121 ( .A(A[10]), .B(n21), .Q(n144) );
  NAND31 U122 ( .A(n3), .B(n53), .C(n54), .Q(n50) );
  XNR21 U123 ( .A(n72), .B(n69), .Q(DIFF[2]) );
  NAND22 U124 ( .A(n43), .B(n44), .Q(n36) );
  NAND22 U125 ( .A(n129), .B(n130), .Q(n44) );
  NOR21 U126 ( .A(n132), .B(n125), .Q(n129) );
  XOR21 U127 ( .A(n59), .B(n60), .Q(DIFF[5]) );
  NAND22 U128 ( .A(n115), .B(n116), .Q(n162) );
  NOR21 U129 ( .A(n155), .B(n156), .Q(n148) );
  NOR21 U130 ( .A(n113), .B(n114), .Q(n111) );
  AOI211 U131 ( .A(n153), .B(n154), .C(n160), .Q(n159) );
  NOR21 U132 ( .A(n108), .B(n125), .Q(n117) );
  NAND22 U133 ( .A(n37), .B(n35), .Q(n160) );
  INV3 U134 ( .A(B[11]), .Q(n22) );
  INV3 U135 ( .A(n14), .Q(n13) );
  NOR21 U136 ( .A(A[4]), .B(n17), .Q(n62) );
  NAND33 U137 ( .A(n172), .B(n49), .C(n48), .Q(n109) );
  NAND22 U138 ( .A(A[7]), .B(n19), .Q(n43) );
  NAND22 U139 ( .A(A[9]), .B(n139), .Q(n38) );
  NAND21 U140 ( .A(B[5]), .B(n175), .Q(n49) );
  INV3 U141 ( .A(A[5]), .Q(n175) );
  NAND22 U142 ( .A(B[9]), .B(n161), .Q(n37) );
  INV3 U143 ( .A(A[9]), .Q(n161) );
  INV3 U144 ( .A(A[7]), .Q(n179) );
  XNR21 U145 ( .A(n9), .B(n47), .Q(DIFF[7]) );
  NAND22 U146 ( .A(n122), .B(n100), .Q(n121) );
  XOR21 U147 ( .A(n76), .B(n77), .Q(DIFF[1]) );
  NAND22 U148 ( .A(n180), .B(n51), .Q(n133) );
  NAND22 U149 ( .A(n91), .B(n87), .Q(n90) );
  INV3 U150 ( .A(n176), .Q(n153) );
  INV3 U151 ( .A(A[12]), .Q(n105) );
  INV3 U152 ( .A(B[2]), .Q(n15) );
  INV3 U153 ( .A(B[14]), .Q(n89) );
  INV3 U154 ( .A(n86), .Q(n83) );
  XNR21 U155 ( .A(n90), .B(n10), .Q(DIFF[14]) );
  XOR20 U156 ( .A(B[14]), .B(A[14]), .Q(n10) );
  INV3 U157 ( .A(n94), .Q(n82) );
  XNR21 U158 ( .A(n67), .B(n68), .Q(DIFF[3]) );
  INV3 U159 ( .A(n92), .Q(n87) );
  NOR21 U160 ( .A(B[13]), .B(n93), .Q(n92) );
  INV1 U161 ( .A(A[13]), .Q(n93) );
  NOR21 U162 ( .A(n6), .B(n123), .Q(n119) );
  OAI2111 U163 ( .A(n6), .B(n177), .C(n43), .D(n46), .Q(n176) );
  NOR20 U164 ( .A(A[14]), .B(n89), .Q(n86) );
  XOR20 U165 ( .A(B[15]), .B(A[15]), .Q(n81) );
  XNR20 U166 ( .A(B[11]), .B(A[11]), .Q(n12) );
  INV3 U167 ( .A(n166), .Q(n163) );
  INV3 U168 ( .A(n110), .Q(n118) );
  NOR21 U169 ( .A(A[13]), .B(n95), .Q(n94) );
  XNR20 U170 ( .A(B[13]), .B(A[13]), .Q(n96) );
  INV2 U171 ( .A(A[6]), .Q(n178) );
  NOR21 U172 ( .A(A[5]), .B(n18), .Q(n180) );
  NOR21 U173 ( .A(A[7]), .B(n19), .Q(n174) );
  CLKIN0 U174 ( .A(A[14]), .Q(n88) );
  XNR20 U175 ( .A(B[3]), .B(A[3]), .Q(n67) );
  NOR21 U176 ( .A(A[9]), .B(n139), .Q(n146) );
  CLKIN3 U177 ( .A(n35), .Q(n34) );
  CLKIN3 U178 ( .A(n36), .Q(n32) );
  CLKIN3 U179 ( .A(n33), .Q(n42) );
  CLKIN3 U180 ( .A(n46), .Q(n30) );
  CLKIN3 U181 ( .A(n54), .Q(n61) );
  OAI212 U182 ( .A(n73), .B(n77), .C(n2), .Q(n69) );
  AOI312 U183 ( .A(n82), .B(n83), .C(n84), .D(n85), .Q(n80) );
  OAI222 U184 ( .A(n86), .B(n87), .C(B[14]), .D(n88), .Q(n85) );
  AOI312 U185 ( .A(n99), .B(n100), .C(n101), .D(n102), .Q(n98) );
  OAI222 U186 ( .A(n103), .B(n104), .C(B[12]), .D(n105), .Q(n102) );
  CLKIN3 U187 ( .A(n115), .Q(n114) );
  CLKIN3 U188 ( .A(n116), .Q(n113) );
  AOI312 U189 ( .A(n117), .B(n118), .C(n119), .D(n120), .Q(n97) );
  CLKIN3 U190 ( .A(n43), .Q(n122) );
  CLKIN3 U191 ( .A(n133), .Q(n125) );
  CLKIN3 U192 ( .A(n124), .Q(n132) );
  OAI212 U193 ( .A(B[8]), .B(n26), .C(n38), .Q(n142) );
  AOI312 U194 ( .A(n148), .B(n35), .C(n149), .D(n150), .Q(n147) );
  CLKIN3 U195 ( .A(n37), .Q(n156) );
  CLKIN3 U196 ( .A(n75), .Q(n71) );
  CLKIN3 U197 ( .A(n79), .Q(n73) );
  CLKIN3 U198 ( .A(n109), .Q(n45) );
  CLKIN3 U199 ( .A(n38), .Q(n152) );
endmodule


module E_alu_DW01_sub_11 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191;

  CLKIN2 U3 ( .A(n139), .Q(n134) );
  CLKIN3 U4 ( .A(A[0]), .Q(n12) );
  INV3 U5 ( .A(n107), .Q(n163) );
  NOR22 U6 ( .A(n112), .B(n113), .Q(n105) );
  NOR24 U7 ( .A(n178), .B(n179), .Q(n177) );
  NAND21 U8 ( .A(n121), .B(n95), .Q(n120) );
  INV3 U9 ( .A(n95), .Q(n102) );
  NAND31 U10 ( .A(n105), .B(n107), .C(n106), .Q(n94) );
  NAND22 U11 ( .A(n50), .B(n35), .Q(n44) );
  NOR21 U12 ( .A(B[3]), .B(n169), .Q(n173) );
  NAND22 U13 ( .A(B[12]), .B(n100), .Q(n95) );
  NAND33 U14 ( .A(n38), .B(n39), .C(n177), .Q(n103) );
  NAND22 U15 ( .A(n34), .B(n35), .Q(n22) );
  INV3 U16 ( .A(n22), .Q(n31) );
  INV3 U17 ( .A(n42), .Q(n41) );
  XOR21 U18 ( .A(n147), .B(n146), .Q(DIFF[11]) );
  XOR21 U19 ( .A(n84), .B(n85), .Q(DIFF[14]) );
  INV3 U20 ( .A(B[8]), .Q(n9) );
  NOR22 U21 ( .A(B[4]), .B(n14), .Q(n188) );
  INV6 U22 ( .A(n175), .Q(n171) );
  NOR22 U23 ( .A(n104), .B(n120), .Q(n119) );
  NOR23 U24 ( .A(n103), .B(n104), .Q(n96) );
  NAND34 U25 ( .A(n134), .B(n135), .C(n136), .Q(n104) );
  NAND32 U26 ( .A(n43), .B(n44), .C(n45), .Q(n40) );
  NAND33 U27 ( .A(n171), .B(n62), .C(n166), .Q(n115) );
  NOR22 U28 ( .A(A[11]), .B(n11), .Q(n139) );
  NOR21 U29 ( .A(A[0]), .B(n3), .Q(n110) );
  INV3 U30 ( .A(B[5]), .Q(n7) );
  INV1 U31 ( .A(A[1]), .Q(n176) );
  NAND22 U32 ( .A(n129), .B(n130), .Q(n33) );
  NAND23 U33 ( .A(n32), .B(n33), .Q(n25) );
  NAND22 U34 ( .A(A[6]), .B(n189), .Q(n42) );
  AOI210 U35 ( .A(n61), .B(n62), .C(n63), .Q(n60) );
  NAND22 U36 ( .A(n185), .B(n42), .Q(n133) );
  INV3 U37 ( .A(n115), .Q(n112) );
  NOR23 U38 ( .A(n137), .B(n145), .Q(n136) );
  INV3 U39 ( .A(n186), .Q(n122) );
  NAND33 U40 ( .A(n43), .B(n42), .C(n187), .Q(n186) );
  INV3 U41 ( .A(B[7]), .Q(n8) );
  INV3 U42 ( .A(B[2]), .Q(n4) );
  NOR21 U43 ( .A(n139), .B(n102), .Q(n101) );
  INV6 U44 ( .A(n162), .Q(n35) );
  NOR21 U45 ( .A(n110), .B(n111), .Q(n164) );
  NAND23 U46 ( .A(B[2]), .B(n13), .Q(n62) );
  IMUX21 U47 ( .A(n28), .B(n29), .S(n30), .Q(DIFF[8]) );
  NOR22 U48 ( .A(n31), .B(n25), .Q(n30) );
  XOR21 U49 ( .A(n46), .B(n47), .Q(DIFF[6]) );
  NAND22 U50 ( .A(A[1]), .B(n167), .Q(n67) );
  NOR22 U51 ( .A(A[3]), .B(n5), .Q(n175) );
  NAND22 U52 ( .A(n153), .B(n154), .Q(n149) );
  INV3 U53 ( .A(B[0]), .Q(n3) );
  INV3 U54 ( .A(A[8]), .Q(n15) );
  INV3 U55 ( .A(A[2]), .Q(n13) );
  INV3 U56 ( .A(A[4]), .Q(n14) );
  INV3 U57 ( .A(n72), .Q(n191) );
  NAND22 U58 ( .A(B[1]), .B(n176), .Q(n73) );
  XOR22 U59 ( .A(n157), .B(n158), .Q(DIFF[10]) );
  CLKIN3 U60 ( .A(n35), .Q(n57) );
  XNR22 U61 ( .A(n2), .B(n126), .Q(DIFF[12]) );
  NOR21 U62 ( .A(n122), .B(n123), .Q(n118) );
  NOR21 U63 ( .A(B[0]), .B(n12), .Q(n72) );
  INV3 U64 ( .A(n38), .Q(n131) );
  OAI222 U65 ( .A(n98), .B(n99), .C(B[12]), .D(n100), .Q(n97) );
  AOI212 U66 ( .A(n48), .B(n39), .C(n49), .Q(n47) );
  INV3 U67 ( .A(n25), .Q(n21) );
  NAND22 U68 ( .A(A[2]), .B(n4), .Q(n68) );
  CLKIN3 U69 ( .A(B[6]), .Q(n189) );
  AOI211 U70 ( .A(n50), .B(n35), .C(n53), .Q(n52) );
  AOI212 U71 ( .A(B[3]), .B(n169), .C(n170), .Q(n168) );
  NAND23 U72 ( .A(n168), .B(n73), .Q(n111) );
  NOR22 U73 ( .A(n152), .B(n159), .Q(n158) );
  AOI212 U74 ( .A(n153), .B(n154), .C(n160), .Q(n159) );
  NAND23 U75 ( .A(n86), .B(n81), .Q(n84) );
  NAND22 U76 ( .A(n76), .B(n78), .Q(n86) );
  OAI2112 U77 ( .A(n57), .B(n103), .C(n33), .D(n32), .Q(n128) );
  AOI312 U78 ( .A(n116), .B(n117), .C(n118), .D(n119), .Q(n92) );
  INV1 U79 ( .A(A[3]), .Q(n169) );
  NAND21 U80 ( .A(A[4]), .B(n6), .Q(n45) );
  INV3 U81 ( .A(B[4]), .Q(n6) );
  NAND24 U82 ( .A(n92), .B(n93), .Q(n78) );
  NAND22 U83 ( .A(A[9]), .B(n138), .Q(n27) );
  XOR22 U84 ( .A(n17), .B(n18), .Q(DIFF[9]) );
  AOI212 U85 ( .A(n21), .B(n22), .C(n23), .Q(n20) );
  XOR22 U86 ( .A(n74), .B(n75), .Q(DIFF[15]) );
  CLKIN2 U87 ( .A(B[10]), .Q(n10) );
  NOR32 U88 ( .A(n163), .B(n164), .C(n165), .Q(n162) );
  NAND20 U89 ( .A(n62), .B(n68), .Q(n64) );
  INV6 U90 ( .A(n62), .Q(n170) );
  INV3 U91 ( .A(B[1]), .Q(n167) );
  NOR23 U92 ( .A(A[8]), .B(n9), .Q(n137) );
  NAND24 U93 ( .A(n34), .B(n35), .Q(n154) );
  OAI2111 U94 ( .A(n122), .B(n182), .C(n32), .D(n36), .Q(n181) );
  NAND31 U95 ( .A(n133), .B(n124), .C(n38), .Q(n182) );
  INV2 U96 ( .A(A[12]), .Q(n100) );
  INV6 U97 ( .A(n67), .Q(n166) );
  NOR21 U98 ( .A(n132), .B(n125), .Q(n129) );
  NOR22 U99 ( .A(n19), .B(n20), .Q(n18) );
  NOR21 U100 ( .A(n131), .B(n122), .Q(n130) );
  NAND22 U101 ( .A(A[5]), .B(n7), .Q(n43) );
  CLKIN2 U102 ( .A(n110), .Q(n109) );
  CLKIN2 U103 ( .A(n45), .Q(n53) );
  INV0 U104 ( .A(B[13]), .Q(n90) );
  INV2 U105 ( .A(n101), .Q(n99) );
  NAND21 U106 ( .A(B[8]), .B(n15), .Q(n24) );
  XOR20 U107 ( .A(B[8]), .B(A[8]), .Q(n29) );
  AOI210 U108 ( .A(B[8]), .B(n15), .C(n19), .Q(n28) );
  NAND20 U109 ( .A(n12), .B(B[0]), .Q(n190) );
  AOI312 U110 ( .A(n135), .B(n140), .C(n141), .D(n142), .Q(n98) );
  NAND20 U111 ( .A(n39), .B(n43), .Q(n51) );
  NAND20 U112 ( .A(n151), .B(n143), .Q(n150) );
  XOR20 U113 ( .A(B[11]), .B(A[11]), .Q(n147) );
  NOR20 U114 ( .A(A[0]), .B(n3), .Q(n71) );
  CLKIN3 U115 ( .A(n54), .Q(n50) );
  CLKIN0 U116 ( .A(n135), .Q(n155) );
  NOR22 U117 ( .A(A[9]), .B(n138), .Q(n145) );
  XNR20 U118 ( .A(B[7]), .B(A[7]), .Q(n1) );
  NAND20 U119 ( .A(n38), .B(n42), .Q(n46) );
  NAND21 U120 ( .A(n124), .B(n38), .Q(n123) );
  NOR20 U121 ( .A(n58), .B(n53), .Q(n55) );
  IMUX20 U122 ( .A(n55), .B(n56), .S(n57), .Q(DIFF[4]) );
  NAND20 U123 ( .A(n73), .B(n67), .Q(n69) );
  XOR20 U124 ( .A(n69), .B(n66), .Q(DIFF[1]) );
  NAND22 U125 ( .A(n190), .B(n191), .Q(DIFF[0]) );
  NAND22 U126 ( .A(n45), .B(n44), .Q(n48) );
  NAND22 U127 ( .A(n152), .B(n135), .Q(n151) );
  INV3 U128 ( .A(n104), .Q(n117) );
  INV3 U129 ( .A(n98), .Q(n127) );
  INV3 U130 ( .A(n145), .Q(n140) );
  NAND22 U131 ( .A(n143), .B(n144), .Q(n142) );
  NAND22 U132 ( .A(B[10]), .B(n16), .Q(n135) );
  INV3 U133 ( .A(A[10]), .Q(n16) );
  NAND22 U134 ( .A(A[10]), .B(n10), .Q(n143) );
  NAND22 U135 ( .A(n26), .B(n27), .Q(n17) );
  XOR21 U136 ( .A(n51), .B(n52), .Q(DIFF[5]) );
  NAND22 U137 ( .A(n191), .B(n71), .Q(n70) );
  NAND22 U138 ( .A(A[8]), .B(n9), .Q(n36) );
  NOR21 U139 ( .A(n155), .B(n156), .Q(n148) );
  XNR21 U140 ( .A(n64), .B(n61), .Q(DIFF[2]) );
  NAND22 U141 ( .A(A[11]), .B(n11), .Q(n144) );
  NAND22 U142 ( .A(n135), .B(n143), .Q(n157) );
  NOR20 U143 ( .A(A[4]), .B(n6), .Q(n58) );
  NOR21 U144 ( .A(A[2]), .B(n4), .Q(n174) );
  NAND22 U145 ( .A(n26), .B(n24), .Q(n160) );
  NOR20 U146 ( .A(A[4]), .B(n6), .Q(n54) );
  NAND22 U147 ( .A(n108), .B(n109), .Q(n106) );
  INV3 U148 ( .A(B[11]), .Q(n11) );
  NOR32 U149 ( .A(n12), .B(B[0]), .C(n174), .Q(n172) );
  NAND22 U150 ( .A(A[7]), .B(n8), .Q(n32) );
  INV3 U151 ( .A(n188), .Q(n187) );
  XNR21 U152 ( .A(n1), .B(n37), .Q(DIFF[7]) );
  NAND22 U153 ( .A(B[5]), .B(n180), .Q(n39) );
  INV3 U154 ( .A(A[5]), .Q(n180) );
  NAND22 U155 ( .A(B[9]), .B(n161), .Q(n26) );
  INV3 U156 ( .A(A[9]), .Q(n161) );
  NAND22 U157 ( .A(B[7]), .B(n184), .Q(n124) );
  INV3 U158 ( .A(A[7]), .Q(n184) );
  NAND22 U159 ( .A(n63), .B(n171), .Q(n114) );
  INV3 U160 ( .A(B[9]), .Q(n138) );
  INV3 U161 ( .A(n181), .Q(n153) );
  INV6 U162 ( .A(B[3]), .Q(n5) );
  INV3 U163 ( .A(B[14]), .Q(n83) );
  NAND22 U164 ( .A(B[6]), .B(n183), .Q(n38) );
  INV3 U165 ( .A(n80), .Q(n77) );
  XNR21 U166 ( .A(n59), .B(n60), .Q(DIFF[3]) );
  INV3 U167 ( .A(n89), .Q(n76) );
  INV3 U168 ( .A(n87), .Q(n81) );
  NOR21 U169 ( .A(B[13]), .B(n88), .Q(n87) );
  INV3 U170 ( .A(A[13]), .Q(n88) );
  NAND22 U171 ( .A(n114), .B(n115), .Q(n165) );
  NOR22 U172 ( .A(A[7]), .B(n8), .Q(n179) );
  NOR20 U173 ( .A(A[14]), .B(n83), .Q(n80) );
  XNR20 U174 ( .A(B[12]), .B(A[12]), .Q(n2) );
  XOR20 U175 ( .A(B[4]), .B(A[4]), .Q(n56) );
  XOR20 U176 ( .A(B[15]), .B(A[15]), .Q(n75) );
  NOR21 U177 ( .A(n102), .B(n125), .Q(n116) );
  XOR20 U178 ( .A(n91), .B(n78), .Q(DIFF[13]) );
  NOR21 U179 ( .A(A[13]), .B(n90), .Q(n89) );
  XNR20 U180 ( .A(B[13]), .B(A[13]), .Q(n91) );
  INV2 U181 ( .A(A[6]), .Q(n183) );
  NOR21 U182 ( .A(A[5]), .B(n7), .Q(n185) );
  XNR20 U183 ( .A(B[14]), .B(A[14]), .Q(n85) );
  CLKIN0 U184 ( .A(A[14]), .Q(n82) );
  XNR20 U185 ( .A(B[3]), .B(A[3]), .Q(n59) );
  CLKIN3 U186 ( .A(n24), .Q(n23) );
  CLKIN3 U187 ( .A(n36), .Q(n19) );
  AOI312 U188 ( .A(n38), .B(n39), .C(n40), .D(n41), .Q(n37) );
  CLKIN3 U189 ( .A(n43), .Q(n49) );
  OAI212 U190 ( .A(n65), .B(n66), .C(n67), .Q(n61) );
  CLKIN3 U191 ( .A(n70), .Q(n66) );
  AOI312 U192 ( .A(n76), .B(n77), .C(n78), .D(n79), .Q(n74) );
  OAI222 U193 ( .A(n80), .B(n81), .C(B[14]), .D(n82), .Q(n79) );
  AOI312 U194 ( .A(n94), .B(n95), .C(n96), .D(n97), .Q(n93) );
  CLKIN3 U195 ( .A(n111), .Q(n108) );
  CLKIN3 U196 ( .A(n114), .Q(n113) );
  CLKIN3 U197 ( .A(n32), .Q(n121) );
  AOI222 U198 ( .A(n127), .B(n134), .C(n117), .D(n128), .Q(n126) );
  CLKIN3 U199 ( .A(n133), .Q(n125) );
  CLKIN3 U200 ( .A(n124), .Q(n132) );
  OAI212 U201 ( .A(B[8]), .B(n15), .C(n27), .Q(n141) );
  AOI312 U202 ( .A(n148), .B(n24), .C(n149), .D(n150), .Q(n146) );
  CLKIN3 U203 ( .A(n26), .Q(n156) );
  CLKIN3 U204 ( .A(n68), .Q(n63) );
  CLKIN3 U205 ( .A(n73), .Q(n65) );
  AOI312 U206 ( .A(n73), .B(n171), .C(n172), .D(n173), .Q(n107) );
  CLKIN3 U207 ( .A(n103), .Q(n34) );
  NOR24 U208 ( .A(A[4]), .B(n6), .Q(n178) );
  CLKIN3 U209 ( .A(n27), .Q(n152) );
endmodule


module E_alu ( o_data_AluRes, i_data_A, i_data_B, i_con_AluCtrl, i_data_shamt
 );
  output [31:0] o_data_AluRes;
  input [31:0] i_data_A;
  input [31:0] i_data_B;
  input [3:0] i_con_AluCtrl;
  input [4:0] i_data_shamt;
  wire   N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N306, n41, n42,
         n139, n161, n169, n176, n183, n190, n198, n218, n219, n220, n221,
         n333, n428, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n162, n163, n164, n165, n166, n167,
         n168, n170, n171, n172, n173, n174, n175, n177, n178, n179, n180,
         n181, n182, n184, n185, n186, n187, n188, n189, n191, n192, n193,
         n194, n195, n196, n197, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545;
  wire   [8:0] sum_1;
  wire   [8:0] pre_sum_2a;
  wire   [8:0] pre_sum_2b;
  wire   [8:0] pre_sum_3a;
  wire   [8:0] pre_sum_3b;
  wire   [7:0] pre_sum_4a;
  wire   [7:0] pre_sum_4b;
  wire   [16:0] half_sub;
  wire   [15:0] pre_suba;
  wire   [15:0] pre_subb;

  E_alu_DW01_sub_3 sub_33 ( .A({n42, i_data_A[15:12], n30, n115, i_data_A[9:4], 
        n46, i_data_A[2:0]}), .B({n42, n79, n77, i_data_B[13:12], n105, n103, 
        n75, n101, i_data_B[7:0]}), .CI(n42), .DIFF(half_sub) );
  E_alu_DW01_add_7 add_25 ( .A({n42, i_data_A[7:4], n46, i_data_A[2:0]}), .B({
        n42, i_data_B[7:0]}), .CI(n42), .SUM(sum_1) );
  E_alu_DW01_add_12 add_1_root_add_31_2 ( .A({n88, i_data_A[30:28], n126, n124, 
        i_data_A[25], n122}), .B({n113, n86, n85, n112, n111, n64, n83, n62}), 
        .CI(n41), .SUM(pre_sum_4b) );
  E_alu_DW01_add_13 add_30 ( .A({n88, i_data_A[30:28], n126, n124, 
        i_data_A[25], n122}), .B({n113, n86, n85, n112, n67, n64, n83, n63}), 
        .CI(n42), .SUM(pre_sum_4a) );
  E_alu_DW01_ash_1 sll_56 ( .A({n113, n86, n85, n112, n67, n65, n83, n62, n61, 
        n81, n60, n56, n55, n110, i_data_B[17], n109, n79, n77, n76, 
        i_data_B[12], n105, n103, n74, n101, i_data_B[7:0]}), .DATA_TC(n42), 
        .SH(i_data_shamt), .SH_TC(n42), .B({N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, 
        N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193}) );
  E_alu_DW01_add_18 add_28 ( .A({n42, i_data_A[23:21], n120, i_data_A[19:17], 
        n117}), .B({n42, n61, n82, n60, n56, n54, n110, i_data_B[17], n109}), 
        .CI(n42), .SUM(pre_sum_3a) );
  E_alu_DW01_add_17 add_1_root_add_29_2 ( .A({n42, i_data_A[23:21], n120, 
        i_data_A[19:17], n117}), .B({n42, n61, n82, n60, n56, n54, n110, 
        i_data_B[17], n109}), .CI(n41), .SUM(pre_sum_3b) );
  E_alu_DW01_cmp2_2 r131 ( .A({n87, i_data_A[30:28], n126, n124, i_data_A[25], 
        n122, i_data_A[23:21], n120, i_data_A[19:17], n117, i_data_A[15:12], 
        n30, n115, i_data_A[9:4], n46, i_data_A[2:0]}), .B({n113, n86, n85, 
        n112, n111, n65, n84, n62, n61, n81, n59, n56, n54, n110, i_data_B[17], 
        n109, n80, n78, n76, i_data_B[12], n105, n103, n75, n101, 
        i_data_B[7:6], n7, i_data_B[4:0]}), .LEQ(n42), .TC(n42), .LT_LE(N306)
         );
  E_alu_DW01_add_15 add_26 ( .A({n42, i_data_A[15:12], n30, n115, 
        i_data_A[9:8]}), .B({n42, n80, n78, i_data_B[13:12], n105, n103, n74, 
        n101}), .CI(n42), .SUM(pre_sum_2a) );
  E_alu_DW01_add_16 add_1_root_add_27_2 ( .A({n42, i_data_A[15:12], n30, n115, 
        i_data_A[9:8]}), .B({n42, n79, n78, i_data_B[13:12], n105, n103, n74, 
        n101}), .CI(n41), .SUM(pre_sum_2b) );
  E_alu_DW_rash_3 r130 ( .A({n113, n86, n85, n112, n66, n65, n84, n62, n61, 
        n81, n59, n56, n54, n110, i_data_B[17], n109, n80, n77, n76, 
        i_data_B[12], n105, n103, n75, n101, i_data_B[7:6], n7, i_data_B[4], 
        n2, i_data_B[2:0]}), .DATA_TC(n42), .SH(i_data_shamt), .SH_TC(n42), 
        .B({N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, 
        N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, 
        N233, N232, N231, N230, N229, N228, N227, N226, N225}) );
  E_alu_DW01_sub_10 sub_1_root_sub_35_2 ( .A({n87, i_data_A[30:28], n126, n124, 
        i_data_A[25], n122, i_data_A[23:21], n120, i_data_A[19:17], n117}), 
        .B({n113, n86, n85, n112, n111, i_data_B[26], n84, n63, n61, n82, n60, 
        n57, n54, n110, i_data_B[17], n109}), .CI(n41), .DIFF(pre_subb) );
  E_alu_DW01_sub_11 sub_34 ( .A({n87, i_data_A[30:28], n126, n124, 
        i_data_A[25], n122, i_data_A[23:21], n120, i_data_A[19:17], n117}), 
        .B({n113, n86, n85, n112, n66, n64, n84, n62, n61, n82, n59, n56, n55, 
        n110, i_data_B[17], n109}), .CI(n42), .DIFF(pre_suba) );
  AOI222 U3 ( .A(pre_subb[11]), .B(n524), .C(n523), .D(pre_suba[11]), .Q(n472)
         );
  NAND24 U4 ( .A(n388), .B(n389), .Q(n5) );
  INV15 U5 ( .A(n305), .Q(n400) );
  INV4 U6 ( .A(i_con_AluCtrl[1]), .Q(n136) );
  AOI212 U7 ( .A(n96), .B(n392), .C(n10), .Q(n36) );
  CLKBU15 U8 ( .A(n111), .Q(n66) );
  BUF6 U9 ( .A(n100), .Q(n97) );
  BUF6 U10 ( .A(i_data_B[9]), .Q(n75) );
  NAND21 U11 ( .A(n232), .B(n231), .Q(n233) );
  IMUX31 U12 ( .A(n526), .B(n96), .C(n174), .S0(i_data_A[4]), .S1(i_data_B[4]), 
        .Q(n175) );
  INV12 U13 ( .A(n536), .Q(n483) );
  INV2 U14 ( .A(n495), .Q(n28) );
  NAND28 U15 ( .A(n411), .B(pre_sum_3b[8]), .Q(n521) );
  CLKIN10 U16 ( .A(n58), .Q(n60) );
  OAI210 U17 ( .A(n11), .B(n295), .C(n117), .Q(n300) );
  IMUX31 U18 ( .A(n526), .B(n96), .C(n195), .S0(i_data_A[7]), .S1(i_data_B[7]), 
        .Q(n199) );
  OAI210 U19 ( .A(n10), .B(n230), .C(n115), .Q(n231) );
  CLKIN12 U20 ( .A(n545), .Q(n100) );
  CLKIN15 U21 ( .A(n51), .Q(n436) );
  AOI222 U22 ( .A(N206), .B(n70), .C(half_sub[13]), .D(n1), .Q(n267) );
  INV12 U23 ( .A(n121), .Q(n120) );
  INV10 U24 ( .A(i_data_A[10]), .Q(n116) );
  NAND24 U25 ( .A(pre_subb[6]), .B(n524), .Q(n389) );
  NAND24 U26 ( .A(pre_subb[4]), .B(n524), .Q(n363) );
  NAND24 U27 ( .A(pre_subb[0]), .B(n524), .Q(n313) );
  NAND24 U28 ( .A(pre_subb[2]), .B(n524), .Q(n338) );
  AOI222 U29 ( .A(pre_subb[8]), .B(n524), .C(pre_suba[8]), .D(n523), .Q(n419)
         );
  CLKIN15 U30 ( .A(n303), .Q(n524) );
  BUF12 U31 ( .A(sum_1[8]), .Q(n51) );
  INV12 U32 ( .A(pre_sum_2b[8]), .Q(n437) );
  AOI221 U33 ( .A(pre_sum_3b[6]), .B(n400), .C(pre_sum_3a[6]), .D(n399), .Q(
        n388) );
  CLKBU12 U34 ( .A(n309), .Q(n1) );
  NAND33 U35 ( .A(n135), .B(n293), .C(n136), .Q(n503) );
  BUF12 U36 ( .A(i_data_B[15]), .Q(n80) );
  INV6 U37 ( .A(i_data_B[11]), .Q(n106) );
  INV12 U38 ( .A(pre_sum_2a[8]), .Q(n422) );
  NAND26 U39 ( .A(n414), .B(n441), .Q(n495) );
  AOI2111 U40 ( .A(N234), .B(n91), .C(n222), .D(n217), .Q(n226) );
  INV3 U41 ( .A(i_data_A[16]), .Q(n118) );
  IMUX21 U42 ( .A(n318), .B(n317), .S(i_data_B[17]), .Q(n319) );
  INV6 U43 ( .A(n118), .Q(n117) );
  BUF8 U44 ( .A(i_data_A[11]), .Q(n30) );
  AOI211 U45 ( .A(N246), .B(n92), .C(n369), .Q(n370) );
  IMUX21 U46 ( .A(n343), .B(n342), .S(n55), .Q(n344) );
  INV3 U47 ( .A(n544), .Q(n527) );
  NAND33 U48 ( .A(n27), .B(n294), .C(n292), .Q(n139) );
  NOR32 U49 ( .A(n47), .B(n48), .C(n26), .Q(n49) );
  INV3 U50 ( .A(n372), .Q(n7) );
  AOI2111 U51 ( .A(N240), .B(n91), .C(n285), .D(n284), .Q(n291) );
  AOI211 U52 ( .A(N203), .B(n71), .C(n233), .Q(n235) );
  AOI311 U53 ( .A(n28), .B(n536), .C(pre_sum_4b[7]), .D(n535), .Q(n538) );
  CLKIN8 U54 ( .A(n503), .Q(n542) );
  INV12 U55 ( .A(n53), .Q(n54) );
  AOI222 U56 ( .A(pre_sum_3b[7]), .B(n400), .C(pre_sum_3a[7]), .D(n399), .Q(
        n402) );
  NAND21 U57 ( .A(n52), .B(n437), .Q(n440) );
  NAND23 U58 ( .A(n142), .B(n293), .Q(n143) );
  NAND23 U59 ( .A(pre_sum_2b[3]), .B(n287), .Q(n240) );
  CLKBU12 U60 ( .A(i_data_B[9]), .Q(n74) );
  NAND34 U61 ( .A(n312), .B(n311), .C(n313), .Q(n19) );
  OAI312 U62 ( .A(n151), .B(n530), .C(n145), .D(n144), .Q(n146) );
  BUF12 U63 ( .A(i_con_AluCtrl[2]), .Q(n27) );
  INV3 U64 ( .A(n137), .Q(n532) );
  NAND22 U65 ( .A(pre_suba[5]), .B(n523), .Q(n374) );
  NAND22 U66 ( .A(pre_suba[3]), .B(n523), .Q(n349) );
  NAND23 U67 ( .A(pre_suba[1]), .B(n523), .Q(n324) );
  AOI221 U68 ( .A(N200), .B(n522), .C(half_sub[7]), .D(n1), .Q(n197) );
  NAND21 U69 ( .A(N201), .B(n522), .Q(n210) );
  NAND21 U70 ( .A(N195), .B(n522), .Q(n166) );
  NAND21 U71 ( .A(N204), .B(n522), .Q(n239) );
  NAND21 U72 ( .A(N193), .B(n522), .Q(n144) );
  BUF6 U73 ( .A(i_data_B[13]), .Q(n76) );
  NAND23 U74 ( .A(n324), .B(n325), .Q(n23) );
  NAND21 U75 ( .A(pre_subb[1]), .B(n524), .Q(n326) );
  NAND21 U76 ( .A(pre_subb[7]), .B(n524), .Q(n403) );
  NAND21 U77 ( .A(pre_subb[3]), .B(n524), .Q(n351) );
  NAND21 U78 ( .A(pre_subb[5]), .B(n524), .Q(n376) );
  OAI2110 U79 ( .A(i_data_A[7]), .B(n21), .C(n14), .D(n161), .Q(n195) );
  NAND20 U80 ( .A(i_data_A[7]), .B(n32), .Q(n161) );
  AOI220 U81 ( .A(sum_1[5]), .B(n441), .C(i_data_A[5]), .D(n90), .Q(n182) );
  OAI210 U82 ( .A(n89), .B(n353), .C(n120), .Q(n358) );
  AOI210 U83 ( .A(n99), .B(n281), .C(n90), .Q(n282) );
  NAND21 U84 ( .A(pre_suba[7]), .B(n523), .Q(n401) );
  NAND21 U85 ( .A(pre_suba[14]), .B(n523), .Q(n518) );
  INV2 U86 ( .A(i_con_AluCtrl[0]), .Q(n292) );
  BUF12 U87 ( .A(i_con_AluCtrl[0]), .Q(n37) );
  INV3 U88 ( .A(i_con_AluCtrl[3]), .Q(n135) );
  CLKIN12 U89 ( .A(n495), .Q(n537) );
  INV8 U90 ( .A(n125), .Q(n124) );
  INV12 U91 ( .A(n127), .Q(n126) );
  NAND22 U92 ( .A(n450), .B(n449), .Q(o_data_AluRes[25]) );
  INV3 U93 ( .A(n138), .Q(n309) );
  IMUX31 U94 ( .A(n139), .B(n22), .C(n130), .S0(i_data_A[0]), .S1(n50), .Q(
        n149) );
  INV12 U95 ( .A(n139), .Q(n526) );
  CLKBU12 U96 ( .A(n503), .Q(n16) );
  BUF6 U97 ( .A(n532), .Q(n92) );
  INV12 U98 ( .A(n143), .Q(n522) );
  NAND31 U99 ( .A(n27), .B(n141), .C(n292), .Q(n138) );
  INV6 U100 ( .A(i_data_B[21]), .Q(n58) );
  INV3 U101 ( .A(i_data_A[20]), .Q(n121) );
  BUF6 U102 ( .A(i_data_B[22]), .Q(n81) );
  INV8 U103 ( .A(i_data_B[8]), .Q(n102) );
  INV3 U104 ( .A(i_data_A[24]), .Q(n123) );
  BUF6 U105 ( .A(i_data_B[24]), .Q(n63) );
  INV6 U106 ( .A(n123), .Q(n122) );
  CLKIN8 U107 ( .A(n128), .Q(n294) );
  INV3 U108 ( .A(i_data_B[12]), .Q(n108) );
  CLKBU12 U109 ( .A(i_data_A[3]), .Q(n46) );
  NAND23 U110 ( .A(n338), .B(n337), .Q(n40) );
  OAI2110 U111 ( .A(i_data_A[6]), .B(n21), .C(n169), .D(n544), .Q(n186) );
  CLKIN4 U112 ( .A(n544), .Q(n12) );
  NAND22 U113 ( .A(half_sub[10]), .B(n1), .Q(n234) );
  INV3 U114 ( .A(n521), .Q(n48) );
  AOI221 U115 ( .A(pre_subb[15]), .B(n524), .C(pre_suba[15]), .D(n523), .Q(
        n539) );
  AOI221 U116 ( .A(pre_subb[9]), .B(n524), .C(pre_suba[9]), .D(n523), .Q(n449)
         );
  NAND42 U117 ( .A(n261), .B(n260), .C(n259), .D(n258), .Q(o_data_AluRes[12])
         );
  INV3 U118 ( .A(i_data_A[27]), .Q(n127) );
  CLKIN6 U119 ( .A(i_data_B[19]), .Q(n53) );
  INV3 U120 ( .A(n38), .Q(n425) );
  INV8 U121 ( .A(pre_sum_3b[8]), .Q(n439) );
  IMUX21 U122 ( .A(n330), .B(n329), .S(n110), .Q(n331) );
  INV8 U123 ( .A(n116), .Q(n115) );
  INV3 U124 ( .A(n98), .Q(n39) );
  IMUX21 U125 ( .A(n368), .B(n367), .S(n60), .Q(n369) );
  INV8 U126 ( .A(n114), .Q(n113) );
  BUF6 U127 ( .A(sum_1[8]), .Q(n52) );
  OAI2111 U128 ( .A(n46), .B(n21), .C(n14), .D(n190), .Q(n168) );
  NAND23 U129 ( .A(n362), .B(n363), .Q(n3) );
  AOI221 U130 ( .A(n400), .B(pre_sum_3b[4]), .C(pre_sum_3a[4]), .D(n399), .Q(
        n362) );
  AOI211 U131 ( .A(n99), .B(n272), .C(n11), .Q(n270) );
  AOI211 U132 ( .A(n280), .B(n15), .C(n281), .Q(n285) );
  AOI211 U133 ( .A(n99), .B(n250), .C(n89), .Q(n251) );
  NAND23 U134 ( .A(half_sub[12]), .B(n1), .Q(n258) );
  AOI221 U135 ( .A(pre_sum_3b[0]), .B(n400), .C(pre_sum_3a[0]), .D(n399), .Q(
        n312) );
  NAND22 U136 ( .A(pre_suba[0]), .B(n523), .Q(n311) );
  AOI211 U137 ( .A(N247), .B(n92), .C(n382), .Q(n383) );
  INV3 U138 ( .A(n40), .Q(n43) );
  AOI211 U139 ( .A(N231), .B(n93), .C(n189), .Q(n194) );
  INV3 U140 ( .A(n17), .Q(n18) );
  NAND42 U141 ( .A(n474), .B(n473), .C(n472), .D(n471), .Q(o_data_AluRes[27])
         );
  NOR22 U142 ( .A(n49), .B(n470), .Q(n471) );
  NAND31 U143 ( .A(pre_sum_4a[7]), .B(n521), .C(n25), .Q(n541) );
  NAND42 U144 ( .A(n520), .B(n519), .C(n518), .D(n517), .Q(o_data_AluRes[30])
         );
  AOI221 U145 ( .A(pre_sum_3b[3]), .B(n400), .C(pre_sum_3a[3]), .D(n399), .Q(
        n350) );
  NOR31 U146 ( .A(pre_sum_2b[8]), .B(pre_sum_3a[8]), .C(n436), .Q(n435) );
  INV12 U147 ( .A(n104), .Q(n103) );
  AOI211 U148 ( .A(N211), .B(n522), .C(n335), .Q(n339) );
  NAND21 U149 ( .A(N202), .B(n522), .Q(n224) );
  NAND21 U150 ( .A(N223), .B(n522), .Q(n519) );
  NAND21 U151 ( .A(N205), .B(n522), .Q(n260) );
  AOI211 U152 ( .A(N212), .B(n522), .C(n348), .Q(n352) );
  CLKBU12 U153 ( .A(i_data_B[20]), .Q(n56) );
  INV6 U154 ( .A(n544), .Q(n11) );
  BUF8 U155 ( .A(i_data_B[24]), .Q(n62) );
  BUF2 U156 ( .A(n527), .Q(n90) );
  CLKBU12 U157 ( .A(i_data_B[30]), .Q(n86) );
  BUF8 U158 ( .A(i_data_B[26]), .Q(n64) );
  BUF6 U159 ( .A(i_data_B[26]), .Q(n65) );
  CLKBU12 U160 ( .A(i_data_B[23]), .Q(n61) );
  INV6 U161 ( .A(n25), .Q(n26) );
  BUF12 U162 ( .A(i_data_B[29]), .Q(n85) );
  NAND23 U163 ( .A(n33), .B(n135), .Q(n131) );
  CLKBU12 U164 ( .A(n111), .Q(n67) );
  BUF2 U165 ( .A(n544), .Q(n68) );
  BUF12 U166 ( .A(i_data_B[14]), .Q(n78) );
  INV6 U167 ( .A(n19), .Q(n20) );
  CLKIN6 U168 ( .A(pre_sum_3a[8]), .Q(n443) );
  CLKIN3 U169 ( .A(n347), .Q(n2) );
  INV3 U170 ( .A(i_data_B[3]), .Q(n347) );
  INV3 U171 ( .A(pre_sum_4b[3]), .Q(n469) );
  INV2 U172 ( .A(n150), .Q(n142) );
  OAI2111 U173 ( .A(i_data_A[4]), .B(n21), .C(n15), .D(n183), .Q(n174) );
  NAND26 U174 ( .A(n1), .B(n308), .Q(n310) );
  AOI212 U175 ( .A(n97), .B(n366), .C(n11), .Q(n367) );
  AOI222 U176 ( .A(N196), .B(n70), .C(N228), .D(n92), .Q(n173) );
  AOI2112 U177 ( .A(N253), .B(n91), .C(n481), .D(n480), .Q(n488) );
  NAND28 U178 ( .A(n415), .B(n439), .Q(n536) );
  IMUX20 U179 ( .A(n97), .B(n32), .S(n80), .Q(n280) );
  CLKIN6 U180 ( .A(n515), .Q(n25) );
  BUF6 U181 ( .A(n100), .Q(n96) );
  CLKIN6 U182 ( .A(n95), .Q(n22) );
  NAND21 U183 ( .A(pre_suba[13]), .B(n523), .Q(n500) );
  CLKBU12 U184 ( .A(i_data_B[25]), .Q(n83) );
  AOI212 U185 ( .A(N248), .B(n92), .C(n394), .Q(n395) );
  AOI212 U186 ( .A(N242), .B(n92), .C(n319), .Q(n320) );
  AOI222 U187 ( .A(pre_sum_3b[1]), .B(n400), .C(pre_sum_3a[1]), .D(n399), .Q(
        n325) );
  IMUX23 U188 ( .A(n422), .B(n437), .S(n51), .Q(n304) );
  NAND22 U189 ( .A(n428), .B(n68), .Q(n129) );
  AOI210 U190 ( .A(n97), .B(n134), .C(n129), .Q(n130) );
  NAND33 U191 ( .A(n364), .B(n361), .C(n4), .Q(o_data_AluRes[20]) );
  INV6 U192 ( .A(n3), .Q(n4) );
  NAND21 U193 ( .A(pre_suba[4]), .B(n523), .Q(n361) );
  AOI312 U194 ( .A(pre_sum_4a[4]), .B(n521), .C(n25), .D(n484), .Q(n485) );
  NAND33 U195 ( .A(n390), .B(n387), .C(n6), .Q(o_data_AluRes[22]) );
  INV6 U196 ( .A(n5), .Q(n6) );
  AOI211 U197 ( .A(N215), .B(n70), .C(n386), .Q(n390) );
  OAI2111 U198 ( .A(n73), .B(n385), .C(n384), .D(n383), .Q(n386) );
  AOI222 U199 ( .A(N225), .B(n92), .C(half_sub[0]), .D(n1), .Q(n140) );
  AOI212 U200 ( .A(n98), .B(n341), .C(n11), .Q(n342) );
  AOI211 U201 ( .A(n99), .B(n116), .C(n10), .Q(n227) );
  AOI212 U202 ( .A(N245), .B(n92), .C(n356), .Q(n357) );
  AOI212 U203 ( .A(N214), .B(n522), .C(n373), .Q(n377) );
  CLKBU4 U204 ( .A(i_data_B[14]), .Q(n77) );
  INV10 U205 ( .A(n544), .Q(n10) );
  NAND24 U206 ( .A(i_con_AluCtrl[3]), .B(n136), .Q(n128) );
  AOI211 U207 ( .A(n213), .B(n15), .C(n214), .Q(n222) );
  AOI2112 U208 ( .A(N236), .B(n91), .C(n247), .D(n246), .Q(n249) );
  CLKIN0 U209 ( .A(i_data_B[1]), .Q(n322) );
  NAND33 U210 ( .A(n327), .B(n326), .C(n24), .Q(o_data_AluRes[17]) );
  AOI212 U211 ( .A(N241), .B(n92), .C(n298), .Q(n299) );
  IMUX21 U212 ( .A(n297), .B(n296), .S(n109), .Q(n298) );
  AOI212 U213 ( .A(N244), .B(n92), .C(n344), .Q(n345) );
  NAND23 U214 ( .A(N306), .B(n153), .Q(n154) );
  AOI222 U215 ( .A(n436), .B(n422), .C(n52), .D(n437), .Q(n411) );
  AOI212 U216 ( .A(n98), .B(n379), .C(n10), .Q(n380) );
  NOR32 U217 ( .A(pre_sum_3a[8]), .B(pre_sum_2a[8]), .C(n51), .Q(n413) );
  AOI221 U218 ( .A(n219), .B(n543), .C(i_data_B[2]), .D(n220), .Q(n218) );
  INV4 U219 ( .A(n23), .Q(n24) );
  OAI2112 U220 ( .A(n73), .B(n301), .C(n300), .D(n299), .Q(n302) );
  AOI211 U221 ( .A(N243), .B(n92), .C(n331), .Q(n332) );
  CLKIN0 U222 ( .A(i_data_B[13]), .Q(n489) );
  NAND24 U223 ( .A(half_sub[16]), .B(n1), .Q(n303) );
  INV2 U224 ( .A(i_data_B[5]), .Q(n372) );
  NAND34 U225 ( .A(n27), .B(n37), .C(n294), .Q(n545) );
  AOI211 U226 ( .A(n98), .B(n316), .C(n11), .Q(n317) );
  AOI212 U227 ( .A(N216), .B(n69), .C(n398), .Q(n404) );
  AOI221 U228 ( .A(sum_1[3]), .B(n441), .C(n46), .D(n10), .Q(n171) );
  AOI220 U229 ( .A(i_data_A[13]), .B(n263), .C(pre_sum_2a[5]), .D(n286), .Q(
        n269) );
  AOI211 U230 ( .A(n98), .B(n121), .C(n12), .Q(n354) );
  CLKIN6 U231 ( .A(half_sub[16]), .Q(n308) );
  INV15 U232 ( .A(n310), .Q(n523) );
  AOI2112 U233 ( .A(N218), .B(n522), .C(n447), .D(n448), .Q(n450) );
  NOR32 U234 ( .A(n446), .B(n445), .C(n444), .Q(n447) );
  MUX21 U235 ( .A(n526), .B(n96), .S(i_data_A[6]), .Q(n8) );
  IMUX21 U236 ( .A(n8), .B(n186), .S(i_data_B[6]), .Q(n187) );
  NAND42 U237 ( .A(n242), .B(n241), .C(n240), .D(n239), .Q(n247) );
  CLKIN6 U238 ( .A(n95), .Q(n21) );
  BUF15 U239 ( .A(n100), .Q(n95) );
  OAI2112 U240 ( .A(n73), .B(n372), .C(n371), .D(n370), .Q(n373) );
  AOI222 U241 ( .A(pre_sum_2b[8]), .B(n52), .C(pre_sum_2a[8]), .D(n436), .Q(
        n306) );
  CLKIN12 U242 ( .A(n307), .Q(n399) );
  NAND24 U243 ( .A(n306), .B(n441), .Q(n307) );
  NAND42 U244 ( .A(n226), .B(n225), .C(n224), .D(n223), .Q(o_data_AluRes[9])
         );
  OAI2112 U245 ( .A(n73), .B(n397), .C(n396), .D(n395), .Q(n398) );
  CLKIN4 U246 ( .A(n58), .Q(n59) );
  NAND24 U247 ( .A(n441), .B(n304), .Q(n305) );
  OAI210 U248 ( .A(n11), .B(n238), .C(n30), .Q(n241) );
  INV12 U249 ( .A(n208), .Q(n286) );
  NAND26 U250 ( .A(n441), .B(n436), .Q(n208) );
  NAND26 U251 ( .A(n537), .B(n536), .Q(n512) );
  NAND33 U252 ( .A(n234), .B(n237), .C(n236), .Q(n17) );
  NOR41 U253 ( .A(n149), .B(n148), .C(n147), .D(n146), .Q(n155) );
  AOI212 U254 ( .A(N210), .B(n522), .C(n323), .Q(n327) );
  OAI2112 U255 ( .A(n73), .B(n322), .C(n321), .D(n320), .Q(n323) );
  IMUX21 U256 ( .A(n355), .B(n354), .S(n57), .Q(n356) );
  CLKBU4 U257 ( .A(i_data_B[20]), .Q(n57) );
  OAI312 U258 ( .A(n435), .B(n433), .C(n434), .D(n432), .Q(n448) );
  OAI2111 U259 ( .A(pre_sum_3b[8]), .B(n438), .C(pre_sum_4b[1]), .D(n441), .Q(
        n433) );
  AOI2112 U260 ( .A(N250), .B(n91), .C(n431), .D(n430), .Q(n432) );
  OAI2112 U261 ( .A(n73), .B(n359), .C(n358), .D(n357), .Q(n360) );
  NAND22 U262 ( .A(n436), .B(n422), .Q(n442) );
  AOI212 U263 ( .A(N213), .B(n522), .C(n360), .Q(n364) );
  OAI2112 U264 ( .A(n73), .B(n347), .C(n346), .D(n345), .Q(n348) );
  AOI222 U265 ( .A(pre_sum_3b[2]), .B(n400), .C(pre_sum_3a[2]), .D(n399), .Q(
        n337) );
  IMUX22 U266 ( .A(n426), .B(n425), .S(n84), .Q(n431) );
  BUF6 U267 ( .A(n132), .Q(n9) );
  CLKIN1 U268 ( .A(n527), .Q(n13) );
  CLKIN2 U269 ( .A(n11), .Q(n14) );
  INV3 U270 ( .A(n11), .Q(n15) );
  BUF6 U271 ( .A(n522), .Q(n70) );
  BUF6 U272 ( .A(n522), .Q(n69) );
  AOI211 U273 ( .A(n99), .B(n118), .C(n12), .Q(n296) );
  AOI211 U274 ( .A(n99), .B(n202), .C(n10), .Q(n203) );
  CLKBU12 U275 ( .A(n95), .Q(n99) );
  OAI211 U276 ( .A(n13), .B(n163), .C(n162), .Q(n164) );
  NAND28 U277 ( .A(n542), .B(n37), .Q(n544) );
  CLKBU4 U278 ( .A(n100), .Q(n98) );
  NAND42 U279 ( .A(n194), .B(n193), .C(n192), .D(n191), .Q(o_data_AluRes[6])
         );
  NAND21 U280 ( .A(sum_1[6]), .B(n441), .Q(n191) );
  NAND22 U281 ( .A(n235), .B(n18), .Q(o_data_AluRes[10]) );
  AOI211 U282 ( .A(pre_sum_2b[2]), .B(n287), .C(n229), .Q(n237) );
  NAND21 U283 ( .A(pre_sum_2a[2]), .B(n286), .Q(n236) );
  NAND22 U284 ( .A(n314), .B(n20), .Q(o_data_AluRes[16]) );
  AOI212 U285 ( .A(N209), .B(n71), .C(n302), .Q(n314) );
  CLKBU15 U286 ( .A(i_data_B[16]), .Q(n109) );
  NAND42 U287 ( .A(n291), .B(n290), .C(n289), .D(n288), .Q(o_data_AluRes[15])
         );
  NAND21 U288 ( .A(pre_suba[6]), .B(n523), .Q(n387) );
  AOI221 U289 ( .A(pre_sum_2a[6]), .B(n286), .C(pre_sum_2b[6]), .D(n287), .Q(
        n277) );
  CLKIN3 U290 ( .A(n95), .Q(n94) );
  CLKIN12 U291 ( .A(n9), .Q(n441) );
  CLKIN0 U292 ( .A(i_data_A[18]), .Q(n119) );
  NAND21 U293 ( .A(pre_sum_2a[8]), .B(n436), .Q(n438) );
  INV15 U294 ( .A(n106), .Q(n105) );
  BUF15 U295 ( .A(i_data_B[27]), .Q(n111) );
  NOR31 U296 ( .A(n495), .B(n483), .C(n416), .Q(n417) );
  BUF2 U297 ( .A(n527), .Q(n89) );
  AOI221 U298 ( .A(pre_sum_3b[5]), .B(n400), .C(pre_sum_3a[5]), .D(n399), .Q(
        n375) );
  IMUX21 U299 ( .A(n454), .B(n453), .S(n65), .Q(n455) );
  AOI211 U300 ( .A(sum_1[2]), .B(n441), .C(n164), .Q(n165) );
  IMUX21 U301 ( .A(n271), .B(n270), .S(n78), .Q(n275) );
  INV15 U302 ( .A(n102), .Q(n101) );
  OAI210 U303 ( .A(n10), .B(n35), .C(i_data_A[29]), .Q(n34) );
  NAND41 U304 ( .A(n185), .B(n184), .C(n182), .D(n181), .Q(o_data_AluRes[5])
         );
  OAI2111 U305 ( .A(n198), .B(n114), .C(n534), .D(n533), .Q(n535) );
  IMUX21 U306 ( .A(n466), .B(n465), .S(n67), .Q(n467) );
  NAND20 U307 ( .A(n526), .B(n121), .Q(n355) );
  CLKIN6 U308 ( .A(n207), .Q(n287) );
  AOI210 U309 ( .A(n201), .B(n15), .C(n202), .Q(n206) );
  AOI210 U310 ( .A(n97), .B(n477), .C(n11), .Q(n478) );
  AOI210 U311 ( .A(n99), .B(n243), .C(n10), .Q(n244) );
  INV0 U312 ( .A(n30), .Q(n243) );
  AOI210 U313 ( .A(n97), .B(n490), .C(n12), .Q(n491) );
  NAND20 U314 ( .A(n526), .B(n123), .Q(n408) );
  AOI210 U315 ( .A(n97), .B(n125), .C(n12), .Q(n453) );
  NOR20 U316 ( .A(n113), .B(n88), .Q(n525) );
  CLKIN3 U317 ( .A(n140), .Q(n147) );
  NAND42 U318 ( .A(n200), .B(n199), .C(n197), .D(n196), .Q(o_data_AluRes[7])
         );
  AOI220 U319 ( .A(N197), .B(n522), .C(N229), .D(n92), .Q(n179) );
  NAND20 U320 ( .A(n526), .B(n116), .Q(n228) );
  AOI210 U321 ( .A(n97), .B(n507), .C(n10), .Q(n508) );
  BUF15 U322 ( .A(i_data_B[18]), .Q(n110) );
  IMUX20 U323 ( .A(n252), .B(n251), .S(n107), .Q(n253) );
  BUF15 U324 ( .A(i_data_B[25]), .Q(n84) );
  OAI210 U325 ( .A(n12), .B(n254), .C(i_data_A[12]), .Q(n255) );
  BUF15 U326 ( .A(i_data_B[28]), .Q(n112) );
  BUF2 U327 ( .A(n522), .Q(n71) );
  BUF2 U328 ( .A(n542), .Q(n31) );
  INV3 U329 ( .A(n16), .Q(n32) );
  AOI2111 U330 ( .A(N233), .B(n91), .C(n206), .D(n205), .Q(n212) );
  BUF6 U331 ( .A(n532), .Q(n91) );
  BUF2 U332 ( .A(n529), .Q(n73) );
  BUF2 U333 ( .A(n532), .Q(n93) );
  AOI210 U334 ( .A(n98), .B(n123), .C(n12), .Q(n407) );
  NAND41 U335 ( .A(n218), .B(n167), .C(n166), .D(n165), .Q(o_data_AluRes[2])
         );
  AOI2111 U336 ( .A(N239), .B(n91), .C(n275), .D(n274), .Q(n279) );
  NAND41 U337 ( .A(n212), .B(n211), .C(n210), .D(n209), .Q(o_data_AluRes[8])
         );
  AOI2111 U338 ( .A(N249), .B(n91), .C(n410), .D(n409), .Q(n421) );
  AOI2111 U339 ( .A(N251), .B(n91), .C(n456), .D(n455), .Q(n462) );
  AOI221 U340 ( .A(pre_subb[10]), .B(n524), .C(pre_suba[10]), .D(n523), .Q(
        n460) );
  AOI211 U341 ( .A(N237), .B(n92), .C(n253), .Q(n261) );
  AOI221 U342 ( .A(pre_subb[12]), .B(n524), .C(n523), .D(pre_suba[12]), .Q(
        n486) );
  INV3 U343 ( .A(n108), .Q(n107) );
  AOI210 U344 ( .A(n97), .B(n127), .C(n10), .Q(n465) );
  IMUX21 U345 ( .A(n393), .B(n36), .S(n61), .Q(n394) );
  IMUX21 U346 ( .A(n94), .B(n16), .S(n84), .Q(n427) );
  NAND22 U347 ( .A(n155), .B(n154), .Q(o_data_AluRes[0]) );
  IMUX21 U348 ( .A(n216), .B(n215), .S(n74), .Q(n217) );
  AOI210 U349 ( .A(n99), .B(n214), .C(n12), .Q(n215) );
  IMUX21 U350 ( .A(n492), .B(n491), .S(n85), .Q(n493) );
  IMUX21 U351 ( .A(n283), .B(n282), .S(n80), .Q(n284) );
  IMUX20 U352 ( .A(n11), .B(n526), .S(n525), .Q(n534) );
  AOI211 U353 ( .A(N256), .B(n93), .C(n531), .Q(n533) );
  NAND41 U354 ( .A(n269), .B(n268), .C(n267), .D(n266), .Q(o_data_AluRes[13])
         );
  IMUX21 U355 ( .A(n265), .B(n264), .S(i_data_B[13]), .Q(n266) );
  NAND41 U356 ( .A(n160), .B(n159), .C(n158), .D(n157), .Q(o_data_AluRes[1])
         );
  NAND22 U357 ( .A(half_sub[1]), .B(n1), .Q(n159) );
  AOI221 U358 ( .A(N194), .B(n69), .C(N226), .D(n92), .Q(n160) );
  NAND41 U359 ( .A(n173), .B(n172), .C(n171), .D(n170), .Q(o_data_AluRes[3])
         );
  NAND22 U360 ( .A(half_sub[3]), .B(n1), .Q(n172) );
  NAND41 U361 ( .A(n179), .B(n178), .C(n177), .D(n175), .Q(o_data_AluRes[4])
         );
  NAND22 U362 ( .A(half_sub[4]), .B(n1), .Q(n178) );
  NAND22 U363 ( .A(half_sub[5]), .B(n1), .Q(n184) );
  AOI221 U364 ( .A(N198), .B(n69), .C(N230), .D(n92), .Q(n185) );
  NAND22 U365 ( .A(sum_1[7]), .B(n441), .Q(n196) );
  IMUX21 U366 ( .A(n479), .B(n478), .S(n112), .Q(n480) );
  IMUX21 U367 ( .A(n509), .B(n508), .S(n86), .Q(n510) );
  BUF12 U368 ( .A(i_data_B[15]), .Q(n79) );
  BUF2 U369 ( .A(i_data_A[31]), .Q(n88) );
  BUF2 U370 ( .A(i_data_A[31]), .Q(n87) );
  INV3 U371 ( .A(i_data_A[26]), .Q(n125) );
  INV6 U372 ( .A(i_data_B[10]), .Q(n104) );
  INV3 U373 ( .A(i_data_B[31]), .Q(n114) );
  LOGIC0 U374 ( .Q(n42) );
  LOGIC1 U375 ( .Q(n41) );
  IMUX20 U376 ( .A(n204), .B(n203), .S(n101), .Q(n205) );
  INV0 U377 ( .A(i_data_A[9]), .Q(n214) );
  INV6 U378 ( .A(n131), .Q(n141) );
  IMUX20 U379 ( .A(n245), .B(n244), .S(n105), .Q(n246) );
  AOI220 U380 ( .A(sum_1[1]), .B(n441), .C(i_data_A[1]), .D(n11), .Q(n158) );
  OAI212 U381 ( .A(n15), .B(n188), .C(n187), .Q(n189) );
  INV0 U382 ( .A(i_data_A[2]), .Q(n163) );
  OAI211 U383 ( .A(n10), .B(n378), .C(i_data_A[22]), .Q(n384) );
  OAI211 U384 ( .A(n10), .B(n340), .C(i_data_A[19]), .Q(n346) );
  OAI211 U385 ( .A(n10), .B(n365), .C(i_data_A[21]), .Q(n371) );
  INV8 U386 ( .A(n27), .Q(n293) );
  NAND21 U387 ( .A(n32), .B(n88), .Q(n198) );
  IMUX20 U388 ( .A(n94), .B(n16), .S(n112), .Q(n475) );
  IMUX20 U389 ( .A(n94), .B(n16), .S(n82), .Q(n378) );
  IMUX20 U390 ( .A(n22), .B(n16), .S(n67), .Q(n463) );
  IMUX20 U391 ( .A(n21), .B(n16), .S(n86), .Q(n504) );
  IMUX20 U392 ( .A(n22), .B(n16), .S(i_data_B[21]), .Q(n365) );
  IMUX20 U393 ( .A(n22), .B(n16), .S(n110), .Q(n328) );
  IMUX20 U394 ( .A(n22), .B(n16), .S(i_data_B[17]), .Q(n315) );
  IMUX20 U395 ( .A(n21), .B(n16), .S(n109), .Q(n295) );
  OAI211 U396 ( .A(n12), .B(n405), .C(n122), .Q(n406) );
  OAI211 U397 ( .A(n12), .B(n328), .C(i_data_A[18]), .Q(n334) );
  IMUX20 U398 ( .A(n95), .B(n32), .S(n75), .Q(n213) );
  CLKIN6 U399 ( .A(n53), .Q(n55) );
  IMUX20 U400 ( .A(n94), .B(n16), .S(n56), .Q(n353) );
  INV0 U401 ( .A(n103), .Q(n29) );
  IMUX20 U402 ( .A(n21), .B(n16), .S(n55), .Q(n340) );
  OAI211 U403 ( .A(n11), .B(n391), .C(i_data_A[23]), .Q(n396) );
  IMUX20 U404 ( .A(n94), .B(n16), .S(i_data_B[23]), .Q(n391) );
  CLKIN0 U405 ( .A(i_data_B[6]), .Q(n385) );
  NAND42 U406 ( .A(n404), .B(n403), .C(n402), .D(n401), .Q(o_data_AluRes[23])
         );
  IMUX30 U407 ( .A(n526), .B(n96), .C(n168), .S0(n46), .S1(n2), .Q(n170) );
  NAND21 U408 ( .A(pre_sum_2b[8]), .B(n52), .Q(n423) );
  INV1 U409 ( .A(n136), .Q(n33) );
  OAI211 U410 ( .A(n72), .B(n29), .C(n452), .Q(n456) );
  AOI221 U411 ( .A(pre_sum_2b[7]), .B(n287), .C(N208), .D(n522), .Q(n289) );
  IMUX20 U412 ( .A(n21), .B(n16), .S(n105), .Q(n238) );
  IMUX20 U413 ( .A(n97), .B(n32), .S(n78), .Q(n273) );
  IMUX20 U414 ( .A(n97), .B(n32), .S(i_data_B[13]), .Q(n262) );
  IMUX30 U415 ( .A(n526), .B(n95), .C(n156), .S0(i_data_A[1]), .S1(i_data_B[1]), .Q(n157) );
  OAI210 U416 ( .A(i_data_A[13]), .B(n94), .C(n68), .Q(n264) );
  NOR20 U417 ( .A(i_data_A[13]), .B(n139), .Q(n265) );
  NAND30 U418 ( .A(n27), .B(n136), .C(n135), .Q(n137) );
  NAND20 U419 ( .A(n46), .B(n31), .Q(n190) );
  NAND20 U420 ( .A(i_data_A[0]), .B(n542), .Q(n428) );
  NAND20 U421 ( .A(i_data_A[2]), .B(n31), .Q(n221) );
  NAND20 U422 ( .A(i_data_A[1]), .B(n31), .Q(n333) );
  NAND20 U423 ( .A(i_data_A[5]), .B(n31), .Q(n176) );
  NAND20 U424 ( .A(i_data_A[4]), .B(n32), .Q(n183) );
  OAI211 U425 ( .A(n11), .B(n475), .C(i_data_A[28]), .Q(n476) );
  OAI211 U426 ( .A(n12), .B(n463), .C(n126), .Q(n464) );
  OAI211 U427 ( .A(n11), .B(n504), .C(i_data_A[30]), .Q(n505) );
  OAI211 U428 ( .A(n10), .B(n315), .C(i_data_A[17]), .Q(n321) );
  AOI211 U429 ( .A(n273), .B(n15), .C(n272), .Q(n274) );
  NAND21 U430 ( .A(n262), .B(n15), .Q(n263) );
  OAI2110 U431 ( .A(i_data_A[1]), .B(n39), .C(n13), .D(n333), .Q(n156) );
  IMUX21 U432 ( .A(n21), .B(n16), .S(n85), .Q(n35) );
  OAI2111 U433 ( .A(n443), .B(n442), .C(pre_sum_4a[1]), .D(n441), .Q(n444) );
  OAI221 U434 ( .A(n443), .B(n440), .C(n439), .D(n438), .Q(n445) );
  INV2 U435 ( .A(i_data_B[4]), .Q(n359) );
  CLKIN0 U436 ( .A(i_data_A[6]), .Q(n188) );
  NAND20 U437 ( .A(i_data_A[6]), .B(n542), .Q(n169) );
  OAI2110 U438 ( .A(i_data_A[5]), .B(n22), .C(n13), .D(n176), .Q(n180) );
  IMUX30 U439 ( .A(n526), .B(n96), .C(n180), .S0(i_data_A[5]), .S1(n7), .Q(
        n181) );
  AOI221 U440 ( .A(N232), .B(n92), .C(i_data_A[7]), .D(n10), .Q(n200) );
  NOR31 U441 ( .A(n495), .B(n483), .C(n469), .Q(n470) );
  NOR31 U442 ( .A(n495), .B(n483), .C(n457), .Q(n458) );
  NOR31 U443 ( .A(n495), .B(n483), .C(n482), .Q(n484) );
  CLKIN0 U444 ( .A(i_data_B[2]), .Q(n543) );
  INV3 U445 ( .A(pre_sum_4b[4]), .Q(n482) );
  NOR31 U446 ( .A(n436), .B(n437), .C(n439), .Q(n446) );
  IMUX21 U447 ( .A(n21), .B(n16), .S(n107), .Q(n254) );
  OAI2110 U448 ( .A(i_data_A[2]), .B(n22), .C(n15), .D(n221), .Q(n220) );
  OAI220 U449 ( .A(n22), .B(n163), .C(i_data_A[2]), .D(n139), .Q(n219) );
  OAI212 U450 ( .A(n39), .B(i_data_A[25]), .C(n68), .Q(n38) );
  IMUX20 U451 ( .A(n97), .B(n32), .S(n101), .Q(n201) );
  NAND33 U452 ( .A(n339), .B(n336), .C(n43), .Q(o_data_AluRes[18]) );
  NAND21 U453 ( .A(pre_suba[2]), .B(n523), .Q(n336) );
  IMUX22 U454 ( .A(n381), .B(n380), .S(n82), .Q(n382) );
  AOI211 U455 ( .A(pre_sum_2b[4]), .B(n287), .C(n257), .Q(n259) );
  AOI220 U456 ( .A(pre_sum_2a[1]), .B(n286), .C(pre_sum_2b[1]), .D(n287), .Q(
        n225) );
  AOI220 U457 ( .A(pre_sum_2b[5]), .B(n287), .C(N238), .D(n91), .Q(n268) );
  AOI220 U458 ( .A(pre_sum_2b[0]), .B(n287), .C(pre_sum_2a[0]), .D(n286), .Q(
        n211) );
  NAND30 U459 ( .A(n37), .B(n294), .C(n293), .Q(n151) );
  NAND21 U460 ( .A(n37), .B(n141), .Q(n150) );
  IMUX20 U461 ( .A(n228), .B(n227), .S(n103), .Q(n229) );
  IMUX20 U462 ( .A(n22), .B(n16), .S(n103), .Q(n230) );
  INV2 U463 ( .A(i_data_A[15]), .Q(n281) );
  IMUX21 U464 ( .A(n408), .B(n407), .S(n63), .Q(n409) );
  NAND22 U465 ( .A(n44), .B(n74), .Q(n45) );
  NAND22 U466 ( .A(n45), .B(n429), .Q(n430) );
  INV3 U467 ( .A(n72), .Q(n44) );
  BUF6 U468 ( .A(n529), .Q(n72) );
  OAI212 U469 ( .A(n11), .B(n427), .C(i_data_A[25]), .Q(n429) );
  INV2 U470 ( .A(i_data_A[29]), .Q(n490) );
  IMUX21 U471 ( .A(n22), .B(n16), .S(n62), .Q(n405) );
  IMUX21 U472 ( .A(n22), .B(n16), .S(n64), .Q(n451) );
  CLKIN0 U473 ( .A(i_data_A[22]), .Q(n379) );
  NAND41 U474 ( .A(n352), .B(n351), .C(n350), .D(n349), .Q(o_data_AluRes[19])
         );
  NAND41 U475 ( .A(n377), .B(n376), .C(n375), .D(n374), .Q(o_data_AluRes[21])
         );
  INV2 U476 ( .A(i_data_A[0]), .Q(n134) );
  INV2 U477 ( .A(i_data_A[21]), .Q(n366) );
  INV2 U478 ( .A(i_data_A[12]), .Q(n250) );
  INV2 U479 ( .A(i_data_A[23]), .Q(n392) );
  AOI311 U480 ( .A(pre_sum_4a[0]), .B(n521), .C(n25), .D(n417), .Q(n418) );
  AOI220 U481 ( .A(sum_1[4]), .B(n441), .C(i_data_A[4]), .D(n12), .Q(n177) );
  AOI311 U482 ( .A(pre_sum_4a[2]), .B(n521), .C(n25), .D(n458), .Q(n459) );
  INV3 U483 ( .A(pre_sum_4a[3]), .Q(n47) );
  CLKIN0 U484 ( .A(i_data_A[30]), .Q(n507) );
  OAI220 U485 ( .A(n152), .B(n151), .C(n293), .D(n150), .Q(n153) );
  NAND31 U486 ( .A(n294), .B(n293), .C(n292), .Q(n529) );
  NAND31 U487 ( .A(n141), .B(n293), .C(n292), .Q(n132) );
  BUF2 U488 ( .A(i_data_B[0]), .Q(n50) );
  OAI220 U489 ( .A(pre_sum_3b[8]), .B(n423), .C(pre_sum_3a[8]), .D(n442), .Q(
        n434) );
  INV2 U490 ( .A(i_data_A[19]), .Q(n341) );
  INV2 U491 ( .A(i_data_A[25]), .Q(n424) );
  BUF15 U492 ( .A(i_data_B[22]), .Q(n82) );
  NAND22 U493 ( .A(sum_1[0]), .B(n441), .Q(n133) );
  OAI212 U494 ( .A(n14), .B(n134), .C(n133), .Q(n148) );
  XNR21 U495 ( .A(n113), .B(n88), .Q(n530) );
  CLKIN3 U496 ( .A(n88), .Q(n145) );
  CLKIN3 U497 ( .A(n530), .Q(n152) );
  NAND22 U498 ( .A(N227), .B(n93), .Q(n167) );
  NAND22 U499 ( .A(half_sub[2]), .B(n1), .Q(n162) );
  NAND22 U500 ( .A(N199), .B(n522), .Q(n193) );
  NAND22 U501 ( .A(half_sub[6]), .B(n1), .Q(n192) );
  CLKIN3 U502 ( .A(i_data_A[8]), .Q(n202) );
  NAND22 U503 ( .A(n526), .B(n202), .Q(n204) );
  NAND22 U504 ( .A(n441), .B(n52), .Q(n207) );
  NAND22 U505 ( .A(half_sub[8]), .B(n1), .Q(n209) );
  NAND22 U506 ( .A(n526), .B(n214), .Q(n216) );
  NAND22 U507 ( .A(half_sub[9]), .B(n1), .Q(n223) );
  NAND22 U508 ( .A(N235), .B(n93), .Q(n232) );
  NAND22 U509 ( .A(pre_sum_2a[3]), .B(n286), .Q(n242) );
  NAND22 U510 ( .A(n526), .B(n243), .Q(n245) );
  NAND22 U511 ( .A(half_sub[11]), .B(n1), .Q(n248) );
  NAND22 U512 ( .A(n249), .B(n248), .Q(o_data_AluRes[11]) );
  NAND22 U513 ( .A(n526), .B(n250), .Q(n252) );
  NAND22 U514 ( .A(pre_sum_2a[4]), .B(n286), .Q(n256) );
  NAND22 U515 ( .A(n256), .B(n255), .Q(n257) );
  CLKIN3 U516 ( .A(i_data_A[14]), .Q(n272) );
  NAND22 U517 ( .A(n526), .B(n272), .Q(n271) );
  NAND22 U518 ( .A(N207), .B(n522), .Q(n278) );
  NAND22 U519 ( .A(half_sub[14]), .B(n1), .Q(n276) );
  NAND42 U520 ( .A(n279), .B(n278), .C(n277), .D(n276), .Q(o_data_AluRes[14])
         );
  NAND22 U521 ( .A(n526), .B(n281), .Q(n283) );
  NAND22 U522 ( .A(pre_sum_2a[7]), .B(n286), .Q(n290) );
  NAND22 U523 ( .A(half_sub[15]), .B(n1), .Q(n288) );
  CLKIN3 U524 ( .A(n50), .Q(n301) );
  NAND22 U525 ( .A(n526), .B(n118), .Q(n297) );
  CLKIN3 U526 ( .A(i_data_A[17]), .Q(n316) );
  NAND22 U527 ( .A(n526), .B(n316), .Q(n318) );
  NAND22 U528 ( .A(n526), .B(n119), .Q(n330) );
  AOI212 U529 ( .A(n98), .B(n119), .C(n10), .Q(n329) );
  OAI2112 U530 ( .A(n543), .B(n73), .C(n334), .D(n332), .Q(n335) );
  NAND22 U531 ( .A(n526), .B(n341), .Q(n343) );
  NAND22 U532 ( .A(n526), .B(n366), .Q(n368) );
  NAND22 U533 ( .A(n526), .B(n379), .Q(n381) );
  CLKIN3 U534 ( .A(i_data_B[7]), .Q(n397) );
  NAND22 U535 ( .A(n526), .B(n392), .Q(n393) );
  OAI212 U536 ( .A(n72), .B(n102), .C(n406), .Q(n410) );
  NAND22 U537 ( .A(N217), .B(n522), .Q(n420) );
  OAI222 U538 ( .A(n436), .B(n437), .C(n51), .D(n422), .Q(n412) );
  OAI212 U539 ( .A(n443), .B(n412), .C(n441), .Q(n515) );
  AOI312 U540 ( .A(n437), .B(n443), .C(n52), .D(n413), .Q(n414) );
  OAI222 U541 ( .A(n52), .B(n422), .C(n436), .D(n437), .Q(n415) );
  CLKIN3 U542 ( .A(pre_sum_4b[0]), .Q(n416) );
  NAND42 U543 ( .A(n421), .B(n420), .C(n419), .D(n418), .Q(o_data_AluRes[24])
         );
  NAND22 U544 ( .A(n526), .B(n424), .Q(n426) );
  OAI212 U545 ( .A(n12), .B(n451), .C(n124), .Q(n452) );
  NAND22 U546 ( .A(n526), .B(n125), .Q(n454) );
  NAND22 U547 ( .A(N219), .B(n522), .Q(n461) );
  CLKIN3 U548 ( .A(pre_sum_4b[2]), .Q(n457) );
  NAND42 U549 ( .A(n462), .B(n461), .C(n460), .D(n459), .Q(o_data_AluRes[26])
         );
  OAI212 U550 ( .A(n72), .B(n106), .C(n464), .Q(n468) );
  NAND22 U551 ( .A(n526), .B(n127), .Q(n466) );
  AOI2112 U552 ( .A(N252), .B(n91), .C(n468), .D(n467), .Q(n474) );
  NAND22 U553 ( .A(N220), .B(n522), .Q(n473) );
  OAI212 U554 ( .A(n72), .B(n108), .C(n476), .Q(n481) );
  CLKIN3 U555 ( .A(i_data_A[28]), .Q(n477) );
  NAND22 U556 ( .A(n526), .B(n477), .Q(n479) );
  NAND22 U557 ( .A(N221), .B(n522), .Q(n487) );
  NAND42 U558 ( .A(n488), .B(n487), .C(n486), .D(n485), .Q(o_data_AluRes[28])
         );
  OAI212 U559 ( .A(n72), .B(n489), .C(n34), .Q(n494) );
  NAND22 U560 ( .A(n526), .B(n490), .Q(n492) );
  AOI2112 U561 ( .A(N254), .B(n91), .C(n494), .D(n493), .Q(n502) );
  NAND22 U562 ( .A(N222), .B(n522), .Q(n501) );
  NAND22 U563 ( .A(pre_sum_4a[5]), .B(n521), .Q(n497) );
  CLKIN3 U564 ( .A(pre_sum_4b[5]), .Q(n496) );
  OAI222 U565 ( .A(n26), .B(n497), .C(n512), .D(n496), .Q(n498) );
  AOI212 U566 ( .A(pre_subb[13]), .B(n524), .C(n498), .Q(n499) );
  NAND42 U567 ( .A(n502), .B(n501), .C(n500), .D(n499), .Q(o_data_AluRes[29])
         );
  CLKIN3 U568 ( .A(n78), .Q(n506) );
  OAI212 U569 ( .A(n72), .B(n506), .C(n505), .Q(n511) );
  NAND22 U570 ( .A(n526), .B(n507), .Q(n509) );
  AOI2112 U571 ( .A(N255), .B(n91), .C(n511), .D(n510), .Q(n520) );
  NAND22 U572 ( .A(pre_sum_4a[6]), .B(n521), .Q(n514) );
  CLKIN3 U573 ( .A(pre_sum_4b[6]), .Q(n513) );
  OAI222 U574 ( .A(n26), .B(n514), .C(n512), .D(n513), .Q(n516) );
  AOI212 U575 ( .A(pre_subb[14]), .B(n524), .C(n516), .Q(n517) );
  NAND22 U576 ( .A(N224), .B(n522), .Q(n540) );
  CLKIN3 U577 ( .A(n80), .Q(n528) );
  OAI222 U578 ( .A(n22), .B(n530), .C(n72), .D(n528), .Q(n531) );
  NAND42 U579 ( .A(n541), .B(n540), .C(n538), .D(n539), .Q(o_data_AluRes[31])
         );
endmodule


module E_alu_control ( o_con_AluCtrl, i_con_AluOp, i_con_FuncCode );
  output [3:0] o_con_AluCtrl;
  input [5:0] i_con_AluOp;
  input [5:0] i_con_FuncCode;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n54, n55, n56, n57, n58;

  OAI2112 U3 ( .A(n15), .B(n22), .C(n23), .D(n24), .Q(o_con_AluCtrl[3]) );
  OAI2112 U7 ( .A(n57), .B(n32), .C(n16), .D(n55), .Q(n26) );
  NOR42 U20 ( .A(n15), .B(n43), .C(n44), .D(n9), .Q(n46) );
  NOR42 U27 ( .A(n25), .B(n35), .C(n31), .D(n51), .Q(n50) );
  NOR24 U35 ( .A(n19), .B(i_con_FuncCode[0]), .Q(n25) );
  NOR42 U36 ( .A(n20), .B(n56), .C(n57), .D(i_con_FuncCode[2]), .Q(n53) );
  AOI211 U4 ( .A(n13), .B(i_con_AluOp[0]), .C(n46), .Q(n38) );
  OAI2111 U5 ( .A(n27), .B(n28), .C(n29), .D(n7), .Q(o_con_AluCtrl[2]) );
  NAND22 U6 ( .A(n38), .B(n45), .Q(n30) );
  INV3 U8 ( .A(n57), .Q(n1) );
  INV6 U9 ( .A(i_con_FuncCode[1]), .Q(n57) );
  OAI2112 U10 ( .A(n41), .B(n28), .C(n24), .D(n42), .Q(o_con_AluCtrl[0]) );
  INV3 U11 ( .A(i_con_AluOp[2]), .Q(n12) );
  CLKIN6 U12 ( .A(i_con_FuncCode[5]), .Q(n20) );
  CLKIN6 U13 ( .A(i_con_FuncCode[3]), .Q(n56) );
  NAND41 U14 ( .A(n36), .B(n29), .C(n11), .D(n37), .Q(o_con_AluCtrl[1]) );
  NOR21 U15 ( .A(n13), .B(n6), .Q(n37) );
  BUF2 U16 ( .A(i_con_FuncCode[5]), .Q(n2) );
  INV3 U17 ( .A(n56), .Q(n3) );
  NOR31 U18 ( .A(n21), .B(n31), .C(n17), .Q(n4) );
  NOR21 U19 ( .A(n5), .B(n26), .Q(n27) );
  INV3 U21 ( .A(n4), .Q(n5) );
  INV0 U22 ( .A(n33), .Q(n21) );
  NAND21 U23 ( .A(n44), .B(i_con_AluOp[0]), .Q(n29) );
  NOR32 U24 ( .A(i_con_FuncCode[3]), .B(i_con_FuncCode[5]), .C(
        i_con_FuncCode[2]), .Q(n47) );
  OAI210 U25 ( .A(n25), .B(n26), .C(n14), .Q(n23) );
  NAND32 U26 ( .A(n58), .B(n57), .C(n47), .Q(n49) );
  NAND33 U28 ( .A(n49), .B(n32), .C(n33), .Q(n51) );
  NOR32 U29 ( .A(n3), .B(i_con_FuncCode[2]), .C(n20), .Q(n35) );
  CLKIN1 U30 ( .A(n30), .Q(n7) );
  NAND22 U31 ( .A(n47), .B(i_con_FuncCode[1]), .Q(n33) );
  NOR41 U32 ( .A(n10), .B(n12), .C(i_con_AluOp[3]), .D(i_con_AluOp[4]), .Q(n44) );
  AOI311 U33 ( .A(n9), .B(n12), .C(i_con_AluOp[0]), .D(n30), .Q(n24) );
  CLKIN3 U34 ( .A(i_con_AluOp[5]), .Q(n10) );
  CLKIN1 U37 ( .A(n29), .Q(n8) );
  AOI310 U38 ( .A(i_con_AluOp[3]), .B(i_con_AluOp[0]), .C(n43), .D(n8), .Q(n42) );
  CLKIN1 U39 ( .A(n32), .Q(n54) );
  NAND21 U40 ( .A(i_con_AluOp[1]), .B(n15), .Q(n28) );
  NOR30 U41 ( .A(i_con_AluOp[2]), .B(i_con_AluOp[3]), .C(n15), .Q(n39) );
  CLKIN3 U42 ( .A(i_con_FuncCode[0]), .Q(n58) );
  NAND40 U43 ( .A(n43), .B(i_con_AluOp[2]), .C(i_con_AluOp[3]), .D(
        i_con_AluOp[0]), .Q(n45) );
  INV2 U44 ( .A(n34), .Q(n17) );
  CLKIN3 U45 ( .A(i_con_AluOp[1]), .Q(n13) );
  INV3 U46 ( .A(n39), .Q(n11) );
  INV3 U47 ( .A(n22), .Q(n9) );
  INV3 U48 ( .A(n38), .Q(n6) );
  INV3 U49 ( .A(n28), .Q(n14) );
  NAND31 U50 ( .A(i_con_AluOp[3]), .B(n10), .C(i_con_AluOp[4]), .Q(n22) );
  NOR21 U51 ( .A(i_con_AluOp[5]), .B(i_con_AluOp[4]), .Q(n43) );
  INV3 U52 ( .A(i_con_AluOp[0]), .Q(n15) );
  INV3 U53 ( .A(i_con_FuncCode[4]), .Q(n55) );
  NAND20 U54 ( .A(i_con_FuncCode[1]), .B(n35), .Q(n34) );
  INV3 U55 ( .A(n31), .Q(n18) );
  OAI212 U56 ( .A(n35), .B(n40), .C(n14), .Q(n36) );
  NAND43 U57 ( .A(n49), .B(n18), .C(n16), .D(n55), .Q(n40) );
  NAND32 U58 ( .A(n2), .B(n56), .C(i_con_FuncCode[2]), .Q(n32) );
  AOI2111 U59 ( .A(n47), .B(i_con_FuncCode[0]), .C(n48), .D(n40), .Q(n41) );
  NOR23 U60 ( .A(n58), .B(n19), .Q(n31) );
  INV6 U61 ( .A(n50), .Q(n16) );
  OAI310 U62 ( .A(n32), .B(n1), .C(n58), .D(n52), .Q(n48) );
  AOI310 U63 ( .A(n1), .B(n58), .C(n54), .D(n25), .Q(n52) );
  CLKIN6 U64 ( .A(n53), .Q(n19) );
endmodule


module E_famux5 ( i_data_rs, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fa, o_data_alusra );
  input [31:0] i_data_rs;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fa;
  output [31:0] o_data_alusra;
  wire   n134, n135, n136, n137, n1, n2, n3, n4, n6, n9, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133;

  AOI221 U1 ( .A(i_data_lwM[22]), .B(n15), .C(i_data_alures[22]), .D(n21), .Q(
        n100) );
  NAND33 U2 ( .A(n45), .B(n44), .C(n43), .Q(o_data_alusra[4]) );
  NAND32 U3 ( .A(i_con_fa[1]), .B(n32), .C(n31), .Q(n26) );
  CLKIN12 U4 ( .A(i_con_fa[0]), .Q(n31) );
  CLKIN6 U5 ( .A(n11), .Q(n13) );
  INV6 U6 ( .A(n128), .Q(n11) );
  NAND34 U7 ( .A(n65), .B(n64), .C(n63), .Q(o_data_alusra[10]) );
  INV12 U8 ( .A(n24), .Q(n12) );
  INV8 U9 ( .A(i_con_fa[1]), .Q(n24) );
  BUF12 U10 ( .A(n129), .Q(n21) );
  CLKIN12 U11 ( .A(n27), .Q(n121) );
  AOI221 U12 ( .A(i_data_writeres[4]), .B(n13), .C(i_data_lwW[4]), .D(n4), .Q(
        n45) );
  AOI221 U13 ( .A(i_data_lwM[30]), .B(n15), .C(i_data_alures[30]), .D(n21), 
        .Q(n126) );
  NAND33 U14 ( .A(n95), .B(n94), .C(n93), .Q(o_data_alusra[20]) );
  NAND22 U15 ( .A(i_data_rs[10]), .B(n121), .Q(n63) );
  NAND22 U16 ( .A(i_data_rs[29]), .B(n121), .Q(n122) );
  CLKIN12 U17 ( .A(n33), .Q(n46) );
  AOI221 U18 ( .A(i_data_writeres[18]), .B(n1), .C(i_data_lwW[18]), .D(n4), 
        .Q(n89) );
  AOI221 U19 ( .A(i_data_rs[1]), .B(n111), .C(i_data_writeres[1]), .D(n13), 
        .Q(n36) );
  NAND22 U20 ( .A(i_data_rs[4]), .B(n111), .Q(n43) );
  CLKIN6 U21 ( .A(n19), .Q(n111) );
  NAND34 U22 ( .A(n42), .B(n41), .C(n40), .Q(o_data_alusra[3]) );
  AOI221 U23 ( .A(i_data_lwM[3]), .B(n15), .C(i_data_alures[3]), .D(n21), .Q(
        n41) );
  INV15 U24 ( .A(n25), .Q(n15) );
  AOI221 U25 ( .A(i_data_rs[28]), .B(n111), .C(i_data_writeres[28]), .D(n13), 
        .Q(n120) );
  NAND22 U26 ( .A(i_data_rs[20]), .B(n111), .Q(n93) );
  AOI221 U27 ( .A(i_data_writeres[8]), .B(n13), .C(i_data_lwW[8]), .D(n17), 
        .Q(n59) );
  AOI221 U28 ( .A(i_data_lwM[1]), .B(n15), .C(i_data_lwW[1]), .D(n4), .Q(n34)
         );
  BUF8 U29 ( .A(n20), .Q(n4) );
  INV12 U30 ( .A(n6), .Q(o_data_alusra[22]) );
  INV6 U31 ( .A(n134), .Q(n6) );
  AOI221 U32 ( .A(i_data_lwM[17]), .B(n15), .C(i_data_alures[17]), .D(n22), 
        .Q(n85) );
  AOI221 U33 ( .A(i_data_lwM[26]), .B(n15), .C(i_data_alures[26]), .D(n21), 
        .Q(n113) );
  INV3 U34 ( .A(n23), .Q(n128) );
  CLKIN12 U35 ( .A(n9), .Q(o_data_alusra[17]) );
  AOI221 U36 ( .A(i_data_writeres[2]), .B(n1), .C(i_data_lwW[2]), .D(n4), .Q(
        n39) );
  NAND22 U37 ( .A(i_data_rs[2]), .B(n111), .Q(n37) );
  AOI221 U38 ( .A(i_data_writeres[19]), .B(n1), .C(i_data_lwW[19]), .D(n18), 
        .Q(n92) );
  INV3 U39 ( .A(n16), .Q(n17) );
  BUF8 U40 ( .A(n129), .Q(n22) );
  NAND22 U41 ( .A(i_data_rs[21]), .B(n130), .Q(n96) );
  INV8 U42 ( .A(n47), .Q(n130) );
  BUF12 U43 ( .A(n137), .Q(o_data_alusra[0]) );
  AOI221 U44 ( .A(i_data_lwM[28]), .B(n15), .C(i_data_lwW[28]), .D(n17), .Q(
        n118) );
  INV3 U45 ( .A(n23), .Q(n1) );
  INV3 U46 ( .A(n11), .Q(n3) );
  NAND32 U47 ( .A(i_con_fa[2]), .B(n31), .C(n24), .Q(n25) );
  INV3 U48 ( .A(n20), .Q(n16) );
  INV6 U49 ( .A(i_con_fa[2]), .Q(n32) );
  NAND26 U50 ( .A(n32), .B(n31), .Q(n33) );
  NAND33 U51 ( .A(n124), .B(n123), .C(n122), .Q(o_data_alusra[29]) );
  NAND22 U52 ( .A(i_data_rs[18]), .B(n111), .Q(n87) );
  NAND22 U53 ( .A(i_data_rs[6]), .B(n121), .Q(n51) );
  AOI221 U54 ( .A(i_data_lwM[19]), .B(n15), .C(i_data_alures[19]), .D(n129), 
        .Q(n91) );
  NOR32 U55 ( .A(n32), .B(n31), .C(i_con_fa[1]), .Q(n20) );
  INV6 U56 ( .A(n26), .Q(n129) );
  AOI221 U57 ( .A(i_data_lwM[20]), .B(n15), .C(i_data_alures[20]), .D(n22), 
        .Q(n94) );
  NAND33 U58 ( .A(i_con_fa[0]), .B(n32), .C(n24), .Q(n23) );
  AOI221 U59 ( .A(n14), .B(i_data_rs[27]), .C(i_data_writeres[27]), .D(n3), 
        .Q(n117) );
  AOI221 U60 ( .A(i_data_lwM[12]), .B(n15), .C(i_data_alures[12]), .D(n22), 
        .Q(n70) );
  AOI221 U61 ( .A(i_data_writeres[16]), .B(n3), .C(i_data_lwW[16]), .D(n4), 
        .Q(n83) );
  INV2 U62 ( .A(n16), .Q(n18) );
  NAND33 U63 ( .A(n30), .B(n29), .C(n28), .Q(n137) );
  NAND22 U64 ( .A(i_data_rs[0]), .B(n121), .Q(n28) );
  AOI221 U65 ( .A(i_data_lwM[0]), .B(n15), .C(i_data_alures[0]), .D(n22), .Q(
        n29) );
  AOI221 U66 ( .A(i_data_rs[13]), .B(n121), .C(i_data_writeres[13]), .D(n13), 
        .Q(n74) );
  AOI221 U67 ( .A(i_data_writeres[23]), .B(n1), .C(i_data_lwW[23]), .D(n4), 
        .Q(n104) );
  NAND33 U68 ( .A(n92), .B(n91), .C(n90), .Q(o_data_alusra[19]) );
  INV3 U69 ( .A(n11), .Q(n2) );
  AOI221 U70 ( .A(i_data_lwM[23]), .B(n15), .C(i_data_alures[23]), .D(n21), 
        .Q(n103) );
  XNR22 U71 ( .A(n33), .B(n12), .Q(n14) );
  NAND32 U72 ( .A(n127), .B(n126), .C(n125), .Q(o_data_alusra[30]) );
  AOI221 U73 ( .A(i_data_lwM[13]), .B(n15), .C(i_data_lwW[13]), .D(n17), .Q(
        n72) );
  NAND21 U74 ( .A(i_data_rs[23]), .B(n130), .Q(n102) );
  AOI221 U75 ( .A(i_data_lwM[5]), .B(n15), .C(i_data_alures[5]), .D(n22), .Q(
        n49) );
  NAND33 U76 ( .A(n71), .B(n70), .C(n69), .Q(o_data_alusra[12]) );
  AOI221 U77 ( .A(i_data_lwM[21]), .B(n15), .C(i_data_alures[21]), .D(n21), 
        .Q(n97) );
  NAND33 U78 ( .A(n86), .B(n85), .C(n84), .Q(n135) );
  BUF15 U79 ( .A(n136), .Q(o_data_alusra[14]) );
  NAND33 U80 ( .A(n77), .B(n76), .C(n75), .Q(n136) );
  NAND22 U81 ( .A(i_data_rs[12]), .B(n130), .Q(n69) );
  XOR22 U82 ( .A(n33), .B(n12), .Q(n19) );
  NAND21 U83 ( .A(n14), .B(i_data_rs[19]), .Q(n90) );
  NAND33 U84 ( .A(n104), .B(n103), .C(n102), .Q(o_data_alusra[23]) );
  CLKIN3 U85 ( .A(n135), .Q(n9) );
  NAND22 U86 ( .A(i_data_rs[22]), .B(n130), .Q(n99) );
  NAND33 U87 ( .A(n101), .B(n100), .C(n99), .Q(n134) );
  AOI221 U88 ( .A(i_data_lwM[8]), .B(n15), .C(i_data_alures[8]), .D(n21), .Q(
        n58) );
  NAND22 U89 ( .A(i_data_rs[3]), .B(n121), .Q(n40) );
  XNR22 U90 ( .A(n12), .B(n46), .Q(n47) );
  AOI221 U91 ( .A(i_data_writeres[3]), .B(n2), .C(i_data_lwW[3]), .D(n17), .Q(
        n42) );
  NAND21 U92 ( .A(i_data_rs[31]), .B(n130), .Q(n131) );
  NAND33 U93 ( .A(n98), .B(n97), .C(n96), .Q(o_data_alusra[21]) );
  NAND22 U94 ( .A(i_data_rs[9]), .B(n121), .Q(n60) );
  AOI221 U95 ( .A(i_data_lwM[9]), .B(n15), .C(i_data_alures[9]), .D(n22), .Q(
        n61) );
  AOI221 U96 ( .A(i_data_lwM[11]), .B(n15), .C(i_data_alures[11]), .D(n21), 
        .Q(n67) );
  NAND33 U97 ( .A(n80), .B(n79), .C(n78), .Q(o_data_alusra[15]) );
  NAND21 U98 ( .A(i_data_alures[25]), .B(n21), .Q(n109) );
  NAND21 U99 ( .A(i_data_alures[13]), .B(n21), .Q(n73) );
  AOI221 U100 ( .A(i_data_lwM[7]), .B(n15), .C(i_data_alures[7]), .D(n22), .Q(
        n55) );
  AOI221 U101 ( .A(i_data_lwM[10]), .B(n15), .C(i_data_alures[10]), .D(n22), 
        .Q(n64) );
  AOI221 U102 ( .A(i_data_lwM[14]), .B(n15), .C(i_data_alures[14]), .D(n22), 
        .Q(n76) );
  NAND33 U103 ( .A(n68), .B(n67), .C(n66), .Q(o_data_alusra[11]) );
  NAND33 U104 ( .A(n83), .B(n82), .C(n81), .Q(o_data_alusra[16]) );
  AOI221 U105 ( .A(i_data_writeres[15]), .B(n2), .C(i_data_lwW[15]), .D(n4), 
        .Q(n80) );
  NAND33 U106 ( .A(n110), .B(n109), .C(n108), .Q(o_data_alusra[25]) );
  NAND33 U107 ( .A(n59), .B(n58), .C(n57), .Q(o_data_alusra[8]) );
  AOI221 U108 ( .A(i_data_lwM[6]), .B(n15), .C(i_data_alures[6]), .D(n21), .Q(
        n52) );
  AOI221 U109 ( .A(i_data_lwM[16]), .B(n15), .C(i_data_alures[16]), .D(n21), 
        .Q(n82) );
  NAND22 U110 ( .A(i_data_rs[16]), .B(n130), .Q(n81) );
  NAND21 U111 ( .A(i_data_rs[15]), .B(n121), .Q(n78) );
  NAND21 U112 ( .A(i_data_alures[28]), .B(n21), .Q(n119) );
  NAND21 U113 ( .A(i_data_alures[27]), .B(n21), .Q(n116) );
  AOI221 U114 ( .A(i_data_lwM[2]), .B(n15), .C(i_data_alures[2]), .D(n22), .Q(
        n38) );
  AOI221 U115 ( .A(i_data_lwM[15]), .B(n15), .C(i_data_alures[15]), .D(n21), 
        .Q(n79) );
  AOI221 U116 ( .A(i_data_lwM[4]), .B(n15), .C(i_data_alures[4]), .D(n22), .Q(
        n44) );
  AOI221 U117 ( .A(i_data_lwM[29]), .B(n15), .C(i_data_alures[29]), .D(n22), 
        .Q(n123) );
  NAND21 U118 ( .A(i_data_rs[26]), .B(n111), .Q(n112) );
  AOI220 U119 ( .A(i_data_rs[25]), .B(n111), .C(i_data_writeres[25]), .D(n1), 
        .Q(n110) );
  NAND34 U120 ( .A(n62), .B(n61), .C(n60), .Q(o_data_alusra[9]) );
  NAND34 U121 ( .A(n74), .B(n73), .C(n72), .Q(o_data_alusra[13]) );
  NAND33 U122 ( .A(n120), .B(n119), .C(n118), .Q(o_data_alusra[28]) );
  NAND34 U123 ( .A(n39), .B(n38), .C(n37), .Q(o_data_alusra[2]) );
  AOI221 U124 ( .A(i_data_writeres[29]), .B(n13), .C(i_data_lwW[29]), .D(n4), 
        .Q(n124) );
  AOI221 U125 ( .A(i_data_writeres[21]), .B(n3), .C(i_data_lwW[21]), .D(n4), 
        .Q(n98) );
  AOI221 U126 ( .A(i_data_writeres[14]), .B(n13), .C(i_data_lwW[14]), .D(n18), 
        .Q(n77) );
  AOI221 U127 ( .A(i_data_writeres[17]), .B(n1), .C(i_data_lwW[17]), .D(n17), 
        .Q(n86) );
  AOI221 U128 ( .A(i_data_writeres[30]), .B(n2), .C(i_data_lwW[30]), .D(n4), 
        .Q(n127) );
  AOI220 U129 ( .A(i_data_writeres[31]), .B(n2), .C(i_data_lwW[31]), .D(n4), 
        .Q(n133) );
  AOI221 U130 ( .A(i_data_writeres[11]), .B(n13), .C(i_data_lwW[11]), .D(n4), 
        .Q(n68) );
  AOI221 U131 ( .A(i_data_writeres[22]), .B(n3), .C(i_data_lwW[22]), .D(n4), 
        .Q(n101) );
  AOI221 U132 ( .A(i_data_writeres[24]), .B(n1), .C(i_data_lwW[24]), .D(n4), 
        .Q(n107) );
  AOI221 U133 ( .A(i_data_writeres[9]), .B(n13), .C(i_data_lwW[9]), .D(n17), 
        .Q(n62) );
  AOI221 U134 ( .A(i_data_writeres[6]), .B(n13), .C(i_data_lwW[6]), .D(n17), 
        .Q(n53) );
  AOI221 U135 ( .A(i_data_writeres[0]), .B(n1), .C(i_data_lwW[0]), .D(n4), .Q(
        n30) );
  AOI221 U136 ( .A(i_data_writeres[7]), .B(n13), .C(i_data_lwW[7]), .D(n4), 
        .Q(n56) );
  AOI221 U137 ( .A(i_data_writeres[5]), .B(n3), .C(i_data_lwW[5]), .D(n17), 
        .Q(n50) );
  AOI221 U138 ( .A(i_data_writeres[10]), .B(n1), .C(i_data_lwW[10]), .D(n18), 
        .Q(n65) );
  AOI221 U139 ( .A(i_data_writeres[26]), .B(n13), .C(i_data_lwW[26]), .D(n18), 
        .Q(n114) );
  AOI221 U140 ( .A(i_data_writeres[20]), .B(n1), .C(i_data_lwW[20]), .D(n4), 
        .Q(n95) );
  AOI221 U141 ( .A(i_data_lwM[25]), .B(n15), .C(i_data_lwW[25]), .D(n4), .Q(
        n108) );
  AOI221 U142 ( .A(i_data_lwM[24]), .B(n15), .C(i_data_alures[24]), .D(n21), 
        .Q(n106) );
  AOI220 U143 ( .A(i_data_lwM[31]), .B(n15), .C(i_data_alures[31]), .D(n21), 
        .Q(n132) );
  AOI221 U144 ( .A(i_data_lwM[27]), .B(n15), .C(i_data_lwW[27]), .D(n17), .Q(
        n115) );
  AOI221 U145 ( .A(i_data_lwM[18]), .B(n15), .C(i_data_alures[18]), .D(n22), 
        .Q(n88) );
  NAND21 U146 ( .A(i_data_rs[8]), .B(n130), .Q(n57) );
  NAND34 U147 ( .A(n50), .B(n49), .C(n48), .Q(o_data_alusra[5]) );
  NAND34 U148 ( .A(n56), .B(n55), .C(n54), .Q(o_data_alusra[7]) );
  AOI221 U149 ( .A(i_data_writeres[12]), .B(n2), .C(i_data_lwW[12]), .D(n4), 
        .Q(n71) );
  NAND22 U150 ( .A(n14), .B(i_data_rs[30]), .Q(n125) );
  NAND34 U151 ( .A(n36), .B(n35), .C(n34), .Q(o_data_alusra[1]) );
  NAND21 U152 ( .A(n14), .B(i_data_rs[24]), .Q(n105) );
  XNR22 U153 ( .A(n46), .B(n12), .Q(n27) );
  NAND22 U154 ( .A(i_data_alures[1]), .B(n21), .Q(n35) );
  NAND22 U155 ( .A(i_data_rs[5]), .B(n130), .Q(n48) );
  NAND33 U156 ( .A(n53), .B(n52), .C(n51), .Q(o_data_alusra[6]) );
  NAND22 U157 ( .A(i_data_rs[7]), .B(n130), .Q(n54) );
  NAND22 U158 ( .A(i_data_rs[11]), .B(n121), .Q(n66) );
  NAND22 U159 ( .A(i_data_rs[14]), .B(n121), .Q(n75) );
  NAND22 U160 ( .A(i_data_rs[17]), .B(n111), .Q(n84) );
  NAND33 U161 ( .A(n89), .B(n88), .C(n87), .Q(o_data_alusra[18]) );
  NAND33 U162 ( .A(n107), .B(n106), .C(n105), .Q(o_data_alusra[24]) );
  NAND33 U163 ( .A(n114), .B(n113), .C(n112), .Q(o_data_alusra[26]) );
  NAND33 U164 ( .A(n117), .B(n116), .C(n115), .Q(o_data_alusra[27]) );
  NAND33 U165 ( .A(n133), .B(n132), .C(n131), .Q(o_data_alusra[31]) );
endmodule


module E_fbmux5 ( i_data_rt, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fb, o_data_alusrb );
  input [31:0] i_data_rt;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fb;
  output [31:0] o_data_alusrb;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135;

  NAND34 U1 ( .A(n32), .B(n31), .C(n30), .Q(o_data_alusrb[1]) );
  NAND26 U2 ( .A(n38), .B(n14), .Q(o_data_alusrb[3]) );
  CLKIN12 U3 ( .A(i_con_fb[1]), .Q(n74) );
  NAND23 U4 ( .A(i_data_rt[11]), .B(n94), .Q(n62) );
  INV4 U5 ( .A(n74), .Q(n9) );
  NAND34 U6 ( .A(n49), .B(n50), .C(n51), .Q(o_data_alusrb[7]) );
  CLKIN8 U7 ( .A(i_con_fb[2]), .Q(n72) );
  AOI222 U8 ( .A(i_data_lwM[25]), .B(n18), .C(i_data_lwW[25]), .D(n21), .Q(
        n111) );
  NAND34 U9 ( .A(n64), .B(n63), .C(n62), .Q(o_data_alusrb[11]) );
  NAND34 U10 ( .A(n42), .B(n41), .C(n40), .Q(o_data_alusrb[4]) );
  AOI222 U11 ( .A(i_data_writeres[1]), .B(n15), .C(i_data_alures[1]), .D(n6), 
        .Q(n32) );
  AOI222 U12 ( .A(i_data_writeres[25]), .B(n16), .C(i_data_alures[25]), .D(n7), 
        .Q(n112) );
  NAND34 U13 ( .A(n112), .B(n111), .C(n110), .Q(o_data_alusrb[25]) );
  INV6 U14 ( .A(n13), .Q(n14) );
  AOI221 U15 ( .A(i_data_lwM[4]), .B(n17), .C(i_data_alures[4]), .D(n7), .Q(
        n41) );
  NAND33 U16 ( .A(n58), .B(n57), .C(n56), .Q(o_data_alusrb[9]) );
  NAND33 U17 ( .A(n70), .B(n69), .C(n68), .Q(o_data_alusrb[13]) );
  NAND33 U18 ( .A(n87), .B(n86), .C(n85), .Q(o_data_alusrb[17]) );
  NAND33 U19 ( .A(n90), .B(n89), .C(n88), .Q(o_data_alusrb[18]) );
  NAND33 U20 ( .A(n100), .B(n99), .C(n98), .Q(o_data_alusrb[21]) );
  NAND33 U21 ( .A(n103), .B(n102), .C(n101), .Q(o_data_alusrb[22]) );
  AOI222 U22 ( .A(i_data_writeres[3]), .B(n15), .C(i_data_lwW[3]), .D(n20), 
        .Q(n39) );
  INV6 U23 ( .A(n26), .Q(n129) );
  NAND24 U24 ( .A(n72), .B(n71), .Q(n19) );
  INV6 U25 ( .A(n19), .Q(n10) );
  NAND22 U26 ( .A(i_data_rt[10]), .B(n94), .Q(n59) );
  NAND24 U27 ( .A(n39), .B(n37), .Q(n13) );
  NAND33 U28 ( .A(n55), .B(n54), .C(n53), .Q(o_data_alusrb[8]) );
  NAND33 U29 ( .A(n65), .B(n66), .C(n67), .Q(o_data_alusrb[12]) );
  NAND33 U30 ( .A(n83), .B(n82), .C(n81), .Q(o_data_alusrb[16]) );
  NAND22 U31 ( .A(i_data_rt[21]), .B(n94), .Q(n98) );
  AOI221 U32 ( .A(i_data_lwM[23]), .B(n17), .C(i_data_lwW[23]), .D(n21), .Q(
        n105) );
  NAND33 U33 ( .A(n115), .B(n114), .C(n113), .Q(o_data_alusrb[26]) );
  NAND23 U34 ( .A(i_data_rt[19]), .B(n84), .Q(n91) );
  CLKBU12 U35 ( .A(n131), .Q(n6) );
  CLKBU12 U36 ( .A(n131), .Q(n7) );
  AOI222 U37 ( .A(i_data_lwM[24]), .B(n18), .C(i_data_lwW[24]), .D(n22), .Q(
        n108) );
  NAND33 U38 ( .A(n61), .B(n60), .C(n59), .Q(o_data_alusrb[10]) );
  NAND33 U39 ( .A(n45), .B(n44), .C(n43), .Q(o_data_alusrb[5]) );
  AOI221 U40 ( .A(i_data_lwM[28]), .B(n18), .C(i_data_alures[28]), .D(n7), .Q(
        n120) );
  AOI220 U41 ( .A(i_data_lwM[31]), .B(n18), .C(i_data_alures[31]), .D(n7), .Q(
        n134) );
  AOI221 U42 ( .A(i_data_lwM[29]), .B(n18), .C(i_data_alures[29]), .D(n7), .Q(
        n123) );
  NAND33 U43 ( .A(n48), .B(n47), .C(n46), .Q(o_data_alusrb[6]) );
  AOI221 U44 ( .A(i_data_lwM[6]), .B(n18), .C(i_data_lwW[6]), .D(n20), .Q(n47)
         );
  NAND21 U45 ( .A(i_data_rt[15]), .B(n3), .Q(n78) );
  INV6 U46 ( .A(n24), .Q(n131) );
  NAND23 U47 ( .A(i_data_rt[18]), .B(n84), .Q(n88) );
  NAND33 U48 ( .A(n135), .B(n134), .C(n133), .Q(o_data_alusrb[31]) );
  AOI222 U49 ( .A(i_data_writeres[24]), .B(n16), .C(i_data_alures[24]), .D(n6), 
        .Q(n109) );
  NAND34 U50 ( .A(n109), .B(n108), .C(n107), .Q(o_data_alusrb[24]) );
  AOI221 U51 ( .A(i_data_writeres[28]), .B(n16), .C(i_data_lwW[28]), .D(n22), 
        .Q(n121) );
  AOI222 U52 ( .A(i_data_writeres[18]), .B(n15), .C(i_data_lwW[18]), .D(n22), 
        .Q(n90) );
  AOI222 U53 ( .A(i_data_writeres[2]), .B(n15), .C(i_data_lwW[2]), .D(n20), 
        .Q(n36) );
  AOI222 U54 ( .A(i_data_writeres[7]), .B(n16), .C(i_data_alures[7]), .D(n7), 
        .Q(n51) );
  AOI221 U55 ( .A(i_data_rt[30]), .B(n8), .C(i_data_writeres[30]), .D(n16), 
        .Q(n128) );
  AOI221 U56 ( .A(i_data_lwM[7]), .B(n18), .C(i_data_lwW[7]), .D(n20), .Q(n50)
         );
  AOI221 U57 ( .A(i_data_lwM[0]), .B(n18), .C(i_data_lwW[0]), .D(n20), .Q(n28)
         );
  AOI221 U58 ( .A(i_data_lwM[22]), .B(n18), .C(i_data_lwW[22]), .D(n20), .Q(
        n102) );
  AOI221 U59 ( .A(i_data_lwM[5]), .B(n18), .C(i_data_lwW[5]), .D(n20), .Q(n44)
         );
  CLKIN3 U60 ( .A(n52), .Q(n3) );
  CLKIN6 U61 ( .A(n52), .Q(n125) );
  AOI222 U62 ( .A(i_data_writeres[8]), .B(n15), .C(i_data_alures[8]), .D(n6), 
        .Q(n55) );
  AOI221 U63 ( .A(i_data_writeres[4]), .B(n15), .C(i_data_lwW[4]), .D(n20), 
        .Q(n42) );
  NAND34 U64 ( .A(n77), .B(n76), .C(n75), .Q(o_data_alusrb[14]) );
  NAND24 U65 ( .A(n80), .B(n2), .Q(o_data_alusrb[15]) );
  AOI221 U66 ( .A(i_data_writeres[15]), .B(n16), .C(i_data_alures[15]), .D(n6), 
        .Q(n80) );
  CLKIN3 U67 ( .A(n52), .Q(n8) );
  CLKIN6 U68 ( .A(n25), .Q(n132) );
  NAND32 U69 ( .A(n71), .B(n74), .C(i_con_fb[2]), .Q(n25) );
  CLKIN6 U70 ( .A(i_con_fb[0]), .Q(n71) );
  AOI222 U71 ( .A(i_data_lwM[17]), .B(n17), .C(i_data_alures[17]), .D(n7), .Q(
        n86) );
  AOI222 U72 ( .A(i_data_writeres[17]), .B(n16), .C(i_data_lwW[17]), .D(n21), 
        .Q(n87) );
  BUF15 U73 ( .A(n132), .Q(n17) );
  BUF15 U74 ( .A(n132), .Q(n18) );
  NAND34 U75 ( .A(n97), .B(n96), .C(n95), .Q(o_data_alusrb[20]) );
  NAND34 U76 ( .A(n106), .B(n105), .C(n104), .Q(o_data_alusrb[23]) );
  AOI221 U77 ( .A(i_data_lwM[30]), .B(n18), .C(i_data_lwW[30]), .D(n22), .Q(
        n126) );
  CLKBU15 U78 ( .A(n129), .Q(n22) );
  NAND22 U79 ( .A(i_data_rt[3]), .B(n84), .Q(n37) );
  CLKBU15 U80 ( .A(n129), .Q(n21) );
  AOI222 U81 ( .A(i_data_lwM[11]), .B(n17), .C(i_data_lwW[11]), .D(n21), .Q(
        n63) );
  AOI221 U82 ( .A(i_data_writeres[5]), .B(n16), .C(i_data_alures[5]), .D(n7), 
        .Q(n45) );
  AOI221 U83 ( .A(i_data_writeres[29]), .B(n16), .C(i_data_lwW[29]), .D(n21), 
        .Q(n124) );
  NAND23 U84 ( .A(n74), .B(n19), .Q(n11) );
  CLKIN15 U85 ( .A(n52), .Q(n94) );
  NAND22 U86 ( .A(n78), .B(n79), .Q(n1) );
  INV3 U87 ( .A(n1), .Q(n2) );
  NAND22 U88 ( .A(i_data_rt[13]), .B(n125), .Q(n68) );
  NAND22 U89 ( .A(i_data_rt[16]), .B(n94), .Q(n81) );
  AOI222 U90 ( .A(i_data_writeres[9]), .B(n15), .C(i_data_alures[9]), .D(n7), 
        .Q(n58) );
  AOI221 U91 ( .A(i_data_writeres[22]), .B(n16), .C(i_data_alures[22]), .D(n6), 
        .Q(n103) );
  BUF15 U92 ( .A(n130), .Q(n16) );
  NAND32 U93 ( .A(i_con_fb[1]), .B(n71), .C(n72), .Q(n24) );
  AOI221 U94 ( .A(i_data_writeres[0]), .B(n16), .C(i_data_alures[0]), .D(n6), 
        .Q(n29) );
  AOI221 U95 ( .A(i_data_lwM[3]), .B(n17), .C(i_data_alures[3]), .D(n7), .Q(
        n38) );
  CLKIN8 U96 ( .A(n33), .Q(n84) );
  XOR22 U97 ( .A(n9), .B(n73), .Q(n33) );
  CLKBU15 U98 ( .A(n129), .Q(n20) );
  NAND21 U99 ( .A(i_con_fb[2]), .B(i_con_fb[0]), .Q(n4) );
  NAND24 U100 ( .A(n74), .B(n5), .Q(n26) );
  INV3 U101 ( .A(n4), .Q(n5) );
  AOI222 U102 ( .A(i_data_lwM[16]), .B(n17), .C(i_data_lwW[16]), .D(n22), .Q(
        n82) );
  NAND26 U103 ( .A(n9), .B(n10), .Q(n12) );
  NAND28 U104 ( .A(n11), .B(n12), .Q(n52) );
  NAND21 U105 ( .A(i_data_rt[7]), .B(n125), .Q(n49) );
  NAND31 U106 ( .A(n74), .B(n72), .C(i_con_fb[0]), .Q(n23) );
  NAND22 U107 ( .A(i_data_rt[1]), .B(n125), .Q(n30) );
  NAND33 U108 ( .A(n29), .B(n28), .C(n27), .Q(o_data_alusrb[0]) );
  NAND21 U109 ( .A(i_data_rt[22]), .B(n94), .Q(n101) );
  NAND22 U110 ( .A(n72), .B(n71), .Q(n73) );
  AOI221 U111 ( .A(i_data_lwM[27]), .B(n18), .C(i_data_lwW[27]), .D(n21), .Q(
        n117) );
  AOI221 U112 ( .A(i_data_writeres[27]), .B(n16), .C(i_data_alures[27]), .D(n6), .Q(n118) );
  AOI220 U113 ( .A(i_data_writeres[31]), .B(n16), .C(i_data_lwW[31]), .D(n21), 
        .Q(n135) );
  BUF15 U114 ( .A(n130), .Q(n15) );
  CLKIN6 U115 ( .A(n23), .Q(n130) );
  NAND22 U116 ( .A(i_data_rt[25]), .B(n125), .Q(n110) );
  NAND22 U117 ( .A(i_data_rt[17]), .B(n84), .Q(n85) );
  NAND22 U118 ( .A(i_data_rt[4]), .B(n84), .Q(n40) );
  NAND34 U119 ( .A(n36), .B(n35), .C(n34), .Q(o_data_alusrb[2]) );
  NAND22 U120 ( .A(i_data_rt[20]), .B(n125), .Q(n95) );
  NAND22 U121 ( .A(i_data_rt[23]), .B(n125), .Q(n104) );
  NAND22 U122 ( .A(i_data_rt[8]), .B(n94), .Q(n53) );
  NAND22 U123 ( .A(i_data_rt[9]), .B(n94), .Q(n56) );
  NAND34 U124 ( .A(n92), .B(n93), .C(n91), .Q(o_data_alusrb[19]) );
  NAND22 U125 ( .A(i_data_rt[0]), .B(n94), .Q(n27) );
  AOI222 U126 ( .A(i_data_lwM[1]), .B(n17), .C(i_data_lwW[1]), .D(n20), .Q(n31) );
  AOI222 U127 ( .A(i_data_lwM[2]), .B(n17), .C(i_data_alures[2]), .D(n6), .Q(
        n35) );
  NAND22 U128 ( .A(i_data_rt[2]), .B(n84), .Q(n34) );
  NAND22 U129 ( .A(i_data_rt[5]), .B(n3), .Q(n43) );
  AOI222 U130 ( .A(i_data_writeres[6]), .B(n16), .C(i_data_alures[6]), .D(n6), 
        .Q(n48) );
  NAND22 U131 ( .A(i_data_rt[6]), .B(n94), .Q(n46) );
  AOI222 U132 ( .A(i_data_lwM[8]), .B(n17), .C(i_data_lwW[8]), .D(n20), .Q(n54) );
  AOI222 U133 ( .A(i_data_lwM[9]), .B(n17), .C(i_data_lwW[9]), .D(n20), .Q(n57) );
  AOI222 U134 ( .A(i_data_writeres[10]), .B(n15), .C(i_data_alures[10]), .D(n7), .Q(n61) );
  AOI222 U135 ( .A(i_data_lwM[10]), .B(n17), .C(i_data_lwW[10]), .D(n20), .Q(
        n60) );
  AOI222 U136 ( .A(i_data_writeres[11]), .B(n15), .C(i_data_alures[11]), .D(n6), .Q(n64) );
  AOI222 U137 ( .A(i_data_writeres[12]), .B(n15), .C(i_data_alures[12]), .D(n6), .Q(n67) );
  AOI222 U138 ( .A(i_data_lwM[12]), .B(n18), .C(i_data_lwW[12]), .D(n22), .Q(
        n66) );
  NAND22 U139 ( .A(i_data_rt[12]), .B(n8), .Q(n65) );
  AOI222 U140 ( .A(i_data_writeres[13]), .B(n16), .C(i_data_alures[13]), .D(n6), .Q(n70) );
  AOI222 U141 ( .A(i_data_lwM[13]), .B(n18), .C(i_data_lwW[13]), .D(n21), .Q(
        n69) );
  AOI222 U142 ( .A(i_data_writeres[14]), .B(n16), .C(i_data_alures[14]), .D(n7), .Q(n77) );
  AOI222 U143 ( .A(i_data_lwM[14]), .B(n18), .C(i_data_lwW[14]), .D(n22), .Q(
        n76) );
  NAND22 U144 ( .A(i_data_rt[14]), .B(n125), .Q(n75) );
  AOI222 U145 ( .A(i_data_lwM[15]), .B(n18), .C(i_data_lwW[15]), .D(n21), .Q(
        n79) );
  AOI222 U146 ( .A(i_data_writeres[16]), .B(n15), .C(i_data_alures[16]), .D(n6), .Q(n83) );
  AOI222 U147 ( .A(i_data_lwM[18]), .B(n17), .C(i_data_alures[18]), .D(n7), 
        .Q(n89) );
  AOI222 U148 ( .A(i_data_writeres[19]), .B(n15), .C(i_data_lwW[19]), .D(n21), 
        .Q(n93) );
  AOI222 U149 ( .A(i_data_lwM[19]), .B(n17), .C(i_data_alures[19]), .D(n7), 
        .Q(n92) );
  AOI222 U150 ( .A(i_data_writeres[20]), .B(n16), .C(i_data_alures[20]), .D(n7), .Q(n97) );
  AOI222 U151 ( .A(i_data_lwM[20]), .B(n18), .C(i_data_lwW[20]), .D(n22), .Q(
        n96) );
  AOI222 U152 ( .A(i_data_writeres[21]), .B(n16), .C(i_data_alures[21]), .D(n7), .Q(n100) );
  AOI222 U153 ( .A(i_data_lwM[21]), .B(n18), .C(i_data_lwW[21]), .D(n21), .Q(
        n99) );
  AOI222 U154 ( .A(i_data_writeres[23]), .B(n16), .C(i_data_alures[23]), .D(n6), .Q(n106) );
  NAND22 U155 ( .A(i_data_rt[24]), .B(n3), .Q(n107) );
  AOI222 U156 ( .A(i_data_writeres[26]), .B(n16), .C(i_data_alures[26]), .D(n6), .Q(n115) );
  AOI222 U157 ( .A(i_data_lwM[26]), .B(n18), .C(i_data_lwW[26]), .D(n22), .Q(
        n114) );
  NAND22 U158 ( .A(i_data_rt[26]), .B(n94), .Q(n113) );
  NAND22 U159 ( .A(i_data_rt[27]), .B(n3), .Q(n116) );
  NAND33 U160 ( .A(n118), .B(n117), .C(n116), .Q(o_data_alusrb[27]) );
  NAND22 U161 ( .A(i_data_rt[28]), .B(n8), .Q(n119) );
  NAND33 U162 ( .A(n121), .B(n120), .C(n119), .Q(o_data_alusrb[28]) );
  NAND22 U163 ( .A(i_data_rt[29]), .B(n8), .Q(n122) );
  NAND33 U164 ( .A(n124), .B(n123), .C(n122), .Q(o_data_alusrb[29]) );
  NAND22 U165 ( .A(i_data_alures[30]), .B(n6), .Q(n127) );
  NAND33 U166 ( .A(n128), .B(n127), .C(n126), .Q(o_data_alusrb[30]) );
  NAND22 U167 ( .A(i_data_rt[31]), .B(n8), .Q(n133) );
endmodule


module E_alubmux ( i_data_fb, i_data_imm, i_con_imm, o_data_alub );
  input [31:0] i_data_fb;
  input [31:0] i_data_imm;
  output [31:0] o_data_alub;
  input i_con_imm;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60;

  INV6 U1 ( .A(n42), .Q(o_data_alub[19]) );
  INV12 U2 ( .A(n14), .Q(o_data_alub[3]) );
  CLKIN6 U3 ( .A(n46), .Q(o_data_alub[21]) );
  CLKIN15 U4 ( .A(n15), .Q(o_data_alub[4]) );
  CLKIN12 U5 ( .A(n38), .Q(o_data_alub[17]) );
  CLKIN12 U6 ( .A(n31), .Q(o_data_alub[12]) );
  CLKIN12 U7 ( .A(n19), .Q(o_data_alub[6]) );
  INV3 U8 ( .A(n50), .Q(o_data_alub[25]) );
  INV3 U9 ( .A(n26), .Q(o_data_alub[9]) );
  INV3 U10 ( .A(n43), .Q(o_data_alub[20]) );
  INV3 U11 ( .A(n37), .Q(o_data_alub[16]) );
  INV8 U12 ( .A(n22), .Q(o_data_alub[7]) );
  CLKIN6 U13 ( .A(n34), .Q(o_data_alub[15]) );
  CLKIN6 U14 ( .A(n49), .Q(o_data_alub[24]) );
  INV4 U15 ( .A(n56), .Q(o_data_alub[27]) );
  INV3 U16 ( .A(n27), .Q(o_data_alub[10]) );
  INV6 U17 ( .A(n18), .Q(o_data_alub[5]) );
  INV3 U18 ( .A(n54), .Q(n55) );
  CLKIN6 U19 ( .A(n28), .Q(o_data_alub[11]) );
  INV3 U20 ( .A(n53), .Q(o_data_alub[26]) );
  INV6 U21 ( .A(n9), .Q(o_data_alub[0]) );
  INV6 U22 ( .A(n47), .Q(o_data_alub[22]) );
  CLKIN6 U23 ( .A(n48), .Q(o_data_alub[23]) );
  CLKIN6 U24 ( .A(n32), .Q(o_data_alub[13]) );
  AOI221 U25 ( .A(i_data_fb[30]), .B(n1), .C(i_data_imm[30]), .D(n4), .Q(n59)
         );
  AOI221 U26 ( .A(i_data_fb[29]), .B(n1), .C(i_data_imm[29]), .D(n4), .Q(n58)
         );
  INV4 U27 ( .A(n33), .Q(o_data_alub[14]) );
  AOI222 U28 ( .A(i_data_fb[25]), .B(n1), .C(i_data_imm[25]), .D(n4), .Q(n50)
         );
  INV6 U29 ( .A(n25), .Q(o_data_alub[8]) );
  AOI222 U30 ( .A(i_data_fb[28]), .B(n1), .C(i_data_imm[28]), .D(n4), .Q(n57)
         );
  INV3 U31 ( .A(n60), .Q(o_data_alub[31]) );
  AOI221 U32 ( .A(i_data_fb[31]), .B(n2), .C(i_data_imm[31]), .D(n6), .Q(n60)
         );
  BUF6 U33 ( .A(i_con_imm), .Q(n6) );
  AOI222 U34 ( .A(i_data_fb[2]), .B(n3), .C(i_data_imm[2]), .D(n6), .Q(n13) );
  CLKIN2 U35 ( .A(i_con_imm), .Q(n3) );
  NAND22 U36 ( .A(i_data_imm[18]), .B(n6), .Q(n39) );
  NAND22 U37 ( .A(i_data_imm[21]), .B(n6), .Q(n44) );
  NAND21 U38 ( .A(i_data_imm[8]), .B(n6), .Q(n23) );
  CLKIN3 U39 ( .A(i_con_imm), .Q(n1) );
  AOI222 U40 ( .A(i_data_fb[24]), .B(n1), .C(i_data_imm[24]), .D(n4), .Q(n49)
         );
  CLKIN3 U41 ( .A(i_con_imm), .Q(n2) );
  NAND20 U42 ( .A(i_data_imm[26]), .B(n6), .Q(n51) );
  AOI222 U43 ( .A(i_data_fb[3]), .B(n2), .C(i_data_imm[3]), .D(n6), .Q(n14) );
  INV2 U44 ( .A(n39), .Q(n40) );
  AOI222 U45 ( .A(i_data_fb[20]), .B(n1), .C(i_data_imm[20]), .D(n4), .Q(n43)
         );
  INV2 U46 ( .A(n44), .Q(n45) );
  NAND20 U47 ( .A(i_data_imm[0]), .B(n6), .Q(n7) );
  NAND20 U48 ( .A(i_data_imm[5]), .B(n6), .Q(n16) );
  NAND20 U49 ( .A(i_data_imm[1]), .B(n6), .Q(n10) );
  NAND20 U50 ( .A(i_data_imm[16]), .B(n6), .Q(n35) );
  INV8 U51 ( .A(n12), .Q(o_data_alub[1]) );
  BUF2 U52 ( .A(i_con_imm), .Q(n5) );
  BUF2 U53 ( .A(i_con_imm), .Q(n4) );
  INV12 U54 ( .A(n13), .Q(o_data_alub[2]) );
  CLKIN3 U55 ( .A(n7), .Q(n8) );
  OAI222 U56 ( .A(n8), .B(n3), .C(i_data_fb[0]), .D(n8), .Q(n9) );
  CLKIN3 U57 ( .A(n10), .Q(n11) );
  OAI222 U58 ( .A(n11), .B(n3), .C(i_data_fb[1]), .D(n11), .Q(n12) );
  AOI222 U59 ( .A(i_data_fb[4]), .B(n2), .C(i_data_imm[4]), .D(n6), .Q(n15) );
  CLKIN3 U60 ( .A(n16), .Q(n17) );
  OAI222 U61 ( .A(i_data_fb[5]), .B(n17), .C(n17), .D(n2), .Q(n18) );
  AOI222 U62 ( .A(i_data_fb[6]), .B(n2), .C(i_data_imm[6]), .D(n6), .Q(n19) );
  NAND22 U63 ( .A(i_data_imm[7]), .B(n5), .Q(n20) );
  CLKIN3 U64 ( .A(n20), .Q(n21) );
  OAI222 U65 ( .A(n21), .B(n3), .C(i_data_fb[7]), .D(n21), .Q(n22) );
  CLKIN3 U66 ( .A(n23), .Q(n24) );
  OAI222 U67 ( .A(n24), .B(n3), .C(i_data_fb[8]), .D(n24), .Q(n25) );
  AOI222 U68 ( .A(i_data_fb[9]), .B(n2), .C(i_data_imm[9]), .D(n5), .Q(n26) );
  AOI222 U69 ( .A(i_data_fb[10]), .B(n2), .C(i_data_imm[10]), .D(n5), .Q(n27)
         );
  AOI222 U70 ( .A(i_data_fb[11]), .B(n2), .C(i_data_imm[11]), .D(n5), .Q(n28)
         );
  NAND22 U71 ( .A(i_data_imm[12]), .B(n6), .Q(n29) );
  CLKIN3 U72 ( .A(n29), .Q(n30) );
  OAI222 U73 ( .A(i_data_fb[12]), .B(n30), .C(n30), .D(n2), .Q(n31) );
  AOI222 U74 ( .A(i_data_fb[13]), .B(n2), .C(i_data_imm[13]), .D(n5), .Q(n32)
         );
  AOI222 U75 ( .A(i_data_fb[14]), .B(n2), .C(i_data_imm[14]), .D(n5), .Q(n33)
         );
  AOI222 U76 ( .A(i_data_fb[15]), .B(n2), .C(i_data_imm[15]), .D(n5), .Q(n34)
         );
  CLKIN3 U77 ( .A(n35), .Q(n36) );
  OAI222 U78 ( .A(n36), .B(n3), .C(i_data_fb[16]), .D(n36), .Q(n37) );
  AOI222 U79 ( .A(i_data_fb[17]), .B(n2), .C(i_data_imm[17]), .D(n5), .Q(n38)
         );
  OAI222 U80 ( .A(i_data_fb[18]), .B(n40), .C(n40), .D(n1), .Q(n41) );
  CLKIN3 U81 ( .A(n41), .Q(o_data_alub[18]) );
  AOI222 U82 ( .A(i_data_fb[19]), .B(n1), .C(i_data_imm[19]), .D(n5), .Q(n42)
         );
  OAI222 U83 ( .A(i_data_fb[21]), .B(n45), .C(n45), .D(n1), .Q(n46) );
  AOI222 U84 ( .A(i_data_fb[22]), .B(n1), .C(i_data_imm[22]), .D(n4), .Q(n47)
         );
  AOI222 U85 ( .A(i_data_fb[23]), .B(n1), .C(i_data_imm[23]), .D(n4), .Q(n48)
         );
  CLKIN3 U86 ( .A(n51), .Q(n52) );
  OAI222 U87 ( .A(i_data_fb[26]), .B(n52), .C(n52), .D(n1), .Q(n53) );
  NAND22 U88 ( .A(i_data_imm[27]), .B(n4), .Q(n54) );
  OAI222 U89 ( .A(i_data_fb[27]), .B(n55), .C(n55), .D(n1), .Q(n56) );
  CLKIN3 U90 ( .A(n57), .Q(o_data_alub[28]) );
  CLKIN3 U91 ( .A(n58), .Q(o_data_alub[29]) );
  CLKIN3 U92 ( .A(n59), .Q(o_data_alub[30]) );
endmodule


module E_rdmux ( i_data_rtE, i_data_rdE, i_con_regdst, i_con_aluPC4, 
        o_data_writeE );
  input [4:0] i_data_rtE;
  input [4:0] i_data_rdE;
  output [4:0] o_data_writeE;
  input i_con_regdst, i_con_aluPC4;
  wire   n7, n8, n9, n10, n11, n1, n2, n3, n4, n5, n6, n12;

  NAND21 U2 ( .A(i_data_rdE[1]), .B(n1), .Q(n10) );
  NAND21 U3 ( .A(i_data_rdE[2]), .B(n1), .Q(n9) );
  OAI2110 U4 ( .A(n1), .B(n2), .C(n12), .D(n7), .Q(o_data_writeE[4]) );
  NAND20 U5 ( .A(i_data_rdE[4]), .B(n1), .Q(n7) );
  OAI2111 U6 ( .A(n1), .B(n6), .C(n12), .D(n11), .Q(o_data_writeE[0]) );
  INV3 U7 ( .A(i_data_rtE[0]), .Q(n6) );
  NAND22 U8 ( .A(i_data_rdE[0]), .B(n1), .Q(n11) );
  OAI2111 U9 ( .A(n1), .B(n5), .C(n12), .D(n10), .Q(o_data_writeE[1]) );
  INV3 U10 ( .A(i_data_rtE[1]), .Q(n5) );
  OAI2111 U11 ( .A(n1), .B(n4), .C(n12), .D(n9), .Q(o_data_writeE[2]) );
  INV3 U12 ( .A(i_data_rtE[2]), .Q(n4) );
  INV3 U13 ( .A(i_data_rtE[4]), .Q(n2) );
  OAI2111 U14 ( .A(n1), .B(n3), .C(n12), .D(n8), .Q(o_data_writeE[3]) );
  INV3 U15 ( .A(i_data_rtE[3]), .Q(n3) );
  NAND22 U16 ( .A(i_data_rdE[3]), .B(n1), .Q(n8) );
  BUF2 U17 ( .A(i_con_regdst), .Q(n1) );
  INV3 U18 ( .A(i_con_aluPC4), .Q(n12) );
endmodule


module D_compare_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172;

  CLKIN2 U1 ( .A(B[27]), .Q(n95) );
  INV6 U2 ( .A(A[6]), .Q(n68) );
  CLKIN3 U3 ( .A(A[4]), .Q(n72) );
  NAND22 U4 ( .A(n107), .B(n108), .Q(n101) );
  NOR21 U5 ( .A(n56), .B(n57), .Q(n48) );
  NOR23 U6 ( .A(n19), .B(n20), .Q(n18) );
  INV3 U7 ( .A(A[19]), .Q(n109) );
  INV3 U8 ( .A(A[0]), .Q(n97) );
  NOR22 U9 ( .A(n31), .B(n32), .Q(n15) );
  NAND23 U10 ( .A(n61), .B(n62), .Q(n44) );
  NOR22 U11 ( .A(n63), .B(n64), .Q(n62) );
  NAND22 U12 ( .A(n65), .B(n66), .Q(n64) );
  NOR22 U13 ( .A(n36), .B(n35), .Q(n11) );
  INV1 U14 ( .A(B[19]), .Q(n171) );
  NAND21 U15 ( .A(n33), .B(n34), .Q(n170) );
  NAND20 U16 ( .A(A[9]), .B(n92), .Q(n37) );
  NAND20 U17 ( .A(B[19]), .B(n109), .Q(n107) );
  NAND34 U18 ( .A(n17), .B(n16), .C(n15), .Q(n3) );
  NOR22 U19 ( .A(n27), .B(n28), .Q(n16) );
  AOI2112 U20 ( .A(A[1]), .B(n91), .C(n130), .D(n131), .Q(n129) );
  INV0 U21 ( .A(A[10]), .Q(n5) );
  INV2 U22 ( .A(B[15]), .Q(n53) );
  CLKIN1 U23 ( .A(A[8]), .Q(n82) );
  NAND22 U24 ( .A(n158), .B(n159), .Q(n19) );
  NAND22 U25 ( .A(n161), .B(n162), .Q(n20) );
  NAND22 U26 ( .A(n151), .B(n152), .Q(n145) );
  NOR23 U27 ( .A(n101), .B(n102), .Q(n100) );
  INV3 U28 ( .A(B[28]), .Q(n96) );
  INV3 U29 ( .A(A[12]), .Q(n78) );
  INV3 U30 ( .A(A[5]), .Q(n81) );
  NAND22 U31 ( .A(n69), .B(n70), .Q(n63) );
  NOR21 U32 ( .A(A[9]), .B(n92), .Q(n89) );
  NAND22 U33 ( .A(n25), .B(n26), .Q(n21) );
  INV3 U34 ( .A(n34), .Q(n31) );
  INV3 U35 ( .A(n35), .Q(n119) );
  NAND22 U36 ( .A(n156), .B(n157), .Q(n155) );
  NAND23 U37 ( .A(n1), .B(n134), .Q(n13) );
  INV3 U38 ( .A(A[2]), .Q(n71) );
  INV2 U39 ( .A(A[21]), .Q(n106) );
  AOI2111 U40 ( .A(n2), .B(A[21]), .C(n145), .D(n146), .Q(n1) );
  NAND22 U41 ( .A(n37), .B(n129), .Q(n36) );
  INV3 U42 ( .A(n129), .Q(n38) );
  NOR21 U43 ( .A(A[1]), .B(n91), .Q(n90) );
  AOI2111 U44 ( .A(B[10]), .B(n5), .C(n89), .D(n90), .Q(n88) );
  NOR31 U45 ( .A(n50), .B(n51), .C(n52), .Q(n49) );
  INV1 U46 ( .A(B[1]), .Q(n91) );
  NAND21 U47 ( .A(n25), .B(n26), .Q(n165) );
  CLKIN1 U48 ( .A(B[25]), .Q(n144) );
  NAND21 U49 ( .A(B[25]), .B(n114), .Q(n112) );
  NOR32 U50 ( .A(n40), .B(n41), .C(n39), .Q(EQ) );
  NAND21 U51 ( .A(B[13]), .B(n60), .Q(n46) );
  NAND22 U52 ( .A(B[6]), .B(n68), .Q(n65) );
  NAND24 U53 ( .A(n99), .B(n100), .Q(n83) );
  NOR24 U54 ( .A(n83), .B(n84), .Q(n42) );
  NOR21 U55 ( .A(A[27]), .B(n95), .Q(n94) );
  CLKIN3 U56 ( .A(A[13]), .Q(n60) );
  NOR21 U57 ( .A(B[12]), .B(n78), .Q(n126) );
  INV3 U58 ( .A(A[23]), .Q(n117) );
  NAND24 U59 ( .A(n18), .B(n4), .Q(n14) );
  NAND21 U60 ( .A(B[3]), .B(n67), .Q(n66) );
  INV2 U61 ( .A(B[3]), .Q(n167) );
  NAND26 U62 ( .A(n42), .B(n43), .Q(n39) );
  NOR24 U63 ( .A(n44), .B(n45), .Q(n43) );
  NAND22 U64 ( .A(B[8]), .B(n82), .Q(n79) );
  NAND22 U65 ( .A(B[26]), .B(n9), .Q(n113) );
  INV6 U66 ( .A(n3), .Q(n4) );
  NAND21 U67 ( .A(B[2]), .B(n71), .Q(n70) );
  NAND22 U68 ( .A(B[4]), .B(n72), .Q(n69) );
  NAND21 U69 ( .A(A[13]), .B(n160), .Q(n158) );
  NAND24 U70 ( .A(n120), .B(n121), .Q(n35) );
  NOR22 U71 ( .A(n73), .B(n74), .Q(n61) );
  NOR23 U72 ( .A(n13), .B(n14), .Q(n12) );
  NAND21 U73 ( .A(B[29]), .B(n98), .Q(n85) );
  NAND21 U74 ( .A(B[5]), .B(n81), .Q(n80) );
  NOR22 U75 ( .A(n21), .B(n22), .Q(n17) );
  NOR22 U76 ( .A(A[17]), .B(n54), .Q(n51) );
  NOR21 U77 ( .A(A[18]), .B(n55), .Q(n50) );
  NOR21 U78 ( .A(B[7]), .B(n77), .Q(n127) );
  NAND21 U79 ( .A(n29), .B(n30), .Q(n169) );
  NAND22 U80 ( .A(A[17]), .B(n54), .Q(n29) );
  CLKIN2 U81 ( .A(A[25]), .Q(n114) );
  NAND22 U82 ( .A(A[25]), .B(n144), .Q(n143) );
  NOR22 U83 ( .A(B[0]), .B(n97), .Q(n130) );
  NOR21 U84 ( .A(A[15]), .B(n53), .Q(n52) );
  NOR21 U85 ( .A(B[2]), .B(n71), .Q(n131) );
  NAND34 U86 ( .A(n10), .B(n11), .C(n12), .Q(NE) );
  NAND43 U87 ( .A(n46), .B(n47), .C(n48), .D(n49), .Q(n45) );
  CLKIN2 U88 ( .A(n29), .Q(n28) );
  AOI2111 U89 ( .A(A[10]), .B(n125), .C(n127), .D(n126), .Q(n120) );
  NAND21 U90 ( .A(A[28]), .B(n96), .Q(n142) );
  NAND22 U91 ( .A(A[15]), .B(n53), .Q(n23) );
  CLKIN2 U92 ( .A(A[24]), .Q(n8) );
  NAND21 U93 ( .A(A[29]), .B(n150), .Q(n147) );
  NAND20 U94 ( .A(B[0]), .B(n97), .Q(n86) );
  NAND22 U95 ( .A(n138), .B(n139), .Q(n137) );
  NOR22 U96 ( .A(n154), .B(n155), .Q(n132) );
  INV3 U97 ( .A(n37), .Q(n128) );
  NAND22 U98 ( .A(A[14]), .B(n58), .Q(n24) );
  CLKIN0 U99 ( .A(B[13]), .Q(n160) );
  CLKIN0 U100 ( .A(B[26]), .Q(n153) );
  NAND20 U101 ( .A(A[23]), .B(n141), .Q(n138) );
  CLKIN0 U102 ( .A(B[29]), .Q(n150) );
  INV6 U103 ( .A(n39), .Q(n10) );
  NAND24 U104 ( .A(n118), .B(n119), .Q(n41) );
  INV6 U105 ( .A(A[7]), .Q(n77) );
  AOI2112 U106 ( .A(A[24]), .B(n135), .C(n136), .D(n137), .Q(n134) );
  NAND22 U107 ( .A(n147), .B(n148), .Q(n146) );
  NAND20 U108 ( .A(A[27]), .B(n95), .Q(n151) );
  NOR21 U109 ( .A(A[28]), .B(n96), .Q(n93) );
  NAND20 U110 ( .A(A[11]), .B(n59), .Q(n159) );
  CLKIN0 U111 ( .A(A[16]), .Q(n6) );
  CLKIN0 U112 ( .A(B[21]), .Q(n2) );
  NAND22 U113 ( .A(n163), .B(n164), .Q(n154) );
  NOR21 U114 ( .A(n169), .B(n170), .Q(n163) );
  NOR21 U115 ( .A(n110), .B(n111), .Q(n99) );
  NAND42 U116 ( .A(n85), .B(n86), .C(n87), .D(n88), .Q(n84) );
  NOR21 U117 ( .A(n165), .B(n166), .Q(n164) );
  NAND22 U118 ( .A(n23), .B(n24), .Q(n166) );
  NAND22 U119 ( .A(n23), .B(n24), .Q(n22) );
  INV3 U120 ( .A(A[3]), .Q(n67) );
  NAND22 U121 ( .A(A[3]), .B(n167), .Q(n26) );
  NAND22 U122 ( .A(n79), .B(n80), .Q(n73) );
  NAND22 U123 ( .A(A[19]), .B(n171), .Q(n33) );
  NAND22 U124 ( .A(A[18]), .B(n55), .Q(n34) );
  XNR21 U125 ( .A(B[31]), .B(A[31]), .Q(n161) );
  NAND22 U126 ( .A(A[16]), .B(n172), .Q(n30) );
  NOR21 U127 ( .A(B[5]), .B(n81), .Q(n122) );
  NAND22 U128 ( .A(n142), .B(n143), .Q(n136) );
  NAND22 U129 ( .A(A[8]), .B(n168), .Q(n25) );
  NOR21 U130 ( .A(A[11]), .B(n59), .Q(n56) );
  NAND22 U131 ( .A(n115), .B(n116), .Q(n110) );
  NOR21 U132 ( .A(A[14]), .B(n58), .Q(n57) );
  NAND22 U133 ( .A(n103), .B(n104), .Q(n102) );
  INV3 U134 ( .A(A[22]), .Q(n105) );
  NAND22 U135 ( .A(n112), .B(n113), .Q(n111) );
  NAND22 U136 ( .A(n75), .B(n76), .Q(n74) );
  NAND22 U137 ( .A(B[7]), .B(n77), .Q(n76) );
  NAND22 U138 ( .A(A[26]), .B(n153), .Q(n152) );
  NOR21 U139 ( .A(n93), .B(n94), .Q(n87) );
  INV3 U140 ( .A(A[26]), .Q(n9) );
  INV3 U141 ( .A(A[29]), .Q(n98) );
  NAND22 U142 ( .A(A[20]), .B(n149), .Q(n148) );
  INV3 U143 ( .A(A[20]), .Q(n7) );
  INV2 U144 ( .A(B[14]), .Q(n58) );
  NAND20 U145 ( .A(n106), .B(B[21]), .Q(n103) );
  INV1 U146 ( .A(B[9]), .Q(n92) );
  NAND22 U147 ( .A(B[22]), .B(n105), .Q(n104) );
  INV1 U148 ( .A(B[22]), .Q(n140) );
  INV1 U149 ( .A(B[11]), .Q(n59) );
  INV0 U150 ( .A(B[10]), .Q(n125) );
  CLKIN1 U151 ( .A(B[20]), .Q(n149) );
  INV2 U152 ( .A(B[18]), .Q(n55) );
  INV1 U153 ( .A(B[8]), .Q(n168) );
  INV2 U154 ( .A(n13), .Q(n133) );
  NAND21 U155 ( .A(B[24]), .B(n8), .Q(n116) );
  INV0 U156 ( .A(B[24]), .Q(n135) );
  NAND21 U157 ( .A(B[23]), .B(n117), .Q(n115) );
  NOR32 U158 ( .A(n122), .B(n123), .C(n124), .Q(n121) );
  INV2 U159 ( .A(B[17]), .Q(n54) );
  NOR21 U160 ( .A(B[6]), .B(n68), .Q(n123) );
  NAND21 U161 ( .A(B[20]), .B(n7), .Q(n108) );
  NAND22 U162 ( .A(B[12]), .B(n78), .Q(n75) );
  CLKIN1 U163 ( .A(B[23]), .Q(n141) );
  CLKIN2 U164 ( .A(B[16]), .Q(n172) );
  NAND21 U165 ( .A(B[16]), .B(n6), .Q(n47) );
  NOR21 U166 ( .A(B[4]), .B(n72), .Q(n124) );
  NAND22 U167 ( .A(A[22]), .B(n140), .Q(n139) );
  NOR21 U168 ( .A(n38), .B(n128), .Q(n118) );
  CLKIN3 U169 ( .A(n30), .Q(n27) );
  CLKIN3 U170 ( .A(n33), .Q(n32) );
  NAND24 U171 ( .A(n132), .B(n133), .Q(n40) );
  CLKIN3 U172 ( .A(n19), .Q(n157) );
  CLKIN3 U173 ( .A(n20), .Q(n156) );
  XNR22 U174 ( .A(B[30]), .B(A[30]), .Q(n162) );
endmodule


module D_compare ( o_con_ifbranch, i_data_rs, i_data_rt, i_con_bop );
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [2:0] i_con_bop;
  output o_con_ifbranch;
  wire   N32, N33, n4, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n1,
         n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n27;

  D_compare_DW01_cmp6_1 r49 ( .A(i_data_rs), .B(i_data_rt), .TC(n4), .EQ(N32), 
        .NE(N33) );
  NAND43 U2 ( .A(n19), .B(n22), .C(n21), .D(n20), .Q(n18) );
  NOR40 U3 ( .A(i_data_rs[9]), .B(i_data_rs[8]), .C(i_data_rs[7]), .D(
        i_data_rs[6]), .Q(n26) );
  NAND42 U4 ( .A(n23), .B(n24), .C(n25), .D(n26), .Q(n17) );
  NOR40 U5 ( .A(i_data_rs[26]), .B(i_data_rs[25]), .C(i_data_rs[24]), .D(
        i_data_rs[23]), .Q(n23) );
  NOR40 U6 ( .A(i_data_rs[2]), .B(i_data_rs[29]), .C(i_data_rs[28]), .D(
        i_data_rs[27]), .Q(n24) );
  NOR30 U7 ( .A(i_data_rs[0]), .B(i_data_rs[11]), .C(i_data_rs[10]), .Q(n19)
         );
  INV3 U8 ( .A(n3), .Q(n7) );
  NOR40 U9 ( .A(i_data_rs[15]), .B(i_data_rs[14]), .C(i_data_rs[13]), .D(
        i_data_rs[12]), .Q(n20) );
  NOR40 U10 ( .A(i_data_rs[5]), .B(i_data_rs[4]), .C(i_data_rs[3]), .D(
        i_data_rs[30]), .Q(n25) );
  NOR40 U11 ( .A(i_data_rs[19]), .B(i_data_rs[18]), .C(i_data_rs[17]), .D(
        i_data_rs[16]), .Q(n21) );
  NOR21 U12 ( .A(n3), .B(n9), .Q(n6) );
  LOGIC0 U13 ( .Q(n4) );
  NOR31 U14 ( .A(n2), .B(i_data_rs[1]), .C(i_data_rs[21]), .Q(n22) );
  OAI211 U15 ( .A(n18), .B(n17), .C(i_con_bop[0]), .Q(n5) );
  NOR21 U16 ( .A(i_data_rs[20]), .B(i_data_rs[22]), .Q(n1) );
  INV3 U17 ( .A(n1), .Q(n2) );
  BUF2 U18 ( .A(i_data_rs[31]), .Q(n3) );
  NOR24 U19 ( .A(i_con_bop[0]), .B(N33), .Q(n27) );
  OAI212 U20 ( .A(n3), .B(n5), .C(i_con_bop[1]), .Q(n16) );
  CLKIN3 U21 ( .A(i_con_bop[2]), .Q(n9) );
  OAI312 U22 ( .A(i_con_bop[1]), .B(n18), .C(n17), .D(n6), .Q(n13) );
  CLKIN3 U23 ( .A(i_con_bop[0]), .Q(n12) );
  NAND22 U24 ( .A(i_con_bop[0]), .B(n7), .Q(n10) );
  CLKIN3 U25 ( .A(i_con_bop[1]), .Q(n8) );
  OAI222 U26 ( .A(n10), .B(n9), .C(n12), .D(n8), .Q(n11) );
  AOI212 U27 ( .A(n13), .B(n12), .C(n11), .Q(n14) );
  OAI212 U28 ( .A(N32), .B(i_con_bop[2]), .C(n14), .Q(n15) );
  OAI312 U29 ( .A(n27), .B(i_con_bop[2]), .C(n16), .D(n15), .Q(o_con_ifbranch)
         );
endmodule


module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Efamux, i_con_Efbmux, 
        i_con_Ealuop, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread, 
        i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_bop, o_data_pc4, o_data_alures, o_data_rt, o_addr_regdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_addr_Erd, o_addr_Mrt, o_con_ifbranch );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [5:0] i_con_Ealuop;
  input [2:0] i_con_bop;
  output [31:0] o_data_pc4;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;
  wire   [31:0] alu_o_data_AluRes;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;

  DFC3 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[0]) );
  DFC3 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC3 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC3 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC3 pipe_rt_reg_28_ ( .D(compare_i_data_rt[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[28]) );
  DFC3 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC3 pipe_rt_reg_25_ ( .D(compare_i_data_rt[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[25]) );
  DFC3 pipe_rt_reg_23_ ( .D(compare_i_data_rt[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[23]) );
  DFC3 pipe_rt_reg_21_ ( .D(compare_i_data_rt[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[21]) );
  DFC3 pipe_rt_reg_20_ ( .D(compare_i_data_rt[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[20]) );
  DFC3 pipe_rt_reg_19_ ( .D(compare_i_data_rt[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[19]) );
  DFC3 pipe_rt_reg_18_ ( .D(compare_i_data_rt[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[18]) );
  DFC3 pipe_rt_reg_17_ ( .D(compare_i_data_rt[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[17]) );
  DFC3 pipe_rt_reg_16_ ( .D(compare_i_data_rt[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[16]) );
  DFC3 pipe_rt_reg_14_ ( .D(compare_i_data_rt[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[14]) );
  DFC3 pipe_rt_reg_13_ ( .D(compare_i_data_rt[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[13]) );
  DFC3 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC3 pipe_rt_reg_11_ ( .D(compare_i_data_rt[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[11]) );
  DFC3 pipe_rt_reg_9_ ( .D(compare_i_data_rt[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[9]) );
  DFC3 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC3 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC3 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC3 pipe_rt_reg_2_ ( .D(compare_i_data_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[2]) );
  DFC3 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC3 pipe_rt_reg_0_ ( .D(n5), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[0]) );
  DFC3 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC3 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Malupc8_reg ( .D(i_con_Malupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Malupc8) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  E_alu u_alu ( .o_data_AluRes(alu_o_data_AluRes), .i_data_A({
        compare_i_data_rs[31], n8, n4, n21, compare_i_data_rs[27:26], n20, 
        compare_i_data_rs[24], n17, compare_i_data_rs[22], n14, 
        compare_i_data_rs[20], n13, n7, compare_i_data_rs[17:16], n15, 
        compare_i_data_rs[14:13], n10, compare_i_data_rs[11:9], n22, 
        compare_i_data_rs[7], n12, compare_i_data_rs[5], n19, 
        compare_i_data_rs[3:0]}), .i_data_B(alu_i_data_B), .i_con_AluCtrl(
        alu_i_con_AluCtrl), .i_data_shamt(i_data_immext[10:6]) );
  E_alu_control u_alu_control ( .o_con_AluCtrl(alu_i_con_AluCtrl), 
        .i_con_AluOp(i_con_Ealuop), .i_con_FuncCode(i_data_immext[5:0]) );
  E_famux5 u_famux5 ( .i_data_rs(i_data_rs), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fa(i_con_Efamux), .o_data_alusra(
        compare_i_data_rs) );
  E_fbmux5 u_fbmux ( .i_data_rt(i_data_rt), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fb(i_con_Efbmux), .o_data_alusrb(
        compare_i_data_rt) );
  E_alubmux u_alubmux ( .i_data_fb(compare_i_data_rt), .i_data_imm(
        i_data_immext), .i_con_imm(i_con_Ealusrc), .o_data_alub(alu_i_data_B)
         );
  E_rdmux u_rdmux ( .i_data_rtE(i_addr_rt), .i_data_rdE(i_addr_rd), 
        .i_con_regdst(i_con_Eregdst), .i_con_aluPC4(i_con_Malupc8), 
        .o_data_writeE(o_addr_Erd) );
  D_compare u_compare ( .o_con_ifbranch(o_con_ifbranch), .i_data_rs({
        compare_i_data_rs[31], n8, compare_i_data_rs[29:20], n13, n7, 
        compare_i_data_rs[17:13], n10, compare_i_data_rs[11:7], n12, 
        compare_i_data_rs[5], n19, compare_i_data_rs[3:0]}), .i_data_rt({
        compare_i_data_rt[31:11], n2, compare_i_data_rt[9:1], n5}), 
        .i_con_bop(i_con_bop) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_rt_reg_10_ ( .D(n2), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_rt_reg_24_ ( .D(compare_i_data_rt[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[24]) );
  DFC1 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC1 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC1 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC1 pipe_rt_reg_5_ ( .D(compare_i_data_rt[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[5]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  DFC1 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC1 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC1 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC1 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC1 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC1 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC1 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC1 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC1 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC1 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC1 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC1 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC1 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC1 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC1 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC1 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC1 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC1 pipe_alures_reg_15_ ( .D(alu_o_data_AluRes[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[15]) );
  DFC1 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC1 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC1 pipe_alures_reg_14_ ( .D(alu_o_data_AluRes[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[14]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC3 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC1 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC1 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC3 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC1 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC1 pipe_rt_reg_15_ ( .D(compare_i_data_rt[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[15]) );
  DFC1 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC1 pipe_alures_reg_13_ ( .D(alu_o_data_AluRes[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[13]) );
  DFC1 pipe_rt_reg_22_ ( .D(n1), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC1 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC1 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  CLKBU12 U3 ( .A(compare_i_data_rs[30]), .Q(n8) );
  CLKBU12 U4 ( .A(compare_i_data_rs[25]), .Q(n20) );
  INV6 U5 ( .A(n11), .Q(n12) );
  INV12 U6 ( .A(n18), .Q(n19) );
  BUF2 U7 ( .A(compare_i_data_rt[22]), .Q(n1) );
  INV8 U8 ( .A(n16), .Q(n17) );
  CLKIN6 U9 ( .A(compare_i_data_rs[12]), .Q(n9) );
  INV3 U10 ( .A(compare_i_data_rs[23]), .Q(n16) );
  BUF8 U11 ( .A(compare_i_data_rs[28]), .Q(n21) );
  BUF8 U12 ( .A(compare_i_data_rs[8]), .Q(n22) );
  BUF12 U13 ( .A(compare_i_data_rs[19]), .Q(n13) );
  BUF2 U14 ( .A(compare_i_data_rt[0]), .Q(n5) );
  BUF12 U15 ( .A(compare_i_data_rs[21]), .Q(n14) );
  INV12 U16 ( .A(n9), .Q(n10) );
  BUF2 U17 ( .A(compare_i_data_rt[10]), .Q(n2) );
  INV3 U18 ( .A(compare_i_data_rs[29]), .Q(n3) );
  INV3 U19 ( .A(n3), .Q(n4) );
  INV6 U20 ( .A(compare_i_data_rs[6]), .Q(n11) );
  INV12 U21 ( .A(n6), .Q(n7) );
  INV6 U22 ( .A(compare_i_data_rs[18]), .Q(n6) );
  CLKIN6 U23 ( .A(compare_i_data_rs[4]), .Q(n18) );
  BUF6 U24 ( .A(compare_i_data_rs[15]), .Q(n15) );
endmodule


module M_resmux ( i_data_alures, i_data_pc8, i_con_pc8, o_data_alu );
  input [31:0] i_data_alures;
  input [31:0] i_data_pc8;
  output [31:0] o_data_alu;
  input i_con_pc8;
  wire   n34, n35, n36, n37, n38, n39, n40, n43, n54, n62, n63, n64, n65, n1;

  INV3 U1 ( .A(n34), .Q(o_data_alu[9]) );
  INV3 U2 ( .A(n62), .Q(o_data_alu[12]) );
  INV3 U3 ( .A(n40), .Q(o_data_alu[3]) );
  INV3 U4 ( .A(n38), .Q(o_data_alu[5]) );
  INV3 U5 ( .A(n36), .Q(o_data_alu[7]) );
  INV3 U6 ( .A(n64), .Q(o_data_alu[10]) );
  MUX22 U7 ( .A(i_data_alures[31]), .B(i_data_pc8[31]), .S(i_con_pc8), .Q(
        o_data_alu[31]) );
  AOI220 U8 ( .A(i_data_alures[11]), .B(n1), .C(i_data_pc8[11]), .D(i_con_pc8), 
        .Q(n63) );
  AOI220 U9 ( .A(i_data_alures[1]), .B(n1), .C(i_data_pc8[1]), .D(i_con_pc8), 
        .Q(n54) );
  AOI220 U10 ( .A(i_data_alures[9]), .B(n1), .C(i_data_pc8[9]), .D(i_con_pc8), 
        .Q(n34) );
  MUX21 U11 ( .A(i_data_alures[18]), .B(i_data_pc8[18]), .S(i_con_pc8), .Q(
        o_data_alu[18]) );
  MUX21 U12 ( .A(i_data_alures[13]), .B(i_data_pc8[13]), .S(i_con_pc8), .Q(
        o_data_alu[13]) );
  MUX21 U13 ( .A(i_data_alures[23]), .B(i_data_pc8[23]), .S(i_con_pc8), .Q(
        o_data_alu[23]) );
  MUX21 U14 ( .A(i_data_alures[24]), .B(i_data_pc8[24]), .S(i_con_pc8), .Q(
        o_data_alu[24]) );
  AOI220 U15 ( .A(i_data_alures[10]), .B(n1), .C(i_data_pc8[10]), .D(i_con_pc8), .Q(n64) );
  MUX21 U16 ( .A(i_data_alures[16]), .B(i_data_pc8[16]), .S(i_con_pc8), .Q(
        o_data_alu[16]) );
  AOI220 U17 ( .A(i_data_alures[2]), .B(n1), .C(i_data_pc8[2]), .D(i_con_pc8), 
        .Q(n43) );
  AOI220 U18 ( .A(i_data_alures[12]), .B(n1), .C(i_data_pc8[12]), .D(i_con_pc8), .Q(n62) );
  MUX21 U19 ( .A(i_data_alures[19]), .B(i_data_pc8[19]), .S(i_con_pc8), .Q(
        o_data_alu[19]) );
  MUX21 U20 ( .A(i_data_alures[30]), .B(i_data_pc8[30]), .S(i_con_pc8), .Q(
        o_data_alu[30]) );
  MUX21 U21 ( .A(i_data_alures[27]), .B(i_data_pc8[27]), .S(i_con_pc8), .Q(
        o_data_alu[27]) );
  MUX21 U22 ( .A(i_data_alures[15]), .B(i_data_pc8[15]), .S(i_con_pc8), .Q(
        o_data_alu[15]) );
  MUX21 U23 ( .A(i_data_alures[20]), .B(i_data_pc8[20]), .S(i_con_pc8), .Q(
        o_data_alu[20]) );
  AOI221 U24 ( .A(i_data_alures[7]), .B(n1), .C(i_data_pc8[7]), .D(i_con_pc8), 
        .Q(n36) );
  AOI220 U25 ( .A(i_data_alures[3]), .B(n1), .C(i_data_pc8[3]), .D(i_con_pc8), 
        .Q(n40) );
  AOI221 U26 ( .A(i_data_alures[5]), .B(n1), .C(i_data_pc8[5]), .D(i_con_pc8), 
        .Q(n38) );
  AOI220 U27 ( .A(i_data_alures[0]), .B(n1), .C(i_data_pc8[0]), .D(i_con_pc8), 
        .Q(n65) );
  AOI220 U28 ( .A(i_data_alures[4]), .B(n1), .C(i_data_pc8[4]), .D(i_con_pc8), 
        .Q(n39) );
  AOI220 U29 ( .A(i_data_alures[8]), .B(n1), .C(i_data_pc8[8]), .D(i_con_pc8), 
        .Q(n35) );
  MUX22 U30 ( .A(i_data_alures[14]), .B(i_data_pc8[14]), .S(i_con_pc8), .Q(
        o_data_alu[14]) );
  INV3 U31 ( .A(n63), .Q(o_data_alu[11]) );
  MUX22 U32 ( .A(i_data_alures[21]), .B(i_data_pc8[21]), .S(i_con_pc8), .Q(
        o_data_alu[21]) );
  MUX22 U33 ( .A(i_data_alures[22]), .B(i_data_pc8[22]), .S(i_con_pc8), .Q(
        o_data_alu[22]) );
  MUX22 U34 ( .A(i_data_alures[17]), .B(i_data_pc8[17]), .S(i_con_pc8), .Q(
        o_data_alu[17]) );
  MUX22 U35 ( .A(i_data_alures[25]), .B(i_data_pc8[25]), .S(i_con_pc8), .Q(
        o_data_alu[25]) );
  MUX22 U36 ( .A(i_data_alures[26]), .B(i_data_pc8[26]), .S(i_con_pc8), .Q(
        o_data_alu[26]) );
  MUX22 U37 ( .A(i_data_alures[29]), .B(i_data_pc8[29]), .S(i_con_pc8), .Q(
        o_data_alu[29]) );
  MUX22 U38 ( .A(i_data_alures[28]), .B(i_data_pc8[28]), .S(i_con_pc8), .Q(
        o_data_alu[28]) );
  INV3 U39 ( .A(n65), .Q(o_data_alu[0]) );
  INV3 U40 ( .A(n54), .Q(o_data_alu[1]) );
  INV3 U41 ( .A(n43), .Q(o_data_alu[2]) );
  INV3 U42 ( .A(n39), .Q(o_data_alu[4]) );
  INV3 U43 ( .A(n37), .Q(o_data_alu[6]) );
  AOI221 U44 ( .A(i_data_alures[6]), .B(n1), .C(i_data_pc8[6]), .D(i_con_pc8), 
        .Q(n37) );
  INV3 U45 ( .A(n35), .Q(o_data_alu[8]) );
  INV3 U46 ( .A(i_con_pc8), .Q(n1) );
endmodule


module mem_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  XNR21 U2 ( .A(n41), .B(n39), .Q(SUM[22]) );
  XNR21 U3 ( .A(n29), .B(n26), .Q(SUM[26]) );
  XNR21 U4 ( .A(A[29]), .B(n17), .Q(SUM[29]) );
  XNR21 U5 ( .A(n72), .B(n65), .Q(SUM[14]) );
  XNR21 U6 ( .A(n55), .B(n50), .Q(SUM[17]) );
  XNR21 U7 ( .A(n31), .B(n27), .Q(SUM[25]) );
  XOR21 U8 ( .A(n7), .B(n6), .Q(SUM[6]) );
  INV3 U9 ( .A(n5), .Q(n7) );
  INV3 U10 ( .A(n85), .Q(n3) );
  NAND22 U11 ( .A(n86), .B(n87), .Q(n85) );
  NOR21 U12 ( .A(SUM[2]), .B(n91), .Q(n86) );
  NOR21 U13 ( .A(n66), .B(n73), .Q(n72) );
  INV3 U14 ( .A(n57), .Q(n19) );
  NAND22 U15 ( .A(n58), .B(n59), .Q(n57) );
  NOR21 U16 ( .A(n61), .B(n62), .Q(n59) );
  NOR31 U17 ( .A(n67), .B(n68), .C(n69), .Q(n58) );
  NAND22 U18 ( .A(n63), .B(A[2]), .Q(n62) );
  NOR21 U19 ( .A(n65), .B(n66), .Q(n63) );
  INV3 U20 ( .A(n18), .Q(n16) );
  NAND22 U21 ( .A(n19), .B(n20), .Q(n18) );
  NOR21 U22 ( .A(n21), .B(n22), .Q(n20) );
  NAND22 U23 ( .A(n23), .B(n24), .Q(n21) );
  NOR21 U24 ( .A(n84), .B(n2), .Q(n83) );
  INV3 U25 ( .A(n54), .Q(n53) );
  NAND22 U26 ( .A(n55), .B(A[17]), .Q(n54) );
  INV3 U27 ( .A(n42), .Q(n41) );
  NAND22 U28 ( .A(n43), .B(A[21]), .Q(n42) );
  INV3 U29 ( .A(n30), .Q(n29) );
  NAND22 U30 ( .A(n31), .B(A[25]), .Q(n30) );
  NOR21 U31 ( .A(n8), .B(n10), .Q(n5) );
  NAND22 U32 ( .A(n76), .B(n3), .Q(n75) );
  INV3 U33 ( .A(n67), .Q(n76) );
  NAND22 U34 ( .A(n5), .B(A[6]), .Q(n4) );
  NOR21 U35 ( .A(n26), .B(n27), .Q(n23) );
  NAND22 U36 ( .A(n77), .B(n78), .Q(n67) );
  NOR21 U37 ( .A(n2), .B(n80), .Q(n77) );
  INV3 U38 ( .A(n79), .Q(n78) );
  NAND22 U39 ( .A(A[11]), .B(A[8]), .Q(n79) );
  NAND22 U40 ( .A(n35), .B(n36), .Q(n22) );
  NOR31 U41 ( .A(n39), .B(n37), .C(n38), .Q(n35) );
  NAND22 U42 ( .A(A[23]), .B(A[20]), .Q(n37) );
  NOR31 U43 ( .A(n68), .B(n85), .C(n67), .Q(n74) );
  NOR21 U44 ( .A(n57), .B(n56), .Q(n55) );
  INV3 U45 ( .A(A[16]), .Q(n56) );
  NOR21 U46 ( .A(n57), .B(n44), .Q(n43) );
  NAND22 U47 ( .A(A[20]), .B(n36), .Q(n44) );
  NOR21 U48 ( .A(n57), .B(n32), .Q(n31) );
  NAND22 U49 ( .A(A[24]), .B(n33), .Q(n32) );
  NAND22 U50 ( .A(n88), .B(n89), .Q(n61) );
  NOR21 U51 ( .A(n60), .B(n90), .Q(n88) );
  NOR21 U52 ( .A(n8), .B(n6), .Q(n89) );
  INV3 U53 ( .A(A[7]), .Q(n90) );
  INV3 U54 ( .A(A[14]), .Q(n65) );
  INV3 U55 ( .A(A[22]), .Q(n39) );
  INV3 U56 ( .A(A[13]), .Q(n66) );
  INV3 U57 ( .A(A[21]), .Q(n38) );
  INV3 U58 ( .A(A[5]), .Q(n8) );
  INV3 U59 ( .A(A[10]), .Q(n80) );
  INV3 U60 ( .A(A[18]), .Q(n51) );
  INV3 U61 ( .A(A[9]), .Q(n2) );
  INV3 U62 ( .A(A[17]), .Q(n50) );
  INV3 U63 ( .A(A[6]), .Q(n6) );
  NAND22 U64 ( .A(A[15]), .B(A[3]), .Q(n69) );
  NAND22 U65 ( .A(A[30]), .B(n14), .Q(n13) );
  XOR21 U66 ( .A(n70), .B(A[15]), .Q(SUM[15]) );
  NOR21 U67 ( .A(n65), .B(n71), .Q(n70) );
  XOR21 U68 ( .A(n40), .B(A[23]), .Q(SUM[23]) );
  NOR21 U69 ( .A(n39), .B(n42), .Q(n40) );
  XOR21 U70 ( .A(n81), .B(A[11]), .Q(SUM[11]) );
  NOR21 U71 ( .A(n80), .B(n82), .Q(n81) );
  INV3 U72 ( .A(n15), .Q(n14) );
  NAND31 U73 ( .A(A[28]), .B(n16), .C(A[29]), .Q(n15) );
  INV3 U74 ( .A(A[2]), .Q(SUM[2]) );
  INV3 U75 ( .A(n84), .Q(n1) );
  NAND22 U76 ( .A(A[8]), .B(n3), .Q(n84) );
  INV3 U77 ( .A(A[4]), .Q(n60) );
  INV3 U78 ( .A(A[12]), .Q(n68) );
  NAND22 U79 ( .A(n47), .B(n48), .Q(n45) );
  NOR21 U80 ( .A(n50), .B(n51), .Q(n47) );
  INV3 U81 ( .A(n49), .Q(n48) );
  NAND22 U82 ( .A(A[19]), .B(A[16]), .Q(n49) );
  INV3 U83 ( .A(n25), .Q(n24) );
  NAND22 U84 ( .A(A[27]), .B(A[24]), .Q(n25) );
  XOR21 U85 ( .A(n43), .B(A[21]), .Q(SUM[21]) );
  XOR21 U86 ( .A(n52), .B(A[19]), .Q(SUM[19]) );
  NOR21 U87 ( .A(n51), .B(n54), .Q(n52) );
  XOR21 U88 ( .A(n14), .B(A[30]), .Q(SUM[30]) );
  XOR21 U89 ( .A(n28), .B(A[27]), .Q(SUM[27]) );
  NOR21 U90 ( .A(n26), .B(n30), .Q(n28) );
  XNR21 U91 ( .A(n13), .B(A[31]), .Q(SUM[31]) );
  XNR21 U92 ( .A(n83), .B(n80), .Q(SUM[10]) );
  XOR21 U93 ( .A(n46), .B(A[20]), .Q(SUM[20]) );
  NOR21 U94 ( .A(n57), .B(n45), .Q(n46) );
  XOR21 U95 ( .A(n34), .B(A[24]), .Q(SUM[24]) );
  NOR21 U96 ( .A(n57), .B(n22), .Q(n34) );
  XOR21 U97 ( .A(n53), .B(A[18]), .Q(SUM[18]) );
  NAND22 U98 ( .A(A[28]), .B(n16), .Q(n17) );
  XNR21 U99 ( .A(n1), .B(n2), .Q(SUM[9]) );
  INV3 U100 ( .A(A[26]), .Q(n26) );
  INV3 U101 ( .A(A[25]), .Q(n27) );
  INV3 U102 ( .A(n12), .Q(n11) );
  NAND22 U103 ( .A(A[3]), .B(A[2]), .Q(n12) );
  INV3 U104 ( .A(n10), .Q(n9) );
  NAND22 U105 ( .A(A[4]), .B(n11), .Q(n10) );
  INV3 U106 ( .A(A[3]), .Q(n91) );
  XOR21 U107 ( .A(n16), .B(A[28]), .Q(SUM[28]) );
  XNR21 U108 ( .A(n9), .B(n8), .Q(SUM[5]) );
  XNR21 U109 ( .A(A[12]), .B(n75), .Q(SUM[12]) );
  XNR21 U110 ( .A(A[3]), .B(SUM[2]), .Q(SUM[3]) );
  XOR21 U111 ( .A(n11), .B(A[4]), .Q(SUM[4]) );
  XNR21 U112 ( .A(A[7]), .B(n4), .Q(SUM[7]) );
  XOR21 U113 ( .A(n3), .B(A[8]), .Q(SUM[8]) );
  XOR21 U114 ( .A(n74), .B(A[13]), .Q(SUM[13]) );
  XOR21 U115 ( .A(n19), .B(A[16]), .Q(SUM[16]) );
  CLKIN3 U116 ( .A(n22), .Q(n33) );
  CLKIN3 U117 ( .A(n45), .Q(n36) );
  CLKIN3 U118 ( .A(n72), .Q(n71) );
  CLKIN3 U119 ( .A(n74), .Q(n73) );
  CLKIN3 U120 ( .A(n83), .Q(n82) );
  CLKIN3 U121 ( .A(n61), .Q(n87) );
endmodule


module mem ( i_clk, i_nrst, i_data_pc4, i_data_alures, i_data_memout, 
        i_addr_regdst, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_FWmemread, i_addr_Mrt, o_data_alures, o_data_memout, 
        o_addr_regdst, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread, 
        o_addr_Wrt );
  input [31:0] i_data_pc4;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [4:0] i_addr_regdst;
  input [4:0] i_addr_Mrt;
  output [31:0] o_data_alures;
  output [31:0] o_data_memout;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Wrt;
  input i_clk, i_nrst, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite,
         i_con_FWmemread;
  output o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread;
  wire   n_Logic1_, n_Logic0_;
  wire   [31:0] pc8;
  wire   [31:0] resmux_o_data_alu;

  DFC3 pipe_rt_reg_4_ ( .D(i_addr_Mrt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(i_addr_Mrt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(i_addr_Mrt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[2]) );
  DFC3 pipe_rt_reg_1_ ( .D(i_addr_Mrt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[1]) );
  DFC3 pipe_rt_reg_0_ ( .D(i_addr_Mrt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[0]) );
  DFC3 pipe_data_alures_reg_31_ ( .D(resmux_o_data_alu[31]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[31]) );
  DFC3 pipe_data_alures_reg_30_ ( .D(resmux_o_data_alu[30]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[30]) );
  DFC3 pipe_data_alures_reg_29_ ( .D(resmux_o_data_alu[29]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[29]) );
  DFC3 pipe_data_alures_reg_28_ ( .D(resmux_o_data_alu[28]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[28]) );
  DFC3 pipe_data_alures_reg_27_ ( .D(resmux_o_data_alu[27]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[27]) );
  DFC3 pipe_data_alures_reg_26_ ( .D(resmux_o_data_alu[26]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[26]) );
  DFC3 pipe_data_alures_reg_25_ ( .D(resmux_o_data_alu[25]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[25]) );
  DFC3 pipe_data_alures_reg_24_ ( .D(resmux_o_data_alu[24]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[24]) );
  DFC3 pipe_data_alures_reg_23_ ( .D(resmux_o_data_alu[23]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[23]) );
  DFC3 pipe_data_alures_reg_22_ ( .D(resmux_o_data_alu[22]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[22]) );
  DFC3 pipe_data_alures_reg_21_ ( .D(resmux_o_data_alu[21]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[21]) );
  DFC3 pipe_data_alures_reg_20_ ( .D(resmux_o_data_alu[20]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[20]) );
  DFC3 pipe_data_alures_reg_19_ ( .D(resmux_o_data_alu[19]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[19]) );
  DFC3 pipe_data_alures_reg_18_ ( .D(resmux_o_data_alu[18]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[18]) );
  DFC3 pipe_data_alures_reg_17_ ( .D(resmux_o_data_alu[17]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[17]) );
  DFC3 pipe_data_alures_reg_16_ ( .D(resmux_o_data_alu[16]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[16]) );
  DFC3 pipe_data_alures_reg_15_ ( .D(resmux_o_data_alu[15]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[15]) );
  DFC3 pipe_data_alures_reg_14_ ( .D(resmux_o_data_alu[14]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[14]) );
  DFC3 pipe_data_alures_reg_13_ ( .D(resmux_o_data_alu[13]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[13]) );
  DFC3 pipe_data_alures_reg_12_ ( .D(resmux_o_data_alu[12]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[12]) );
  DFC3 pipe_data_alures_reg_11_ ( .D(resmux_o_data_alu[11]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[11]) );
  DFC3 pipe_data_alures_reg_10_ ( .D(resmux_o_data_alu[10]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[10]) );
  DFC3 pipe_data_alures_reg_9_ ( .D(resmux_o_data_alu[9]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[9]) );
  DFC3 pipe_data_alures_reg_8_ ( .D(resmux_o_data_alu[8]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[8]) );
  DFC3 pipe_data_alures_reg_7_ ( .D(resmux_o_data_alu[7]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[7]) );
  DFC3 pipe_data_alures_reg_6_ ( .D(resmux_o_data_alu[6]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[6]) );
  DFC3 pipe_data_alures_reg_5_ ( .D(resmux_o_data_alu[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[5]) );
  DFC3 pipe_data_alures_reg_4_ ( .D(resmux_o_data_alu[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[4]) );
  DFC3 pipe_data_alures_reg_3_ ( .D(resmux_o_data_alu[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[3]) );
  DFC3 pipe_data_alures_reg_2_ ( .D(resmux_o_data_alu[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[2]) );
  DFC3 pipe_data_alures_reg_1_ ( .D(resmux_o_data_alu[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[1]) );
  DFC3 pipe_data_alures_reg_0_ ( .D(resmux_o_data_alu[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[0]) );
  DFC3 pipe_data_memout_reg_31_ ( .D(i_data_memout[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[31]) );
  DFC3 pipe_data_memout_reg_30_ ( .D(i_data_memout[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[30]) );
  DFC3 pipe_data_memout_reg_29_ ( .D(i_data_memout[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[29]) );
  DFC3 pipe_data_memout_reg_28_ ( .D(i_data_memout[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[28]) );
  DFC3 pipe_data_memout_reg_27_ ( .D(i_data_memout[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[27]) );
  DFC3 pipe_data_memout_reg_26_ ( .D(i_data_memout[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[26]) );
  DFC3 pipe_data_memout_reg_25_ ( .D(i_data_memout[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[25]) );
  DFC3 pipe_data_memout_reg_24_ ( .D(i_data_memout[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[24]) );
  DFC3 pipe_data_memout_reg_23_ ( .D(i_data_memout[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[23]) );
  DFC3 pipe_data_memout_reg_22_ ( .D(i_data_memout[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[22]) );
  DFC3 pipe_data_memout_reg_21_ ( .D(i_data_memout[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[21]) );
  DFC3 pipe_data_memout_reg_20_ ( .D(i_data_memout[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[20]) );
  DFC3 pipe_data_memout_reg_19_ ( .D(i_data_memout[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[19]) );
  DFC3 pipe_data_memout_reg_18_ ( .D(i_data_memout[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[18]) );
  DFC3 pipe_data_memout_reg_17_ ( .D(i_data_memout[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[17]) );
  DFC3 pipe_data_memout_reg_16_ ( .D(i_data_memout[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[16]) );
  DFC3 pipe_data_memout_reg_15_ ( .D(i_data_memout[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[15]) );
  DFC3 pipe_data_memout_reg_14_ ( .D(i_data_memout[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[14]) );
  DFC3 pipe_data_memout_reg_13_ ( .D(i_data_memout[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[13]) );
  DFC3 pipe_data_memout_reg_12_ ( .D(i_data_memout[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[12]) );
  DFC3 pipe_data_memout_reg_11_ ( .D(i_data_memout[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[11]) );
  DFC3 pipe_data_memout_reg_10_ ( .D(i_data_memout[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[10]) );
  DFC3 pipe_data_memout_reg_9_ ( .D(i_data_memout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[9]) );
  DFC3 pipe_data_memout_reg_8_ ( .D(i_data_memout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[8]) );
  DFC3 pipe_data_memout_reg_7_ ( .D(i_data_memout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[7]) );
  DFC3 pipe_data_memout_reg_6_ ( .D(i_data_memout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[6]) );
  DFC3 pipe_data_memout_reg_5_ ( .D(i_data_memout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[5]) );
  DFC3 pipe_data_memout_reg_4_ ( .D(i_data_memout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[4]) );
  DFC3 pipe_data_memout_reg_3_ ( .D(i_data_memout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[3]) );
  DFC3 pipe_data_memout_reg_2_ ( .D(i_data_memout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[2]) );
  DFC3 pipe_data_memout_reg_1_ ( .D(i_data_memout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[1]) );
  DFC3 pipe_data_memout_reg_0_ ( .D(i_data_memout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[0]) );
  DFC3 pipe_addr_regdst_reg_4_ ( .D(i_addr_regdst[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[4]) );
  DFC3 pipe_addr_regdst_reg_3_ ( .D(i_addr_regdst[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[3]) );
  DFC3 pipe_addr_regdst_reg_2_ ( .D(i_addr_regdst[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[2]) );
  DFC3 pipe_addr_regdst_reg_1_ ( .D(i_addr_regdst[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[1]) );
  DFC3 pipe_addr_regdst_reg_0_ ( .D(i_addr_regdst[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[0]) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_con_FWmemread_reg ( .D(i_con_FWmemread), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_FWmemread) );
  M_resmux u_resmux ( .i_data_alures(i_data_alures), .i_data_pc8(pc8), 
        .i_con_pc8(i_con_Malupc8), .o_data_alu(resmux_o_data_alu) );
  mem_DW01_add_1 add_27 ( .A(i_data_pc4), .B({n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic1_, n_Logic0_, n_Logic0_}), .CI(n_Logic0_), .SUM(pc8) );
  LOGIC0 U3 ( .Q(n_Logic0_) );
  LOGIC1 U4 ( .Q(n_Logic1_) );
endmodule


module W_datamux ( i_data_alu, i_data_load, i_con_memtoreg, o_data_toreg );
  input [31:0] i_data_alu;
  input [31:0] i_data_load;
  output [31:0] o_data_toreg;
  input i_con_memtoreg;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n1;

  AOI220 U1 ( .A(i_data_alu[16]), .B(n1), .C(i_data_load[16]), .D(
        i_con_memtoreg), .Q(n58) );
  AOI220 U2 ( .A(i_data_alu[24]), .B(n1), .C(i_data_load[24]), .D(
        i_con_memtoreg), .Q(n49) );
  AOI220 U3 ( .A(i_data_alu[9]), .B(n1), .C(i_data_load[9]), .D(i_con_memtoreg), .Q(n34) );
  AOI220 U4 ( .A(i_data_alu[0]), .B(n1), .C(i_data_load[0]), .D(i_con_memtoreg), .Q(n65) );
  AOI220 U5 ( .A(i_data_alu[2]), .B(n1), .C(i_data_load[2]), .D(i_con_memtoreg), .Q(n43) );
  AOI220 U6 ( .A(i_data_alu[3]), .B(n1), .C(i_data_load[3]), .D(i_con_memtoreg), .Q(n40) );
  AOI220 U7 ( .A(i_data_alu[10]), .B(n1), .C(i_data_load[10]), .D(
        i_con_memtoreg), .Q(n64) );
  AOI220 U8 ( .A(i_data_alu[11]), .B(n1), .C(i_data_load[11]), .D(
        i_con_memtoreg), .Q(n63) );
  AOI220 U9 ( .A(i_data_alu[12]), .B(n1), .C(i_data_load[12]), .D(
        i_con_memtoreg), .Q(n62) );
  AOI220 U10 ( .A(i_data_alu[13]), .B(n1), .C(i_data_load[13]), .D(
        i_con_memtoreg), .Q(n61) );
  AOI220 U11 ( .A(i_data_alu[14]), .B(n1), .C(i_data_load[14]), .D(
        i_con_memtoreg), .Q(n60) );
  AOI220 U12 ( .A(i_data_alu[15]), .B(n1), .C(i_data_load[15]), .D(
        i_con_memtoreg), .Q(n59) );
  AOI220 U13 ( .A(i_data_alu[17]), .B(n1), .C(i_data_load[17]), .D(
        i_con_memtoreg), .Q(n57) );
  AOI220 U14 ( .A(i_data_alu[18]), .B(n1), .C(i_data_load[18]), .D(
        i_con_memtoreg), .Q(n56) );
  AOI220 U15 ( .A(i_data_alu[19]), .B(n1), .C(i_data_load[19]), .D(
        i_con_memtoreg), .Q(n55) );
  AOI220 U16 ( .A(i_data_alu[20]), .B(n1), .C(i_data_load[20]), .D(
        i_con_memtoreg), .Q(n53) );
  AOI220 U17 ( .A(i_data_alu[23]), .B(n1), .C(i_data_load[23]), .D(
        i_con_memtoreg), .Q(n50) );
  AOI220 U18 ( .A(i_data_alu[25]), .B(n1), .C(i_data_load[25]), .D(
        i_con_memtoreg), .Q(n48) );
  AOI220 U19 ( .A(i_data_alu[26]), .B(n1), .C(i_data_load[26]), .D(
        i_con_memtoreg), .Q(n47) );
  AOI220 U20 ( .A(i_data_alu[27]), .B(n1), .C(i_data_load[27]), .D(
        i_con_memtoreg), .Q(n46) );
  AOI220 U21 ( .A(i_data_alu[28]), .B(n1), .C(i_data_load[28]), .D(
        i_con_memtoreg), .Q(n45) );
  AOI220 U22 ( .A(i_data_alu[29]), .B(n1), .C(i_data_load[29]), .D(
        i_con_memtoreg), .Q(n44) );
  AOI220 U23 ( .A(i_data_alu[30]), .B(n1), .C(i_data_load[30]), .D(
        i_con_memtoreg), .Q(n42) );
  AOI220 U24 ( .A(i_data_alu[4]), .B(n1), .C(i_data_load[4]), .D(
        i_con_memtoreg), .Q(n39) );
  AOI220 U25 ( .A(i_data_alu[6]), .B(n1), .C(i_data_load[6]), .D(
        i_con_memtoreg), .Q(n37) );
  AOI220 U26 ( .A(i_data_alu[7]), .B(n1), .C(i_data_load[7]), .D(
        i_con_memtoreg), .Q(n36) );
  AOI220 U27 ( .A(i_data_alu[8]), .B(n1), .C(i_data_load[8]), .D(
        i_con_memtoreg), .Q(n35) );
  INV3 U28 ( .A(n54), .Q(o_data_toreg[1]) );
  AOI221 U29 ( .A(i_data_alu[1]), .B(n1), .C(i_data_load[1]), .D(
        i_con_memtoreg), .Q(n54) );
  INV3 U30 ( .A(n55), .Q(o_data_toreg[19]) );
  INV3 U31 ( .A(n65), .Q(o_data_toreg[0]) );
  INV3 U32 ( .A(n43), .Q(o_data_toreg[2]) );
  INV3 U33 ( .A(n40), .Q(o_data_toreg[3]) );
  INV3 U34 ( .A(n39), .Q(o_data_toreg[4]) );
  INV3 U35 ( .A(n38), .Q(o_data_toreg[5]) );
  AOI221 U36 ( .A(i_data_alu[5]), .B(n1), .C(i_data_load[5]), .D(
        i_con_memtoreg), .Q(n38) );
  INV3 U37 ( .A(n37), .Q(o_data_toreg[6]) );
  INV3 U38 ( .A(n36), .Q(o_data_toreg[7]) );
  INV3 U39 ( .A(n34), .Q(o_data_toreg[9]) );
  INV3 U40 ( .A(n64), .Q(o_data_toreg[10]) );
  INV3 U41 ( .A(n63), .Q(o_data_toreg[11]) );
  INV3 U42 ( .A(n62), .Q(o_data_toreg[12]) );
  INV3 U43 ( .A(n60), .Q(o_data_toreg[14]) );
  INV3 U44 ( .A(n59), .Q(o_data_toreg[15]) );
  INV3 U45 ( .A(n57), .Q(o_data_toreg[17]) );
  INV3 U46 ( .A(n56), .Q(o_data_toreg[18]) );
  INV3 U47 ( .A(n53), .Q(o_data_toreg[20]) );
  INV3 U48 ( .A(n52), .Q(o_data_toreg[21]) );
  AOI221 U49 ( .A(i_data_alu[21]), .B(n1), .C(i_data_load[21]), .D(
        i_con_memtoreg), .Q(n52) );
  INV3 U50 ( .A(n51), .Q(o_data_toreg[22]) );
  AOI221 U51 ( .A(i_data_alu[22]), .B(n1), .C(i_data_load[22]), .D(
        i_con_memtoreg), .Q(n51) );
  INV3 U52 ( .A(n49), .Q(o_data_toreg[24]) );
  INV3 U53 ( .A(n47), .Q(o_data_toreg[26]) );
  INV3 U54 ( .A(n44), .Q(o_data_toreg[29]) );
  INV3 U55 ( .A(n35), .Q(o_data_toreg[8]) );
  INV3 U56 ( .A(n61), .Q(o_data_toreg[13]) );
  INV3 U57 ( .A(n58), .Q(o_data_toreg[16]) );
  INV3 U58 ( .A(n50), .Q(o_data_toreg[23]) );
  INV3 U59 ( .A(n48), .Q(o_data_toreg[25]) );
  INV3 U60 ( .A(n46), .Q(o_data_toreg[27]) );
  INV3 U61 ( .A(n45), .Q(o_data_toreg[28]) );
  INV3 U62 ( .A(n41), .Q(o_data_toreg[31]) );
  AOI221 U63 ( .A(i_data_alu[31]), .B(n1), .C(i_data_load[31]), .D(
        i_con_memtoreg), .Q(n41) );
  INV3 U64 ( .A(n42), .Q(o_data_toreg[30]) );
  INV3 U65 ( .A(i_con_memtoreg), .Q(n1) );
endmodule


module writeback ( i_data_alures, i_data_memout, i_con_Wmemtoreg, 
        o_data_regwrite );
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  output [31:0] o_data_regwrite;
  input i_con_Wmemtoreg;


  W_datamux u_datamux ( .i_data_alu(i_data_alures), .i_data_load(i_data_memout), .i_con_memtoreg(i_con_Wmemtoreg), .o_data_toreg(o_data_regwrite) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Mmemread, ex_con_Mmemwrite, ex_con_Malupc8, ex_con_Wmemtoreg,
         mem_con_Malupc8, mem_con_Wmemtoreg, wb_con_Wmemtoreg, n1,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2;
  wire   [31:0] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [31:0] id_addr_pc4;
  wire   [31:0] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] wb_data_memout;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] mem_data_alures;
  wire   [31:0] mem_data_pc4;

  fetch u_fetch ( .i_clk(clk), .i_nrst(rst_n), .i_addr_b(if_addr_b), 
        .i_addr_j({if_addr_j, n1, n1}), .i_addr_jr(id_data_jr), .i_con_b(
        if_con_b), .i_con_j(if_con_j), .i_data_instr(read_instruction), 
        .i_con_ifstall(if_con_ifstall), .o_addr_pc(instruction_address), 
        .o_addr_pc4(id_addr_pc4), .o_data_instr(id_data_instr) );
  decode u_decode ( .i_clk(clk), .i_nrst(rst_n), .i_addr_pc4(id_addr_pc4), 
        .i_data_instr(id_data_instr), .i_con_Wregwrite(id_con_Wregwrite), 
        .i_data_Wregwrite(id_data_Wregwrite), .i_addr_Wregwrite(
        id_addr_Wregwrite), .i_addr_Erd(for_o_addr_Erd), .i_addr_Mrd(
        mem_addr_regdst), .i_con_Eregwrite(ex_con_Wregwrite), 
        .i_con_Mregwrite(mem_con_Wregwrite), .i_addr_rtM(for_addr_rtM), 
        .i_addr_rtW(for_addr_rtW), .i_con_memreadM(mem_read), .i_con_memreadW(
        for_FWmemread), .i_data_Wmemout(wb_data_memout), .o_data_rs(id_data_rs), .o_data_rt(ex_data_rt), .o_addr_rd(ex_addr_rd), .o_addr_rt(ex_addr_rt), 
        .o_data_jr(id_data_jr), .o_con_jump(if_con_j), .o_addr_pc4(ex_data_pc4), .o_addr_branch(if_addr_b), .o_addr_jump({if_addr_j, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .o_con_Ealuop(ex_con_Ealuop), 
        .o_con_Ealusrc(ex_con_Ealusrc), .o_con_Eregdst(ex_con_Eregdst), 
        .o_con_Mmemread(ex_con_Mmemread), .o_con_Mmemwrite(ex_con_Mmemwrite), 
        .o_con_Malupc8(ex_con_Malupc8), .o_con_Wmemtoreg(ex_con_Wmemtoreg), 
        .o_con_Wregwrite(ex_con_Wregwrite), .o_con_ifstall(if_con_ifstall), 
        .o_con_Ebop(ex_con_bop), .o_data_signext(ex_data_immext), 
        .o_con_Efamux(for_o_con_Efamux), .o_con_Efbmux(for_o_con_Efbmux), 
        .o_data_Fmemout(for_memout) );
  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext(
        ex_data_immext), .i_addr_rt(ex_addr_rt), .i_addr_rd(ex_addr_rd), 
        .i_data_FEalures(data_address), .i_data_FMalures(mem_data_alures), 
        .i_data_FMmemout(wb_data_memout), .i_data_FWmemout(for_memout), 
        .i_con_Efamux(for_o_con_Efamux), .i_con_Efbmux(for_o_con_Efbmux), 
        .i_con_Ealuop(ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), 
        .i_con_Mmemwrite(ex_con_Mmemwrite), .i_con_Malupc8(ex_con_Malupc8), 
        .i_con_Wmemtoreg(ex_con_Wmemtoreg), .i_con_Wregwrite(ex_con_Wregwrite), 
        .i_con_bop(ex_con_bop), .o_data_pc4(mem_data_pc4), .o_data_alures(
        data_address), .o_data_rt(write_data), .o_addr_regdst(mem_addr_regdst), 
        .o_con_Mmemread(mem_read), .o_con_Mmemwrite(mem_write), 
        .o_con_Malupc8(mem_con_Malupc8), .o_con_Wmemtoreg(mem_con_Wmemtoreg), 
        .o_con_Wregwrite(mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), 
        .o_addr_Mrt(for_addr_rtM), .o_con_ifbranch(if_con_b) );
  mem u_mem ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(mem_data_pc4), 
        .i_data_alures(data_address), .i_data_memout(read_data), 
        .i_addr_regdst(mem_addr_regdst), .i_con_Malupc8(mem_con_Malupc8), 
        .i_con_Wmemtoreg(mem_con_Wmemtoreg), .i_con_Wregwrite(
        mem_con_Wregwrite), .i_con_FWmemread(ex_con_Mmemread), .i_addr_Mrt(
        for_addr_rtM), .o_data_alures(mem_data_alures), .o_data_memout(
        wb_data_memout), .o_addr_regdst(id_addr_Wregwrite), .o_con_Wmemtoreg(
        wb_con_Wmemtoreg), .o_con_Wregwrite(id_con_Wregwrite), 
        .o_con_FWmemread(for_FWmemread), .o_addr_Wrt(for_addr_rtW) );
  writeback u_writeback ( .i_data_alures(mem_data_alures), .i_data_memout(
        wb_data_memout), .i_con_Wmemtoreg(wb_con_Wmemtoreg), .o_data_regwrite(
        id_data_Wregwrite) );
  LOGIC0 U1 ( .Q(n1) );
endmodule

