module W_imm_extend