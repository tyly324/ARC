
module F_jumpmux ( i_addr_j, i_addr_jr, i_addr_pc4, i_con_jump, o_addr_jumpmux
 );
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [31:0] i_addr_pc4;
  input [1:0] i_con_jump;
  output [31:0] o_addr_jumpmux;
  wire   n3, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n23,
         n24, n45, n46, n61, n62, n63, n64, n65, n66, n67, n68, n1, n2, n5, n6,
         n19, n20, n21, n22, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n69, n70, n71, n72,
         n73;

  BUF2 U1 ( .A(n72), .Q(n1) );
  BUF2 U2 ( .A(n72), .Q(n2) );
  INV3 U3 ( .A(n20), .Q(n71) );
  AOI221 U4 ( .A(i_addr_j[13]), .B(n73), .C(i_addr_pc4[13]), .D(n1), .Q(n22)
         );
  AOI221 U5 ( .A(i_addr_j[14]), .B(n73), .C(i_addr_pc4[14]), .D(n1), .Q(n26)
         );
  AOI221 U6 ( .A(i_addr_j[15]), .B(n73), .C(i_addr_pc4[15]), .D(n1), .Q(n28)
         );
  AOI221 U7 ( .A(i_addr_j[16]), .B(n73), .C(i_addr_pc4[16]), .D(n1), .Q(n30)
         );
  AOI221 U8 ( .A(i_addr_j[17]), .B(n73), .C(i_addr_pc4[17]), .D(n1), .Q(n32)
         );
  AOI221 U9 ( .A(i_addr_j[18]), .B(n73), .C(i_addr_pc4[18]), .D(n1), .Q(n34)
         );
  AOI221 U10 ( .A(i_addr_j[19]), .B(n73), .C(i_addr_pc4[19]), .D(n1), .Q(n36)
         );
  AOI221 U11 ( .A(i_addr_j[20]), .B(n73), .C(i_addr_pc4[20]), .D(n1), .Q(n38)
         );
  AOI221 U12 ( .A(i_addr_j[21]), .B(n73), .C(i_addr_pc4[21]), .D(n1), .Q(n40)
         );
  AOI221 U13 ( .A(i_addr_j[22]), .B(n73), .C(i_addr_pc4[22]), .D(n1), .Q(n42)
         );
  AOI221 U14 ( .A(i_addr_j[23]), .B(n73), .C(i_addr_pc4[23]), .D(n1), .Q(n44)
         );
  AOI221 U15 ( .A(i_addr_j[24]), .B(n73), .C(i_addr_pc4[24]), .D(n1), .Q(n48)
         );
  AOI221 U16 ( .A(i_addr_j[25]), .B(n73), .C(i_addr_pc4[25]), .D(n1), .Q(n50)
         );
  AOI221 U17 ( .A(i_addr_j[26]), .B(n73), .C(i_addr_pc4[26]), .D(n2), .Q(n52)
         );
  AOI221 U18 ( .A(i_addr_j[27]), .B(n73), .C(i_addr_pc4[27]), .D(n2), .Q(n54)
         );
  AOI221 U19 ( .A(i_addr_j[28]), .B(n73), .C(i_addr_pc4[28]), .D(n2), .Q(n56)
         );
  AOI221 U20 ( .A(i_addr_j[29]), .B(n73), .C(i_addr_pc4[29]), .D(n2), .Q(n58)
         );
  AOI221 U21 ( .A(i_addr_j[30]), .B(n73), .C(i_addr_pc4[30]), .D(n2), .Q(n60)
         );
  AOI221 U22 ( .A(i_addr_j[31]), .B(n73), .C(i_addr_pc4[31]), .D(n2), .Q(n70)
         );
  NAND22 U23 ( .A(n67), .B(n68), .Q(o_addr_jumpmux[0]) );
  NAND22 U24 ( .A(i_addr_j[0]), .B(n73), .Q(n68) );
  AOI221 U25 ( .A(i_addr_pc4[0]), .B(n2), .C(i_addr_jr[0]), .D(n71), .Q(n67)
         );
  NAND22 U26 ( .A(n45), .B(n46), .Q(o_addr_jumpmux[1]) );
  NAND22 U27 ( .A(i_addr_j[1]), .B(n73), .Q(n46) );
  AOI221 U28 ( .A(i_addr_pc4[1]), .B(n2), .C(i_addr_jr[1]), .D(n71), .Q(n45)
         );
  NAND22 U29 ( .A(n23), .B(n24), .Q(o_addr_jumpmux[2]) );
  NAND22 U30 ( .A(i_addr_j[2]), .B(n73), .Q(n24) );
  AOI221 U31 ( .A(i_addr_pc4[2]), .B(n2), .C(i_addr_jr[2]), .D(n71), .Q(n23)
         );
  NAND22 U32 ( .A(n17), .B(n18), .Q(o_addr_jumpmux[3]) );
  NAND22 U33 ( .A(i_addr_j[3]), .B(n73), .Q(n18) );
  AOI221 U34 ( .A(i_addr_pc4[3]), .B(n2), .C(i_addr_jr[3]), .D(n71), .Q(n17)
         );
  NAND22 U35 ( .A(n15), .B(n16), .Q(o_addr_jumpmux[4]) );
  NAND22 U36 ( .A(i_addr_j[4]), .B(n73), .Q(n16) );
  AOI221 U37 ( .A(i_addr_pc4[4]), .B(n1), .C(i_addr_jr[4]), .D(n71), .Q(n15)
         );
  NAND22 U38 ( .A(n13), .B(n14), .Q(o_addr_jumpmux[5]) );
  NAND22 U39 ( .A(i_addr_j[5]), .B(n73), .Q(n14) );
  AOI221 U40 ( .A(i_addr_pc4[5]), .B(n2), .C(i_addr_jr[5]), .D(n71), .Q(n13)
         );
  NAND22 U41 ( .A(n11), .B(n12), .Q(o_addr_jumpmux[6]) );
  NAND22 U42 ( .A(i_addr_j[6]), .B(n73), .Q(n12) );
  AOI221 U43 ( .A(i_addr_pc4[6]), .B(n72), .C(i_addr_jr[6]), .D(n71), .Q(n11)
         );
  NAND22 U44 ( .A(n9), .B(n10), .Q(o_addr_jumpmux[7]) );
  NAND22 U45 ( .A(i_addr_j[7]), .B(n73), .Q(n10) );
  AOI221 U46 ( .A(i_addr_pc4[7]), .B(n72), .C(i_addr_jr[7]), .D(n71), .Q(n9)
         );
  NAND22 U47 ( .A(n7), .B(n8), .Q(o_addr_jumpmux[8]) );
  NAND22 U48 ( .A(i_addr_j[8]), .B(n73), .Q(n8) );
  AOI221 U49 ( .A(i_addr_pc4[8]), .B(n72), .C(i_addr_jr[8]), .D(n71), .Q(n7)
         );
  NAND22 U50 ( .A(n3), .B(n4), .Q(o_addr_jumpmux[9]) );
  NAND22 U51 ( .A(i_addr_j[9]), .B(n73), .Q(n4) );
  AOI221 U52 ( .A(i_addr_pc4[9]), .B(n72), .C(i_addr_jr[9]), .D(n71), .Q(n3)
         );
  NAND22 U53 ( .A(n65), .B(n66), .Q(o_addr_jumpmux[10]) );
  NAND22 U54 ( .A(i_addr_j[10]), .B(n73), .Q(n66) );
  AOI221 U55 ( .A(i_addr_pc4[10]), .B(n2), .C(i_addr_jr[10]), .D(n71), .Q(n65)
         );
  NAND22 U56 ( .A(n63), .B(n64), .Q(o_addr_jumpmux[11]) );
  NAND22 U57 ( .A(i_addr_j[11]), .B(n73), .Q(n64) );
  AOI221 U58 ( .A(i_addr_pc4[11]), .B(n2), .C(i_addr_jr[11]), .D(n71), .Q(n63)
         );
  NAND22 U59 ( .A(n61), .B(n62), .Q(o_addr_jumpmux[12]) );
  NAND22 U60 ( .A(i_addr_j[12]), .B(n73), .Q(n62) );
  AOI221 U61 ( .A(i_addr_pc4[12]), .B(n2), .C(i_addr_jr[12]), .D(n71), .Q(n61)
         );
  CLKIN3 U62 ( .A(i_con_jump[1]), .Q(n5) );
  NAND22 U63 ( .A(i_con_jump[0]), .B(n5), .Q(n6) );
  CLKIN3 U64 ( .A(n6), .Q(n73) );
  XNR21 U65 ( .A(i_con_jump[0]), .B(i_con_jump[1]), .Q(n72) );
  CLKIN3 U66 ( .A(i_con_jump[0]), .Q(n19) );
  NAND22 U67 ( .A(i_con_jump[1]), .B(n19), .Q(n20) );
  NAND22 U68 ( .A(i_addr_jr[13]), .B(n71), .Q(n21) );
  NAND22 U69 ( .A(n22), .B(n21), .Q(o_addr_jumpmux[13]) );
  NAND22 U70 ( .A(i_addr_jr[14]), .B(n71), .Q(n25) );
  NAND22 U71 ( .A(n26), .B(n25), .Q(o_addr_jumpmux[14]) );
  NAND22 U72 ( .A(i_addr_jr[15]), .B(n71), .Q(n27) );
  NAND22 U73 ( .A(n28), .B(n27), .Q(o_addr_jumpmux[15]) );
  NAND22 U74 ( .A(i_addr_jr[16]), .B(n71), .Q(n29) );
  NAND22 U75 ( .A(n30), .B(n29), .Q(o_addr_jumpmux[16]) );
  NAND22 U76 ( .A(i_addr_jr[17]), .B(n71), .Q(n31) );
  NAND22 U77 ( .A(n32), .B(n31), .Q(o_addr_jumpmux[17]) );
  NAND22 U78 ( .A(i_addr_jr[18]), .B(n71), .Q(n33) );
  NAND22 U79 ( .A(n34), .B(n33), .Q(o_addr_jumpmux[18]) );
  NAND22 U80 ( .A(i_addr_jr[19]), .B(n71), .Q(n35) );
  NAND22 U81 ( .A(n36), .B(n35), .Q(o_addr_jumpmux[19]) );
  NAND22 U82 ( .A(i_addr_jr[20]), .B(n71), .Q(n37) );
  NAND22 U83 ( .A(n38), .B(n37), .Q(o_addr_jumpmux[20]) );
  NAND22 U84 ( .A(i_addr_jr[21]), .B(n71), .Q(n39) );
  NAND22 U85 ( .A(n40), .B(n39), .Q(o_addr_jumpmux[21]) );
  NAND22 U86 ( .A(i_addr_jr[22]), .B(n71), .Q(n41) );
  NAND22 U87 ( .A(n42), .B(n41), .Q(o_addr_jumpmux[22]) );
  NAND22 U88 ( .A(i_addr_jr[23]), .B(n71), .Q(n43) );
  NAND22 U89 ( .A(n44), .B(n43), .Q(o_addr_jumpmux[23]) );
  NAND22 U90 ( .A(i_addr_jr[24]), .B(n71), .Q(n47) );
  NAND22 U91 ( .A(n48), .B(n47), .Q(o_addr_jumpmux[24]) );
  NAND22 U92 ( .A(i_addr_jr[25]), .B(n71), .Q(n49) );
  NAND22 U93 ( .A(n50), .B(n49), .Q(o_addr_jumpmux[25]) );
  NAND22 U94 ( .A(i_addr_jr[26]), .B(n71), .Q(n51) );
  NAND22 U95 ( .A(n52), .B(n51), .Q(o_addr_jumpmux[26]) );
  NAND22 U96 ( .A(i_addr_jr[27]), .B(n71), .Q(n53) );
  NAND22 U97 ( .A(n54), .B(n53), .Q(o_addr_jumpmux[27]) );
  NAND22 U98 ( .A(i_addr_jr[28]), .B(n71), .Q(n55) );
  NAND22 U99 ( .A(n56), .B(n55), .Q(o_addr_jumpmux[28]) );
  NAND22 U100 ( .A(i_addr_jr[29]), .B(n71), .Q(n57) );
  NAND22 U101 ( .A(n58), .B(n57), .Q(o_addr_jumpmux[29]) );
  NAND22 U102 ( .A(i_addr_jr[30]), .B(n71), .Q(n59) );
  NAND22 U103 ( .A(n60), .B(n59), .Q(o_addr_jumpmux[30]) );
  NAND22 U104 ( .A(i_addr_jr[31]), .B(n71), .Q(n69) );
  NAND22 U105 ( .A(n70), .B(n69), .Q(o_addr_jumpmux[31]) );
endmodule


module F_branchmux ( i_addr_jumpmux, i_addr_b, i_con_ifbranch, o_addr_nextpc
 );
  input [31:0] i_addr_jumpmux;
  input [31:0] i_addr_b;
  output [31:0] o_addr_nextpc;
  input i_con_ifbranch;
  wire   n1, n2;

  CLKBU15 U1 ( .A(i_con_ifbranch), .Q(n1) );
  CLKBU15 U2 ( .A(i_con_ifbranch), .Q(n2) );
  MUX21 U3 ( .A(i_addr_jumpmux[0]), .B(i_addr_b[0]), .S(n2), .Q(
        o_addr_nextpc[0]) );
  MUX21 U4 ( .A(i_addr_jumpmux[2]), .B(i_addr_b[2]), .S(n1), .Q(
        o_addr_nextpc[2]) );
  MUX21 U5 ( .A(i_addr_jumpmux[4]), .B(i_addr_b[4]), .S(n2), .Q(
        o_addr_nextpc[4]) );
  MUX21 U6 ( .A(i_addr_jumpmux[6]), .B(i_addr_b[6]), .S(n2), .Q(
        o_addr_nextpc[6]) );
  MUX21 U7 ( .A(i_addr_jumpmux[8]), .B(i_addr_b[8]), .S(n1), .Q(
        o_addr_nextpc[8]) );
  MUX21 U8 ( .A(i_addr_jumpmux[10]), .B(i_addr_b[10]), .S(n2), .Q(
        o_addr_nextpc[10]) );
  MUX21 U9 ( .A(i_addr_jumpmux[12]), .B(i_addr_b[12]), .S(n1), .Q(
        o_addr_nextpc[12]) );
  MUX21 U10 ( .A(i_addr_jumpmux[14]), .B(i_addr_b[14]), .S(n1), .Q(
        o_addr_nextpc[14]) );
  MUX21 U11 ( .A(i_addr_jumpmux[15]), .B(i_addr_b[15]), .S(n1), .Q(
        o_addr_nextpc[15]) );
  MUX21 U12 ( .A(i_addr_jumpmux[16]), .B(i_addr_b[16]), .S(n2), .Q(
        o_addr_nextpc[16]) );
  MUX21 U13 ( .A(i_addr_jumpmux[17]), .B(i_addr_b[17]), .S(n1), .Q(
        o_addr_nextpc[17]) );
  MUX21 U14 ( .A(i_addr_jumpmux[18]), .B(i_addr_b[18]), .S(n2), .Q(
        o_addr_nextpc[18]) );
  MUX21 U15 ( .A(i_addr_jumpmux[19]), .B(i_addr_b[19]), .S(n1), .Q(
        o_addr_nextpc[19]) );
  MUX21 U16 ( .A(i_addr_jumpmux[20]), .B(i_addr_b[20]), .S(n2), .Q(
        o_addr_nextpc[20]) );
  MUX21 U17 ( .A(i_addr_jumpmux[21]), .B(i_addr_b[21]), .S(n1), .Q(
        o_addr_nextpc[21]) );
  MUX21 U18 ( .A(i_addr_jumpmux[22]), .B(i_addr_b[22]), .S(n2), .Q(
        o_addr_nextpc[22]) );
  MUX21 U19 ( .A(i_addr_jumpmux[23]), .B(i_addr_b[23]), .S(n1), .Q(
        o_addr_nextpc[23]) );
  MUX21 U20 ( .A(i_addr_jumpmux[24]), .B(i_addr_b[24]), .S(n2), .Q(
        o_addr_nextpc[24]) );
  MUX21 U21 ( .A(i_addr_jumpmux[25]), .B(i_addr_b[25]), .S(n1), .Q(
        o_addr_nextpc[25]) );
  MUX21 U22 ( .A(i_addr_jumpmux[26]), .B(i_addr_b[26]), .S(n2), .Q(
        o_addr_nextpc[26]) );
  MUX21 U23 ( .A(i_addr_jumpmux[28]), .B(i_addr_b[28]), .S(n1), .Q(
        o_addr_nextpc[28]) );
  MUX21 U24 ( .A(i_addr_jumpmux[30]), .B(i_addr_b[30]), .S(n2), .Q(
        o_addr_nextpc[30]) );
  MUX21 U25 ( .A(i_addr_jumpmux[1]), .B(i_addr_b[1]), .S(n2), .Q(
        o_addr_nextpc[1]) );
  MUX21 U26 ( .A(i_addr_jumpmux[3]), .B(i_addr_b[3]), .S(n1), .Q(
        o_addr_nextpc[3]) );
  MUX21 U27 ( .A(i_addr_jumpmux[5]), .B(i_addr_b[5]), .S(n2), .Q(
        o_addr_nextpc[5]) );
  MUX21 U28 ( .A(i_addr_jumpmux[7]), .B(i_addr_b[7]), .S(n1), .Q(
        o_addr_nextpc[7]) );
  MUX21 U29 ( .A(i_addr_jumpmux[9]), .B(i_addr_b[9]), .S(n1), .Q(
        o_addr_nextpc[9]) );
  MUX21 U30 ( .A(i_addr_jumpmux[11]), .B(i_addr_b[11]), .S(n2), .Q(
        o_addr_nextpc[11]) );
  MUX21 U31 ( .A(i_addr_jumpmux[13]), .B(i_addr_b[13]), .S(n1), .Q(
        o_addr_nextpc[13]) );
  MUX21 U32 ( .A(i_addr_jumpmux[27]), .B(i_addr_b[27]), .S(n2), .Q(
        o_addr_nextpc[27]) );
  MUX21 U33 ( .A(i_addr_jumpmux[29]), .B(i_addr_b[29]), .S(n2), .Q(
        o_addr_nextpc[29]) );
  MUX21 U34 ( .A(i_addr_jumpmux[31]), .B(i_addr_b[31]), .S(n1), .Q(
        o_addr_nextpc[31]) );
endmodule


module F_pc ( i_clk, i_rst_n, i_con_stall, i_addr_next_pc, o_addr_pc );
  input [31:0] i_addr_next_pc;
  output [31:0] o_addr_pc;
  input i_clk, i_rst_n, i_con_stall;


  DFEC1 program_counter_reg_31_ ( .D(i_addr_next_pc[31]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[31]) );
  DFEC1 program_counter_reg_1_ ( .D(i_addr_next_pc[1]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[1]) );
  DFEC1 program_counter_reg_0_ ( .D(i_addr_next_pc[0]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[0]) );
  DFEC1 program_counter_reg_30_ ( .D(i_addr_next_pc[30]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[30]) );
  DFEC1 program_counter_reg_26_ ( .D(i_addr_next_pc[26]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[26]) );
  DFEC1 program_counter_reg_25_ ( .D(i_addr_next_pc[25]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[25]) );
  DFEC1 program_counter_reg_22_ ( .D(i_addr_next_pc[22]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[22]) );
  DFEC1 program_counter_reg_21_ ( .D(i_addr_next_pc[21]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[21]) );
  DFEC1 program_counter_reg_17_ ( .D(i_addr_next_pc[17]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[17]) );
  DFEC1 program_counter_reg_27_ ( .D(i_addr_next_pc[27]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[27]) );
  DFEC1 program_counter_reg_23_ ( .D(i_addr_next_pc[23]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[23]) );
  DFEC1 program_counter_reg_29_ ( .D(i_addr_next_pc[29]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[29]) );
  DFEC1 program_counter_reg_28_ ( .D(i_addr_next_pc[28]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[28]) );
  DFEC1 program_counter_reg_24_ ( .D(i_addr_next_pc[24]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[24]) );
  DFEC1 program_counter_reg_18_ ( .D(i_addr_next_pc[18]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[18]) );
  DFEC1 program_counter_reg_14_ ( .D(i_addr_next_pc[14]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[14]) );
  DFEC1 program_counter_reg_13_ ( .D(i_addr_next_pc[13]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[13]) );
  DFEC1 program_counter_reg_10_ ( .D(i_addr_next_pc[10]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[10]) );
  DFEC1 program_counter_reg_9_ ( .D(i_addr_next_pc[9]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[9]) );
  DFEC1 program_counter_reg_6_ ( .D(i_addr_next_pc[6]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[6]) );
  DFEC1 program_counter_reg_5_ ( .D(i_addr_next_pc[5]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[5]) );
  DFEC1 program_counter_reg_2_ ( .D(i_addr_next_pc[2]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[2]) );
  DFEC1 program_counter_reg_15_ ( .D(i_addr_next_pc[15]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[15]) );
  DFEC1 program_counter_reg_19_ ( .D(i_addr_next_pc[19]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[19]) );
  DFEC1 program_counter_reg_7_ ( .D(i_addr_next_pc[7]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[7]) );
  DFEC1 program_counter_reg_11_ ( .D(i_addr_next_pc[11]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[11]) );
  DFEC1 program_counter_reg_12_ ( .D(i_addr_next_pc[12]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[12]) );
  DFEC1 program_counter_reg_16_ ( .D(i_addr_next_pc[16]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[16]) );
  DFEC1 program_counter_reg_20_ ( .D(i_addr_next_pc[20]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[20]) );
  DFEC1 program_counter_reg_8_ ( .D(i_addr_next_pc[8]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[8]) );
  DFEC1 program_counter_reg_4_ ( .D(i_addr_next_pc[4]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[4]) );
  DFEC1 program_counter_reg_3_ ( .D(i_addr_next_pc[3]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[3]) );
endmodule


module F_add4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  XNR21 U2 ( .A(n48), .B(n42), .Q(SUM[21]) );
  XNR21 U3 ( .A(n34), .B(n28), .Q(SUM[25]) );
  XNR21 U4 ( .A(n71), .B(n68), .Q(SUM[14]) );
  XNR21 U5 ( .A(n57), .B(n54), .Q(SUM[18]) );
  XNR21 U6 ( .A(n46), .B(n43), .Q(SUM[22]) );
  XNR21 U7 ( .A(n32), .B(n29), .Q(SUM[26]) );
  INV3 U8 ( .A(n61), .Q(n23) );
  NAND41 U9 ( .A(n62), .B(n63), .C(n64), .D(n65), .Q(n61) );
  NOR21 U10 ( .A(n67), .B(n68), .Q(n62) );
  NOR21 U11 ( .A(n66), .B(SUM[2]), .Q(n64) );
  NOR21 U12 ( .A(n82), .B(n2), .Q(n81) );
  INV3 U13 ( .A(n21), .Q(n17) );
  NAND22 U14 ( .A(n22), .B(n23), .Q(n21) );
  NOR21 U15 ( .A(n24), .B(n25), .Q(n22) );
  INV3 U16 ( .A(n51), .Q(n50) );
  NAND22 U17 ( .A(n40), .B(n23), .Q(n51) );
  INV3 U18 ( .A(n37), .Q(n36) );
  NAND22 U19 ( .A(n38), .B(n23), .Q(n37) );
  INV3 U20 ( .A(n76), .Q(n75) );
  NAND22 U21 ( .A(n65), .B(n3), .Q(n76) );
  INV3 U22 ( .A(n47), .Q(n46) );
  NAND22 U23 ( .A(n48), .B(A[21]), .Q(n47) );
  INV3 U24 ( .A(n33), .Q(n32) );
  NAND22 U25 ( .A(n34), .B(A[25]), .Q(n33) );
  INV3 U26 ( .A(n58), .Q(n57) );
  NAND22 U27 ( .A(n59), .B(A[17]), .Q(n58) );
  INV3 U28 ( .A(n72), .Q(n71) );
  NAND22 U29 ( .A(n73), .B(A[13]), .Q(n72) );
  XNR21 U30 ( .A(n73), .B(n67), .Q(SUM[13]) );
  XNR21 U31 ( .A(n59), .B(n53), .Q(SUM[17]) );
  XNR21 U32 ( .A(n81), .B(n78), .Q(SUM[10]) );
  XNR21 U33 ( .A(n9), .B(n8), .Q(SUM[5]) );
  XNR21 U34 ( .A(n1), .B(n2), .Q(SUM[9]) );
  NOR21 U35 ( .A(n8), .B(n10), .Q(n6) );
  XNR21 U36 ( .A(n6), .B(n7), .Q(SUM[6]) );
  NAND31 U37 ( .A(A[15]), .B(A[12]), .C(A[3]), .Q(n66) );
  XOR21 U38 ( .A(n15), .B(A[30]), .Q(SUM[30]) );
  XOR21 U39 ( .A(n19), .B(n20), .Q(SUM[29]) );
  INV3 U40 ( .A(A[29]), .Q(n19) );
  NAND22 U41 ( .A(A[28]), .B(n17), .Q(n20) );
  XOR21 U42 ( .A(n69), .B(n70), .Q(SUM[15]) );
  INV3 U43 ( .A(A[15]), .Q(n69) );
  NAND22 U44 ( .A(n71), .B(A[14]), .Q(n70) );
  XOR21 U45 ( .A(n55), .B(n56), .Q(SUM[19]) );
  INV3 U46 ( .A(A[19]), .Q(n55) );
  NAND22 U47 ( .A(n57), .B(A[18]), .Q(n56) );
  XOR21 U48 ( .A(n44), .B(n45), .Q(SUM[23]) );
  INV3 U49 ( .A(A[23]), .Q(n44) );
  NAND22 U50 ( .A(n46), .B(A[22]), .Q(n45) );
  XOR21 U51 ( .A(n30), .B(n31), .Q(SUM[27]) );
  INV3 U52 ( .A(A[27]), .Q(n30) );
  NAND22 U53 ( .A(n32), .B(A[26]), .Q(n31) );
  XOR21 U54 ( .A(n13), .B(n14), .Q(SUM[31]) );
  INV3 U55 ( .A(A[31]), .Q(n13) );
  NAND22 U56 ( .A(A[30]), .B(n15), .Q(n14) );
  NOR31 U57 ( .A(n54), .B(n52), .C(n53), .Q(n40) );
  NAND22 U58 ( .A(A[19]), .B(A[16]), .Q(n52) );
  NOR31 U59 ( .A(n78), .B(n77), .C(n2), .Q(n65) );
  NAND22 U60 ( .A(A[11]), .B(A[8]), .Q(n77) );
  NAND22 U61 ( .A(n39), .B(n40), .Q(n24) );
  NOR31 U62 ( .A(n43), .B(n41), .C(n42), .Q(n39) );
  NAND22 U63 ( .A(A[23]), .B(A[20]), .Q(n41) );
  INV3 U64 ( .A(A[5]), .Q(n8) );
  INV3 U65 ( .A(A[10]), .Q(n78) );
  INV3 U66 ( .A(A[9]), .Q(n2) );
  INV3 U67 ( .A(A[18]), .Q(n54) );
  INV3 U68 ( .A(A[6]), .Q(n7) );
  INV3 U69 ( .A(n83), .Q(n3) );
  NAND22 U70 ( .A(n84), .B(n63), .Q(n83) );
  NOR21 U71 ( .A(n88), .B(SUM[2]), .Q(n84) );
  INV3 U72 ( .A(A[3]), .Q(n88) );
  INV3 U73 ( .A(A[13]), .Q(n67) );
  INV3 U74 ( .A(A[14]), .Q(n68) );
  INV3 U75 ( .A(A[2]), .Q(SUM[2]) );
  XOR21 U76 ( .A(n79), .B(A[11]), .Q(SUM[11]) );
  NOR21 U77 ( .A(n78), .B(n80), .Q(n79) );
  INV3 U78 ( .A(n16), .Q(n15) );
  NAND31 U79 ( .A(A[28]), .B(n17), .C(A[29]), .Q(n16) );
  INV3 U80 ( .A(n49), .Q(n48) );
  NAND22 U81 ( .A(A[20]), .B(n50), .Q(n49) );
  INV3 U82 ( .A(n35), .Q(n34) );
  NAND22 U83 ( .A(A[24]), .B(n36), .Q(n35) );
  INV3 U84 ( .A(n60), .Q(n59) );
  NAND22 U85 ( .A(A[16]), .B(n23), .Q(n60) );
  INV3 U86 ( .A(n74), .Q(n73) );
  NAND22 U87 ( .A(A[12]), .B(n75), .Q(n74) );
  INV3 U88 ( .A(n82), .Q(n1) );
  NAND22 U89 ( .A(A[8]), .B(n3), .Q(n82) );
  NOR21 U90 ( .A(n85), .B(n86), .Q(n63) );
  NAND22 U91 ( .A(A[7]), .B(A[4]), .Q(n86) );
  INV3 U92 ( .A(n87), .Q(n85) );
  NOR21 U93 ( .A(n8), .B(n7), .Q(n87) );
  XOR21 U94 ( .A(n17), .B(A[28]), .Q(SUM[28]) );
  XOR21 U95 ( .A(n50), .B(A[20]), .Q(SUM[20]) );
  XOR21 U96 ( .A(n36), .B(A[24]), .Q(SUM[24]) );
  XOR21 U97 ( .A(A[16]), .B(n23), .Q(SUM[16]) );
  XOR21 U98 ( .A(n3), .B(A[8]), .Q(SUM[8]) );
  XOR21 U99 ( .A(n11), .B(A[4]), .Q(SUM[4]) );
  XOR21 U100 ( .A(n75), .B(A[12]), .Q(SUM[12]) );
  XOR21 U101 ( .A(A[3]), .B(A[2]), .Q(SUM[3]) );
  XOR21 U102 ( .A(n4), .B(n5), .Q(SUM[7]) );
  INV3 U103 ( .A(A[7]), .Q(n4) );
  NAND22 U104 ( .A(n6), .B(A[6]), .Q(n5) );
  INV3 U105 ( .A(A[22]), .Q(n43) );
  INV3 U106 ( .A(A[26]), .Q(n29) );
  INV3 U107 ( .A(A[17]), .Q(n53) );
  INV3 U108 ( .A(A[21]), .Q(n42) );
  INV3 U109 ( .A(A[25]), .Q(n28) );
  NOR31 U110 ( .A(n29), .B(n27), .C(n28), .Q(n26) );
  NAND22 U111 ( .A(A[27]), .B(A[24]), .Q(n27) );
  INV3 U112 ( .A(n12), .Q(n11) );
  NAND22 U113 ( .A(A[3]), .B(A[2]), .Q(n12) );
  INV3 U114 ( .A(n10), .Q(n9) );
  NAND22 U115 ( .A(A[4]), .B(n11), .Q(n10) );
  CLKIN3 U116 ( .A(n26), .Q(n25) );
  CLKIN3 U117 ( .A(n24), .Q(n38) );
  CLKIN3 U118 ( .A(n81), .Q(n80) );
endmodule


module F_add4 ( i_addr_pc, o_addr_pcadd4 );
  input [31:0] i_addr_pc;
  output [31:0] o_addr_pcadd4;
  wire   n2, n1;

  F_add4_DW01_add_1 add_5 ( .A(i_addr_pc), .B({n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n2, n1, n1}), .CI(n1), .SUM(o_addr_pcadd4) );
  LOGIC0 U3 ( .Q(n1) );
  LOGIC1 U4 ( .Q(n2) );
endmodule


module fetch ( i_clk, i_nrst, i_addr_b, i_addr_j, i_addr_jr, i_con_b, i_con_j, 
        i_data_instr, i_con_ifstall, o_addr_pc, o_addr_pc4, o_data_instr );
  input [31:0] i_addr_b;
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [1:0] i_con_j;
  input [31:0] i_data_instr;
  output [31:0] o_addr_pc;
  output [31:0] o_addr_pc4;
  output [31:0] o_data_instr;
  input i_clk, i_nrst, i_con_b, i_con_ifstall;

  wire   [31:0] jmux_i_addr_pc4;
  wire   [31:0] bmux_i_addr_jumpmux;
  wire   [31:0] pc_i_addr_next_pc;

  DFC3 pipe_instr_reg_31_ ( .D(i_data_instr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[31]) );
  DFC3 pipe_instr_reg_30_ ( .D(i_data_instr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[30]) );
  DFC3 pipe_instr_reg_29_ ( .D(i_data_instr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[29]) );
  DFC3 pipe_instr_reg_28_ ( .D(i_data_instr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[28]) );
  DFC3 pipe_instr_reg_27_ ( .D(i_data_instr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[27]) );
  DFC3 pipe_instr_reg_26_ ( .D(i_data_instr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[26]) );
  DFC3 pipe_instr_reg_25_ ( .D(i_data_instr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[25]) );
  DFC3 pipe_instr_reg_24_ ( .D(i_data_instr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[24]) );
  DFC3 pipe_instr_reg_23_ ( .D(i_data_instr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[23]) );
  DFC3 pipe_instr_reg_22_ ( .D(i_data_instr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[22]) );
  DFC3 pipe_instr_reg_21_ ( .D(i_data_instr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[21]) );
  DFC3 pipe_instr_reg_20_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[20]) );
  DFC3 pipe_instr_reg_19_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[19]) );
  DFC3 pipe_instr_reg_18_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[18]) );
  DFC3 pipe_instr_reg_17_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[17]) );
  DFC3 pipe_instr_reg_16_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[16]) );
  DFC3 pipe_instr_reg_15_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[15]) );
  DFC3 pipe_instr_reg_14_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[14]) );
  DFC3 pipe_instr_reg_13_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[13]) );
  DFC3 pipe_instr_reg_12_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[12]) );
  DFC3 pipe_instr_reg_11_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[11]) );
  DFC3 pipe_instr_reg_10_ ( .D(i_data_instr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[10]) );
  DFC3 pipe_instr_reg_9_ ( .D(i_data_instr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[9]) );
  DFC3 pipe_instr_reg_8_ ( .D(i_data_instr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[8]) );
  DFC3 pipe_instr_reg_7_ ( .D(i_data_instr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[7]) );
  DFC3 pipe_instr_reg_6_ ( .D(i_data_instr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[6]) );
  DFC3 pipe_instr_reg_5_ ( .D(i_data_instr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[5]) );
  DFC3 pipe_instr_reg_4_ ( .D(i_data_instr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[4]) );
  DFC3 pipe_instr_reg_3_ ( .D(i_data_instr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[3]) );
  DFC3 pipe_instr_reg_2_ ( .D(i_data_instr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[2]) );
  DFC3 pipe_instr_reg_1_ ( .D(i_data_instr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[1]) );
  DFC3 pipe_instr_reg_0_ ( .D(i_data_instr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(jmux_i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(jmux_i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(jmux_i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(jmux_i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(jmux_i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(jmux_i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(jmux_i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(jmux_i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(jmux_i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(jmux_i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(jmux_i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(jmux_i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(jmux_i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(jmux_i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(jmux_i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(jmux_i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(jmux_i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(jmux_i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(jmux_i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(jmux_i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(jmux_i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(jmux_i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(jmux_i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(jmux_i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(jmux_i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(jmux_i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(jmux_i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(jmux_i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(jmux_i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(jmux_i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(jmux_i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(jmux_i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  F_jumpmux u_jumpmux ( .i_addr_j(i_addr_j), .i_addr_jr(i_addr_jr), 
        .i_addr_pc4(jmux_i_addr_pc4), .i_con_jump(i_con_j), .o_addr_jumpmux(
        bmux_i_addr_jumpmux) );
  F_branchmux u_branchmux ( .i_addr_jumpmux(bmux_i_addr_jumpmux), .i_addr_b(
        i_addr_b), .i_con_ifbranch(i_con_b), .o_addr_nextpc(pc_i_addr_next_pc)
         );
  F_pc u_pc ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_con_stall(i_con_ifstall), 
        .i_addr_next_pc(pc_i_addr_next_pc), .o_addr_pc(o_addr_pc) );
  F_add4 u_add4 ( .i_addr_pc(o_addr_pc), .o_addr_pcadd4(jmux_i_addr_pc4) );
endmodule


module D_control ( o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite, 
        o_con_alusrc, o_con_regwrite, o_con_ifsign, o_con_aluop, i_con_instru
 );
  output [5:0] o_con_aluop;
  input [5:0] i_con_instru;
  output o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite,
         o_con_alusrc, o_con_regwrite, o_con_ifsign;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n1, n2, n3, n5, n6, n7, n8, n9, n10;

  OAI212 U2 ( .A(i_con_instru[3]), .B(n11), .C(n12), .Q(o_con_regwrite) );
  OAI212 U3 ( .A(n5), .B(n13), .C(n3), .Q(n12) );
  OAI222 U6 ( .A(i_con_instru[3]), .B(n15), .C(i_con_instru[4]), .D(n17), .Q(
        o_con_memread) );
  OAI212 U23 ( .A(i_con_instru[5]), .B(n20), .C(n14), .Q(o_con_aluop[1]) );
  NAND31 U4 ( .A(n24), .B(n3), .C(n13), .Q(n14) );
  NAND22 U5 ( .A(n9), .B(n13), .Q(n11) );
  AOI211 U7 ( .A(n5), .B(n8), .C(o_con_memwrite), .Q(n18) );
  INV3 U8 ( .A(n20), .Q(n5) );
  INV3 U9 ( .A(n24), .Q(n9) );
  NAND22 U10 ( .A(n20), .B(n15), .Q(o_con_alusrc) );
  NAND22 U11 ( .A(n15), .B(n16), .Q(o_con_memtoreg) );
  NOR21 U12 ( .A(n11), .B(n21), .Q(o_con_aluop[5]) );
  INV3 U13 ( .A(n16), .Q(o_con_memwrite) );
  INV3 U14 ( .A(n21), .Q(n2) );
  NOR31 U15 ( .A(i_con_instru[2]), .B(i_con_instru[4]), .C(n27), .Q(n13) );
  XNR21 U16 ( .A(i_con_instru[1]), .B(n10), .Q(n27) );
  OAI2111 U17 ( .A(n9), .B(n18), .C(n19), .D(n15), .Q(o_con_ifsign) );
  NAND31 U18 ( .A(n9), .B(n5), .C(i_con_instru[2]), .Q(n19) );
  NAND22 U19 ( .A(i_con_instru[0]), .B(i_con_instru[1]), .Q(n24) );
  NAND22 U20 ( .A(i_con_instru[3]), .B(n6), .Q(n20) );
  INV3 U21 ( .A(i_con_instru[4]), .Q(n6) );
  NAND22 U22 ( .A(i_con_instru[5]), .B(n5), .Q(n16) );
  INV3 U24 ( .A(i_con_instru[0]), .Q(n10) );
  NOR21 U25 ( .A(i_con_instru[3]), .B(n14), .Q(o_con_regdst) );
  NAND22 U26 ( .A(i_con_instru[5]), .B(n7), .Q(n15) );
  INV3 U27 ( .A(n11), .Q(n7) );
  NAND22 U28 ( .A(i_con_instru[3]), .B(n3), .Q(n21) );
  NAND31 U29 ( .A(n2), .B(n9), .C(i_con_instru[2]), .Q(n17) );
  NAND31 U30 ( .A(i_con_instru[1]), .B(n10), .C(n2), .Q(n23) );
  INV3 U31 ( .A(i_con_instru[2]), .Q(n8) );
  AOI2111 U32 ( .A(n24), .B(n26), .C(n21), .D(i_con_instru[4]), .Q(
        o_con_aluop[2]) );
  NAND22 U33 ( .A(i_con_instru[2]), .B(n10), .Q(n26) );
  NOR21 U34 ( .A(i_con_instru[4]), .B(n21), .Q(o_con_aluop[0]) );
  AOI211 U35 ( .A(n23), .B(n25), .C(i_con_instru[4]), .Q(o_con_aluop[3]) );
  NAND31 U36 ( .A(n2), .B(i_con_instru[0]), .C(i_con_instru[2]), .Q(n25) );
  INV3 U37 ( .A(i_con_instru[5]), .Q(n3) );
  AOI211 U38 ( .A(n17), .B(n22), .C(i_con_instru[4]), .Q(o_con_aluop[4]) );
  NAND22 U39 ( .A(n1), .B(n8), .Q(n22) );
  INV3 U40 ( .A(n23), .Q(n1) );
endmodule


module D_jb_control ( o_con_jump, o_con_bop, o_con_aluPC4, o_con_ifstall, 
        i_con_instru, i_con_func, i_con_rt );
  output [1:0] o_con_jump;
  output [2:0] o_con_bop;
  input [5:0] i_con_instru;
  input [5:0] i_con_func;
  input i_con_rt;
  output o_con_aluPC4, o_con_ifstall;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n2, n3, n4,
         n5, n6;

  OAI222 U13 ( .A(n5), .B(n16), .C(n14), .D(n17), .Q(o_con_bop[1]) );
  NAND31 U3 ( .A(n5), .B(n3), .C(n6), .Q(n8) );
  NAND22 U4 ( .A(n7), .B(n8), .Q(o_con_jump[1]) );
  INV3 U5 ( .A(n7), .Q(n2) );
  INV3 U6 ( .A(n13), .Q(o_con_ifstall) );
  AOI211 U7 ( .A(n3), .B(n14), .C(n2), .Q(n13) );
  NAND22 U8 ( .A(n7), .B(n4), .Q(n17) );
  OAI311 U9 ( .A(n4), .B(n2), .C(n14), .D(n16), .Q(o_con_bop[0]) );
  OAI2111 U10 ( .A(n9), .B(n8), .C(n10), .D(n7), .Q(o_con_jump[0]) );
  NOR40 U11 ( .A(n11), .B(i_con_func[2]), .C(i_con_func[5]), .D(i_con_func[4]), 
        .Q(n9) );
  NAND22 U12 ( .A(i_con_instru[1]), .B(n3), .Q(n10) );
  NAND22 U14 ( .A(n12), .B(i_con_func[3]), .Q(n11) );
  NOR31 U15 ( .A(i_con_instru[3]), .B(i_con_instru[5]), .C(i_con_instru[4]), 
        .Q(n7) );
  INV3 U16 ( .A(i_con_instru[2]), .Q(n3) );
  INV3 U17 ( .A(i_con_instru[1]), .Q(n5) );
  INV3 U18 ( .A(i_con_instru[0]), .Q(n6) );
  NOR21 U19 ( .A(i_con_func[1]), .B(i_con_func[0]), .Q(n12) );
  NAND22 U20 ( .A(i_con_instru[0]), .B(n5), .Q(n14) );
  NOR40 U21 ( .A(i_con_instru[2]), .B(n2), .C(n5), .D(n6), .Q(o_con_aluPC4) );
  NAND31 U22 ( .A(n7), .B(n6), .C(i_con_instru[2]), .Q(n16) );
  NOR31 U23 ( .A(n15), .B(n2), .C(n6), .Q(o_con_bop[2]) );
  XNR21 U24 ( .A(n5), .B(i_con_instru[2]), .Q(n15) );
  INV3 U25 ( .A(n18), .Q(n4) );
  NOR21 U26 ( .A(i_con_instru[2]), .B(i_con_rt), .Q(n18) );
endmodule


module D_pcadd_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274;

  NAND22 U2 ( .A(n29), .B(n26), .Q(n31) );
  NAND22 U3 ( .A(n23), .B(n30), .Q(n25) );
  NAND22 U4 ( .A(n224), .B(n233), .Q(n234) );
  NAND22 U5 ( .A(n192), .B(n191), .Q(n207) );
  NAND22 U6 ( .A(n187), .B(n201), .Q(n202) );
  NAND22 U7 ( .A(n153), .B(n152), .Q(n170) );
  NAND22 U8 ( .A(n148), .B(n165), .Q(n166) );
  NAND22 U9 ( .A(n115), .B(n117), .Q(n131) );
  NAND22 U10 ( .A(n86), .B(n85), .Q(n98) );
  NAND22 U11 ( .A(n81), .B(n93), .Q(n94) );
  MUX22 U12 ( .A(B[0]), .B(n274), .S(A[0]), .Q(SUM[0]) );
  INV3 U13 ( .A(B[30]), .Q(n9) );
  NAND31 U14 ( .A(n244), .B(n245), .C(n243), .Q(n37) );
  INV3 U15 ( .A(n252), .Q(n244) );
  AOI211 U16 ( .A(n246), .B(n247), .C(n248), .Q(n245) );
  INV3 U17 ( .A(n255), .Q(n243) );
  NOR31 U18 ( .A(n65), .B(n66), .C(n67), .Q(n54) );
  INV3 U19 ( .A(n70), .Q(n66) );
  NOR21 U20 ( .A(n69), .B(n71), .Q(n65) );
  NOR31 U21 ( .A(n103), .B(n68), .C(n69), .Q(n67) );
  OAI311 U22 ( .A(n261), .B(n262), .C(n263), .D(n264), .Q(n260) );
  INV3 U23 ( .A(n29), .Q(n263) );
  AOI211 U24 ( .A(n265), .B(n23), .C(n24), .Q(n264) );
  INV3 U25 ( .A(n23), .Q(n261) );
  AOI2111 U26 ( .A(n19), .B(n13), .C(n222), .D(n223), .Q(n218) );
  AOI211 U27 ( .A(n114), .B(n115), .C(n116), .Q(n106) );
  INV3 U28 ( .A(n117), .Q(n116) );
  NAND22 U29 ( .A(n175), .B(n176), .Q(n111) );
  AOI211 U30 ( .A(n180), .B(n181), .C(n182), .Q(n175) );
  NAND22 U31 ( .A(n177), .B(n16), .Q(n176) );
  XNR21 U32 ( .A(n98), .B(n96), .Q(SUM[25]) );
  XOR21 U33 ( .A(n134), .B(n132), .Q(SUM[21]) );
  NAND22 U34 ( .A(n121), .B(n120), .Q(n134) );
  XNR21 U35 ( .A(n166), .B(n164), .Q(SUM[18]) );
  XNR21 U36 ( .A(n94), .B(n92), .Q(SUM[26]) );
  NAND22 U37 ( .A(n152), .B(n167), .Q(n164) );
  NAND22 U38 ( .A(n168), .B(n153), .Q(n167) );
  NAND22 U39 ( .A(n85), .B(n95), .Q(n92) );
  NAND22 U40 ( .A(n96), .B(n86), .Q(n95) );
  XNR21 U41 ( .A(n131), .B(n130), .Q(SUM[22]) );
  NAND22 U42 ( .A(n110), .B(n111), .Q(n109) );
  NOR21 U43 ( .A(n112), .B(n113), .Q(n110) );
  NOR21 U44 ( .A(n178), .B(n179), .Q(n177) );
  NOR21 U45 ( .A(n249), .B(n250), .Q(n248) );
  INV3 U46 ( .A(n72), .Q(n71) );
  INV3 U47 ( .A(n103), .Q(n76) );
  NOR21 U48 ( .A(n104), .B(n105), .Q(n103) );
  OAI2111 U49 ( .A(n106), .B(n107), .C(n108), .D(n109), .Q(n105) );
  NOR21 U50 ( .A(n143), .B(n113), .Q(n104) );
  INV3 U51 ( .A(n26), .Q(n265) );
  AOI211 U52 ( .A(n215), .B(n16), .C(n181), .Q(n208) );
  INV3 U53 ( .A(n178), .Q(n215) );
  NAND22 U54 ( .A(n19), .B(n238), .Q(n237) );
  NAND22 U55 ( .A(n239), .B(n16), .Q(n238) );
  INV3 U56 ( .A(n271), .Q(n239) );
  XNR21 U57 ( .A(n31), .B(n28), .Q(SUM[5]) );
  XOR21 U58 ( .A(n10), .B(n11), .Q(SUM[9]) );
  NAND22 U59 ( .A(n12), .B(n13), .Q(n10) );
  XNR21 U60 ( .A(n207), .B(n204), .Q(SUM[13]) );
  XNR21 U61 ( .A(n170), .B(n168), .Q(SUM[17]) );
  XNR21 U62 ( .A(n234), .B(n232), .Q(SUM[10]) );
  XNR21 U63 ( .A(n202), .B(n200), .Q(SUM[14]) );
  NAND22 U64 ( .A(n26), .B(n27), .Q(n22) );
  NAND22 U65 ( .A(n28), .B(n29), .Q(n27) );
  NAND22 U66 ( .A(n191), .B(n203), .Q(n200) );
  NAND22 U67 ( .A(n204), .B(n192), .Q(n203) );
  XNR21 U68 ( .A(n25), .B(n22), .Q(SUM[6]) );
  XOR21 U69 ( .A(n44), .B(n57), .Q(SUM[2]) );
  NOR21 U70 ( .A(n58), .B(n46), .Q(n57) );
  XOR21 U71 ( .A(n61), .B(n159), .Q(SUM[1]) );
  NOR21 U72 ( .A(n160), .B(n63), .Q(n159) );
  INV3 U73 ( .A(n19), .Q(n18) );
  NAND22 U74 ( .A(n59), .B(n60), .Q(n44) );
  NAND22 U75 ( .A(n61), .B(n62), .Q(n60) );
  INV3 U76 ( .A(n63), .Q(n62) );
  AOI211 U77 ( .A(n250), .B(n249), .C(n63), .Q(n246) );
  INV3 U78 ( .A(n46), .Q(n45) );
  NAND31 U79 ( .A(n115), .B(n121), .C(n122), .Q(n113) );
  NOR21 U80 ( .A(n123), .B(n124), .Q(n122) );
  NOR21 U81 ( .A(B[23]), .B(A[23]), .Q(n124) );
  NOR21 U82 ( .A(B[20]), .B(A[20]), .Q(n123) );
  NAND31 U83 ( .A(n224), .B(n12), .C(n225), .Q(n178) );
  NOR21 U84 ( .A(n226), .B(n227), .Q(n225) );
  NOR21 U85 ( .A(B[11]), .B(A[11]), .Q(n226) );
  NOR21 U86 ( .A(B[8]), .B(A[8]), .Q(n227) );
  NAND22 U87 ( .A(n266), .B(n267), .Q(n29) );
  INV3 U88 ( .A(A[5]), .Q(n267) );
  INV3 U89 ( .A(B[5]), .Q(n266) );
  NAND31 U90 ( .A(n148), .B(n153), .C(n154), .Q(n112) );
  NOR21 U91 ( .A(n155), .B(n156), .Q(n154) );
  NOR21 U92 ( .A(B[16]), .B(A[16]), .Q(n155) );
  NOR21 U93 ( .A(B[19]), .B(A[19]), .Q(n156) );
  NOR21 U94 ( .A(A[24]), .B(B[24]), .Q(n99) );
  NOR21 U95 ( .A(A[16]), .B(B[16]), .Q(n171) );
  NAND22 U96 ( .A(B[29]), .B(A[29]), .Q(n56) );
  NOR21 U97 ( .A(A[29]), .B(B[29]), .Q(n55) );
  NAND31 U98 ( .A(n187), .B(n192), .C(n193), .Q(n179) );
  NOR21 U99 ( .A(n194), .B(n195), .Q(n193) );
  NOR21 U100 ( .A(B[15]), .B(A[15]), .Q(n195) );
  NOR21 U101 ( .A(B[12]), .B(A[12]), .Q(n194) );
  NAND22 U102 ( .A(n4), .B(n169), .Q(n148) );
  INV3 U103 ( .A(A[18]), .Q(n169) );
  INV3 U104 ( .A(B[18]), .Q(n4) );
  NAND22 U105 ( .A(n6), .B(n133), .Q(n115) );
  INV3 U106 ( .A(A[22]), .Q(n133) );
  INV3 U107 ( .A(B[22]), .Q(n6) );
  NAND22 U108 ( .A(B[5]), .B(A[5]), .Q(n26) );
  NAND22 U109 ( .A(B[8]), .B(A[8]), .Q(n19) );
  NAND22 U110 ( .A(B[22]), .B(A[22]), .Q(n117) );
  XOR21 U111 ( .A(n47), .B(n48), .Q(SUM[31]) );
  XNR21 U112 ( .A(B[31]), .B(A[31]), .Q(n47) );
  AOI211 U113 ( .A(n49), .B(n50), .C(n51), .Q(n48) );
  NOR21 U114 ( .A(n52), .B(n9), .Q(n51) );
  NAND22 U115 ( .A(B[9]), .B(A[9]), .Q(n13) );
  NAND22 U116 ( .A(n240), .B(n241), .Q(n16) );
  AOI221 U117 ( .A(A[7]), .B(B[7]), .C(n259), .D(n260), .Q(n240) );
  NAND31 U118 ( .A(n242), .B(n23), .C(n37), .Q(n241) );
  INV3 U119 ( .A(n270), .Q(n259) );
  NAND22 U120 ( .A(B[13]), .B(A[13]), .Q(n191) );
  NAND22 U121 ( .A(B[17]), .B(A[17]), .Q(n152) );
  NAND22 U122 ( .A(B[25]), .B(A[25]), .Q(n85) );
  NAND22 U123 ( .A(B[16]), .B(A[16]), .Q(n151) );
  NAND22 U124 ( .A(B[20]), .B(A[20]), .Q(n119) );
  NAND22 U125 ( .A(B[24]), .B(A[24]), .Q(n84) );
  NAND22 U126 ( .A(B[21]), .B(A[21]), .Q(n120) );
  NOR21 U127 ( .A(A[3]), .B(B[3]), .Q(n254) );
  NAND22 U128 ( .A(B[19]), .B(A[19]), .Q(n146) );
  NOR21 U129 ( .A(A[19]), .B(B[19]), .Q(n145) );
  AOI211 U130 ( .A(n147), .B(n148), .C(n149), .Q(n144) );
  NAND22 U131 ( .A(B[27]), .B(A[27]), .Q(n79) );
  NOR21 U132 ( .A(A[27]), .B(B[27]), .Q(n78) );
  AOI211 U133 ( .A(n80), .B(n81), .C(n82), .Q(n77) );
  NOR21 U134 ( .A(A[20]), .B(B[20]), .Q(n137) );
  NAND22 U135 ( .A(B[6]), .B(A[6]), .Q(n30) );
  NAND22 U136 ( .A(B[18]), .B(A[18]), .Q(n165) );
  NAND22 U137 ( .A(B[10]), .B(A[10]), .Q(n233) );
  NAND22 U138 ( .A(B[14]), .B(A[14]), .Q(n201) );
  NAND22 U139 ( .A(B[26]), .B(A[26]), .Q(n93) );
  NAND22 U140 ( .A(A[4]), .B(B[4]), .Q(n262) );
  NAND22 U141 ( .A(n216), .B(n217), .Q(n181) );
  NAND22 U142 ( .A(B[11]), .B(A[11]), .Q(n216) );
  INV3 U143 ( .A(n221), .Q(n220) );
  NOR31 U144 ( .A(n263), .B(n257), .C(n258), .Q(n242) );
  NOR21 U145 ( .A(B[7]), .B(A[7]), .Q(n258) );
  NOR21 U146 ( .A(B[4]), .B(A[4]), .Q(n257) );
  NOR21 U147 ( .A(n254), .B(n256), .Q(n255) );
  NAND22 U148 ( .A(A[2]), .B(B[2]), .Q(n256) );
  XOR21 U149 ( .A(n162), .B(n163), .Q(SUM[19]) );
  XNR21 U150 ( .A(B[19]), .B(A[19]), .Q(n162) );
  AOI211 U151 ( .A(n164), .B(n148), .C(n149), .Q(n163) );
  XOR21 U152 ( .A(n128), .B(n129), .Q(SUM[23]) );
  XNR21 U153 ( .A(B[23]), .B(A[23]), .Q(n128) );
  AOI211 U154 ( .A(n130), .B(n115), .C(n116), .Q(n129) );
  XOR21 U155 ( .A(n90), .B(n91), .Q(SUM[27]) );
  XNR21 U156 ( .A(B[27]), .B(A[27]), .Q(n90) );
  AOI211 U157 ( .A(n92), .B(n81), .C(n82), .Q(n91) );
  XOR21 U158 ( .A(n64), .B(n54), .Q(SUM[29]) );
  XNR21 U159 ( .A(B[29]), .B(A[29]), .Q(n64) );
  NOR21 U160 ( .A(A[11]), .B(B[11]), .Q(n221) );
  NOR21 U161 ( .A(A[7]), .B(B[7]), .Q(n270) );
  INV3 U162 ( .A(B[3]), .Q(n250) );
  NOR21 U163 ( .A(A[15]), .B(B[15]), .Q(n184) );
  XOR21 U164 ( .A(n2), .B(n50), .Q(SUM[30]) );
  XOR21 U165 ( .A(B[30]), .B(A[30]), .Q(n2) );
  IMUX21 U166 ( .A(n101), .B(n102), .S(n103), .Q(SUM[24]) );
  XNR21 U167 ( .A(B[24]), .B(A[24]), .Q(n102) );
  NOR21 U168 ( .A(n126), .B(n127), .Q(n101) );
  NOR21 U169 ( .A(B[24]), .B(A[24]), .Q(n126) );
  NOR21 U170 ( .A(A[23]), .B(B[23]), .Q(n107) );
  INV3 U171 ( .A(A[3]), .Q(n249) );
  NAND22 U172 ( .A(B[15]), .B(A[15]), .Q(n185) );
  NAND22 U173 ( .A(A[23]), .B(B[23]), .Q(n108) );
  AOI211 U174 ( .A(n186), .B(n187), .C(n188), .Q(n183) );
  NAND22 U175 ( .A(A[12]), .B(B[12]), .Q(n190) );
  NAND22 U176 ( .A(n268), .B(n269), .Q(n23) );
  INV3 U177 ( .A(A[6]), .Q(n269) );
  INV3 U178 ( .A(B[6]), .Q(n268) );
  NAND22 U179 ( .A(n211), .B(n212), .Q(n192) );
  INV3 U180 ( .A(A[13]), .Q(n212) );
  INV3 U181 ( .A(B[13]), .Q(n211) );
  NAND22 U182 ( .A(n205), .B(n206), .Q(n187) );
  INV3 U183 ( .A(A[14]), .Q(n206) );
  INV3 U184 ( .A(B[14]), .Q(n205) );
  NAND22 U185 ( .A(n235), .B(n236), .Q(n12) );
  INV3 U186 ( .A(A[9]), .Q(n236) );
  INV3 U187 ( .A(B[9]), .Q(n235) );
  NAND22 U188 ( .A(n272), .B(n273), .Q(n224) );
  INV3 U189 ( .A(A[10]), .Q(n273) );
  INV3 U190 ( .A(B[10]), .Q(n272) );
  NAND22 U191 ( .A(n3), .B(n172), .Q(n153) );
  INV3 U192 ( .A(A[17]), .Q(n172) );
  INV3 U193 ( .A(B[17]), .Q(n3) );
  NAND22 U194 ( .A(n5), .B(n138), .Q(n121) );
  INV3 U195 ( .A(A[21]), .Q(n138) );
  INV3 U196 ( .A(B[21]), .Q(n5) );
  NAND22 U197 ( .A(n7), .B(n100), .Q(n86) );
  INV3 U198 ( .A(A[25]), .Q(n100) );
  INV3 U199 ( .A(B[25]), .Q(n7) );
  NAND31 U200 ( .A(n81), .B(n86), .C(n87), .Q(n68) );
  NOR21 U201 ( .A(n88), .B(n89), .Q(n87) );
  NOR21 U202 ( .A(B[27]), .B(A[27]), .Q(n89) );
  NOR21 U203 ( .A(B[24]), .B(A[24]), .Q(n88) );
  NOR21 U204 ( .A(A[12]), .B(B[12]), .Q(n209) );
  NOR21 U205 ( .A(A[4]), .B(B[4]), .Q(n33) );
  NOR21 U206 ( .A(A[28]), .B(B[28]), .Q(n69) );
  NAND22 U207 ( .A(B[4]), .B(A[4]), .Q(n34) );
  NOR21 U208 ( .A(A[8]), .B(B[8]), .Q(n271) );
  NAND22 U209 ( .A(B[12]), .B(A[12]), .Q(n210) );
  XOR21 U210 ( .A(n20), .B(n21), .Q(SUM[7]) );
  XNR21 U211 ( .A(B[7]), .B(A[7]), .Q(n20) );
  AOI211 U212 ( .A(n22), .B(n23), .C(n24), .Q(n21) );
  XOR21 U213 ( .A(n230), .B(n231), .Q(SUM[11]) );
  XNR21 U214 ( .A(B[11]), .B(A[11]), .Q(n230) );
  AOI211 U215 ( .A(n232), .B(n224), .C(n219), .Q(n231) );
  XOR21 U216 ( .A(n198), .B(n199), .Q(SUM[15]) );
  XNR21 U217 ( .A(B[15]), .B(A[15]), .Q(n198) );
  AOI211 U218 ( .A(n200), .B(n187), .C(n188), .Q(n199) );
  XOR21 U219 ( .A(n73), .B(n74), .Q(SUM[28]) );
  XNR21 U220 ( .A(B[28]), .B(A[28]), .Q(n73) );
  AOI211 U221 ( .A(n75), .B(n76), .C(n72), .Q(n74) );
  NAND22 U222 ( .A(B[28]), .B(A[28]), .Q(n70) );
  IMUX21 U223 ( .A(n14), .B(n15), .S(n16), .Q(SUM[8]) );
  NOR21 U224 ( .A(n17), .B(n18), .Q(n15) );
  XNR21 U225 ( .A(B[8]), .B(A[8]), .Q(n14) );
  NOR21 U226 ( .A(B[8]), .B(A[8]), .Q(n17) );
  IMUX21 U227 ( .A(n213), .B(n214), .S(n208), .Q(SUM[12]) );
  NOR21 U228 ( .A(n228), .B(n229), .Q(n213) );
  XNR21 U229 ( .A(B[12]), .B(A[12]), .Q(n214) );
  NOR21 U230 ( .A(B[12]), .B(A[12]), .Q(n228) );
  IMUX21 U231 ( .A(n173), .B(n174), .S(n142), .Q(SUM[16]) );
  NOR21 U232 ( .A(n196), .B(n197), .Q(n173) );
  XNR21 U233 ( .A(B[16]), .B(A[16]), .Q(n174) );
  NOR21 U234 ( .A(B[16]), .B(A[16]), .Q(n196) );
  IMUX21 U235 ( .A(n139), .B(n140), .S(n136), .Q(SUM[20]) );
  XNR21 U236 ( .A(B[20]), .B(A[20]), .Q(n140) );
  NOR21 U237 ( .A(n157), .B(n158), .Q(n139) );
  NOR21 U238 ( .A(B[20]), .B(A[20]), .Q(n157) );
  NAND22 U239 ( .A(n8), .B(n97), .Q(n81) );
  INV3 U240 ( .A(A[26]), .Q(n97) );
  INV3 U241 ( .A(B[26]), .Q(n8) );
  INV3 U242 ( .A(n53), .Q(n49) );
  NOR21 U243 ( .A(A[30]), .B(B[30]), .Q(n53) );
  NOR21 U244 ( .A(A[2]), .B(B[2]), .Q(n46) );
  NOR21 U245 ( .A(A[1]), .B(B[1]), .Q(n63) );
  NAND22 U246 ( .A(B[2]), .B(A[2]), .Q(n42) );
  XOR21 U247 ( .A(n40), .B(n41), .Q(SUM[3]) );
  NAND22 U248 ( .A(n42), .B(n43), .Q(n40) );
  XOR21 U249 ( .A(B[3]), .B(A[3]), .Q(n41) );
  NAND22 U250 ( .A(n44), .B(n45), .Q(n43) );
  IMUX21 U251 ( .A(n35), .B(n36), .S(n32), .Q(SUM[4]) );
  NOR21 U252 ( .A(n38), .B(n39), .Q(n35) );
  XNR21 U253 ( .A(B[4]), .B(A[4]), .Q(n36) );
  NOR21 U254 ( .A(B[4]), .B(A[4]), .Q(n38) );
  INV3 U255 ( .A(A[30]), .Q(n52) );
  INV3 U256 ( .A(B[0]), .Q(n274) );
  NOR31 U257 ( .A(n253), .B(n46), .C(n254), .Q(n252) );
  NAND22 U258 ( .A(B[1]), .B(A[1]), .Q(n253) );
  NAND22 U259 ( .A(B[1]), .B(A[1]), .Q(n59) );
  NOR21 U260 ( .A(n46), .B(n251), .Q(n247) );
  NAND22 U261 ( .A(B[0]), .B(A[0]), .Q(n251) );
  INV3 U262 ( .A(n161), .Q(n61) );
  NAND22 U263 ( .A(B[0]), .B(A[0]), .Q(n161) );
  OAI212 U264 ( .A(n32), .B(n33), .C(n34), .Q(n28) );
  CLKIN3 U265 ( .A(n37), .Q(n32) );
  CLKIN3 U266 ( .A(n34), .Q(n39) );
  OAI212 U267 ( .A(n54), .B(n55), .C(n56), .Q(n50) );
  CLKIN3 U268 ( .A(n42), .Q(n58) );
  OAI212 U269 ( .A(n77), .B(n78), .C(n79), .Q(n72) );
  OAI212 U270 ( .A(n83), .B(n84), .C(n85), .Q(n80) );
  CLKIN3 U271 ( .A(n86), .Q(n83) );
  CLKIN3 U272 ( .A(n68), .Q(n75) );
  CLKIN3 U273 ( .A(n93), .Q(n82) );
  OAI212 U274 ( .A(n103), .B(n99), .C(n84), .Q(n96) );
  OAI212 U275 ( .A(n118), .B(n119), .C(n120), .Q(n114) );
  CLKIN3 U276 ( .A(n84), .Q(n127) );
  OAI212 U277 ( .A(n118), .B(n132), .C(n120), .Q(n130) );
  CLKIN3 U278 ( .A(n121), .Q(n118) );
  CLKIN3 U279 ( .A(n135), .Q(n132) );
  OAI212 U280 ( .A(n136), .B(n137), .C(n119), .Q(n135) );
  CLKIN3 U281 ( .A(n141), .Q(n136) );
  OAI212 U282 ( .A(n142), .B(n112), .C(n143), .Q(n141) );
  CLKIN3 U283 ( .A(n125), .Q(n143) );
  OAI212 U284 ( .A(n144), .B(n145), .C(n146), .Q(n125) );
  OAI212 U285 ( .A(n150), .B(n151), .C(n152), .Q(n147) );
  CLKIN3 U286 ( .A(n153), .Q(n150) );
  CLKIN3 U287 ( .A(n119), .Q(n158) );
  CLKIN3 U288 ( .A(n59), .Q(n160) );
  CLKIN3 U289 ( .A(n165), .Q(n149) );
  OAI212 U290 ( .A(n142), .B(n171), .C(n151), .Q(n168) );
  CLKIN3 U291 ( .A(n111), .Q(n142) );
  OAI212 U292 ( .A(n183), .B(n184), .C(n185), .Q(n182) );
  OAI212 U293 ( .A(n189), .B(n190), .C(n191), .Q(n186) );
  CLKIN3 U294 ( .A(n192), .Q(n189) );
  CLKIN3 U295 ( .A(n179), .Q(n180) );
  CLKIN3 U296 ( .A(n151), .Q(n197) );
  CLKIN3 U297 ( .A(n201), .Q(n188) );
  OAI212 U298 ( .A(n208), .B(n209), .C(n210), .Q(n204) );
  OAI212 U299 ( .A(n218), .B(n219), .C(n220), .Q(n217) );
  CLKIN3 U300 ( .A(n224), .Q(n223) );
  CLKIN3 U301 ( .A(n210), .Q(n229) );
  CLKIN3 U302 ( .A(n233), .Q(n219) );
  OAI212 U303 ( .A(n11), .B(n222), .C(n13), .Q(n232) );
  CLKIN3 U304 ( .A(n12), .Q(n222) );
  CLKIN3 U305 ( .A(n237), .Q(n11) );
  CLKIN3 U306 ( .A(n30), .Q(n24) );
endmodule


module D_pcadd ( i_addr_pcadd4E, i_data_immshiftl, o_addr_pcbranchE );
  input [31:0] i_addr_pcadd4E;
  input [31:0] i_data_immshiftl;
  output [31:0] o_addr_pcbranchE;
  wire   n1;

  D_pcadd_DW01_add_1 add_5 ( .A(i_addr_pcadd4E), .B(i_data_immshiftl), .CI(n1), 
        .SUM(o_addr_pcbranchE) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_addr_Rt, i_con_RegWr, 
        i_addr_Rd, i_data_Rd, o_data_Rs, o_data_Rt );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rt;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr;
  wire   n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812;
  wire   [1023:0] regs;

  DFEC1 regs_reg_30__27_ ( .D(i_data_Rd[27]), .E(n776), .C(i_clk), .RN(n768), 
        .Q(regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(i_data_Rd[26]), .E(n776), .C(i_clk), .RN(n768), 
        .Q(regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(i_data_Rd[25]), .E(n776), .C(i_clk), .RN(n768), 
        .Q(regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(i_data_Rd[24]), .E(n776), .C(i_clk), .RN(n768), 
        .Q(regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(i_data_Rd[23]), .E(n776), .C(i_clk), .RN(n768), 
        .Q(regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(i_data_Rd[22]), .E(n776), .C(i_clk), .RN(n768), 
        .Q(regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(i_data_Rd[21]), .E(n776), .C(i_clk), .RN(n768), 
        .Q(regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(i_data_Rd[20]), .E(n776), .C(i_clk), .RN(n768), 
        .Q(regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n776), .C(i_clk), .RN(n768), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(i_data_Rd[18]), .E(n776), .C(i_clk), .RN(n769), 
        .Q(regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(i_data_Rd[17]), .E(n776), .C(i_clk), .RN(n769), 
        .Q(regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(i_data_Rd[16]), .E(n776), .C(i_clk), .RN(n769), 
        .Q(regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(i_data_Rd[15]), .E(n776), .C(i_clk), .RN(n769), 
        .Q(regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(i_data_Rd[14]), .E(n776), .C(i_clk), .RN(n769), 
        .Q(regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(i_data_Rd[13]), .E(n776), .C(i_clk), .RN(n769), 
        .Q(regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(i_data_Rd[12]), .E(n776), .C(i_clk), .RN(n769), 
        .Q(regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(i_data_Rd[11]), .E(n776), .C(i_clk), .RN(n769), 
        .Q(regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(i_data_Rd[10]), .E(n776), .C(i_clk), .RN(n769), 
        .Q(regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(i_data_Rd[9]), .E(n776), .C(i_clk), .RN(n770), 
        .Q(regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(i_data_Rd[8]), .E(n776), .C(i_clk), .RN(n770), 
        .Q(regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(i_data_Rd[7]), .E(n776), .C(i_clk), .RN(n770), 
        .Q(regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n776), .C(i_clk), .RN(n770), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(i_data_Rd[5]), .E(n776), .C(i_clk), .RN(n770), 
        .Q(regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(i_data_Rd[4]), .E(n776), .C(i_clk), .RN(n770), 
        .Q(regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(i_data_Rd[3]), .E(n776), .C(i_clk), .RN(n770), 
        .Q(regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(i_data_Rd[2]), .E(n776), .C(i_clk), .RN(n770), 
        .Q(regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n776), .C(i_clk), .RN(n770), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(i_data_Rd[0]), .E(n776), .C(i_clk), .RN(n771), 
        .Q(regs[960]) );
  DFEC1 regs_reg_26__31_ ( .D(i_data_Rd[31]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(i_data_Rd[30]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(i_data_Rd[29]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(i_data_Rd[28]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(i_data_Rd[27]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(i_data_Rd[26]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(i_data_Rd[25]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(i_data_Rd[24]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(i_data_Rd[23]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(i_data_Rd[22]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(i_data_Rd[21]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(i_data_Rd[20]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(i_data_Rd[18]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(i_data_Rd[17]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(i_data_Rd[16]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(i_data_Rd[15]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(i_data_Rd[14]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(i_data_Rd[13]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(i_data_Rd[12]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(i_data_Rd[11]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(i_data_Rd[10]), .E(n780), .C(i_clk), .RN(i_rst_n), .Q(regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(i_data_Rd[9]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(i_data_Rd[8]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(i_data_Rd[7]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(i_data_Rd[5]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(i_data_Rd[4]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(i_data_Rd[3]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(i_data_Rd[2]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(i_data_Rd[0]), .E(n780), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[832]) );
  DFEC1 regs_reg_22__31_ ( .D(i_data_Rd[31]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(i_data_Rd[30]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(i_data_Rd[29]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(i_data_Rd[28]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(i_data_Rd[27]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(i_data_Rd[26]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(i_data_Rd[25]), .E(n789), .C(i_clk), .RN(n774), 
        .Q(regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(i_data_Rd[24]), .E(n789), .C(i_clk), .RN(n769), 
        .Q(regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(i_data_Rd[23]), .E(n789), .C(i_clk), .RN(n766), 
        .Q(regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(i_data_Rd[22]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(i_data_Rd[21]), .E(n789), .C(i_clk), .RN(n772), 
        .Q(regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(i_data_Rd[20]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(i_data_Rd[19]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(i_data_Rd[18]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(i_data_Rd[17]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(i_data_Rd[16]), .E(n789), .C(i_clk), .RN(n771), 
        .Q(regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(i_data_Rd[15]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(i_data_Rd[14]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(i_data_Rd[13]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(i_data_Rd[12]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(i_data_Rd[11]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(i_data_Rd[10]), .E(n789), .C(i_clk), .RN(i_rst_n), .Q(regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(i_data_Rd[9]), .E(n789), .C(i_clk), .RN(n774), 
        .Q(regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(i_data_Rd[8]), .E(n789), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(i_data_Rd[7]), .E(n789), .C(i_clk), .RN(n766), 
        .Q(regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(i_data_Rd[6]), .E(n789), .C(i_clk), .RN(n767), 
        .Q(regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(i_data_Rd[5]), .E(n789), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(i_data_Rd[4]), .E(n789), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(i_data_Rd[3]), .E(n789), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(i_data_Rd[2]), .E(n789), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(i_data_Rd[1]), .E(n789), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(i_data_Rd[0]), .E(n789), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[704]) );
  DFEC1 regs_reg_18__31_ ( .D(i_data_Rd[31]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(i_data_Rd[30]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(i_data_Rd[29]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(i_data_Rd[28]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(i_data_Rd[27]), .E(n785), .C(i_clk), .RN(n768), 
        .Q(regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(i_data_Rd[26]), .E(n785), .C(i_clk), .RN(n773), 
        .Q(regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(i_data_Rd[25]), .E(n785), .C(i_clk), .RN(n766), 
        .Q(regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(i_data_Rd[24]), .E(n785), .C(i_clk), .RN(n768), 
        .Q(regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(i_data_Rd[23]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(i_data_Rd[22]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(i_data_Rd[21]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(i_data_Rd[20]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(i_data_Rd[19]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(i_data_Rd[18]), .E(n785), .C(i_clk), .RN(n770), 
        .Q(regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(i_data_Rd[17]), .E(n785), .C(i_clk), .RN(n771), 
        .Q(regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(i_data_Rd[16]), .E(n785), .C(i_clk), .RN(n767), 
        .Q(regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(i_data_Rd[15]), .E(n785), .C(i_clk), .RN(n774), 
        .Q(regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(i_data_Rd[14]), .E(n785), .C(i_clk), .RN(n770), 
        .Q(regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(i_data_Rd[13]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(i_data_Rd[12]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(i_data_Rd[11]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(i_data_Rd[10]), .E(n785), .C(i_clk), .RN(i_rst_n), .Q(regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(i_data_Rd[9]), .E(n785), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(i_data_Rd[8]), .E(n785), .C(i_clk), .RN(n770), 
        .Q(regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(i_data_Rd[7]), .E(n785), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(i_data_Rd[6]), .E(n785), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(i_data_Rd[5]), .E(n785), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(i_data_Rd[4]), .E(n785), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(i_data_Rd[3]), .E(n785), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(i_data_Rd[2]), .E(n785), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(i_data_Rd[1]), .E(n785), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(i_data_Rd[0]), .E(n785), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[576]) );
  DFEC1 regs_reg_14__21_ ( .D(i_data_Rd[21]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[469]) );
  DFEC1 regs_reg_14__19_ ( .D(i_data_Rd[19]), .E(n793), .C(i_clk), .RN(n772), 
        .Q(regs[467]) );
  DFEC1 regs_reg_14__13_ ( .D(i_data_Rd[13]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(i_data_Rd[12]), .E(n793), .C(i_clk), .RN(n773), 
        .Q(regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(i_data_Rd[11]), .E(n793), .C(i_clk), .RN(n768), 
        .Q(regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n793), .C(i_clk), .RN(n769), 
        .Q(regs[458]) );
  DFEC1 regs_reg_14__3_ ( .D(i_data_Rd[3]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(i_data_Rd[2]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(i_data_Rd[1]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[449]) );
  DFEC1 regs_reg_10__27_ ( .D(i_data_Rd[27]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(i_data_Rd[26]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(i_data_Rd[25]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(i_data_Rd[24]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(i_data_Rd[23]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(i_data_Rd[22]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(i_data_Rd[21]), .E(n797), .C(i_clk), .RN(n768), 
        .Q(regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(i_data_Rd[20]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(i_data_Rd[19]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(i_data_Rd[18]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(i_data_Rd[17]), .E(n797), .C(i_clk), .RN(n770), 
        .Q(regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(i_data_Rd[16]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(i_data_Rd[15]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(i_data_Rd[13]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(i_data_Rd[12]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(i_data_Rd[11]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n797), .C(i_clk), .RN(n766), 
        .Q(regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(i_data_Rd[9]), .E(n797), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(i_data_Rd[8]), .E(n797), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(i_data_Rd[7]), .E(n797), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(i_data_Rd[6]), .E(n797), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(i_data_Rd[5]), .E(n797), .C(i_clk), .RN(n774), 
        .Q(regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(i_data_Rd[4]), .E(n797), .C(i_clk), .RN(n773), 
        .Q(regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(i_data_Rd[3]), .E(n797), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(i_data_Rd[2]), .E(n797), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(i_data_Rd[1]), .E(n797), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(i_data_Rd[0]), .E(n797), .C(i_clk), .RN(n772), 
        .Q(regs[320]) );
  DFEC1 regs_reg_6__27_ ( .D(i_data_Rd[27]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(i_data_Rd[26]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(i_data_Rd[25]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(i_data_Rd[24]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(i_data_Rd[23]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(i_data_Rd[22]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(i_data_Rd[21]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(i_data_Rd[20]), .E(n801), .C(i_clk), .RN(n773), 
        .Q(regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(i_data_Rd[19]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(i_data_Rd[18]), .E(n801), .C(i_clk), .RN(n768), 
        .Q(regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(i_data_Rd[17]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(i_data_Rd[16]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(i_data_Rd[15]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(i_data_Rd[14]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(i_data_Rd[13]), .E(n801), .C(i_clk), .RN(n774), 
        .Q(regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(i_data_Rd[12]), .E(n801), .C(i_clk), .RN(n766), 
        .Q(regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(i_data_Rd[11]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(i_data_Rd[10]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(i_data_Rd[9]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(i_data_Rd[8]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(i_data_Rd[7]), .E(n801), .C(i_clk), .RN(n772), .Q(
        regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(i_data_Rd[6]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(i_data_Rd[5]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(i_data_Rd[4]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(i_data_Rd[3]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(i_data_Rd[2]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(i_data_Rd[1]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(i_data_Rd[0]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[192]) );
  DFEC1 regs_reg_2__27_ ( .D(i_data_Rd[27]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(i_data_Rd[26]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(i_data_Rd[25]), .E(n805), .C(i_clk), .RN(n766), 
        .Q(regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(i_data_Rd[24]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(i_data_Rd[23]), .E(n805), .C(i_clk), .RN(n771), 
        .Q(regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(i_data_Rd[22]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(i_data_Rd[21]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(i_data_Rd[20]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(i_data_Rd[19]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(i_data_Rd[18]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(i_data_Rd[17]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(i_data_Rd[16]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(i_data_Rd[15]), .E(n805), .C(i_clk), .RN(n774), 
        .Q(regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(i_data_Rd[14]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(i_data_Rd[13]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(i_data_Rd[12]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(i_data_Rd[11]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(i_data_Rd[10]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(i_data_Rd[9]), .E(n805), .C(i_clk), .RN(n767), .Q(
        regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(i_data_Rd[8]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(i_data_Rd[7]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(i_data_Rd[6]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(i_data_Rd[5]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(i_data_Rd[4]), .E(n805), .C(i_clk), .RN(n772), .Q(
        regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(i_data_Rd[3]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(i_data_Rd[2]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(i_data_Rd[1]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(i_data_Rd[0]), .E(n805), .C(i_clk), .RN(n774), .Q(
        regs[64]) );
  DFEC1 regs_reg_31__27_ ( .D(i_data_Rd[27]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(i_data_Rd[26]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(i_data_Rd[25]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(i_data_Rd[24]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(i_data_Rd[23]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(i_data_Rd[22]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(i_data_Rd[21]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(i_data_Rd[20]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(i_data_Rd[18]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(i_data_Rd[17]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(i_data_Rd[16]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(i_data_Rd[15]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(i_data_Rd[14]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(i_data_Rd[13]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(i_data_Rd[12]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(i_data_Rd[11]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(i_data_Rd[10]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(i_data_Rd[9]), .E(n775), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(i_data_Rd[8]), .E(n775), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(i_data_Rd[7]), .E(n775), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n775), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(i_data_Rd[5]), .E(n775), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(i_data_Rd[4]), .E(n775), .C(i_clk), .RN(n767), 
        .Q(regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(i_data_Rd[3]), .E(n775), .C(i_clk), .RN(n767), 
        .Q(regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(i_data_Rd[2]), .E(n775), .C(i_clk), .RN(n767), 
        .Q(regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n775), .C(i_clk), .RN(n767), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(i_data_Rd[0]), .E(n775), .C(i_clk), .RN(n767), 
        .Q(regs[992]) );
  DFEC1 regs_reg_29__27_ ( .D(i_data_Rd[27]), .E(n777), .C(i_clk), .RN(n771), 
        .Q(regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(i_data_Rd[26]), .E(n777), .C(i_clk), .RN(n771), 
        .Q(regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(i_data_Rd[25]), .E(n777), .C(i_clk), .RN(n771), 
        .Q(regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(i_data_Rd[24]), .E(n777), .C(i_clk), .RN(n771), 
        .Q(regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(i_data_Rd[23]), .E(n777), .C(i_clk), .RN(n772), 
        .Q(regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(i_data_Rd[22]), .E(n777), .C(i_clk), .RN(n772), 
        .Q(regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(i_data_Rd[21]), .E(n777), .C(i_clk), .RN(n772), 
        .Q(regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(i_data_Rd[20]), .E(n777), .C(i_clk), .RN(n772), 
        .Q(regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n777), .C(i_clk), .RN(n772), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(i_data_Rd[18]), .E(n777), .C(i_clk), .RN(n772), 
        .Q(regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(i_data_Rd[17]), .E(n777), .C(i_clk), .RN(n772), 
        .Q(regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(i_data_Rd[16]), .E(n777), .C(i_clk), .RN(n772), 
        .Q(regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(i_data_Rd[15]), .E(n777), .C(i_clk), .RN(n772), 
        .Q(regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(i_data_Rd[14]), .E(n777), .C(i_clk), .RN(i_rst_n), .Q(regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(i_data_Rd[13]), .E(n777), .C(i_clk), .RN(i_rst_n), .Q(regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(i_data_Rd[12]), .E(n777), .C(i_clk), .RN(i_rst_n), .Q(regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(i_data_Rd[11]), .E(n777), .C(i_clk), .RN(i_rst_n), .Q(regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(i_data_Rd[10]), .E(n777), .C(i_clk), .RN(i_rst_n), .Q(regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(i_data_Rd[9]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(i_data_Rd[8]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(i_data_Rd[7]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(i_data_Rd[5]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(i_data_Rd[4]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(i_data_Rd[3]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(i_data_Rd[2]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(i_data_Rd[0]), .E(n777), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[928]) );
  DFEC1 regs_reg_28__27_ ( .D(i_data_Rd[27]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(i_data_Rd[26]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(i_data_Rd[25]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(i_data_Rd[24]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(i_data_Rd[23]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(i_data_Rd[22]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(i_data_Rd[21]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(i_data_Rd[20]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(i_data_Rd[18]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(i_data_Rd[17]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(i_data_Rd[16]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(i_data_Rd[15]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(i_data_Rd[14]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(i_data_Rd[13]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(i_data_Rd[12]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(i_data_Rd[11]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(i_data_Rd[10]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(i_data_Rd[9]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(i_data_Rd[8]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(i_data_Rd[7]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(i_data_Rd[5]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(i_data_Rd[4]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(i_data_Rd[3]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(i_data_Rd[2]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(i_data_Rd[0]), .E(n778), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(i_data_Rd[31]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(i_data_Rd[30]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(i_data_Rd[29]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(i_data_Rd[28]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(i_data_Rd[27]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(i_data_Rd[26]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(i_data_Rd[25]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(i_data_Rd[24]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(i_data_Rd[23]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(i_data_Rd[22]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(i_data_Rd[21]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(i_data_Rd[20]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(i_data_Rd[18]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(i_data_Rd[17]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(i_data_Rd[16]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(i_data_Rd[15]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(i_data_Rd[14]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(i_data_Rd[13]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(i_data_Rd[12]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(i_data_Rd[11]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(i_data_Rd[10]), .E(n779), .C(i_clk), .RN(i_rst_n), .Q(regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(i_data_Rd[9]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(i_data_Rd[8]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(i_data_Rd[7]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(i_data_Rd[5]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(i_data_Rd[4]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(i_data_Rd[3]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(i_data_Rd[2]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(i_data_Rd[1]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(i_data_Rd[0]), .E(n779), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[864]) );
  DFEC1 regs_reg_25__31_ ( .D(i_data_Rd[31]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(i_data_Rd[30]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(i_data_Rd[29]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(i_data_Rd[28]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(i_data_Rd[27]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(i_data_Rd[26]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(i_data_Rd[25]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(i_data_Rd[24]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(i_data_Rd[23]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(i_data_Rd[22]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(i_data_Rd[21]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(i_data_Rd[20]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(i_data_Rd[19]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(i_data_Rd[18]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(i_data_Rd[17]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(i_data_Rd[16]), .E(n781), .C(i_clk), .RN(n768), 
        .Q(regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(i_data_Rd[15]), .E(n781), .C(i_clk), .RN(n769), 
        .Q(regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(i_data_Rd[14]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(i_data_Rd[13]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(i_data_Rd[12]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(i_data_Rd[11]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(i_data_Rd[10]), .E(n781), .C(i_clk), .RN(i_rst_n), .Q(regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(i_data_Rd[9]), .E(n781), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(i_data_Rd[8]), .E(n781), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(i_data_Rd[7]), .E(n781), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(i_data_Rd[6]), .E(n781), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(i_data_Rd[5]), .E(n781), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(i_data_Rd[4]), .E(n781), .C(i_clk), .RN(n773), 
        .Q(regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(i_data_Rd[3]), .E(n781), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(i_data_Rd[2]), .E(n781), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(i_data_Rd[1]), .E(n781), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(i_data_Rd[0]), .E(n781), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[800]) );
  DFEC1 regs_reg_24__27_ ( .D(i_data_Rd[27]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(i_data_Rd[26]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(i_data_Rd[25]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(i_data_Rd[24]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(i_data_Rd[23]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(i_data_Rd[22]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(i_data_Rd[21]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(i_data_Rd[20]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(i_data_Rd[19]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(i_data_Rd[18]), .E(n782), .C(i_clk), .RN(n774), 
        .Q(regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(i_data_Rd[17]), .E(n782), .C(i_clk), .RN(n772), 
        .Q(regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(i_data_Rd[16]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(i_data_Rd[15]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(i_data_Rd[14]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(i_data_Rd[13]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(i_data_Rd[12]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(i_data_Rd[11]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(i_data_Rd[10]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(i_data_Rd[9]), .E(n782), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(i_data_Rd[8]), .E(n782), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(i_data_Rd[7]), .E(n782), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(i_data_Rd[6]), .E(n782), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(i_data_Rd[5]), .E(n782), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(i_data_Rd[4]), .E(n782), .C(i_clk), .RN(n774), 
        .Q(regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(i_data_Rd[3]), .E(n782), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(i_data_Rd[2]), .E(n782), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(i_data_Rd[1]), .E(n782), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(i_data_Rd[0]), .E(n782), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(i_data_Rd[31]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(i_data_Rd[30]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(i_data_Rd[29]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(i_data_Rd[28]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(i_data_Rd[27]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(i_data_Rd[26]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(i_data_Rd[25]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(i_data_Rd[24]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(i_data_Rd[23]), .E(n788), .C(i_clk), .RN(n766), 
        .Q(regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(i_data_Rd[22]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(i_data_Rd[21]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(i_data_Rd[20]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(i_data_Rd[19]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(i_data_Rd[18]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(i_data_Rd[17]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(i_data_Rd[16]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(i_data_Rd[15]), .E(n788), .C(i_clk), .RN(n774), 
        .Q(regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(i_data_Rd[14]), .E(n788), .C(i_clk), .RN(n773), 
        .Q(regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(i_data_Rd[13]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(i_data_Rd[12]), .E(n788), .C(i_clk), .RN(n773), 
        .Q(regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(i_data_Rd[11]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(i_data_Rd[10]), .E(n788), .C(i_clk), .RN(i_rst_n), .Q(regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(i_data_Rd[9]), .E(n788), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(i_data_Rd[8]), .E(n788), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(i_data_Rd[7]), .E(n788), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(i_data_Rd[6]), .E(n788), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(i_data_Rd[5]), .E(n788), .C(i_clk), .RN(n767), 
        .Q(regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(i_data_Rd[4]), .E(n788), .C(i_clk), .RN(n768), 
        .Q(regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(i_data_Rd[3]), .E(n788), .C(i_clk), .RN(n769), 
        .Q(regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(i_data_Rd[2]), .E(n788), .C(i_clk), .RN(n770), 
        .Q(regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(i_data_Rd[1]), .E(n788), .C(i_clk), .RN(n771), 
        .Q(regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(i_data_Rd[0]), .E(n788), .C(i_clk), .RN(n772), 
        .Q(regs[736]) );
  DFEC1 regs_reg_21__31_ ( .D(i_data_Rd[31]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(i_data_Rd[30]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(i_data_Rd[29]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(i_data_Rd[28]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(i_data_Rd[27]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(i_data_Rd[26]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(i_data_Rd[25]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(i_data_Rd[24]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(i_data_Rd[23]), .E(n790), .C(i_clk), .RN(n766), 
        .Q(regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(i_data_Rd[22]), .E(n790), .C(i_clk), .RN(n774), 
        .Q(regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(i_data_Rd[21]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(i_data_Rd[20]), .E(n790), .C(i_clk), .RN(n766), 
        .Q(regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(i_data_Rd[19]), .E(n790), .C(i_clk), .RN(n767), 
        .Q(regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(i_data_Rd[18]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(i_data_Rd[17]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(i_data_Rd[16]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(i_data_Rd[15]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(i_data_Rd[14]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(i_data_Rd[13]), .E(n790), .C(i_clk), .RN(n771), 
        .Q(regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(i_data_Rd[12]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(i_data_Rd[11]), .E(n790), .C(i_clk), .RN(n773), 
        .Q(regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(i_data_Rd[10]), .E(n790), .C(i_clk), .RN(i_rst_n), .Q(regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(i_data_Rd[9]), .E(n790), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(i_data_Rd[8]), .E(n790), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(i_data_Rd[7]), .E(n790), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(i_data_Rd[6]), .E(n790), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(i_data_Rd[5]), .E(n790), .C(i_clk), .RN(n769), 
        .Q(regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(i_data_Rd[4]), .E(n790), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(i_data_Rd[3]), .E(n790), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(i_data_Rd[2]), .E(n790), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(i_data_Rd[1]), .E(n790), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(i_data_Rd[0]), .E(n790), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[672]) );
  DFEC1 regs_reg_20__31_ ( .D(i_data_Rd[31]), .E(n783), .C(i_clk), .RN(n767), 
        .Q(regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(i_data_Rd[30]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(i_data_Rd[29]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(i_data_Rd[28]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(i_data_Rd[27]), .E(n783), .C(i_clk), .RN(n773), 
        .Q(regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(i_data_Rd[26]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(i_data_Rd[25]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(i_data_Rd[24]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(i_data_Rd[23]), .E(n783), .C(i_clk), .RN(n766), 
        .Q(regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(i_data_Rd[22]), .E(n783), .C(i_clk), .RN(n772), 
        .Q(regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(i_data_Rd[21]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(i_data_Rd[20]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(i_data_Rd[19]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(i_data_Rd[18]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(i_data_Rd[17]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(i_data_Rd[16]), .E(n783), .C(i_clk), .RN(n774), 
        .Q(regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(i_data_Rd[15]), .E(n783), .C(i_clk), .RN(n773), 
        .Q(regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(i_data_Rd[14]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(i_data_Rd[13]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(i_data_Rd[12]), .E(n783), .C(i_clk), .RN(n768), 
        .Q(regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(i_data_Rd[11]), .E(n783), .C(i_clk), .RN(n766), 
        .Q(regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(i_data_Rd[10]), .E(n783), .C(i_clk), .RN(i_rst_n), .Q(regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(i_data_Rd[9]), .E(n783), .C(i_clk), .RN(n773), 
        .Q(regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(i_data_Rd[8]), .E(n783), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(i_data_Rd[7]), .E(n783), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(i_data_Rd[6]), .E(n783), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(i_data_Rd[5]), .E(n783), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(i_data_Rd[4]), .E(n783), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(i_data_Rd[3]), .E(n783), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(i_data_Rd[2]), .E(n783), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(i_data_Rd[1]), .E(n783), .C(i_clk), .RN(n772), 
        .Q(regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(i_data_Rd[0]), .E(n783), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(i_data_Rd[31]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(i_data_Rd[30]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(i_data_Rd[29]), .E(n784), .C(i_clk), .RN(n769), 
        .Q(regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(i_data_Rd[28]), .E(n784), .C(i_clk), .RN(n767), 
        .Q(regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(i_data_Rd[27]), .E(n784), .C(i_clk), .RN(n766), 
        .Q(regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(i_data_Rd[26]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(i_data_Rd[25]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(i_data_Rd[24]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(i_data_Rd[23]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(i_data_Rd[22]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(i_data_Rd[21]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(i_data_Rd[20]), .E(n784), .C(i_clk), .RN(n766), 
        .Q(regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(i_data_Rd[19]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(i_data_Rd[18]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(i_data_Rd[17]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(i_data_Rd[16]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(i_data_Rd[15]), .E(n784), .C(i_clk), .RN(n774), 
        .Q(regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(i_data_Rd[14]), .E(n784), .C(i_clk), .RN(n773), 
        .Q(regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(i_data_Rd[13]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(i_data_Rd[12]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(i_data_Rd[11]), .E(n784), .C(i_clk), .RN(i_rst_n), .Q(regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(i_data_Rd[10]), .E(n784), .C(i_clk), .RN(n769), 
        .Q(regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(i_data_Rd[9]), .E(n784), .C(i_clk), .RN(n770), 
        .Q(regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(i_data_Rd[8]), .E(n784), .C(i_clk), .RN(n771), 
        .Q(regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(i_data_Rd[7]), .E(n784), .C(i_clk), .RN(n772), 
        .Q(regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(i_data_Rd[6]), .E(n784), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(i_data_Rd[5]), .E(n784), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(i_data_Rd[4]), .E(n784), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(i_data_Rd[3]), .E(n784), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(i_data_Rd[2]), .E(n784), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(i_data_Rd[1]), .E(n784), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(i_data_Rd[0]), .E(n784), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[608]) );
  DFEC1 regs_reg_17__31_ ( .D(i_data_Rd[31]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(i_data_Rd[30]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(i_data_Rd[29]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(i_data_Rd[28]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(i_data_Rd[27]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(i_data_Rd[26]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(i_data_Rd[25]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(i_data_Rd[24]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(i_data_Rd[23]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(i_data_Rd[22]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(i_data_Rd[21]), .E(n786), .C(i_clk), .RN(n774), 
        .Q(regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(i_data_Rd[20]), .E(n786), .C(i_clk), .RN(n766), 
        .Q(regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(i_data_Rd[19]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(i_data_Rd[18]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(i_data_Rd[17]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(i_data_Rd[16]), .E(n786), .C(i_clk), .RN(n771), 
        .Q(regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(i_data_Rd[15]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(i_data_Rd[14]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(i_data_Rd[13]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(i_data_Rd[12]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(i_data_Rd[11]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(i_data_Rd[10]), .E(n786), .C(i_clk), .RN(i_rst_n), .Q(regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(i_data_Rd[9]), .E(n786), .C(i_clk), .RN(n771), 
        .Q(regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(i_data_Rd[8]), .E(n786), .C(i_clk), .RN(n770), 
        .Q(regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(i_data_Rd[7]), .E(n786), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(i_data_Rd[6]), .E(n786), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(i_data_Rd[5]), .E(n786), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(i_data_Rd[4]), .E(n786), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(i_data_Rd[3]), .E(n786), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(i_data_Rd[2]), .E(n786), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(i_data_Rd[1]), .E(n786), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(i_data_Rd[0]), .E(n786), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(i_data_Rd[31]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(i_data_Rd[30]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(i_data_Rd[29]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(i_data_Rd[28]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(i_data_Rd[27]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(i_data_Rd[26]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(i_data_Rd[25]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(i_data_Rd[24]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(i_data_Rd[23]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(i_data_Rd[22]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(i_data_Rd[21]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(i_data_Rd[20]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(i_data_Rd[19]), .E(n787), .C(i_clk), .RN(n774), 
        .Q(regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(i_data_Rd[18]), .E(n787), .C(i_clk), .RN(n773), 
        .Q(regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(i_data_Rd[17]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(i_data_Rd[16]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(i_data_Rd[15]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(i_data_Rd[14]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(i_data_Rd[13]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(i_data_Rd[12]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(i_data_Rd[11]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(i_data_Rd[10]), .E(n787), .C(i_clk), .RN(i_rst_n), .Q(regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(i_data_Rd[9]), .E(n787), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(i_data_Rd[8]), .E(n787), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(i_data_Rd[7]), .E(n787), .C(i_clk), .RN(n770), 
        .Q(regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(i_data_Rd[6]), .E(n787), .C(i_clk), .RN(n771), 
        .Q(regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(i_data_Rd[5]), .E(n787), .C(i_clk), .RN(n772), 
        .Q(regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(i_data_Rd[4]), .E(n787), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(i_data_Rd[3]), .E(n787), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(i_data_Rd[2]), .E(n787), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(i_data_Rd[1]), .E(n787), .C(i_clk), .RN(n773), 
        .Q(regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(i_data_Rd[0]), .E(n787), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[512]) );
  DFEC1 regs_reg_15__21_ ( .D(i_data_Rd[21]), .E(n792), .C(i_clk), .RN(n771), 
        .Q(regs[501]) );
  DFEC1 regs_reg_15__19_ ( .D(i_data_Rd[19]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[499]) );
  DFEC1 regs_reg_15__13_ ( .D(i_data_Rd[13]), .E(n792), .C(i_clk), .RN(n769), 
        .Q(regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(i_data_Rd[12]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(i_data_Rd[11]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[490]) );
  DFEC1 regs_reg_15__3_ ( .D(i_data_Rd[3]), .E(n792), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(i_data_Rd[2]), .E(n792), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(i_data_Rd[1]), .E(n792), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[481]) );
  DFEC1 regs_reg_13__21_ ( .D(i_data_Rd[21]), .E(n794), .C(i_clk), .RN(n770), 
        .Q(regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(i_data_Rd[20]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(i_data_Rd[19]), .E(n794), .C(i_clk), .RN(n768), 
        .Q(regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(i_data_Rd[18]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(i_data_Rd[17]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(i_data_Rd[16]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(i_data_Rd[15]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(i_data_Rd[13]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(i_data_Rd[12]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(i_data_Rd[11]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(i_data_Rd[9]), .E(n794), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(i_data_Rd[8]), .E(n794), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(i_data_Rd[7]), .E(n794), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(i_data_Rd[6]), .E(n794), .C(i_clk), .RN(n773), 
        .Q(regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(i_data_Rd[5]), .E(n794), .C(i_clk), .RN(n774), 
        .Q(regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(i_data_Rd[4]), .E(n794), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(i_data_Rd[3]), .E(n794), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(i_data_Rd[2]), .E(n794), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(i_data_Rd[1]), .E(n794), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(i_data_Rd[0]), .E(n794), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[416]) );
  DFEC1 regs_reg_12__27_ ( .D(i_data_Rd[27]), .E(n795), .C(i_clk), .RN(n770), 
        .Q(regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(i_data_Rd[26]), .E(n795), .C(i_clk), .RN(n769), 
        .Q(regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(i_data_Rd[25]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(i_data_Rd[24]), .E(n795), .C(i_clk), .RN(n770), 
        .Q(regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(i_data_Rd[23]), .E(n795), .C(i_clk), .RN(n772), 
        .Q(regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(i_data_Rd[22]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(i_data_Rd[21]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(i_data_Rd[20]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(i_data_Rd[19]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(i_data_Rd[18]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(i_data_Rd[17]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(i_data_Rd[16]), .E(n795), .C(i_clk), .RN(n773), 
        .Q(regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(i_data_Rd[15]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(i_data_Rd[13]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(i_data_Rd[12]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(i_data_Rd[11]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(i_data_Rd[9]), .E(n795), .C(i_clk), .RN(n767), 
        .Q(regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(i_data_Rd[8]), .E(n795), .C(i_clk), .RN(n773), 
        .Q(regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(i_data_Rd[7]), .E(n795), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(i_data_Rd[6]), .E(n795), .C(i_clk), .RN(n770), 
        .Q(regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(i_data_Rd[5]), .E(n795), .C(i_clk), .RN(n774), 
        .Q(regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(i_data_Rd[4]), .E(n795), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(i_data_Rd[3]), .E(n795), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(i_data_Rd[2]), .E(n795), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(i_data_Rd[1]), .E(n795), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(i_data_Rd[0]), .E(n795), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[384]) );
  DFEC1 regs_reg_11__27_ ( .D(i_data_Rd[27]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(i_data_Rd[26]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(i_data_Rd[25]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(i_data_Rd[24]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(i_data_Rd[23]), .E(n796), .C(i_clk), .RN(n766), 
        .Q(regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(i_data_Rd[22]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(i_data_Rd[21]), .E(n796), .C(i_clk), .RN(n772), 
        .Q(regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(i_data_Rd[20]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(i_data_Rd[19]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(i_data_Rd[18]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(i_data_Rd[17]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(i_data_Rd[16]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(i_data_Rd[15]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(i_data_Rd[13]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(i_data_Rd[12]), .E(n796), .C(i_clk), .RN(n767), 
        .Q(regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(i_data_Rd[11]), .E(n796), .C(i_clk), .RN(n774), 
        .Q(regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(i_data_Rd[10]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(i_data_Rd[9]), .E(n796), .C(i_clk), .RN(n768), 
        .Q(regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(i_data_Rd[8]), .E(n796), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(i_data_Rd[7]), .E(n796), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(i_data_Rd[6]), .E(n796), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(i_data_Rd[5]), .E(n796), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(i_data_Rd[4]), .E(n796), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(i_data_Rd[3]), .E(n796), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(i_data_Rd[2]), .E(n796), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(i_data_Rd[1]), .E(n796), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(i_data_Rd[0]), .E(n796), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[352]) );
  DFEC1 regs_reg_9__27_ ( .D(i_data_Rd[27]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(i_data_Rd[26]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(i_data_Rd[25]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(i_data_Rd[24]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(i_data_Rd[23]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(i_data_Rd[22]), .E(n798), .C(i_clk), .RN(n769), 
        .Q(regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(i_data_Rd[21]), .E(n798), .C(i_clk), .RN(n767), 
        .Q(regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(i_data_Rd[20]), .E(n798), .C(i_clk), .RN(n768), 
        .Q(regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(i_data_Rd[19]), .E(n798), .C(i_clk), .RN(n766), 
        .Q(regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(i_data_Rd[18]), .E(n798), .C(i_clk), .RN(n767), 
        .Q(regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(i_data_Rd[17]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(i_data_Rd[16]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(i_data_Rd[15]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(i_data_Rd[14]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(i_data_Rd[13]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(i_data_Rd[12]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(i_data_Rd[11]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(i_data_Rd[10]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(i_data_Rd[9]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(i_data_Rd[8]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(i_data_Rd[7]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(i_data_Rd[6]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(i_data_Rd[5]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(i_data_Rd[4]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(i_data_Rd[3]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(i_data_Rd[2]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(i_data_Rd[1]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(i_data_Rd[0]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[288]) );
  DFEC1 regs_reg_8__27_ ( .D(i_data_Rd[27]), .E(n799), .C(i_clk), .RN(n767), 
        .Q(regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(i_data_Rd[26]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(i_data_Rd[25]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(i_data_Rd[24]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(i_data_Rd[23]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(i_data_Rd[22]), .E(n799), .C(i_clk), .RN(n771), 
        .Q(regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(i_data_Rd[21]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(i_data_Rd[20]), .E(n799), .C(i_clk), .RN(n766), 
        .Q(regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(i_data_Rd[19]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(i_data_Rd[18]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(i_data_Rd[17]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(i_data_Rd[16]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(i_data_Rd[15]), .E(n799), .C(i_clk), .RN(n766), 
        .Q(regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(i_data_Rd[14]), .E(n799), .C(i_clk), .RN(n768), 
        .Q(regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(i_data_Rd[13]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(i_data_Rd[12]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(i_data_Rd[11]), .E(n799), .C(i_clk), .RN(n774), 
        .Q(regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(i_data_Rd[10]), .E(n799), .C(i_clk), .RN(n771), 
        .Q(regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(i_data_Rd[9]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(i_data_Rd[8]), .E(n799), .C(i_clk), .RN(n767), .Q(
        regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(i_data_Rd[7]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(i_data_Rd[6]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(i_data_Rd[5]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(i_data_Rd[4]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(i_data_Rd[3]), .E(n799), .C(i_clk), .RN(n766), .Q(
        regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(i_data_Rd[2]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(i_data_Rd[1]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(i_data_Rd[0]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[256]) );
  DFEC1 regs_reg_7__27_ ( .D(i_data_Rd[27]), .E(n800), .C(i_clk), .RN(n769), 
        .Q(regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(i_data_Rd[26]), .E(n800), .C(i_clk), .RN(n773), 
        .Q(regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(i_data_Rd[25]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(i_data_Rd[24]), .E(n800), .C(i_clk), .RN(n774), 
        .Q(regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(i_data_Rd[23]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(i_data_Rd[22]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(i_data_Rd[21]), .E(n800), .C(i_clk), .RN(n772), 
        .Q(regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(i_data_Rd[20]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(i_data_Rd[19]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(i_data_Rd[18]), .E(n800), .C(i_clk), .RN(n774), 
        .Q(regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(i_data_Rd[17]), .E(n800), .C(i_clk), .RN(n773), 
        .Q(regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(i_data_Rd[16]), .E(n800), .C(i_clk), .RN(n767), 
        .Q(regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(i_data_Rd[15]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(i_data_Rd[14]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(i_data_Rd[13]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(i_data_Rd[12]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(i_data_Rd[11]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(i_data_Rd[10]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(i_data_Rd[9]), .E(n800), .C(i_clk), .RN(n770), .Q(
        regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(i_data_Rd[8]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(i_data_Rd[7]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(i_data_Rd[6]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(i_data_Rd[5]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(i_data_Rd[4]), .E(n800), .C(i_clk), .RN(n770), .Q(
        regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(i_data_Rd[3]), .E(n800), .C(i_clk), .RN(n774), .Q(
        regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(i_data_Rd[2]), .E(n800), .C(i_clk), .RN(n773), .Q(
        regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(i_data_Rd[1]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(i_data_Rd[0]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[224]) );
  DFEC1 regs_reg_5__27_ ( .D(i_data_Rd[27]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(i_data_Rd[26]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(i_data_Rd[25]), .E(n802), .C(i_clk), .RN(n774), 
        .Q(regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(i_data_Rd[24]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(i_data_Rd[23]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(i_data_Rd[22]), .E(n802), .C(i_clk), .RN(n768), 
        .Q(regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(i_data_Rd[21]), .E(n802), .C(i_clk), .RN(n774), 
        .Q(regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(i_data_Rd[20]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(i_data_Rd[19]), .E(n802), .C(i_clk), .RN(n774), 
        .Q(regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(i_data_Rd[18]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(i_data_Rd[17]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(i_data_Rd[16]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(i_data_Rd[15]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(i_data_Rd[14]), .E(n802), .C(i_clk), .RN(n768), 
        .Q(regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(i_data_Rd[13]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(i_data_Rd[12]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(i_data_Rd[11]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(i_data_Rd[10]), .E(n802), .C(i_clk), .RN(n769), 
        .Q(regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(i_data_Rd[9]), .E(n802), .C(i_clk), .RN(n766), .Q(
        regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(i_data_Rd[8]), .E(n802), .C(i_clk), .RN(n773), .Q(
        regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(i_data_Rd[7]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(i_data_Rd[6]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(i_data_Rd[5]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(i_data_Rd[4]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(i_data_Rd[3]), .E(n802), .C(i_clk), .RN(n772), .Q(
        regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(i_data_Rd[2]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(i_data_Rd[1]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(i_data_Rd[0]), .E(n802), .C(i_clk), .RN(n770), .Q(
        regs[160]) );
  DFEC1 regs_reg_4__27_ ( .D(i_data_Rd[27]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(i_data_Rd[26]), .E(n803), .C(i_clk), .RN(n772), 
        .Q(regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(i_data_Rd[25]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(i_data_Rd[24]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(i_data_Rd[23]), .E(n803), .C(i_clk), .RN(n770), 
        .Q(regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(i_data_Rd[22]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(i_data_Rd[21]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(i_data_Rd[20]), .E(n803), .C(i_clk), .RN(n771), 
        .Q(regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(i_data_Rd[19]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(i_data_Rd[18]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(i_data_Rd[17]), .E(n803), .C(i_clk), .RN(n768), 
        .Q(regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(i_data_Rd[16]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(i_data_Rd[15]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(i_data_Rd[14]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(i_data_Rd[13]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(i_data_Rd[12]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(i_data_Rd[11]), .E(n803), .C(i_clk), .RN(n774), 
        .Q(regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(i_data_Rd[10]), .E(n803), .C(i_clk), .RN(n773), 
        .Q(regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(i_data_Rd[9]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(i_data_Rd[8]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(i_data_Rd[7]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(i_data_Rd[6]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(i_data_Rd[5]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(i_data_Rd[4]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(i_data_Rd[3]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(i_data_Rd[2]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(i_data_Rd[1]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(i_data_Rd[0]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[128]) );
  DFEC1 regs_reg_3__27_ ( .D(i_data_Rd[27]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(i_data_Rd[26]), .E(n804), .C(i_clk), .RN(n768), 
        .Q(regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(i_data_Rd[25]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(i_data_Rd[24]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(i_data_Rd[23]), .E(n804), .C(i_clk), .RN(n769), 
        .Q(regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(i_data_Rd[22]), .E(n804), .C(i_clk), .RN(n767), 
        .Q(regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(i_data_Rd[21]), .E(n804), .C(i_clk), .RN(n771), 
        .Q(regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(i_data_Rd[20]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(i_data_Rd[19]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(i_data_Rd[18]), .E(n804), .C(i_clk), .RN(n773), 
        .Q(regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(i_data_Rd[17]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(i_data_Rd[16]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(i_data_Rd[15]), .E(n804), .C(i_clk), .RN(n766), 
        .Q(regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(i_data_Rd[14]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(i_data_Rd[13]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(i_data_Rd[12]), .E(n804), .C(i_clk), .RN(n773), 
        .Q(regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(i_data_Rd[11]), .E(n804), .C(i_clk), .RN(n771), 
        .Q(regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(i_data_Rd[10]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(i_data_Rd[9]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(i_data_Rd[8]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(i_data_Rd[7]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(i_data_Rd[6]), .E(n804), .C(i_clk), .RN(n767), .Q(
        regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(i_data_Rd[5]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(i_data_Rd[4]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(i_data_Rd[3]), .E(n804), .C(i_clk), .RN(n769), .Q(
        regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(i_data_Rd[2]), .E(n804), .C(i_clk), .RN(n774), .Q(
        regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(i_data_Rd[1]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(i_data_Rd[0]), .E(n804), .C(i_clk), .RN(n772), .Q(
        regs[96]) );
  DFEC1 regs_reg_1__27_ ( .D(i_data_Rd[27]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(i_data_Rd[26]), .E(n806), .C(i_clk), .RN(n771), 
        .Q(regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(i_data_Rd[25]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(i_data_Rd[24]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(i_data_Rd[23]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(i_data_Rd[22]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(i_data_Rd[21]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(i_data_Rd[20]), .E(n806), .C(i_clk), .RN(n773), 
        .Q(regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(i_data_Rd[19]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(i_data_Rd[18]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(i_data_Rd[17]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(i_data_Rd[16]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(i_data_Rd[15]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(i_data_Rd[14]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(i_data_Rd[13]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(i_data_Rd[12]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(i_data_Rd[11]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(i_data_Rd[10]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(i_data_Rd[9]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(i_data_Rd[8]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(i_data_Rd[7]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(i_data_Rd[6]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(i_data_Rd[5]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(i_data_Rd[4]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(i_data_Rd[3]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(i_data_Rd[2]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(i_data_Rd[1]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(i_data_Rd[0]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[32]) );
  DFEC1 regs_reg_0__27_ ( .D(i_data_Rd[27]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(i_data_Rd[26]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(i_data_Rd[25]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(i_data_Rd[24]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(i_data_Rd[23]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(i_data_Rd[22]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(i_data_Rd[21]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(i_data_Rd[20]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(i_data_Rd[19]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(i_data_Rd[18]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(i_data_Rd[17]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(i_data_Rd[16]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(i_data_Rd[15]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(i_data_Rd[14]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(i_data_Rd[13]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(i_data_Rd[12]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(i_data_Rd[11]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(i_data_Rd[10]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(i_data_Rd[9]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(i_data_Rd[8]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(i_data_Rd[7]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(i_data_Rd[6]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(i_data_Rd[5]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(i_data_Rd[4]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(i_data_Rd[3]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(i_data_Rd[2]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(i_data_Rd[1]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(i_data_Rd[0]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[0]) );
  DFEC1 regs_reg_15__31_ ( .D(i_data_Rd[31]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[511]) );
  DFEC1 regs_reg_14__31_ ( .D(i_data_Rd[31]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[479]) );
  DFEC1 regs_reg_13__31_ ( .D(i_data_Rd[31]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[447]) );
  DFEC1 regs_reg_12__31_ ( .D(i_data_Rd[31]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[415]) );
  DFEC1 regs_reg_11__31_ ( .D(i_data_Rd[31]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[383]) );
  DFEC1 regs_reg_10__31_ ( .D(i_data_Rd[31]), .E(n797), .C(i_clk), .RN(i_rst_n), .Q(regs[351]) );
  DFEC1 regs_reg_9__31_ ( .D(i_data_Rd[31]), .E(n798), .C(i_clk), .RN(n766), 
        .Q(regs[319]) );
  DFEC1 regs_reg_8__31_ ( .D(i_data_Rd[31]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[287]) );
  DFEC1 regs_reg_7__31_ ( .D(i_data_Rd[31]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[255]) );
  DFEC1 regs_reg_6__31_ ( .D(i_data_Rd[31]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[223]) );
  DFEC1 regs_reg_5__31_ ( .D(i_data_Rd[31]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[191]) );
  DFEC1 regs_reg_4__31_ ( .D(i_data_Rd[31]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[159]) );
  DFEC1 regs_reg_3__31_ ( .D(i_data_Rd[31]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[127]) );
  DFEC1 regs_reg_2__31_ ( .D(i_data_Rd[31]), .E(n805), .C(i_clk), .RN(n766), 
        .Q(regs[95]) );
  DFEC1 regs_reg_1__31_ ( .D(i_data_Rd[31]), .E(n806), .C(i_clk), .RN(n773), 
        .Q(regs[63]) );
  DFEC1 regs_reg_0__31_ ( .D(i_data_Rd[31]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[31]) );
  DFEC1 regs_reg_15__30_ ( .D(i_data_Rd[30]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(i_data_Rd[29]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(i_data_Rd[28]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[508]) );
  DFEC1 regs_reg_14__30_ ( .D(i_data_Rd[30]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(i_data_Rd[29]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(i_data_Rd[28]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[476]) );
  DFEC1 regs_reg_13__30_ ( .D(i_data_Rd[30]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(i_data_Rd[29]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(i_data_Rd[28]), .E(n794), .C(i_clk), .RN(n767), 
        .Q(regs[444]) );
  DFEC1 regs_reg_12__30_ ( .D(i_data_Rd[30]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(i_data_Rd[29]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(i_data_Rd[28]), .E(n795), .C(i_clk), .RN(i_rst_n), .Q(regs[412]) );
  DFEC1 regs_reg_11__30_ ( .D(i_data_Rd[30]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(i_data_Rd[29]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(i_data_Rd[28]), .E(n796), .C(i_clk), .RN(i_rst_n), .Q(regs[380]) );
  DFEC1 regs_reg_10__30_ ( .D(i_data_Rd[30]), .E(n797), .C(i_clk), .RN(n771), 
        .Q(regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(i_data_Rd[29]), .E(n797), .C(i_clk), .RN(n769), 
        .Q(regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(i_data_Rd[28]), .E(n797), .C(i_clk), .RN(n769), 
        .Q(regs[348]) );
  DFEC1 regs_reg_9__30_ ( .D(i_data_Rd[30]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(i_data_Rd[29]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(i_data_Rd[28]), .E(n798), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[316]) );
  DFEC1 regs_reg_8__30_ ( .D(i_data_Rd[30]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(i_data_Rd[29]), .E(n799), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(i_data_Rd[28]), .E(n799), .C(i_clk), .RN(n766), 
        .Q(regs[284]) );
  DFEC1 regs_reg_7__30_ ( .D(i_data_Rd[30]), .E(n800), .C(i_clk), .RN(n773), 
        .Q(regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(i_data_Rd[29]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(i_data_Rd[28]), .E(n800), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[252]) );
  DFEC1 regs_reg_6__30_ ( .D(i_data_Rd[30]), .E(n801), .C(i_clk), .RN(n766), 
        .Q(regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(i_data_Rd[29]), .E(n801), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(i_data_Rd[28]), .E(n801), .C(i_clk), .RN(n768), 
        .Q(regs[220]) );
  DFEC1 regs_reg_5__30_ ( .D(i_data_Rd[30]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(i_data_Rd[29]), .E(n802), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(i_data_Rd[28]), .E(n802), .C(i_clk), .RN(n770), 
        .Q(regs[188]) );
  DFEC1 regs_reg_4__30_ ( .D(i_data_Rd[30]), .E(n803), .C(i_clk), .RN(n766), 
        .Q(regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(i_data_Rd[29]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(i_data_Rd[28]), .E(n803), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[156]) );
  DFEC1 regs_reg_3__30_ ( .D(i_data_Rd[30]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(i_data_Rd[29]), .E(n804), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(i_data_Rd[28]), .E(n804), .C(i_clk), .RN(n767), 
        .Q(regs[124]) );
  DFEC1 regs_reg_2__30_ ( .D(i_data_Rd[30]), .E(n805), .C(i_clk), .RN(n770), 
        .Q(regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(i_data_Rd[29]), .E(n805), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(i_data_Rd[28]), .E(n805), .C(i_clk), .RN(n766), 
        .Q(regs[92]) );
  DFEC1 regs_reg_1__30_ ( .D(i_data_Rd[30]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(i_data_Rd[29]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(i_data_Rd[28]), .E(n806), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[60]) );
  DFEC1 regs_reg_0__30_ ( .D(i_data_Rd[30]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(i_data_Rd[29]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(i_data_Rd[28]), .E(n807), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[28]) );
  DFEC1 regs_reg_31__31_ ( .D(i_data_Rd[31]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1023]) );
  DFEC1 regs_reg_31__30_ ( .D(i_data_Rd[30]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(i_data_Rd[29]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(i_data_Rd[28]), .E(n775), .C(i_clk), .RN(i_rst_n), .Q(regs[1020]) );
  DFEC1 regs_reg_30__31_ ( .D(i_data_Rd[31]), .E(n776), .C(i_clk), .RN(n767), 
        .Q(regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(i_data_Rd[30]), .E(n776), .C(i_clk), .RN(n767), 
        .Q(regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(i_data_Rd[29]), .E(n776), .C(i_clk), .RN(n767), 
        .Q(regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(i_data_Rd[28]), .E(n776), .C(i_clk), .RN(n767), 
        .Q(regs[988]) );
  DFEC1 regs_reg_29__31_ ( .D(i_data_Rd[31]), .E(n777), .C(i_clk), .RN(n771), 
        .Q(regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(i_data_Rd[30]), .E(n777), .C(i_clk), .RN(n771), 
        .Q(regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(i_data_Rd[29]), .E(n777), .C(i_clk), .RN(n771), 
        .Q(regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(i_data_Rd[28]), .E(n777), .C(i_clk), .RN(n771), 
        .Q(regs[956]) );
  DFEC1 regs_reg_28__31_ ( .D(i_data_Rd[31]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(i_data_Rd[30]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(i_data_Rd[29]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(i_data_Rd[28]), .E(n778), .C(i_clk), .RN(i_rst_n), .Q(regs[924]) );
  DFEC1 regs_reg_24__31_ ( .D(i_data_Rd[31]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(i_data_Rd[30]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(i_data_Rd[29]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(i_data_Rd[28]), .E(n782), .C(i_clk), .RN(i_rst_n), .Q(regs[796]) );
  DFEC1 regs_reg_15__27_ ( .D(i_data_Rd[27]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(i_data_Rd[26]), .E(n792), .C(i_clk), .RN(n767), 
        .Q(regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(i_data_Rd[25]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(i_data_Rd[24]), .E(n792), .C(i_clk), .RN(n772), 
        .Q(regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(i_data_Rd[23]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(i_data_Rd[22]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[502]) );
  DFEC1 regs_reg_15__20_ ( .D(i_data_Rd[20]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[500]) );
  DFEC1 regs_reg_15__18_ ( .D(i_data_Rd[18]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(i_data_Rd[17]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(i_data_Rd[16]), .E(n792), .C(i_clk), .RN(n771), 
        .Q(regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(i_data_Rd[15]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n792), .C(i_clk), .RN(i_rst_n), .Q(regs[494]) );
  DFEC1 regs_reg_15__9_ ( .D(i_data_Rd[9]), .E(n792), .C(i_clk), .RN(n769), 
        .Q(regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(i_data_Rd[8]), .E(n792), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(i_data_Rd[7]), .E(n792), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(i_data_Rd[6]), .E(n792), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(i_data_Rd[5]), .E(n792), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(i_data_Rd[4]), .E(n792), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[484]) );
  DFEC1 regs_reg_15__0_ ( .D(i_data_Rd[0]), .E(n792), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[480]) );
  DFEC1 regs_reg_14__27_ ( .D(i_data_Rd[27]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(i_data_Rd[26]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(i_data_Rd[25]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(i_data_Rd[24]), .E(n793), .C(i_clk), .RN(n768), 
        .Q(regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(i_data_Rd[23]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(i_data_Rd[22]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[470]) );
  DFEC1 regs_reg_14__20_ ( .D(i_data_Rd[20]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[468]) );
  DFEC1 regs_reg_14__18_ ( .D(i_data_Rd[18]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(i_data_Rd[17]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(i_data_Rd[16]), .E(n793), .C(i_clk), .RN(n769), 
        .Q(regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(i_data_Rd[15]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n793), .C(i_clk), .RN(i_rst_n), .Q(regs[462]) );
  DFEC1 regs_reg_14__9_ ( .D(i_data_Rd[9]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(i_data_Rd[8]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(i_data_Rd[7]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(i_data_Rd[6]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(i_data_Rd[5]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(i_data_Rd[4]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[452]) );
  DFEC1 regs_reg_14__0_ ( .D(i_data_Rd[0]), .E(n793), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[448]) );
  DFEC1 regs_reg_13__27_ ( .D(i_data_Rd[27]), .E(n794), .C(i_clk), .RN(n768), 
        .Q(regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(i_data_Rd[26]), .E(n794), .C(i_clk), .RN(n769), 
        .Q(regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(i_data_Rd[25]), .E(n794), .C(i_clk), .RN(n770), 
        .Q(regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(i_data_Rd[24]), .E(n794), .C(i_clk), .RN(n771), 
        .Q(regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(i_data_Rd[23]), .E(n794), .C(i_clk), .RN(n772), 
        .Q(regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(i_data_Rd[22]), .E(n794), .C(i_clk), .RN(i_rst_n), .Q(regs[438]) );
  BUF2 U2 ( .A(n773), .Q(n772) );
  BUF2 U3 ( .A(n773), .Q(n771) );
  BUF2 U4 ( .A(n773), .Q(n770) );
  BUF2 U5 ( .A(n774), .Q(n769) );
  BUF2 U6 ( .A(n774), .Q(n768) );
  BUF2 U7 ( .A(n774), .Q(n767) );
  BUF2 U8 ( .A(n766), .Q(n773) );
  BUF2 U9 ( .A(n766), .Q(n774) );
  BUF2 U10 ( .A(n399), .Q(n385) );
  BUF2 U11 ( .A(n399), .Q(n386) );
  BUF2 U12 ( .A(n399), .Q(n387) );
  BUF2 U13 ( .A(n400), .Q(n388) );
  BUF2 U14 ( .A(n400), .Q(n389) );
  BUF2 U15 ( .A(n400), .Q(n390) );
  BUF2 U16 ( .A(n399), .Q(n391) );
  BUF2 U17 ( .A(i_addr_Rt[0]), .Q(n392) );
  BUF2 U18 ( .A(i_addr_Rt[0]), .Q(n393) );
  BUF2 U19 ( .A(i_addr_Rt[0]), .Q(n394) );
  BUF2 U20 ( .A(i_addr_Rt[0]), .Q(n395) );
  BUF2 U21 ( .A(n400), .Q(n396) );
  BUF2 U22 ( .A(n399), .Q(n397) );
  BUF2 U23 ( .A(i_addr_Rt[0]), .Q(n398) );
  BUF2 U24 ( .A(i_addr_Rs[0]), .Q(n749) );
  BUF2 U25 ( .A(i_addr_Rs[0]), .Q(n750) );
  BUF2 U26 ( .A(i_addr_Rs[0]), .Q(n751) );
  BUF2 U27 ( .A(n763), .Q(n752) );
  BUF2 U28 ( .A(n763), .Q(n753) );
  BUF2 U29 ( .A(n763), .Q(n754) );
  BUF2 U30 ( .A(n763), .Q(n755) );
  BUF2 U31 ( .A(n763), .Q(n756) );
  BUF2 U32 ( .A(i_addr_Rs[0]), .Q(n757) );
  BUF2 U33 ( .A(n765), .Q(n758) );
  BUF2 U34 ( .A(n765), .Q(n759) );
  BUF2 U35 ( .A(n765), .Q(n760) );
  BUF2 U36 ( .A(n765), .Q(n761) );
  BUF2 U37 ( .A(n765), .Q(n762) );
  INV3 U38 ( .A(n60), .Q(n775) );
  NAND22 U39 ( .A(n48), .B(n46), .Q(n60) );
  BUF2 U40 ( .A(i_addr_Rt[1]), .Q(n377) );
  BUF2 U41 ( .A(n375), .Q(n378) );
  BUF2 U42 ( .A(n376), .Q(n379) );
  BUF2 U43 ( .A(n376), .Q(n380) );
  BUF2 U44 ( .A(n376), .Q(n381) );
  BUF2 U45 ( .A(n375), .Q(n382) );
  BUF2 U46 ( .A(n375), .Q(n383) );
  BUF2 U47 ( .A(i_addr_Rs[1]), .Q(n733) );
  BUF2 U48 ( .A(i_addr_Rs[1]), .Q(n734) );
  BUF2 U49 ( .A(n732), .Q(n735) );
  BUF2 U50 ( .A(n732), .Q(n736) );
  BUF2 U51 ( .A(n748), .Q(n737) );
  BUF2 U52 ( .A(i_addr_Rs[1]), .Q(n738) );
  BUF2 U53 ( .A(n732), .Q(n739) );
  BUF2 U54 ( .A(n731), .Q(n740) );
  BUF2 U55 ( .A(n731), .Q(n741) );
  BUF2 U56 ( .A(n731), .Q(n742) );
  BUF2 U57 ( .A(n730), .Q(n743) );
  BUF2 U58 ( .A(n730), .Q(n744) );
  BUF2 U59 ( .A(n730), .Q(n745) );
  BUF2 U60 ( .A(i_rst_n), .Q(n766) );
  NOR31 U61 ( .A(n812), .B(n791), .C(n808), .Q(n48) );
  NOR31 U62 ( .A(n811), .B(n809), .C(n810), .Q(n46) );
  INV3 U63 ( .A(n39), .Q(n783) );
  NAND22 U64 ( .A(n42), .B(n57), .Q(n39) );
  INV3 U65 ( .A(n79), .Q(n787) );
  NAND22 U66 ( .A(n49), .B(n42), .Q(n79) );
  INV3 U67 ( .A(n80), .Q(n786) );
  NAND22 U68 ( .A(n51), .B(n42), .Q(n80) );
  INV3 U69 ( .A(n81), .Q(n785) );
  NAND22 U70 ( .A(n53), .B(n42), .Q(n81) );
  INV3 U71 ( .A(n82), .Q(n784) );
  NAND22 U72 ( .A(n55), .B(n42), .Q(n82) );
  INV3 U73 ( .A(n40), .Q(n790) );
  NAND22 U74 ( .A(n41), .B(n42), .Q(n40) );
  INV3 U75 ( .A(n43), .Q(n789) );
  NAND22 U76 ( .A(n44), .B(n42), .Q(n43) );
  INV3 U77 ( .A(n45), .Q(n788) );
  NAND22 U78 ( .A(n46), .B(n42), .Q(n45) );
  INV3 U79 ( .A(n47), .Q(n782) );
  NAND22 U80 ( .A(n48), .B(n49), .Q(n47) );
  INV3 U81 ( .A(n56), .Q(n778) );
  NAND22 U82 ( .A(n48), .B(n57), .Q(n56) );
  INV3 U83 ( .A(n58), .Q(n777) );
  NAND22 U84 ( .A(n48), .B(n41), .Q(n58) );
  INV3 U85 ( .A(n59), .Q(n776) );
  NAND22 U86 ( .A(n48), .B(n44), .Q(n59) );
  INV3 U87 ( .A(n50), .Q(n781) );
  NAND22 U88 ( .A(n51), .B(n48), .Q(n50) );
  INV3 U89 ( .A(n52), .Q(n780) );
  NAND22 U90 ( .A(n53), .B(n48), .Q(n52) );
  INV3 U91 ( .A(n54), .Q(n779) );
  NAND22 U92 ( .A(n55), .B(n48), .Q(n54) );
  INV3 U93 ( .A(n61), .Q(n807) );
  NAND22 U94 ( .A(n62), .B(n49), .Q(n61) );
  INV3 U95 ( .A(n63), .Q(n806) );
  NAND22 U96 ( .A(n62), .B(n51), .Q(n63) );
  INV3 U97 ( .A(n64), .Q(n805) );
  NAND22 U98 ( .A(n62), .B(n53), .Q(n64) );
  INV3 U99 ( .A(n65), .Q(n804) );
  NAND22 U100 ( .A(n62), .B(n55), .Q(n65) );
  INV3 U101 ( .A(n66), .Q(n803) );
  NAND22 U102 ( .A(n62), .B(n57), .Q(n66) );
  INV3 U103 ( .A(n67), .Q(n802) );
  NAND22 U104 ( .A(n62), .B(n41), .Q(n67) );
  INV3 U105 ( .A(n68), .Q(n801) );
  NAND22 U106 ( .A(n62), .B(n44), .Q(n68) );
  INV3 U107 ( .A(n69), .Q(n800) );
  NAND22 U108 ( .A(n62), .B(n46), .Q(n69) );
  INV3 U109 ( .A(n70), .Q(n799) );
  NAND22 U110 ( .A(n71), .B(n49), .Q(n70) );
  INV3 U111 ( .A(n72), .Q(n798) );
  NAND22 U112 ( .A(n71), .B(n51), .Q(n72) );
  INV3 U113 ( .A(n73), .Q(n797) );
  NAND22 U114 ( .A(n71), .B(n53), .Q(n73) );
  INV3 U115 ( .A(n74), .Q(n796) );
  NAND22 U116 ( .A(n71), .B(n55), .Q(n74) );
  INV3 U117 ( .A(n75), .Q(n795) );
  NAND22 U118 ( .A(n71), .B(n57), .Q(n75) );
  INV3 U119 ( .A(n76), .Q(n794) );
  NAND22 U120 ( .A(n71), .B(n41), .Q(n76) );
  INV3 U121 ( .A(n77), .Q(n793) );
  NAND22 U122 ( .A(n71), .B(n44), .Q(n77) );
  INV3 U123 ( .A(n78), .Q(n792) );
  NAND22 U124 ( .A(n71), .B(n46), .Q(n78) );
  BUF2 U125 ( .A(n748), .Q(n746) );
  BUF2 U126 ( .A(n748), .Q(n747) );
  BUF2 U127 ( .A(i_addr_Rt[0]), .Q(n399) );
  BUF2 U128 ( .A(i_addr_Rt[0]), .Q(n400) );
  BUF2 U129 ( .A(i_addr_Rt[0]), .Q(n401) );
  BUF2 U130 ( .A(i_addr_Rs[0]), .Q(n763) );
  BUF2 U131 ( .A(i_addr_Rs[0]), .Q(n764) );
  BUF2 U132 ( .A(i_addr_Rs[0]), .Q(n765) );
  BUF2 U133 ( .A(i_addr_Rt[1]), .Q(n376) );
  BUF2 U134 ( .A(i_addr_Rt[1]), .Q(n375) );
  BUF2 U135 ( .A(i_addr_Rt[1]), .Q(n374) );
  BUF2 U136 ( .A(i_addr_Rs[1]), .Q(n732) );
  BUF2 U137 ( .A(i_addr_Rs[1]), .Q(n731) );
  BUF2 U138 ( .A(i_addr_Rs[1]), .Q(n730) );
  NOR31 U139 ( .A(n791), .B(i_addr_Rd[3]), .C(n812), .Q(n42) );
  NOR31 U140 ( .A(i_addr_Rd[3]), .B(i_addr_Rd[4]), .C(n812), .Q(n62) );
  NOR31 U141 ( .A(n812), .B(i_addr_Rd[4]), .C(n808), .Q(n71) );
  MUX22 U142 ( .A(n407), .B(n402), .S(n722), .Q(o_data_Rs[0]) );
  IMUX40 U143 ( .A(n403), .B(n404), .C(n405), .D(n406), .S0(n723), .S1(
        i_addr_Rs[2]), .Q(n402) );
  IMUX40 U144 ( .A(n408), .B(n409), .C(n410), .D(n411), .S0(n723), .S1(n727), 
        .Q(n407) );
  MUX22 U145 ( .A(n16), .B(n11), .S(n365), .Q(o_data_Rt[1]) );
  IMUX40 U146 ( .A(n17), .B(n18), .C(n19), .D(n20), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n16) );
  IMUX40 U147 ( .A(n12), .B(n13), .C(n14), .D(n15), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n11) );
  IMUX40 U148 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n385), .S1(n381), .Q(n17) );
  MUX22 U149 ( .A(n26), .B(n21), .S(n365), .Q(o_data_Rt[2]) );
  IMUX40 U150 ( .A(n27), .B(n28), .C(n29), .D(n30), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n26) );
  IMUX40 U151 ( .A(n22), .B(n23), .C(n24), .D(n25), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n21) );
  IMUX40 U152 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n386), .S1(i_addr_Rt[1]), .Q(n27) );
  MUX22 U153 ( .A(n36), .B(n31), .S(n365), .Q(o_data_Rt[3]) );
  IMUX40 U154 ( .A(n37), .B(n38), .C(n83), .D(n84), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n36) );
  IMUX40 U155 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n31) );
  IMUX40 U156 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n387), .S1(n381), .Q(n37) );
  MUX22 U157 ( .A(n90), .B(n85), .S(n365), .Q(o_data_Rt[4]) );
  IMUX40 U158 ( .A(n91), .B(n92), .C(n93), .D(n94), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n90) );
  IMUX40 U159 ( .A(n86), .B(n87), .C(n88), .D(n89), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n85) );
  IMUX40 U160 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n387), .S1(n382), .Q(n91) );
  MUX22 U161 ( .A(n100), .B(n95), .S(n365), .Q(o_data_Rt[5]) );
  IMUX40 U162 ( .A(n101), .B(n102), .C(n103), .D(n104), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n100) );
  IMUX40 U163 ( .A(n96), .B(n97), .C(n98), .D(n99), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n95) );
  IMUX40 U164 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n388), .S1(n384), .Q(n101) );
  MUX22 U165 ( .A(n110), .B(n105), .S(i_addr_Rt[4]), .Q(o_data_Rt[6]) );
  IMUX40 U166 ( .A(n111), .B(n112), .C(n113), .D(n114), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n110) );
  IMUX40 U167 ( .A(n106), .B(n107), .C(n108), .D(n109), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n105) );
  IMUX40 U168 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n389), .S1(n377), .Q(n111) );
  MUX22 U169 ( .A(n120), .B(n115), .S(i_addr_Rt[4]), .Q(o_data_Rt[7]) );
  IMUX40 U170 ( .A(n121), .B(n122), .C(n123), .D(n124), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n120) );
  IMUX40 U171 ( .A(n116), .B(n117), .C(n118), .D(n119), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n115) );
  IMUX40 U172 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n389), .S1(n378), .Q(n121) );
  MUX22 U173 ( .A(n130), .B(n125), .S(i_addr_Rt[4]), .Q(o_data_Rt[8]) );
  IMUX40 U174 ( .A(n131), .B(n132), .C(n133), .D(n134), .S0(n368), .S1(
        i_addr_Rt[2]), .Q(n130) );
  IMUX40 U175 ( .A(n126), .B(n127), .C(n128), .D(n129), .S0(n368), .S1(
        i_addr_Rt[2]), .Q(n125) );
  IMUX40 U176 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n390), .S1(i_addr_Rt[1]), .Q(n131) );
  MUX22 U177 ( .A(n140), .B(n135), .S(i_addr_Rt[4]), .Q(o_data_Rt[9]) );
  IMUX40 U178 ( .A(n141), .B(n142), .C(n143), .D(n144), .S0(n368), .S1(n370), 
        .Q(n140) );
  IMUX40 U179 ( .A(n136), .B(n137), .C(n138), .D(n139), .S0(n368), .S1(
        i_addr_Rt[2]), .Q(n135) );
  IMUX40 U180 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n391), .S1(n379), .Q(n141) );
  MUX22 U181 ( .A(n150), .B(n145), .S(i_addr_Rt[4]), .Q(o_data_Rt[10]) );
  IMUX40 U182 ( .A(n151), .B(n152), .C(n153), .D(n154), .S0(n368), .S1(n370), 
        .Q(n150) );
  IMUX40 U183 ( .A(n146), .B(n147), .C(n148), .D(n149), .S0(n368), .S1(n370), 
        .Q(n145) );
  IMUX40 U184 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n391), .S1(n380), .Q(n151) );
  MUX22 U185 ( .A(n160), .B(n155), .S(i_addr_Rt[4]), .Q(o_data_Rt[11]) );
  IMUX40 U186 ( .A(n161), .B(n162), .C(n163), .D(n164), .S0(n368), .S1(n370), 
        .Q(n160) );
  IMUX40 U187 ( .A(n156), .B(n157), .C(n158), .D(n159), .S0(n368), .S1(n370), 
        .Q(n155) );
  IMUX40 U188 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n394), .S1(n381), .Q(n161) );
  MUX22 U189 ( .A(n170), .B(n165), .S(i_addr_Rt[4]), .Q(o_data_Rt[12]) );
  IMUX40 U190 ( .A(n171), .B(n172), .C(n173), .D(n174), .S0(n368), .S1(n370), 
        .Q(n170) );
  IMUX40 U191 ( .A(n166), .B(n167), .C(n168), .D(n169), .S0(n368), .S1(n370), 
        .Q(n165) );
  IMUX40 U192 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        i_addr_Rt[0]), .S1(n382), .Q(n171) );
  MUX22 U193 ( .A(n180), .B(n175), .S(i_addr_Rt[4]), .Q(o_data_Rt[13]) );
  IMUX40 U194 ( .A(n181), .B(n182), .C(n183), .D(n184), .S0(n368), .S1(n370), 
        .Q(n180) );
  IMUX40 U195 ( .A(n176), .B(n177), .C(n178), .D(n179), .S0(n368), .S1(n370), 
        .Q(n175) );
  IMUX40 U196 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        i_addr_Rt[0]), .S1(n382), .Q(n181) );
  MUX22 U197 ( .A(n190), .B(n185), .S(i_addr_Rt[4]), .Q(o_data_Rt[14]) );
  IMUX40 U198 ( .A(n191), .B(n192), .C(n193), .D(n194), .S0(n369), .S1(n371), 
        .Q(n190) );
  IMUX40 U199 ( .A(n186), .B(n187), .C(n188), .D(n189), .S0(n369), .S1(n371), 
        .Q(n185) );
  IMUX40 U200 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n392), .S1(n374), .Q(n191) );
  MUX22 U201 ( .A(n200), .B(n195), .S(i_addr_Rt[4]), .Q(o_data_Rt[15]) );
  IMUX40 U202 ( .A(n201), .B(n202), .C(n203), .D(n204), .S0(n369), .S1(n371), 
        .Q(n200) );
  IMUX40 U203 ( .A(n196), .B(n197), .C(n198), .D(n199), .S0(n369), .S1(n371), 
        .Q(n195) );
  IMUX40 U204 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n393), .S1(n384), .Q(n201) );
  MUX22 U205 ( .A(n210), .B(n205), .S(i_addr_Rt[4]), .Q(o_data_Rt[16]) );
  IMUX40 U206 ( .A(n211), .B(n212), .C(n213), .D(n214), .S0(n369), .S1(n371), 
        .Q(n210) );
  IMUX40 U207 ( .A(n206), .B(n207), .C(n208), .D(n209), .S0(n369), .S1(n371), 
        .Q(n205) );
  IMUX40 U208 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n393), .S1(n378), .Q(n211) );
  MUX22 U209 ( .A(n220), .B(n215), .S(i_addr_Rt[4]), .Q(o_data_Rt[17]) );
  IMUX40 U210 ( .A(n221), .B(n222), .C(n223), .D(n224), .S0(n369), .S1(n371), 
        .Q(n220) );
  IMUX40 U211 ( .A(n216), .B(n217), .C(n218), .D(n219), .S0(n369), .S1(n371), 
        .Q(n215) );
  IMUX40 U212 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n394), .S1(n384), .Q(n221) );
  MUX22 U213 ( .A(n230), .B(n225), .S(i_addr_Rt[4]), .Q(o_data_Rt[18]) );
  IMUX40 U214 ( .A(n231), .B(n232), .C(n233), .D(n234), .S0(n369), .S1(n372), 
        .Q(n230) );
  IMUX40 U215 ( .A(n226), .B(n227), .C(n228), .D(n229), .S0(n369), .S1(n371), 
        .Q(n225) );
  IMUX40 U216 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n401), .S1(n383), .Q(n231) );
  MUX22 U217 ( .A(n240), .B(n235), .S(n365), .Q(o_data_Rt[19]) );
  IMUX40 U218 ( .A(n241), .B(n242), .C(n243), .D(n244), .S0(n369), .S1(n372), 
        .Q(n240) );
  IMUX40 U219 ( .A(n236), .B(n237), .C(n238), .D(n239), .S0(n369), .S1(n372), 
        .Q(n235) );
  IMUX40 U220 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n401), .S1(n380), .Q(n241) );
  MUX22 U221 ( .A(n250), .B(n245), .S(n365), .Q(o_data_Rt[20]) );
  IMUX40 U222 ( .A(n251), .B(n252), .C(n253), .D(n254), .S0(i_addr_Rt[3]), 
        .S1(n372), .Q(n250) );
  IMUX40 U223 ( .A(n246), .B(n247), .C(n248), .D(n249), .S0(i_addr_Rt[3]), 
        .S1(n372), .Q(n245) );
  IMUX40 U224 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n394), .S1(n376), .Q(n251) );
  MUX22 U225 ( .A(n260), .B(n255), .S(n365), .Q(o_data_Rt[21]) );
  IMUX40 U226 ( .A(n261), .B(n262), .C(n263), .D(n264), .S0(i_addr_Rt[3]), 
        .S1(n372), .Q(n260) );
  IMUX40 U227 ( .A(n256), .B(n257), .C(n258), .D(n259), .S0(i_addr_Rt[3]), 
        .S1(n372), .Q(n255) );
  IMUX40 U228 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n394), .S1(n383), .Q(n261) );
  MUX22 U229 ( .A(n270), .B(n265), .S(n365), .Q(o_data_Rt[22]) );
  IMUX40 U230 ( .A(n271), .B(n272), .C(n273), .D(n274), .S0(i_addr_Rt[3]), 
        .S1(n372), .Q(n270) );
  IMUX40 U231 ( .A(n266), .B(n267), .C(n268), .D(n269), .S0(i_addr_Rt[3]), 
        .S1(n372), .Q(n265) );
  IMUX40 U232 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n390), .S1(n383), .Q(n271) );
  MUX22 U233 ( .A(n280), .B(n275), .S(n365), .Q(o_data_Rt[23]) );
  IMUX40 U234 ( .A(n281), .B(n282), .C(n283), .D(n284), .S0(i_addr_Rt[3]), 
        .S1(n373), .Q(n280) );
  IMUX40 U235 ( .A(n276), .B(n277), .C(n278), .D(n279), .S0(i_addr_Rt[3]), 
        .S1(n373), .Q(n275) );
  IMUX40 U236 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n398), .S1(n379), .Q(n281) );
  MUX22 U237 ( .A(n290), .B(n285), .S(n365), .Q(o_data_Rt[24]) );
  IMUX40 U238 ( .A(n291), .B(n292), .C(n293), .D(n294), .S0(i_addr_Rt[3]), 
        .S1(n373), .Q(n290) );
  IMUX40 U239 ( .A(n286), .B(n287), .C(n288), .D(n289), .S0(i_addr_Rt[3]), 
        .S1(n373), .Q(n285) );
  IMUX40 U240 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n395), .S1(n381), .Q(n291) );
  MUX22 U241 ( .A(n300), .B(n295), .S(n365), .Q(o_data_Rt[25]) );
  IMUX40 U242 ( .A(n301), .B(n302), .C(n303), .D(n304), .S0(i_addr_Rt[3]), 
        .S1(n373), .Q(n300) );
  IMUX40 U243 ( .A(n296), .B(n297), .C(n298), .D(n299), .S0(i_addr_Rt[3]), 
        .S1(n373), .Q(n295) );
  IMUX40 U244 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n395), .S1(n384), .Q(n301) );
  MUX22 U245 ( .A(n310), .B(n305), .S(i_addr_Rt[4]), .Q(o_data_Rt[26]) );
  IMUX40 U246 ( .A(n311), .B(n312), .C(n313), .D(n314), .S0(n366), .S1(n373), 
        .Q(n310) );
  IMUX40 U247 ( .A(n306), .B(n307), .C(n308), .D(n309), .S0(n366), .S1(n373), 
        .Q(n305) );
  IMUX40 U248 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n401), .S1(n384), .Q(n311) );
  MUX22 U249 ( .A(n320), .B(n315), .S(i_addr_Rt[4]), .Q(o_data_Rt[27]) );
  IMUX40 U250 ( .A(n321), .B(n322), .C(n323), .D(n324), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n320) );
  IMUX40 U251 ( .A(n316), .B(n317), .C(n318), .D(n319), .S0(n366), .S1(n373), 
        .Q(n315) );
  IMUX40 U252 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n396), .S1(n379), .Q(n321) );
  MUX22 U253 ( .A(n330), .B(n325), .S(i_addr_Rt[4]), .Q(o_data_Rt[28]) );
  IMUX40 U254 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n330) );
  IMUX40 U255 ( .A(n326), .B(n327), .C(n328), .D(n329), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n325) );
  IMUX40 U256 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n396), .S1(n380), .Q(n331) );
  MUX22 U257 ( .A(n340), .B(n335), .S(i_addr_Rt[4]), .Q(o_data_Rt[29]) );
  IMUX40 U258 ( .A(n341), .B(n342), .C(n343), .D(n344), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n340) );
  IMUX40 U259 ( .A(n336), .B(n337), .C(n338), .D(n339), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n335) );
  IMUX40 U260 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n397), .S1(i_addr_Rt[1]), .Q(n341) );
  MUX22 U261 ( .A(n350), .B(n345), .S(i_addr_Rt[4]), .Q(o_data_Rt[30]) );
  IMUX40 U262 ( .A(n351), .B(n352), .C(n353), .D(n354), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n350) );
  IMUX40 U263 ( .A(n346), .B(n347), .C(n348), .D(n349), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n345) );
  IMUX40 U264 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n398), .S1(n381), .Q(n351) );
  MUX22 U265 ( .A(n360), .B(n355), .S(i_addr_Rt[4]), .Q(o_data_Rt[31]) );
  IMUX40 U266 ( .A(n361), .B(n362), .C(n363), .D(n364), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n360) );
  IMUX40 U267 ( .A(n356), .B(n357), .C(n358), .D(n359), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n355) );
  IMUX40 U268 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n398), .S1(n380), .Q(n361) );
  MUX22 U269 ( .A(n537), .B(n532), .S(i_addr_Rs[4]), .Q(o_data_Rs[13]) );
  IMUX40 U270 ( .A(n538), .B(n539), .C(n540), .D(n541), .S0(n725), .S1(n729), 
        .Q(n537) );
  IMUX40 U271 ( .A(n533), .B(n534), .C(n535), .D(n536), .S0(n724), .S1(n729), 
        .Q(n532) );
  IMUX40 U272 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n749), .S1(i_addr_Rs[1]), .Q(n538) );
  MUX22 U273 ( .A(n547), .B(n542), .S(i_addr_Rs[4]), .Q(o_data_Rs[14]) );
  IMUX40 U274 ( .A(n548), .B(n549), .C(n550), .D(n551), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n547) );
  IMUX40 U275 ( .A(n543), .B(n544), .C(n545), .D(n546), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n542) );
  IMUX40 U276 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n755), .S1(n733), .Q(n548) );
  MUX22 U277 ( .A(n557), .B(n552), .S(i_addr_Rs[4]), .Q(o_data_Rs[15]) );
  IMUX40 U278 ( .A(n558), .B(n559), .C(n560), .D(n561), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n557) );
  IMUX40 U279 ( .A(n553), .B(n554), .C(n555), .D(n556), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n552) );
  IMUX40 U280 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n756), .S1(n734), .Q(n558) );
  MUX22 U281 ( .A(n567), .B(n562), .S(i_addr_Rs[4]), .Q(o_data_Rs[16]) );
  IMUX40 U282 ( .A(n568), .B(n569), .C(n570), .D(n571), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n567) );
  IMUX40 U283 ( .A(n563), .B(n564), .C(n565), .D(n566), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n562) );
  IMUX40 U284 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n756), .S1(n735), .Q(n568) );
  MUX22 U285 ( .A(n577), .B(n572), .S(i_addr_Rs[4]), .Q(o_data_Rs[17]) );
  IMUX40 U286 ( .A(n578), .B(n579), .C(n580), .D(n581), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n577) );
  IMUX40 U287 ( .A(n573), .B(n574), .C(n575), .D(n576), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n572) );
  IMUX40 U288 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n755), .S1(n736), .Q(n578) );
  MUX22 U289 ( .A(n587), .B(n582), .S(i_addr_Rs[4]), .Q(o_data_Rs[18]) );
  IMUX40 U290 ( .A(n588), .B(n589), .C(n590), .D(n591), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n587) );
  IMUX40 U291 ( .A(n583), .B(n584), .C(n585), .D(n586), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n582) );
  IMUX40 U292 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n757), .S1(n737), .Q(n588) );
  MUX22 U293 ( .A(n597), .B(n592), .S(i_addr_Rs[4]), .Q(o_data_Rs[19]) );
  IMUX40 U294 ( .A(n598), .B(n599), .C(n600), .D(n601), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n597) );
  IMUX40 U295 ( .A(n593), .B(n594), .C(n595), .D(n596), .S0(n724), .S1(
        i_addr_Rs[2]), .Q(n592) );
  IMUX40 U296 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n757), .S1(n737), .Q(n598) );
  MUX22 U297 ( .A(n607), .B(n602), .S(i_addr_Rs[4]), .Q(o_data_Rs[20]) );
  IMUX40 U298 ( .A(n608), .B(n609), .C(n610), .D(n611), .S0(n725), .S1(
        i_addr_Rs[2]), .Q(n607) );
  IMUX40 U299 ( .A(n603), .B(n604), .C(n605), .D(n606), .S0(n725), .S1(
        i_addr_Rs[2]), .Q(n602) );
  IMUX40 U300 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n758), .S1(n738), .Q(n608) );
  MUX22 U301 ( .A(n617), .B(n612), .S(i_addr_Rs[4]), .Q(o_data_Rs[21]) );
  IMUX40 U302 ( .A(n618), .B(n619), .C(n620), .D(n621), .S0(n725), .S1(
        i_addr_Rs[2]), .Q(n617) );
  IMUX40 U303 ( .A(n613), .B(n614), .C(n615), .D(n616), .S0(n725), .S1(
        i_addr_Rs[2]), .Q(n612) );
  IMUX40 U304 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n759), .S1(n739), .Q(n618) );
  MUX22 U305 ( .A(n627), .B(n622), .S(i_addr_Rs[4]), .Q(o_data_Rs[22]) );
  IMUX40 U306 ( .A(n628), .B(n629), .C(n630), .D(n631), .S0(n725), .S1(
        i_addr_Rs[2]), .Q(n627) );
  IMUX40 U307 ( .A(n623), .B(n624), .C(n625), .D(n626), .S0(n725), .S1(
        i_addr_Rs[2]), .Q(n622) );
  IMUX40 U308 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n759), .S1(n739), .Q(n628) );
  MUX22 U309 ( .A(n637), .B(n632), .S(i_addr_Rs[4]), .Q(o_data_Rs[23]) );
  IMUX40 U310 ( .A(n638), .B(n639), .C(n640), .D(n641), .S0(n725), .S1(
        i_addr_Rs[2]), .Q(n637) );
  IMUX40 U311 ( .A(n633), .B(n634), .C(n635), .D(n636), .S0(n725), .S1(n727), 
        .Q(n632) );
  IMUX40 U312 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n764), .S1(n740), .Q(n638) );
  MUX22 U313 ( .A(n647), .B(n642), .S(i_addr_Rs[4]), .Q(o_data_Rs[24]) );
  IMUX40 U314 ( .A(n648), .B(n649), .C(n650), .D(n651), .S0(n725), .S1(
        i_addr_Rs[2]), .Q(n647) );
  IMUX40 U315 ( .A(n643), .B(n644), .C(n645), .D(n646), .S0(n725), .S1(n728), 
        .Q(n642) );
  IMUX40 U316 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n761), .S1(n741), .Q(n648) );
  MUX22 U317 ( .A(n657), .B(n652), .S(i_addr_Rs[4]), .Q(o_data_Rs[25]) );
  IMUX40 U318 ( .A(n658), .B(n659), .C(n660), .D(n661), .S0(n725), .S1(
        i_addr_Rs[2]), .Q(n657) );
  IMUX40 U319 ( .A(n653), .B(n654), .C(n655), .D(n656), .S0(n725), .S1(n729), 
        .Q(n652) );
  IMUX40 U320 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n757), .S1(n742), .Q(n658) );
  MUX22 U321 ( .A(n667), .B(n662), .S(i_addr_Rs[4]), .Q(o_data_Rs[26]) );
  IMUX40 U322 ( .A(n668), .B(n669), .C(n670), .D(n671), .S0(n726), .S1(
        i_addr_Rs[2]), .Q(n667) );
  IMUX40 U323 ( .A(n663), .B(n664), .C(n665), .D(n666), .S0(n726), .S1(
        i_addr_Rs[2]), .Q(n662) );
  IMUX40 U324 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n751), .S1(n743), .Q(n668) );
  MUX22 U325 ( .A(n677), .B(n672), .S(i_addr_Rs[4]), .Q(o_data_Rs[27]) );
  IMUX40 U326 ( .A(n678), .B(n679), .C(n680), .D(n681), .S0(n726), .S1(n727), 
        .Q(n677) );
  IMUX40 U327 ( .A(n673), .B(n674), .C(n675), .D(n676), .S0(n726), .S1(n727), 
        .Q(n672) );
  IMUX40 U328 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n760), .S1(n744), .Q(n678) );
  MUX22 U329 ( .A(n687), .B(n682), .S(i_addr_Rs[4]), .Q(o_data_Rs[28]) );
  IMUX40 U330 ( .A(n688), .B(n689), .C(n690), .D(n691), .S0(n726), .S1(n728), 
        .Q(n687) );
  IMUX40 U331 ( .A(n683), .B(n684), .C(n685), .D(n686), .S0(n726), .S1(
        i_addr_Rs[2]), .Q(n682) );
  IMUX40 U332 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n760), .S1(n745), .Q(n688) );
  MUX22 U333 ( .A(n697), .B(n692), .S(i_addr_Rs[4]), .Q(o_data_Rs[29]) );
  IMUX40 U334 ( .A(n698), .B(n699), .C(n700), .D(n701), .S0(n726), .S1(n729), 
        .Q(n697) );
  IMUX40 U335 ( .A(n693), .B(n694), .C(n695), .D(n696), .S0(n726), .S1(n728), 
        .Q(n692) );
  IMUX40 U336 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n761), .S1(n746), .Q(n700) );
  MUX22 U337 ( .A(n707), .B(n702), .S(i_addr_Rs[4]), .Q(o_data_Rs[30]) );
  IMUX40 U338 ( .A(n708), .B(n709), .C(n710), .D(n711), .S0(n726), .S1(
        i_addr_Rs[2]), .Q(n707) );
  IMUX40 U339 ( .A(n703), .B(n704), .C(n705), .D(n706), .S0(n726), .S1(
        i_addr_Rs[2]), .Q(n702) );
  IMUX40 U340 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n762), .S1(n746), .Q(n710) );
  MUX22 U341 ( .A(n717), .B(n712), .S(i_addr_Rs[4]), .Q(o_data_Rs[31]) );
  IMUX40 U342 ( .A(n718), .B(n719), .C(n720), .D(n721), .S0(n726), .S1(
        i_addr_Rs[2]), .Q(n717) );
  IMUX40 U343 ( .A(n713), .B(n714), .C(n715), .D(n716), .S0(n726), .S1(n729), 
        .Q(n712) );
  IMUX40 U344 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n762), .S1(n747), .Q(n720) );
  NOR31 U345 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n809), .Q(n57) );
  NOR31 U346 ( .A(n809), .B(i_addr_Rd[1]), .C(n811), .Q(n41) );
  NOR31 U347 ( .A(n809), .B(i_addr_Rd[0]), .C(n810), .Q(n44) );
  NOR31 U348 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(i_addr_Rd[0]), .Q(n49)
         );
  NOR31 U349 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(n811), .Q(n51) );
  NOR31 U350 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[2]), .C(n810), .Q(n53) );
  NOR31 U351 ( .A(n811), .B(i_addr_Rd[2]), .C(n810), .Q(n55) );
  IMUX40 U352 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n385), .S1(n374), .Q(n10) );
  IMUX40 U353 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n8) );
  IMUX40 U354 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n385), .S1(i_addr_Rt[1]), .Q(n7) );
  IMUX40 U355 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(i_addr_Rt[0]), .S1(n384), .Q(n5) );
  IMUX40 U356 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(i_addr_Rt[0]), .S1(n383), .Q(n3) );
  IMUX40 U357 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(i_addr_Rt[0]), .S1(n384), .Q(n2) );
  IMUX40 U358 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n385), .S1(n383), .Q(n15) );
  IMUX40 U359 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n13) );
  IMUX40 U360 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n12) );
  IMUX40 U361 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n385), .S1(n384), .Q(n20) );
  IMUX40 U362 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n18) );
  IMUX40 U363 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n386), .S1(n382), .Q(n25) );
  IMUX40 U364 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n386), .S1(n384), .Q(n23) );
  IMUX40 U365 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n386), .S1(n380), .Q(n22) );
  IMUX40 U366 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n386), .S1(n379), .Q(n30) );
  IMUX40 U367 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n386), .S1(n379), .Q(n28) );
  IMUX40 U368 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n386), .S1(n378), .Q(n35) );
  IMUX40 U369 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n386), .S1(i_addr_Rt[1]), .Q(n33) );
  IMUX40 U370 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n386), .S1(i_addr_Rt[1]), .Q(n32) );
  IMUX40 U371 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n387), .S1(i_addr_Rt[1]), .Q(n84) );
  IMUX40 U372 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n387), .S1(i_addr_Rt[1]), .Q(n38) );
  IMUX40 U373 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n387), .S1(n380), .Q(n89) );
  IMUX40 U374 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n387), .S1(n374), .Q(n87) );
  IMUX40 U375 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n387), .S1(n380), .Q(n86) );
  IMUX40 U376 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n387), .S1(n374), .Q(n94) );
  IMUX40 U377 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n387), .S1(n379), .Q(n92) );
  IMUX40 U378 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n388), .S1(n381), .Q(n99) );
  IMUX40 U379 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n388), .S1(n374), .Q(n97) );
  IMUX40 U380 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n388), .S1(n377), .Q(n96) );
  IMUX40 U381 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n388), .S1(n384), .Q(n104) );
  IMUX40 U382 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n388), .S1(n375), .Q(n102) );
  IMUX40 U383 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n388), .S1(n384), .Q(n109) );
  IMUX40 U384 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n388), .S1(n377), .Q(n107) );
  IMUX40 U385 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n388), .S1(n377), .Q(n106) );
  IMUX40 U386 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n389), .S1(n377), .Q(n114) );
  IMUX40 U387 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n389), .S1(n377), .Q(n112) );
  IMUX40 U388 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n389), .S1(n377), .Q(n119) );
  IMUX40 U389 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n389), .S1(n377), .Q(n117) );
  IMUX40 U390 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n389), .S1(n378), .Q(n116) );
  IMUX40 U391 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n389), .S1(n378), .Q(n124) );
  IMUX40 U392 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n389), .S1(n378), .Q(n122) );
  IMUX40 U393 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n390), .S1(n378), .Q(n129) );
  IMUX40 U394 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n390), .S1(n378), .Q(n127) );
  IMUX40 U395 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n390), .S1(i_addr_Rt[1]), .Q(n126) );
  IMUX40 U396 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n390), .S1(i_addr_Rt[1]), .Q(n134) );
  IMUX40 U397 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n390), .S1(i_addr_Rt[1]), .Q(n132) );
  IMUX40 U398 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n390), .S1(n375), .Q(n139) );
  IMUX40 U399 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n390), .S1(i_addr_Rt[1]), .Q(n137) );
  IMUX40 U400 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n390), .S1(i_addr_Rt[1]), .Q(n136) );
  IMUX40 U401 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n391), .S1(n379), .Q(n144) );
  IMUX40 U402 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n391), .S1(n379), .Q(n142) );
  IMUX40 U403 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n391), .S1(n379), .Q(n149) );
  IMUX40 U404 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n391), .S1(n379), .Q(n147) );
  IMUX40 U405 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n391), .S1(n379), .Q(n146) );
  IMUX40 U406 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n391), .S1(n379), .Q(n154) );
  IMUX40 U407 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n391), .S1(n380), .Q(n152) );
  IMUX40 U408 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n401), .S1(n380), .Q(n159) );
  IMUX40 U409 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n393), .S1(n380), .Q(n157) );
  IMUX40 U410 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n401), .S1(n380), .Q(n156) );
  IMUX40 U411 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n394), .S1(n380), .Q(n164) );
  IMUX40 U412 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n393), .S1(n380), .Q(n162) );
  IMUX40 U413 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n392), .S1(n381), .Q(n169) );
  IMUX40 U414 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n401), .S1(n381), .Q(n167) );
  IMUX40 U415 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n392), .S1(n381), .Q(n166) );
  IMUX40 U416 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(i_addr_Rt[0]), .S1(n381), .Q(n174) );
  IMUX40 U417 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(i_addr_Rt[0]), .S1(n381), .Q(n172) );
  IMUX40 U418 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n394), .S1(n382), .Q(n179) );
  IMUX40 U419 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n388), .S1(n382), .Q(n177) );
  IMUX40 U420 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(i_addr_Rt[0]), .S1(n382), .Q(n176) );
  IMUX40 U421 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(i_addr_Rt[0]), .S1(n382), .Q(n184) );
  IMUX40 U422 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(i_addr_Rt[0]), .S1(n382), .Q(n182) );
  IMUX40 U423 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n392), .S1(n374), .Q(n189) );
  IMUX40 U424 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n392), .S1(n374), .Q(n187) );
  IMUX40 U425 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n392), .S1(n374), .Q(n186) );
  IMUX40 U426 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n392), .S1(n374), .Q(n194) );
  IMUX40 U427 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n392), .S1(n374), .Q(n192) );
  IMUX40 U428 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n392), .S1(n374), .Q(n199) );
  IMUX40 U429 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n392), .S1(n377), .Q(n197) );
  IMUX40 U430 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n392), .S1(n379), .Q(n196) );
  IMUX40 U431 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n393), .S1(n374), .Q(n204) );
  IMUX40 U432 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n393), .S1(n380), .Q(n202) );
  IMUX40 U433 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n393), .S1(n377), .Q(n209) );
  IMUX40 U434 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n393), .S1(n377), .Q(n207) );
  IMUX40 U435 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n393), .S1(n382), .Q(n206) );
  IMUX40 U436 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n393), .S1(n384), .Q(n214) );
  IMUX40 U437 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n393), .S1(n374), .Q(n212) );
  IMUX40 U438 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n394), .S1(n376), .Q(n219) );
  IMUX40 U439 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n394), .S1(n377), .Q(n217) );
  IMUX40 U440 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n394), .S1(n375), .Q(n216) );
  IMUX40 U441 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n394), .S1(n377), .Q(n224) );
  IMUX40 U442 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n394), .S1(n381), .Q(n222) );
  IMUX40 U443 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n394), .S1(n384), .Q(n229) );
  IMUX40 U444 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n394), .S1(n384), .Q(n227) );
  IMUX40 U445 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n394), .S1(i_addr_Rt[1]), .Q(n226) );
  IMUX40 U446 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n401), .S1(n380), .Q(n234) );
  IMUX40 U447 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n401), .S1(n376), .Q(n232) );
  IMUX40 U448 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n401), .S1(n379), .Q(n239) );
  IMUX40 U449 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n401), .S1(n383), .Q(n237) );
  IMUX40 U450 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n401), .S1(n375), .Q(n236) );
  IMUX40 U451 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n401), .S1(n384), .Q(n244) );
  IMUX40 U452 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n401), .S1(n376), .Q(n242) );
  IMUX40 U453 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n398), .S1(n378), .Q(n249) );
  IMUX40 U454 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n388), .S1(n377), .Q(n247) );
  IMUX40 U455 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n393), .S1(n381), .Q(n246) );
  IMUX40 U456 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n400), .S1(n374), .Q(n254) );
  IMUX40 U457 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n386), .S1(n377), .Q(n252) );
  IMUX40 U458 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n392), .S1(n377), .Q(n259) );
  IMUX40 U459 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n393), .S1(i_addr_Rt[1]), .Q(n257) );
  IMUX40 U460 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n392), .S1(n379), .Q(n256) );
  IMUX40 U461 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n387), .S1(n384), .Q(n264) );
  IMUX40 U462 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n396), .S1(n382), .Q(n262) );
  IMUX40 U463 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n389), .S1(n383), .Q(n269) );
  IMUX40 U464 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n401), .S1(n383), .Q(n267) );
  IMUX40 U465 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n385), .S1(n383), .Q(n266) );
  IMUX40 U466 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n390), .S1(n383), .Q(n274) );
  IMUX40 U467 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n397), .S1(n383), .Q(n272) );
  IMUX40 U468 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n398), .S1(n379), .Q(n279) );
  IMUX40 U469 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n398), .S1(n382), .Q(n277) );
  IMUX40 U470 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n393), .S1(n377), .Q(n276) );
  IMUX40 U471 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n395), .S1(n384), .Q(n284) );
  IMUX40 U472 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n395), .S1(n384), .Q(n282) );
  IMUX40 U473 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n395), .S1(n374), .Q(n289) );
  IMUX40 U474 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n398), .S1(n377), .Q(n287) );
  IMUX40 U475 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n395), .S1(n375), .Q(n286) );
  IMUX40 U476 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n395), .S1(n382), .Q(n294) );
  IMUX40 U477 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n395), .S1(n378), .Q(n292) );
  IMUX40 U478 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n395), .S1(n380), .Q(n299) );
  IMUX40 U479 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n395), .S1(i_addr_Rt[1]), .Q(n297) );
  IMUX40 U480 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n395), .S1(n384), .Q(n296) );
  IMUX40 U481 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n395), .S1(n384), .Q(n304) );
  IMUX40 U482 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n395), .S1(n384), .Q(n302) );
  IMUX40 U483 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n396), .S1(n384), .Q(n309) );
  IMUX40 U484 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n385), .S1(n384), .Q(n307) );
  IMUX40 U485 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n394), .S1(n376), .Q(n306) );
  IMUX40 U486 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n399), .S1(n384), .Q(n314) );
  IMUX40 U487 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n400), .S1(n380), .Q(n312) );
  IMUX40 U488 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n392), .S1(n384), .Q(n319) );
  IMUX40 U489 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n397), .S1(n374), .Q(n317) );
  IMUX40 U490 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n393), .S1(n374), .Q(n316) );
  IMUX40 U491 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n396), .S1(n375), .Q(n324) );
  IMUX40 U492 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n396), .S1(n377), .Q(n322) );
  IMUX40 U493 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n396), .S1(n381), .Q(n329) );
  IMUX40 U494 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n396), .S1(n378), .Q(n327) );
  IMUX40 U495 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n396), .S1(n381), .Q(n326) );
  IMUX40 U496 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n396), .S1(i_addr_Rt[1]), .Q(n334) );
  IMUX40 U497 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n396), .S1(n374), .Q(n332) );
  IMUX40 U498 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n397), .S1(n374), .Q(n339) );
  IMUX40 U499 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n397), .S1(n374), .Q(n337) );
  IMUX40 U500 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n397), .S1(n374), .Q(n336) );
  IMUX40 U501 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n397), .S1(n374), .Q(n344) );
  IMUX40 U502 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n397), .S1(n374), .Q(n342) );
  IMUX40 U503 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n397), .S1(n382), .Q(n349) );
  IMUX40 U504 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n397), .S1(n374), .Q(n347) );
  IMUX40 U505 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n397), .S1(i_addr_Rt[1]), .Q(n346) );
  IMUX40 U506 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n398), .S1(n384), .Q(n354) );
  IMUX40 U507 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n398), .S1(i_addr_Rt[1]), .Q(n352) );
  IMUX40 U508 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n398), .S1(n374), .Q(n359) );
  IMUX40 U509 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n398), .S1(n374), .Q(n357) );
  IMUX40 U510 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n398), .S1(n374), .Q(n356) );
  IMUX40 U511 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n398), .S1(n382), .Q(n364) );
  IMUX40 U512 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n398), .S1(n378), .Q(n362) );
  IMUX40 U513 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n749), .S1(n747), .Q(n411) );
  IMUX40 U514 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n749), .S1(n748), .Q(n408) );
  IMUX40 U515 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n749), .S1(n731), .Q(n409) );
  IMUX40 U516 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(n759), .S1(n746), .Q(n406) );
  IMUX40 U517 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(n760), .S1(n732), .Q(n404) );
  IMUX40 U518 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(n755), .S1(n733), .Q(n403) );
  IMUX40 U519 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n749), .S1(i_addr_Rs[1]), .Q(n416) );
  IMUX40 U520 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n749), .S1(i_addr_Rs[1]), .Q(n414) );
  IMUX40 U521 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n749), .S1(n732), .Q(n413) );
  IMUX40 U522 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n749), .S1(i_addr_Rs[1]), .Q(n421) );
  IMUX40 U523 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n749), .S1(n748), .Q(n418) );
  IMUX40 U524 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n749), .S1(n732), .Q(n419) );
  IMUX40 U525 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n750), .S1(i_addr_Rs[1]), .Q(n426) );
  IMUX40 U526 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n750), .S1(n732), .Q(n424) );
  IMUX40 U527 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n750), .S1(n732), .Q(n423) );
  IMUX40 U528 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n750), .S1(n734), .Q(n431) );
  IMUX40 U529 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n750), .S1(i_addr_Rs[1]), .Q(n428) );
  IMUX40 U530 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n750), .S1(n734), .Q(n429) );
  IMUX40 U531 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n750), .S1(i_addr_Rs[1]), .Q(n436) );
  IMUX40 U532 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n750), .S1(i_addr_Rs[1]), .Q(n434) );
  IMUX40 U533 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n750), .S1(i_addr_Rs[1]), .Q(n433) );
  IMUX40 U534 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n751), .S1(n731), .Q(n441) );
  IMUX40 U535 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n751), .S1(n731), .Q(n439) );
  IMUX40 U536 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n751), .S1(n733), .Q(n438) );
  IMUX40 U537 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n751), .S1(n732), .Q(n446) );
  IMUX40 U538 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n751), .S1(n730), .Q(n444) );
  IMUX40 U539 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n751), .S1(n746), .Q(n443) );
  IMUX40 U540 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n751), .S1(n731), .Q(n451) );
  IMUX40 U541 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n751), .S1(n748), .Q(n449) );
  IMUX40 U542 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n751), .S1(n734), .Q(n448) );
  IMUX40 U543 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n752), .S1(n748), .Q(n456) );
  IMUX40 U544 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n752), .S1(n734), .Q(n454) );
  IMUX40 U545 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n752), .S1(n748), .Q(n453) );
  IMUX40 U546 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n752), .S1(n748), .Q(n461) );
  IMUX40 U547 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n752), .S1(n748), .Q(n459) );
  IMUX40 U548 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n752), .S1(i_addr_Rs[1]), .Q(n458) );
  IMUX40 U549 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n752), .S1(n748), .Q(n466) );
  IMUX40 U550 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n752), .S1(n731), .Q(n464) );
  IMUX40 U551 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n752), .S1(n731), .Q(n463) );
  IMUX40 U552 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n753), .S1(n738), .Q(n471) );
  IMUX40 U553 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n753), .S1(n738), .Q(n469) );
  IMUX40 U554 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n753), .S1(n730), .Q(n468) );
  IMUX40 U555 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n753), .S1(n730), .Q(n476) );
  IMUX40 U556 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n753), .S1(n738), .Q(n474) );
  IMUX40 U557 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n753), .S1(n733), .Q(n473) );
  IMUX40 U558 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n753), .S1(n734), .Q(n481) );
  IMUX40 U559 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n753), .S1(n733), .Q(n479) );
  IMUX40 U560 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n753), .S1(n733), .Q(n478) );
  IMUX40 U561 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n751), .S1(n732), .Q(n486) );
  IMUX40 U562 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n757), .S1(n733), .Q(n484) );
  IMUX40 U563 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n749), .S1(i_addr_Rs[1]), .Q(n483) );
  IMUX40 U564 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n758), .S1(i_addr_Rs[1]), .Q(n491) );
  IMUX40 U565 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n750), .S1(i_addr_Rs[1]), .Q(n489) );
  IMUX40 U566 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n764), .S1(i_addr_Rs[1]), .Q(n488) );
  IMUX40 U567 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n760), .S1(i_addr_Rs[1]), .Q(n496) );
  IMUX40 U568 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n753), .S1(i_addr_Rs[1]), .Q(n494) );
  IMUX40 U569 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n752), .S1(i_addr_Rs[1]), .Q(n493) );
  IMUX40 U570 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n760), .S1(n733), .Q(n501) );
  IMUX40 U571 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n751), .S1(i_addr_Rs[1]), .Q(n499) );
  IMUX40 U572 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n750), .S1(n734), .Q(n498) );
  IMUX40 U573 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n758), .S1(n731), .Q(n506) );
  IMUX40 U574 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n762), .S1(n733), .Q(n504) );
  IMUX40 U575 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n763), .S1(n730), .Q(n503) );
  IMUX40 U576 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n761), .S1(n732), .Q(n511) );
  IMUX40 U577 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n756), .S1(n730), .Q(n509) );
  IMUX40 U578 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n749), .S1(n734), .Q(n508) );
  IMUX40 U579 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n754), .S1(n734), .Q(n516) );
  IMUX40 U580 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n754), .S1(i_addr_Rs[1]), .Q(n514) );
  IMUX40 U581 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n754), .S1(n732), .Q(n513) );
  IMUX40 U582 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n754), .S1(n733), .Q(n521) );
  IMUX40 U583 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n754), .S1(i_addr_Rs[1]), .Q(n519) );
  IMUX40 U584 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n754), .S1(n738), .Q(n518) );
  IMUX40 U585 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n754), .S1(n733), .Q(n526) );
  IMUX40 U586 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n754), .S1(n734), .Q(n524) );
  IMUX40 U587 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n754), .S1(n734), .Q(n523) );
  IMUX40 U588 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n759), .S1(n730), .Q(n531) );
  IMUX40 U589 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n754), .S1(i_addr_Rs[1]), .Q(n529) );
  IMUX40 U590 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n757), .S1(i_addr_Rs[1]), .Q(n528) );
  IMUX40 U591 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n757), .S1(i_addr_Rs[1]), .Q(n536) );
  IMUX40 U592 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n758), .S1(i_addr_Rs[1]), .Q(n534) );
  IMUX40 U593 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n760), .S1(n730), .Q(n533) );
  IMUX40 U594 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n762), .S1(i_addr_Rs[1]), .Q(n541) );
  IMUX40 U595 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n753), .S1(n732), .Q(n539) );
  IMUX40 U596 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n755), .S1(n733), .Q(n546) );
  IMUX40 U597 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n755), .S1(n733), .Q(n544) );
  IMUX40 U598 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n755), .S1(n733), .Q(n543) );
  IMUX40 U599 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n755), .S1(n733), .Q(n551) );
  IMUX40 U600 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n755), .S1(n733), .Q(n549) );
  IMUX40 U601 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n755), .S1(n733), .Q(n556) );
  IMUX40 U602 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n755), .S1(n734), .Q(n554) );
  IMUX40 U603 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n755), .S1(n734), .Q(n553) );
  IMUX40 U604 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n756), .S1(n734), .Q(n561) );
  IMUX40 U605 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n756), .S1(n734), .Q(n559) );
  IMUX40 U606 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n756), .S1(n734), .Q(n566) );
  IMUX40 U607 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n756), .S1(n734), .Q(n564) );
  IMUX40 U608 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n756), .S1(n735), .Q(n563) );
  IMUX40 U609 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n756), .S1(n735), .Q(n571) );
  IMUX40 U610 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n756), .S1(n735), .Q(n569) );
  IMUX40 U611 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n749), .S1(n735), .Q(n576) );
  IMUX40 U612 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n750), .S1(n735), .Q(n574) );
  IMUX40 U613 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n754), .S1(n736), .Q(n573) );
  IMUX40 U614 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n764), .S1(n736), .Q(n581) );
  IMUX40 U615 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n762), .S1(n736), .Q(n579) );
  IMUX40 U616 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n750), .S1(n736), .Q(n586) );
  IMUX40 U617 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n751), .S1(n736), .Q(n584) );
  IMUX40 U618 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n758), .S1(n736), .Q(n583) );
  IMUX40 U619 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n757), .S1(n737), .Q(n591) );
  IMUX40 U620 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n757), .S1(n737), .Q(n589) );
  IMUX40 U621 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n757), .S1(n738), .Q(n596) );
  IMUX40 U622 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n757), .S1(n738), .Q(n594) );
  IMUX40 U623 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n757), .S1(n738), .Q(n593) );
  IMUX40 U624 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n757), .S1(n738), .Q(n601) );
  IMUX40 U625 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n757), .S1(n737), .Q(n599) );
  IMUX40 U626 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n758), .S1(n737), .Q(n606) );
  IMUX40 U627 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n758), .S1(n737), .Q(n604) );
  IMUX40 U628 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n758), .S1(n737), .Q(n603) );
  IMUX40 U629 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n758), .S1(n737), .Q(n611) );
  IMUX40 U630 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n758), .S1(n737), .Q(n609) );
  IMUX40 U631 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n758), .S1(n738), .Q(n616) );
  IMUX40 U632 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n758), .S1(n738), .Q(n614) );
  IMUX40 U633 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n758), .S1(n738), .Q(n613) );
  IMUX40 U634 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n759), .S1(n738), .Q(n621) );
  IMUX40 U635 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n759), .S1(n738), .Q(n619) );
  IMUX40 U636 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n759), .S1(n739), .Q(n626) );
  IMUX40 U637 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n759), .S1(n739), .Q(n624) );
  IMUX40 U638 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n759), .S1(n739), .Q(n623) );
  IMUX40 U639 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n759), .S1(n739), .Q(n631) );
  IMUX40 U640 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n759), .S1(n739), .Q(n629) );
  IMUX40 U641 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n764), .S1(n740), .Q(n636) );
  IMUX40 U642 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n764), .S1(n740), .Q(n634) );
  IMUX40 U643 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n764), .S1(n740), .Q(n633) );
  IMUX40 U644 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n764), .S1(n740), .Q(n641) );
  IMUX40 U645 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n764), .S1(n740), .Q(n639) );
  IMUX40 U646 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n764), .S1(n740), .Q(n646) );
  IMUX40 U647 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n764), .S1(n741), .Q(n644) );
  IMUX40 U648 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n764), .S1(n741), .Q(n643) );
  IMUX40 U649 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n749), .S1(n741), .Q(n651) );
  IMUX40 U650 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n761), .S1(n741), .Q(n649) );
  IMUX40 U651 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n759), .S1(n741), .Q(n656) );
  IMUX40 U652 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n755), .S1(n741), .Q(n654) );
  IMUX40 U653 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n764), .S1(n742), .Q(n653) );
  IMUX40 U654 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n756), .S1(n742), .Q(n661) );
  IMUX40 U655 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n752), .S1(n742), .Q(n659) );
  IMUX40 U656 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n752), .S1(n742), .Q(n666) );
  IMUX40 U657 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n761), .S1(n742), .Q(n664) );
  IMUX40 U658 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n750), .S1(n743), .Q(n663) );
  IMUX40 U659 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n754), .S1(n743), .Q(n671) );
  IMUX40 U660 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n758), .S1(n743), .Q(n669) );
  IMUX40 U661 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n751), .S1(n743), .Q(n676) );
  IMUX40 U662 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n757), .S1(n743), .Q(n674) );
  IMUX40 U663 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n764), .S1(n743), .Q(n673) );
  IMUX40 U664 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n760), .S1(n744), .Q(n681) );
  IMUX40 U665 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n760), .S1(n744), .Q(n679) );
  IMUX40 U666 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n760), .S1(n744), .Q(n686) );
  IMUX40 U667 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n760), .S1(n744), .Q(n684) );
  IMUX40 U668 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n760), .S1(n744), .Q(n683) );
  IMUX40 U669 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n760), .S1(n744), .Q(n691) );
  IMUX40 U670 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n760), .S1(n745), .Q(n689) );
  IMUX40 U671 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n761), .S1(n745), .Q(n696) );
  IMUX40 U672 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n761), .S1(n745), .Q(n694) );
  IMUX40 U673 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n761), .S1(n745), .Q(n693) );
  IMUX40 U674 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n761), .S1(n745), .Q(n701) );
  IMUX40 U675 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n761), .S1(n745), .Q(n699) );
  IMUX40 U676 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n761), .S1(n746), .Q(n698) );
  IMUX40 U677 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n761), .S1(n746), .Q(n706) );
  IMUX40 U678 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n761), .S1(n746), .Q(n704) );
  IMUX40 U679 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n761), .S1(n746), .Q(n703) );
  IMUX40 U680 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n762), .S1(n746), .Q(n711) );
  IMUX40 U681 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n762), .S1(n747), .Q(n708) );
  IMUX40 U682 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n762), .S1(n746), .Q(n709) );
  IMUX40 U683 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n762), .S1(n747), .Q(n716) );
  IMUX40 U684 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n762), .S1(n747), .Q(n714) );
  IMUX40 U685 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n762), .S1(n747), .Q(n713) );
  IMUX40 U686 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n762), .S1(n747), .Q(n721) );
  IMUX40 U687 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n762), .S1(n747), .Q(n718) );
  IMUX40 U688 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n762), .S1(n747), .Q(n719) );
  IMUX40 U689 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n385), .S1(n375), .Q(n9) );
  IMUX40 U690 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(i_addr_Rt[0]), .S1(n377), .Q(n4) );
  IMUX40 U691 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n385), .S1(n384), .Q(n14) );
  IMUX40 U692 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n385), .S1(n375), .Q(n19) );
  IMUX40 U693 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n386), .S1(n383), .Q(n24) );
  IMUX40 U694 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n386), .S1(n375), .Q(n29) );
  IMUX40 U695 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n386), .S1(n377), .Q(n34) );
  IMUX40 U696 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n387), .S1(n378), .Q(n83) );
  IMUX40 U697 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n387), .S1(n377), .Q(n88) );
  IMUX40 U698 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n387), .S1(n376), .Q(n93) );
  IMUX40 U699 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n388), .S1(n377), .Q(n98) );
  IMUX40 U700 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n388), .S1(n380), .Q(n103) );
  IMUX40 U701 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n388), .S1(n377), .Q(n108) );
  IMUX40 U702 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n389), .S1(n377), .Q(n113) );
  IMUX40 U703 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n389), .S1(n378), .Q(n118) );
  IMUX40 U704 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n389), .S1(n378), .Q(n123) );
  IMUX40 U705 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n390), .S1(n378), .Q(n128) );
  IMUX40 U706 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n390), .S1(i_addr_Rt[1]), .Q(n133) );
  IMUX40 U707 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n390), .S1(n384), .Q(n138) );
  IMUX40 U708 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n391), .S1(n379), .Q(n143) );
  IMUX40 U709 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n391), .S1(n379), .Q(n148) );
  IMUX40 U710 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n391), .S1(n380), .Q(n153) );
  IMUX40 U711 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n394), .S1(n380), .Q(n158) );
  IMUX40 U712 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n392), .S1(n381), .Q(n163) );
  IMUX40 U713 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n393), .S1(n381), .Q(n168) );
  IMUX40 U714 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(i_addr_Rt[0]), .S1(n381), .Q(n173) );
  IMUX40 U715 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n391), .S1(n382), .Q(n178) );
  IMUX40 U716 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(i_addr_Rt[0]), .S1(n382), .Q(n183) );
  IMUX40 U717 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n392), .S1(n374), .Q(n188) );
  IMUX40 U718 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n392), .S1(n374), .Q(n193) );
  IMUX40 U719 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n392), .S1(n377), .Q(n198) );
  IMUX40 U720 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n393), .S1(n377), .Q(n203) );
  IMUX40 U721 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n393), .S1(n381), .Q(n208) );
  IMUX40 U722 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n393), .S1(n378), .Q(n213) );
  IMUX40 U723 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n394), .S1(n380), .Q(n218) );
  IMUX40 U724 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n394), .S1(n377), .Q(n223) );
  IMUX40 U725 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n394), .S1(n375), .Q(n228) );
  IMUX40 U726 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n401), .S1(n379), .Q(n233) );
  IMUX40 U727 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n401), .S1(n374), .Q(n238) );
  IMUX40 U728 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n401), .S1(n384), .Q(n243) );
  IMUX40 U729 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n387), .S1(n377), .Q(n248) );
  IMUX40 U730 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n399), .S1(i_addr_Rt[1]), .Q(n253) );
  IMUX40 U731 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n386), .S1(n384), .Q(n258) );
  IMUX40 U732 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n398), .S1(i_addr_Rt[1]), .Q(n263) );
  IMUX40 U733 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n401), .S1(n383), .Q(n268) );
  IMUX40 U734 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n395), .S1(n383), .Q(n273) );
  IMUX40 U735 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n395), .S1(n379), .Q(n278) );
  IMUX40 U736 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n395), .S1(n374), .Q(n283) );
  IMUX40 U737 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n398), .S1(n381), .Q(n288) );
  IMUX40 U738 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n395), .S1(n383), .Q(n293) );
  IMUX40 U739 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n395), .S1(n384), .Q(n298) );
  IMUX40 U740 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n395), .S1(n384), .Q(n303) );
  IMUX40 U741 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n395), .S1(n384), .Q(n308) );
  IMUX40 U742 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n389), .S1(n374), .Q(n313) );
  IMUX40 U743 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n398), .S1(n384), .Q(n318) );
  IMUX40 U744 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n396), .S1(n383), .Q(n323) );
  IMUX40 U745 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n396), .S1(n377), .Q(n328) );
  IMUX40 U746 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n396), .S1(n374), .Q(n333) );
  IMUX40 U747 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n397), .S1(n374), .Q(n338) );
  IMUX40 U748 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n397), .S1(n383), .Q(n343) );
  IMUX40 U749 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n397), .S1(n384), .Q(n348) );
  IMUX40 U750 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n398), .S1(n375), .Q(n353) );
  IMUX40 U751 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n398), .S1(n374), .Q(n358) );
  IMUX40 U752 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n398), .S1(n381), .Q(n363) );
  IMUX40 U753 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n749), .S1(n731), .Q(n410) );
  IMUX40 U754 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(n756), .S1(n748), .Q(n405) );
  IMUX40 U755 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n749), .S1(i_addr_Rs[1]), .Q(n415) );
  IMUX40 U756 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n750), .S1(n732), .Q(n425) );
  IMUX40 U757 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n750), .S1(n730), .Q(n435) );
  IMUX40 U758 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n751), .S1(n730), .Q(n445) );
  IMUX40 U759 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n752), .S1(n747), .Q(n455) );
  IMUX40 U760 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n752), .S1(n730), .Q(n465) );
  IMUX40 U761 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n753), .S1(n732), .Q(n475) );
  IMUX40 U762 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n754), .S1(n733), .Q(n485) );
  IMUX40 U763 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n759), .S1(n734), .Q(n495) );
  IMUX40 U764 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n764), .S1(n733), .Q(n505) );
  IMUX40 U765 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n754), .S1(n730), .Q(n515) );
  IMUX40 U766 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n754), .S1(n731), .Q(n525) );
  IMUX40 U767 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n750), .S1(n731), .Q(n535) );
  IMUX40 U768 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n761), .S1(n738), .Q(n540) );
  IMUX40 U769 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n755), .S1(n733), .Q(n545) );
  IMUX40 U770 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n755), .S1(n733), .Q(n550) );
  IMUX40 U771 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n755), .S1(n734), .Q(n555) );
  IMUX40 U772 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n756), .S1(n734), .Q(n560) );
  IMUX40 U773 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n756), .S1(n735), .Q(n565) );
  IMUX40 U774 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n756), .S1(n735), .Q(n570) );
  IMUX40 U775 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n751), .S1(n735), .Q(n575) );
  IMUX40 U776 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n749), .S1(n736), .Q(n580) );
  IMUX40 U777 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n749), .S1(n736), .Q(n585) );
  IMUX40 U778 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n757), .S1(n738), .Q(n590) );
  IMUX40 U779 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n757), .S1(n738), .Q(n595) );
  IMUX40 U780 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n757), .S1(n737), .Q(n600) );
  IMUX40 U781 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n758), .S1(n737), .Q(n605) );
  IMUX40 U782 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n758), .S1(n738), .Q(n610) );
  IMUX40 U783 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n758), .S1(n738), .Q(n615) );
  IMUX40 U784 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n759), .S1(n738), .Q(n620) );
  IMUX40 U785 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n759), .S1(n739), .Q(n625) );
  IMUX40 U786 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n759), .S1(n739), .Q(n630) );
  IMUX40 U787 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n764), .S1(n740), .Q(n635) );
  IMUX40 U788 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n764), .S1(n740), .Q(n640) );
  IMUX40 U789 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n764), .S1(n741), .Q(n645) );
  IMUX40 U790 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n759), .S1(n741), .Q(n650) );
  IMUX40 U791 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n753), .S1(n742), .Q(n655) );
  IMUX40 U792 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n760), .S1(n742), .Q(n660) );
  IMUX40 U793 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n750), .S1(n742), .Q(n665) );
  IMUX40 U794 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n762), .S1(n743), .Q(n670) );
  IMUX40 U795 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n764), .S1(n743), .Q(n675) );
  IMUX40 U796 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n760), .S1(n744), .Q(n680) );
  IMUX40 U797 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n760), .S1(n744), .Q(n685) );
  IMUX40 U798 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n760), .S1(n745), .Q(n690) );
  IMUX40 U799 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n761), .S1(n745), .Q(n695) );
  IMUX40 U800 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n761), .S1(n746), .Q(n705) );
  IMUX40 U801 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n762), .S1(n747), .Q(n715) );
  BUF2 U802 ( .A(i_addr_Rt[3]), .Q(n367) );
  BUF2 U803 ( .A(i_addr_Rt[3]), .Q(n368) );
  BUF2 U804 ( .A(i_addr_Rt[3]), .Q(n369) );
  BUF2 U805 ( .A(i_addr_Rs[3]), .Q(n724) );
  BUF2 U806 ( .A(i_addr_Rs[3]), .Q(n725) );
  BUF2 U807 ( .A(i_addr_Rs[3]), .Q(n726) );
  INV3 U808 ( .A(i_addr_Rd[2]), .Q(n809) );
  INV3 U809 ( .A(i_addr_Rd[0]), .Q(n811) );
  INV3 U810 ( .A(i_addr_Rd[1]), .Q(n810) );
  INV3 U811 ( .A(i_con_RegWr), .Q(n812) );
  BUF2 U812 ( .A(i_addr_Rs[4]), .Q(n722) );
  BUF2 U813 ( .A(i_addr_Rs[2]), .Q(n727) );
  BUF2 U814 ( .A(i_addr_Rs[2]), .Q(n728) );
  BUF2 U815 ( .A(i_addr_Rs[2]), .Q(n729) );
  INV3 U816 ( .A(i_addr_Rd[4]), .Q(n791) );
  INV3 U817 ( .A(i_addr_Rd[3]), .Q(n808) );
  BUF2 U818 ( .A(i_addr_Rs[3]), .Q(n723) );
  MUX22 U819 ( .A(n417), .B(n412), .S(n722), .Q(o_data_Rs[1]) );
  IMUX40 U820 ( .A(n418), .B(n419), .C(n420), .D(n421), .S0(n723), .S1(n727), 
        .Q(n417) );
  IMUX40 U821 ( .A(n413), .B(n414), .C(n415), .D(n416), .S0(n723), .S1(n727), 
        .Q(n412) );
  IMUX40 U822 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n749), .S1(n733), .Q(n420) );
  MUX22 U823 ( .A(n427), .B(n422), .S(n722), .Q(o_data_Rs[2]) );
  IMUX40 U824 ( .A(n428), .B(n429), .C(n430), .D(n431), .S0(i_addr_Rs[3]), 
        .S1(n727), .Q(n427) );
  IMUX40 U825 ( .A(n423), .B(n424), .C(n425), .D(n426), .S0(n723), .S1(n727), 
        .Q(n422) );
  IMUX40 U826 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n750), .S1(n734), .Q(n430) );
  MUX22 U827 ( .A(n437), .B(n432), .S(n722), .Q(o_data_Rs[3]) );
  IMUX40 U828 ( .A(n438), .B(n439), .C(n440), .D(n441), .S0(i_addr_Rs[3]), 
        .S1(n727), .Q(n437) );
  IMUX40 U829 ( .A(n433), .B(n434), .C(n435), .D(n436), .S0(n726), .S1(n727), 
        .Q(n432) );
  IMUX40 U830 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n751), .S1(i_addr_Rs[1]), .Q(n440) );
  MUX22 U831 ( .A(n447), .B(n442), .S(n722), .Q(o_data_Rs[4]) );
  IMUX40 U832 ( .A(n448), .B(n449), .C(n450), .D(n451), .S0(i_addr_Rs[3]), 
        .S1(n727), .Q(n447) );
  IMUX40 U833 ( .A(n443), .B(n444), .C(n445), .D(n446), .S0(i_addr_Rs[3]), 
        .S1(n727), .Q(n442) );
  IMUX40 U834 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n751), .S1(n732), .Q(n450) );
  MUX22 U835 ( .A(n457), .B(n452), .S(n722), .Q(o_data_Rs[5]) );
  IMUX40 U836 ( .A(n458), .B(n459), .C(n460), .D(n461), .S0(i_addr_Rs[3]), 
        .S1(n728), .Q(n457) );
  IMUX40 U837 ( .A(n453), .B(n454), .C(n455), .D(n456), .S0(i_addr_Rs[3]), 
        .S1(n728), .Q(n452) );
  IMUX40 U838 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n752), .S1(n731), .Q(n460) );
  MUX22 U839 ( .A(n467), .B(n462), .S(n722), .Q(o_data_Rs[6]) );
  IMUX40 U840 ( .A(n468), .B(n469), .C(n470), .D(n471), .S0(i_addr_Rs[3]), 
        .S1(n728), .Q(n467) );
  IMUX40 U841 ( .A(n463), .B(n464), .C(n465), .D(n466), .S0(i_addr_Rs[3]), 
        .S1(n728), .Q(n462) );
  IMUX40 U842 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n753), .S1(n738), .Q(n470) );
  MUX22 U843 ( .A(n477), .B(n472), .S(n722), .Q(o_data_Rs[7]) );
  IMUX40 U844 ( .A(n478), .B(n479), .C(n480), .D(n481), .S0(i_addr_Rs[3]), 
        .S1(n728), .Q(n477) );
  IMUX40 U845 ( .A(n473), .B(n474), .C(n475), .D(n476), .S0(i_addr_Rs[3]), 
        .S1(n728), .Q(n472) );
  IMUX40 U846 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n753), .S1(n733), .Q(n480) );
  MUX22 U847 ( .A(n487), .B(n482), .S(n722), .Q(o_data_Rs[8]) );
  IMUX40 U848 ( .A(n488), .B(n489), .C(n490), .D(n491), .S0(n723), .S1(n728), 
        .Q(n487) );
  IMUX40 U849 ( .A(n483), .B(n484), .C(n485), .D(n486), .S0(n723), .S1(n728), 
        .Q(n482) );
  IMUX40 U850 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n762), .S1(i_addr_Rs[1]), .Q(n490) );
  MUX22 U851 ( .A(n497), .B(n492), .S(i_addr_Rs[4]), .Q(o_data_Rs[9]) );
  IMUX40 U852 ( .A(n498), .B(n499), .C(n500), .D(n501), .S0(n723), .S1(n729), 
        .Q(n497) );
  IMUX40 U853 ( .A(n493), .B(n494), .C(n495), .D(n496), .S0(n723), .S1(n728), 
        .Q(n492) );
  IMUX40 U854 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n751), .S1(n730), .Q(n500) );
  MUX22 U855 ( .A(n507), .B(n502), .S(n722), .Q(o_data_Rs[10]) );
  IMUX40 U856 ( .A(n508), .B(n509), .C(n510), .D(n511), .S0(n723), .S1(n729), 
        .Q(n507) );
  IMUX40 U857 ( .A(n503), .B(n504), .C(n505), .D(n506), .S0(n723), .S1(n729), 
        .Q(n502) );
  IMUX40 U858 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n755), .S1(n734), .Q(n510) );
  MUX22 U859 ( .A(n517), .B(n512), .S(n722), .Q(o_data_Rs[11]) );
  IMUX40 U860 ( .A(n518), .B(n519), .C(n520), .D(n521), .S0(i_addr_Rs[3]), 
        .S1(n729), .Q(n517) );
  IMUX40 U861 ( .A(n513), .B(n514), .C(n515), .D(n516), .S0(n723), .S1(n729), 
        .Q(n512) );
  IMUX40 U862 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n754), .S1(i_addr_Rs[1]), .Q(n520) );
  MUX22 U863 ( .A(n527), .B(n522), .S(n722), .Q(o_data_Rs[12]) );
  IMUX40 U864 ( .A(n528), .B(n529), .C(n530), .D(n531), .S0(i_addr_Rs[3]), 
        .S1(n729), .Q(n527) );
  IMUX40 U865 ( .A(n523), .B(n524), .C(n525), .D(n526), .S0(n723), .S1(n729), 
        .Q(n522) );
  IMUX40 U866 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n764), .S1(n734), .Q(n530) );
  BUF2 U867 ( .A(i_addr_Rt[1]), .Q(n384) );
  BUF2 U868 ( .A(i_addr_Rs[1]), .Q(n748) );
  MUX22 U869 ( .A(n6), .B(n1), .S(n365), .Q(o_data_Rt[0]) );
  IMUX40 U870 ( .A(n2), .B(n3), .C(n4), .D(n5), .S0(n366), .S1(i_addr_Rt[2]), 
        .Q(n1) );
  IMUX40 U871 ( .A(n7), .B(n8), .C(n9), .D(n10), .S0(n366), .S1(i_addr_Rt[2]), 
        .Q(n6) );
  BUF2 U872 ( .A(i_addr_Rt[4]), .Q(n365) );
  BUF2 U873 ( .A(i_addr_Rt[2]), .Q(n370) );
  BUF2 U874 ( .A(i_addr_Rt[2]), .Q(n371) );
  BUF2 U875 ( .A(i_addr_Rt[2]), .Q(n372) );
  BUF2 U876 ( .A(i_addr_Rt[2]), .Q(n373) );
  BUF2 U877 ( .A(i_addr_Rt[3]), .Q(n366) );
endmodule


module D_shiftleft ( i_data_immE, o_data_immshiftl );
  input [15:0] i_data_immE;
  output [31:0] o_data_immshiftl;
  wire   n1;
  assign o_data_immshiftl[0] = o_data_immshiftl[1];
  assign o_data_immshiftl[20] = o_data_immshiftl[31];
  assign o_data_immshiftl[19] = o_data_immshiftl[31];
  assign o_data_immshiftl[29] = o_data_immshiftl[31];
  assign o_data_immshiftl[26] = o_data_immshiftl[31];
  assign o_data_immshiftl[25] = o_data_immshiftl[31];
  assign o_data_immshiftl[21] = o_data_immshiftl[31];
  assign o_data_immshiftl[23] = o_data_immshiftl[30];
  assign o_data_immshiftl[27] = o_data_immshiftl[30];
  assign o_data_immshiftl[28] = o_data_immshiftl[30];
  assign o_data_immshiftl[17] = o_data_immshiftl[30];
  assign o_data_immshiftl[22] = o_data_immshiftl[30];
  assign o_data_immshiftl[18] = o_data_immshiftl[30];
  assign o_data_immshiftl[24] = i_data_immE[15];
  assign o_data_immshiftl[16] = i_data_immE[14];
  assign o_data_immshiftl[15] = i_data_immE[13];
  assign o_data_immshiftl[14] = i_data_immE[12];
  assign o_data_immshiftl[13] = i_data_immE[11];
  assign o_data_immshiftl[12] = i_data_immE[10];
  assign o_data_immshiftl[11] = i_data_immE[9];
  assign o_data_immshiftl[10] = i_data_immE[8];
  assign o_data_immshiftl[9] = i_data_immE[7];
  assign o_data_immshiftl[8] = i_data_immE[6];
  assign o_data_immshiftl[7] = i_data_immE[5];
  assign o_data_immshiftl[6] = i_data_immE[4];
  assign o_data_immshiftl[5] = i_data_immE[3];
  assign o_data_immshiftl[4] = i_data_immE[2];
  assign o_data_immshiftl[3] = i_data_immE[1];
  assign o_data_immshiftl[2] = i_data_immE[0];

  INV3 U2 ( .A(n1), .Q(o_data_immshiftl[30]) );
  INV3 U3 ( .A(n1), .Q(o_data_immshiftl[31]) );
  INV3 U4 ( .A(i_data_immE[15]), .Q(n1) );
  LOGIC0 U5 ( .Q(o_data_immshiftl[1]) );
endmodule


module D_sign_extend ( i_data_immD, i_con_signext, o_data_immD );
  input [15:0] i_data_immD;
  output [31:0] o_data_immD;
  input i_con_signext;
  wire   n2;
  assign o_data_immD[15] = i_data_immD[15];
  assign o_data_immD[14] = i_data_immD[14];
  assign o_data_immD[13] = i_data_immD[13];
  assign o_data_immD[12] = i_data_immD[12];
  assign o_data_immD[11] = i_data_immD[11];
  assign o_data_immD[10] = i_data_immD[10];
  assign o_data_immD[9] = i_data_immD[9];
  assign o_data_immD[8] = i_data_immD[8];
  assign o_data_immD[7] = i_data_immD[7];
  assign o_data_immD[6] = i_data_immD[6];
  assign o_data_immD[5] = i_data_immD[5];
  assign o_data_immD[4] = i_data_immD[4];
  assign o_data_immD[3] = i_data_immD[3];
  assign o_data_immD[2] = i_data_immD[2];
  assign o_data_immD[1] = i_data_immD[1];
  assign o_data_immD[0] = i_data_immD[0];
  assign o_data_immD[16] = o_data_immD[31];
  assign o_data_immD[17] = o_data_immD[31];
  assign o_data_immD[18] = o_data_immD[31];
  assign o_data_immD[19] = o_data_immD[31];
  assign o_data_immD[20] = o_data_immD[31];
  assign o_data_immD[21] = o_data_immD[31];
  assign o_data_immD[22] = o_data_immD[31];
  assign o_data_immD[23] = o_data_immD[31];
  assign o_data_immD[24] = o_data_immD[31];
  assign o_data_immD[25] = o_data_immD[31];
  assign o_data_immD[26] = o_data_immD[31];
  assign o_data_immD[27] = o_data_immD[31];
  assign o_data_immD[28] = o_data_immD[31];
  assign o_data_immD[29] = o_data_immD[31];
  assign o_data_immD[30] = o_data_immD[31];

  INV3 U2 ( .A(n2), .Q(o_data_immD[31]) );
  NAND22 U3 ( .A(i_con_signext), .B(i_data_immD[15]), .Q(n2) );
endmodule


module D_jump_ext ( i_addr_j, i_PC4_j, o_addr_j );
  input [25:0] i_addr_j;
  input [3:0] i_PC4_j;
  output [31:0] o_addr_j;

  assign o_addr_j[0] = o_addr_j[1];
  assign o_addr_j[31] = i_PC4_j[3];
  assign o_addr_j[30] = i_PC4_j[2];
  assign o_addr_j[29] = i_PC4_j[1];
  assign o_addr_j[28] = i_PC4_j[0];
  assign o_addr_j[27] = i_addr_j[25];
  assign o_addr_j[26] = i_addr_j[24];
  assign o_addr_j[25] = i_addr_j[23];
  assign o_addr_j[24] = i_addr_j[22];
  assign o_addr_j[23] = i_addr_j[21];
  assign o_addr_j[22] = i_addr_j[20];
  assign o_addr_j[21] = i_addr_j[19];
  assign o_addr_j[20] = i_addr_j[18];
  assign o_addr_j[19] = i_addr_j[17];
  assign o_addr_j[18] = i_addr_j[16];
  assign o_addr_j[17] = i_addr_j[15];
  assign o_addr_j[16] = i_addr_j[14];
  assign o_addr_j[15] = i_addr_j[13];
  assign o_addr_j[14] = i_addr_j[12];
  assign o_addr_j[13] = i_addr_j[11];
  assign o_addr_j[12] = i_addr_j[10];
  assign o_addr_j[11] = i_addr_j[9];
  assign o_addr_j[10] = i_addr_j[8];
  assign o_addr_j[9] = i_addr_j[7];
  assign o_addr_j[8] = i_addr_j[6];
  assign o_addr_j[7] = i_addr_j[5];
  assign o_addr_j[6] = i_addr_j[4];
  assign o_addr_j[5] = i_addr_j[3];
  assign o_addr_j[4] = i_addr_j[2];
  assign o_addr_j[3] = i_addr_j[1];
  assign o_addr_j[2] = i_addr_j[0];

  LOGIC0 U2 ( .Q(o_addr_j[1]) );
endmodule


module D_forward ( i_addr_rs, i_addr_rt, i_addr_rdE, i_addr_rdM, i_addr_rtM, 
        i_addr_rtW, i_con_regwriteE, i_con_regwriteM, i_con_memreadM, 
        i_con_memreadW, o_con_fa, o_con_fb );
  input [4:0] i_addr_rs;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rdE;
  input [4:0] i_addr_rdM;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  output [2:0] o_con_fa;
  output [2:0] o_con_fb;
  input i_con_regwriteE, i_con_regwriteM, i_con_memreadM, i_con_memreadW;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;

  NOR31 U1 ( .A(i_addr_rs[2]), .B(i_addr_rs[4]), .C(i_addr_rs[3]), .Q(n85) );
  OAI310 U2 ( .A(n1), .B(n2), .C(n3), .D(n4), .Q(o_con_fb[2]) );
  NOR40 U3 ( .A(n5), .B(n6), .C(n7), .D(n8), .Q(o_con_fb[1]) );
  CLKIN0 U4 ( .A(n9), .Q(n6) );
  NAND20 U5 ( .A(n4), .B(n10), .Q(o_con_fb[0]) );
  NAND40 U6 ( .A(n11), .B(i_con_regwriteM), .C(n12), .D(n13), .Q(n10) );
  NOR40 U7 ( .A(n14), .B(n15), .C(n16), .D(n17), .Q(n13) );
  XOR20 U8 ( .A(i_addr_rdM[4]), .B(i_addr_rt[4]), .Q(n17) );
  XNR20 U9 ( .A(n18), .B(i_addr_rt[2]), .Q(n16) );
  XNR20 U10 ( .A(n19), .B(i_addr_rt[1]), .Q(n15) );
  XNR20 U11 ( .A(n20), .B(i_addr_rt[0]), .Q(n14) );
  CLKIN0 U12 ( .A(n21), .Q(n12) );
  OAI210 U13 ( .A(n8), .B(n7), .C(n9), .Q(n21) );
  NAND40 U14 ( .A(n22), .B(n23), .C(n24), .D(n25), .Q(n7) );
  XNR20 U15 ( .A(i_addr_rt[0]), .B(i_addr_rdE[0]), .Q(n25) );
  NOR20 U16 ( .A(n26), .B(n27), .Q(n24) );
  XNR20 U17 ( .A(n28), .B(i_addr_rt[3]), .Q(n27) );
  XOR20 U18 ( .A(i_addr_rdE[1]), .B(i_addr_rt[1]), .Q(n26) );
  XNR20 U19 ( .A(i_addr_rt[2]), .B(i_addr_rdE[2]), .Q(n23) );
  XNR20 U20 ( .A(i_addr_rt[4]), .B(i_addr_rdE[4]), .Q(n22) );
  CLKIN0 U21 ( .A(i_con_regwriteE), .Q(n8) );
  XNR20 U22 ( .A(i_addr_rt[3]), .B(i_addr_rdM[3]), .Q(n11) );
  NAND20 U23 ( .A(n9), .B(n5), .Q(n4) );
  CLKIN0 U24 ( .A(n29), .Q(n5) );
  NAND40 U25 ( .A(n30), .B(i_con_memreadW), .C(n31), .D(n32), .Q(n29) );
  NOR30 U26 ( .A(n33), .B(n34), .C(n35), .Q(n32) );
  XOR20 U27 ( .A(i_addr_rtW[2]), .B(i_addr_rt[2]), .Q(n35) );
  XOR20 U28 ( .A(i_addr_rtW[4]), .B(i_addr_rt[4]), .Q(n34) );
  XOR20 U29 ( .A(i_addr_rtW[3]), .B(i_addr_rt[3]), .Q(n33) );
  XNR20 U30 ( .A(i_addr_rt[0]), .B(i_addr_rtW[0]), .Q(n31) );
  XNR20 U31 ( .A(i_addr_rt[1]), .B(i_addr_rtW[1]), .Q(n30) );
  AOI210 U32 ( .A(n36), .B(i_con_memreadM), .C(n2), .Q(n9) );
  NOR30 U33 ( .A(i_addr_rt[0]), .B(i_addr_rt[1]), .C(n37), .Q(n2) );
  CLKIN0 U34 ( .A(n38), .Q(n37) );
  NOR30 U35 ( .A(i_addr_rt[2]), .B(i_addr_rt[4]), .C(i_addr_rt[3]), .Q(n38) );
  CLKIN0 U36 ( .A(n3), .Q(n36) );
  NAND40 U37 ( .A(n39), .B(n40), .C(n41), .D(n42), .Q(n3) );
  XNR20 U38 ( .A(i_addr_rt[0]), .B(i_addr_rtM[0]), .Q(n42) );
  NOR20 U39 ( .A(n43), .B(n44), .Q(n41) );
  XOR20 U40 ( .A(i_addr_rtM[3]), .B(i_addr_rt[3]), .Q(n44) );
  XNR20 U41 ( .A(n45), .B(i_addr_rt[1]), .Q(n43) );
  XNR20 U42 ( .A(i_addr_rt[2]), .B(i_addr_rtM[2]), .Q(n40) );
  XNR20 U43 ( .A(i_addr_rt[4]), .B(i_addr_rtM[4]), .Q(n39) );
  NOR20 U44 ( .A(o_con_fa[2]), .B(n46), .Q(o_con_fa[1]) );
  OAI210 U45 ( .A(n47), .B(n48), .C(n49), .Q(o_con_fa[0]) );
  NAND20 U46 ( .A(n50), .B(n51), .Q(n49) );
  NOR40 U47 ( .A(o_con_fa[2]), .B(n52), .C(n53), .D(n54), .Q(n51) );
  XNR20 U48 ( .A(n20), .B(i_addr_rs[0]), .Q(n54) );
  CLKIN0 U49 ( .A(i_addr_rdM[0]), .Q(n20) );
  CLKIN0 U50 ( .A(i_con_regwriteM), .Q(n53) );
  CLKIN0 U51 ( .A(n46), .Q(n52) );
  NAND40 U52 ( .A(n55), .B(i_con_regwriteE), .C(n56), .D(n57), .Q(n46) );
  NOR30 U53 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  XNR20 U54 ( .A(n28), .B(i_addr_rs[3]), .Q(n60) );
  CLKIN0 U55 ( .A(i_addr_rdE[3]), .Q(n28) );
  XOR20 U56 ( .A(i_addr_rdE[2]), .B(i_addr_rs[2]), .Q(n59) );
  IMUX20 U57 ( .A(n61), .B(i_addr_rs[4]), .S(i_addr_rdE[4]), .Q(n58) );
  NOR20 U58 ( .A(n62), .B(i_addr_rs[4]), .Q(n61) );
  NOR40 U59 ( .A(i_addr_rdE[3]), .B(i_addr_rdE[2]), .C(i_addr_rdE[1]), .D(
        i_addr_rdE[0]), .Q(n62) );
  XNR20 U60 ( .A(i_addr_rs[0]), .B(i_addr_rdE[0]), .Q(n56) );
  XNR20 U61 ( .A(i_addr_rs[1]), .B(i_addr_rdE[1]), .Q(n55) );
  NAND20 U62 ( .A(n63), .B(n48), .Q(o_con_fa[2]) );
  NOR40 U63 ( .A(n64), .B(n65), .C(n66), .D(n67), .Q(n50) );
  IMUX20 U64 ( .A(n68), .B(i_addr_rs[4]), .S(i_addr_rdM[4]), .Q(n67) );
  NOR20 U65 ( .A(n69), .B(i_addr_rs[4]), .Q(n68) );
  NOR40 U66 ( .A(i_addr_rdM[3]), .B(i_addr_rdM[2]), .C(i_addr_rdM[1]), .D(
        i_addr_rdM[0]), .Q(n69) );
  XOR20 U67 ( .A(i_addr_rdM[3]), .B(i_addr_rs[3]), .Q(n66) );
  XNR20 U68 ( .A(n18), .B(i_addr_rs[2]), .Q(n65) );
  CLKIN0 U69 ( .A(i_addr_rdM[2]), .Q(n18) );
  XNR20 U70 ( .A(n19), .B(i_addr_rs[1]), .Q(n64) );
  CLKIN0 U71 ( .A(i_addr_rdM[1]), .Q(n19) );
  NAND40 U72 ( .A(n70), .B(n71), .C(n72), .D(n73), .Q(n48) );
  NOR40 U73 ( .A(n74), .B(n75), .C(n76), .D(n77), .Q(n73) );
  XOR20 U74 ( .A(i_addr_rtW[1]), .B(i_addr_rs[1]), .Q(n77) );
  XOR20 U75 ( .A(i_addr_rtW[0]), .B(i_addr_rs[0]), .Q(n76) );
  CLKIN0 U76 ( .A(i_con_memreadW), .Q(n75) );
  XNR20 U77 ( .A(i_addr_rtW[3]), .B(i_addr_rs[3]), .Q(n72) );
  XNR20 U78 ( .A(i_addr_rtW[4]), .B(i_addr_rs[4]), .Q(n71) );
  XNR20 U79 ( .A(i_addr_rtW[2]), .B(i_addr_rs[2]), .Q(n70) );
  CLKIN0 U80 ( .A(n63), .Q(n47) );
  NAND40 U81 ( .A(n78), .B(n79), .C(n80), .D(n81), .Q(n63) );
  NOR40 U82 ( .A(n74), .B(n1), .C(n82), .D(n83), .Q(n81) );
  XNR20 U83 ( .A(n45), .B(i_addr_rs[1]), .Q(n83) );
  CLKIN0 U84 ( .A(i_addr_rtM[1]), .Q(n45) );
  XOR20 U85 ( .A(i_addr_rtM[0]), .B(i_addr_rs[0]), .Q(n82) );
  CLKIN0 U86 ( .A(i_con_memreadM), .Q(n1) );
  NOR30 U87 ( .A(i_addr_rs[0]), .B(i_addr_rs[1]), .C(n84), .Q(n74) );
  CLKIN0 U88 ( .A(n85), .Q(n84) );
  XNR20 U89 ( .A(i_addr_rtM[3]), .B(i_addr_rs[3]), .Q(n80) );
  XNR20 U90 ( .A(i_addr_rtM[4]), .B(i_addr_rs[4]), .Q(n79) );
  XNR20 U91 ( .A(i_addr_rtM[2]), .B(i_addr_rs[2]), .Q(n78) );
endmodule


module decode ( i_clk, i_nrst, i_addr_pc4, i_data_instr, i_con_Wregwrite, 
        i_data_Wregwrite, i_addr_Wregwrite, i_addr_Erd, i_addr_Mrd, 
        i_con_Eregwrite, i_con_Mregwrite, i_addr_rtM, i_addr_rtW, 
        i_con_memreadM, i_con_memreadW, i_data_Wmemout, o_data_rs, o_data_rt, 
        o_addr_rd, o_addr_rt, o_data_jr, o_con_jump, o_addr_pc4, o_addr_branch, 
        o_addr_jump, o_con_Ealuop, o_con_Ealusrc, o_con_Eregdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_con_ifstall, o_con_Ebop, o_data_signext, 
        o_con_Efamux, o_con_Efbmux, o_data_Fmemout );
  input [31:0] i_addr_pc4;
  input [31:0] i_data_instr;
  input [31:0] i_data_Wregwrite;
  input [4:0] i_addr_Wregwrite;
  input [4:0] i_addr_Erd;
  input [4:0] i_addr_Mrd;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  input [31:0] i_data_Wmemout;
  output [31:0] o_data_rs;
  output [31:0] o_data_rt;
  output [4:0] o_addr_rd;
  output [4:0] o_addr_rt;
  output [31:0] o_data_jr;
  output [1:0] o_con_jump;
  output [31:0] o_addr_pc4;
  output [31:0] o_addr_branch;
  output [31:0] o_addr_jump;
  output [5:0] o_con_Ealuop;
  output [2:0] o_con_Ebop;
  output [31:0] o_data_signext;
  output [2:0] o_con_Efamux;
  output [2:0] o_con_Efbmux;
  output [31:0] o_data_Fmemout;
  input i_clk, i_nrst, i_con_Wregwrite, i_con_Eregwrite, i_con_Mregwrite,
         i_con_memreadM, i_con_memreadW;
  output o_con_Ealusrc, o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite,
         o_con_Malupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall;
  wire   control_o_con_alusrc, control_o_con_regdst, jbcon_o_con_aluPC4,
         control_o_con_memread, control_o_con_memwrite, control_o_con_memtoreg,
         control_o_con_regwrite, signext_i_con_signext, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;
  wire   [31:0] regbank_o_data_Rt;
  wire   [5:0] control_o_con_aluop;
  wire   [31:0] signext_o_data_immD;
  wire   [2:0] for_o_con_fa;
  wire   [2:0] for_o_con_fb;
  wire   [31:0] pcadd_o_addr_pcbranchE;
  wire   [2:0] jbcon_o_con_bop;
  wire   [31:2] pcadd_i_data_immshiftl;
  assign o_addr_jump[1] = o_addr_jump[0];

  DFC3 pipe_bop_reg_2_ ( .D(jbcon_o_con_bop[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[2]) );
  DFC3 pipe_bop_reg_1_ ( .D(jbcon_o_con_bop[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[1]) );
  DFC3 pipe_bop_reg_0_ ( .D(jbcon_o_con_bop[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[0]) );
  DFC3 pipe_data_rs_reg_31_ ( .D(o_data_jr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[31]) );
  DFC3 pipe_data_rs_reg_30_ ( .D(o_data_jr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[30]) );
  DFC3 pipe_data_rs_reg_29_ ( .D(o_data_jr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[29]) );
  DFC3 pipe_data_rs_reg_28_ ( .D(o_data_jr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[28]) );
  DFC3 pipe_data_rs_reg_27_ ( .D(o_data_jr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[27]) );
  DFC3 pipe_data_rs_reg_26_ ( .D(o_data_jr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[26]) );
  DFC3 pipe_data_rs_reg_25_ ( .D(o_data_jr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[25]) );
  DFC3 pipe_data_rs_reg_24_ ( .D(o_data_jr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[24]) );
  DFC3 pipe_data_rs_reg_23_ ( .D(o_data_jr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[23]) );
  DFC3 pipe_data_rs_reg_22_ ( .D(o_data_jr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[22]) );
  DFC3 pipe_data_rs_reg_21_ ( .D(o_data_jr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[21]) );
  DFC3 pipe_data_rs_reg_20_ ( .D(o_data_jr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[20]) );
  DFC3 pipe_data_rs_reg_19_ ( .D(o_data_jr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[19]) );
  DFC3 pipe_data_rs_reg_18_ ( .D(o_data_jr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[18]) );
  DFC3 pipe_data_rs_reg_17_ ( .D(o_data_jr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[17]) );
  DFC3 pipe_data_rs_reg_16_ ( .D(o_data_jr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[16]) );
  DFC3 pipe_data_rs_reg_15_ ( .D(o_data_jr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[15]) );
  DFC3 pipe_data_rs_reg_14_ ( .D(o_data_jr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[14]) );
  DFC3 pipe_data_rs_reg_13_ ( .D(o_data_jr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[13]) );
  DFC3 pipe_data_rs_reg_12_ ( .D(o_data_jr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[12]) );
  DFC3 pipe_data_rs_reg_11_ ( .D(o_data_jr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[11]) );
  DFC3 pipe_data_rs_reg_10_ ( .D(o_data_jr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[10]) );
  DFC3 pipe_data_rs_reg_9_ ( .D(o_data_jr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[9]) );
  DFC3 pipe_data_rs_reg_8_ ( .D(o_data_jr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[8]) );
  DFC3 pipe_data_rs_reg_7_ ( .D(o_data_jr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[7]) );
  DFC3 pipe_data_rs_reg_6_ ( .D(o_data_jr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[6]) );
  DFC3 pipe_data_rs_reg_5_ ( .D(o_data_jr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[5]) );
  DFC3 pipe_data_rs_reg_4_ ( .D(o_data_jr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[4]) );
  DFC3 pipe_data_rs_reg_3_ ( .D(o_data_jr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[3]) );
  DFC3 pipe_data_rs_reg_2_ ( .D(o_data_jr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[2]) );
  DFC3 pipe_data_rs_reg_1_ ( .D(o_data_jr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[1]) );
  DFC3 pipe_data_rs_reg_0_ ( .D(o_data_jr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[0]) );
  DFC3 pipe_data_rt_reg_31_ ( .D(regbank_o_data_Rt[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[31]) );
  DFC3 pipe_data_rt_reg_30_ ( .D(regbank_o_data_Rt[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC3 pipe_data_rt_reg_29_ ( .D(regbank_o_data_Rt[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[29]) );
  DFC3 pipe_data_rt_reg_28_ ( .D(regbank_o_data_Rt[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28]) );
  DFC3 pipe_data_rt_reg_27_ ( .D(regbank_o_data_Rt[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27]) );
  DFC3 pipe_data_rt_reg_26_ ( .D(regbank_o_data_Rt[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26]) );
  DFC3 pipe_data_rt_reg_25_ ( .D(regbank_o_data_Rt[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25]) );
  DFC3 pipe_data_rt_reg_24_ ( .D(regbank_o_data_Rt[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24]) );
  DFC3 pipe_data_rt_reg_23_ ( .D(regbank_o_data_Rt[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23]) );
  DFC3 pipe_data_rt_reg_22_ ( .D(regbank_o_data_Rt[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC3 pipe_data_rt_reg_21_ ( .D(regbank_o_data_Rt[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21]) );
  DFC3 pipe_data_rt_reg_20_ ( .D(regbank_o_data_Rt[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20]) );
  DFC3 pipe_data_rt_reg_19_ ( .D(regbank_o_data_Rt[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19]) );
  DFC3 pipe_data_rt_reg_18_ ( .D(regbank_o_data_Rt[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18]) );
  DFC3 pipe_data_rt_reg_17_ ( .D(regbank_o_data_Rt[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17]) );
  DFC3 pipe_data_rt_reg_16_ ( .D(regbank_o_data_Rt[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC3 pipe_data_rt_reg_15_ ( .D(regbank_o_data_Rt[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15]) );
  DFC3 pipe_data_rt_reg_14_ ( .D(regbank_o_data_Rt[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14]) );
  DFC3 pipe_data_rt_reg_13_ ( .D(regbank_o_data_Rt[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC3 pipe_data_rt_reg_12_ ( .D(regbank_o_data_Rt[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12]) );
  DFC3 pipe_data_rt_reg_11_ ( .D(regbank_o_data_Rt[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11]) );
  DFC3 pipe_data_rt_reg_10_ ( .D(regbank_o_data_Rt[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC3 pipe_data_rt_reg_9_ ( .D(regbank_o_data_Rt[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[9]) );
  DFC3 pipe_data_rt_reg_8_ ( .D(regbank_o_data_Rt[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[8]) );
  DFC3 pipe_data_rt_reg_7_ ( .D(regbank_o_data_Rt[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[7]) );
  DFC3 pipe_data_rt_reg_6_ ( .D(regbank_o_data_Rt[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[6]) );
  DFC3 pipe_data_rt_reg_5_ ( .D(regbank_o_data_Rt[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[5]) );
  DFC3 pipe_data_rt_reg_4_ ( .D(regbank_o_data_Rt[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[4]) );
  DFC3 pipe_data_rt_reg_3_ ( .D(regbank_o_data_Rt[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[3]) );
  DFC3 pipe_data_rt_reg_2_ ( .D(regbank_o_data_Rt[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[2]) );
  DFC3 pipe_data_rt_reg_1_ ( .D(regbank_o_data_Rt[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[1]) );
  DFC3 pipe_data_rt_reg_0_ ( .D(regbank_o_data_Rt[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[0]) );
  DFC3 pipe_addr_rd_reg_4_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[4]) );
  DFC3 pipe_addr_rd_reg_3_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[3]) );
  DFC3 pipe_addr_rd_reg_2_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[2]) );
  DFC3 pipe_addr_rd_reg_1_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[1]) );
  DFC3 pipe_addr_rd_reg_0_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[0]) );
  DFC3 pipe_addr_rt_reg_4_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[0]) );
  DFC3 pipe_addr_pc4_reg_31_ ( .D(i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_addr_pc4_reg_30_ ( .D(i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_addr_pc4_reg_29_ ( .D(i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_addr_pc4_reg_28_ ( .D(i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_addr_pc4_reg_27_ ( .D(i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_addr_pc4_reg_26_ ( .D(i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_addr_pc4_reg_25_ ( .D(i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_addr_pc4_reg_24_ ( .D(i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_addr_pc4_reg_23_ ( .D(i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_addr_pc4_reg_22_ ( .D(i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_addr_pc4_reg_21_ ( .D(i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_addr_pc4_reg_20_ ( .D(i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_addr_pc4_reg_19_ ( .D(i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_addr_pc4_reg_18_ ( .D(i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_addr_pc4_reg_17_ ( .D(i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_addr_pc4_reg_16_ ( .D(i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_addr_pc4_reg_15_ ( .D(i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_addr_pc4_reg_14_ ( .D(i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_addr_pc4_reg_13_ ( .D(i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_addr_pc4_reg_12_ ( .D(i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_addr_pc4_reg_11_ ( .D(i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_addr_pc4_reg_10_ ( .D(i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_addr_pc4_reg_9_ ( .D(i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_addr_pc4_reg_8_ ( .D(i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_addr_pc4_reg_7_ ( .D(i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_addr_pc4_reg_6_ ( .D(i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_addr_pc4_reg_5_ ( .D(i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_addr_pc4_reg_4_ ( .D(i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_addr_pc4_reg_3_ ( .D(i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_addr_pc4_reg_2_ ( .D(i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_addr_pc4_reg_1_ ( .D(i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_addr_pc4_reg_0_ ( .D(i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  DFC3 pipe_con_Ealuop_reg_5_ ( .D(control_o_con_aluop[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[5]) );
  DFC3 pipe_con_Ealuop_reg_4_ ( .D(control_o_con_aluop[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[4]) );
  DFC3 pipe_con_Ealuop_reg_3_ ( .D(control_o_con_aluop[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[3]) );
  DFC3 pipe_con_Ealuop_reg_2_ ( .D(control_o_con_aluop[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[2]) );
  DFC3 pipe_con_Ealuop_reg_1_ ( .D(control_o_con_aluop[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[1]) );
  DFC3 pipe_con_Ealuop_reg_0_ ( .D(control_o_con_aluop[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[0]) );
  DFC3 pipe_con_Ealusrc_reg ( .D(control_o_con_alusrc), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Ealusrc) );
  DFC3 pipe_con_Eregdst_reg ( .D(control_o_con_regdst), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Eregdst) );
  DFC3 pipe_con_MaluPC4_reg ( .D(jbcon_o_con_aluPC4), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Malupc8) );
  DFC3 pipe_con_Mmemread_reg ( .D(control_o_con_memread), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(control_o_con_memwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(control_o_con_memtoreg), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(control_o_con_regwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wregwrite) );
  DFC3 pipe_signext_o_data_immD_reg_31_ ( .D(signext_o_data_immD[31]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[31]) );
  DFC3 pipe_signext_o_data_immD_reg_30_ ( .D(signext_o_data_immD[30]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[30]) );
  DFC3 pipe_signext_o_data_immD_reg_29_ ( .D(signext_o_data_immD[29]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[29]) );
  DFC3 pipe_signext_o_data_immD_reg_28_ ( .D(signext_o_data_immD[28]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[28]) );
  DFC3 pipe_signext_o_data_immD_reg_27_ ( .D(signext_o_data_immD[27]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[27]) );
  DFC3 pipe_signext_o_data_immD_reg_26_ ( .D(signext_o_data_immD[26]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[26]) );
  DFC3 pipe_signext_o_data_immD_reg_25_ ( .D(signext_o_data_immD[25]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[25]) );
  DFC3 pipe_signext_o_data_immD_reg_24_ ( .D(signext_o_data_immD[24]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[24]) );
  DFC3 pipe_signext_o_data_immD_reg_23_ ( .D(signext_o_data_immD[23]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[23]) );
  DFC3 pipe_signext_o_data_immD_reg_22_ ( .D(signext_o_data_immD[22]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[22]) );
  DFC3 pipe_signext_o_data_immD_reg_21_ ( .D(signext_o_data_immD[21]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[21]) );
  DFC3 pipe_signext_o_data_immD_reg_20_ ( .D(signext_o_data_immD[20]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[20]) );
  DFC3 pipe_signext_o_data_immD_reg_19_ ( .D(signext_o_data_immD[19]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[19]) );
  DFC3 pipe_signext_o_data_immD_reg_18_ ( .D(signext_o_data_immD[18]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[18]) );
  DFC3 pipe_signext_o_data_immD_reg_17_ ( .D(signext_o_data_immD[17]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[17]) );
  DFC3 pipe_signext_o_data_immD_reg_16_ ( .D(signext_o_data_immD[16]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[16]) );
  DFC3 pipe_signext_o_data_immD_reg_15_ ( .D(signext_o_data_immD[15]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[15]) );
  DFC3 pipe_signext_o_data_immD_reg_14_ ( .D(signext_o_data_immD[14]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[14]) );
  DFC3 pipe_signext_o_data_immD_reg_13_ ( .D(signext_o_data_immD[13]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[13]) );
  DFC3 pipe_signext_o_data_immD_reg_12_ ( .D(signext_o_data_immD[12]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[12]) );
  DFC3 pipe_signext_o_data_immD_reg_11_ ( .D(signext_o_data_immD[11]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[11]) );
  DFC3 pipe_signext_o_data_immD_reg_10_ ( .D(signext_o_data_immD[10]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[10]) );
  DFC3 pipe_signext_o_data_immD_reg_9_ ( .D(signext_o_data_immD[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[9]) );
  DFC3 pipe_signext_o_data_immD_reg_8_ ( .D(signext_o_data_immD[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[8]) );
  DFC3 pipe_signext_o_data_immD_reg_7_ ( .D(signext_o_data_immD[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[7]) );
  DFC3 pipe_signext_o_data_immD_reg_6_ ( .D(signext_o_data_immD[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[6]) );
  DFC3 pipe_signext_o_data_immD_reg_5_ ( .D(signext_o_data_immD[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[5]) );
  DFC3 pipe_signext_o_data_immD_reg_4_ ( .D(signext_o_data_immD[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[4]) );
  DFC3 pipe_signext_o_data_immD_reg_3_ ( .D(signext_o_data_immD[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[3]) );
  DFC3 pipe_signext_o_data_immD_reg_2_ ( .D(signext_o_data_immD[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[2]) );
  DFC3 pipe_signext_o_data_immD_reg_1_ ( .D(signext_o_data_immD[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[1]) );
  DFC3 pipe_signext_o_data_immD_reg_0_ ( .D(signext_o_data_immD[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[0]) );
  DFC3 pipe_con_Efamux_reg_2_ ( .D(for_o_con_fa[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[2]) );
  DFC3 pipe_con_Efamux_reg_1_ ( .D(for_o_con_fa[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[1]) );
  DFC3 pipe_con_Efamux_reg_0_ ( .D(for_o_con_fa[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[0]) );
  DFC3 pipe_con_Efbmux_reg_2_ ( .D(for_o_con_fb[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[2]) );
  DFC3 pipe_con_Efbmux_reg_1_ ( .D(for_o_con_fb[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[1]) );
  DFC3 pipe_con_Efbmux_reg_0_ ( .D(for_o_con_fb[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[0]) );
  DFC3 pipe_FWmemout_reg_31_ ( .D(i_data_Wmemout[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[31]) );
  DFC3 pipe_FWmemout_reg_30_ ( .D(i_data_Wmemout[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[30]) );
  DFC3 pipe_FWmemout_reg_29_ ( .D(i_data_Wmemout[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[29]) );
  DFC3 pipe_FWmemout_reg_28_ ( .D(i_data_Wmemout[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[28]) );
  DFC3 pipe_FWmemout_reg_27_ ( .D(i_data_Wmemout[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[27]) );
  DFC3 pipe_FWmemout_reg_26_ ( .D(i_data_Wmemout[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[26]) );
  DFC3 pipe_FWmemout_reg_25_ ( .D(i_data_Wmemout[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[25]) );
  DFC3 pipe_FWmemout_reg_24_ ( .D(i_data_Wmemout[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[24]) );
  DFC3 pipe_FWmemout_reg_23_ ( .D(i_data_Wmemout[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[23]) );
  DFC3 pipe_FWmemout_reg_22_ ( .D(i_data_Wmemout[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[22]) );
  DFC3 pipe_FWmemout_reg_21_ ( .D(i_data_Wmemout[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[21]) );
  DFC3 pipe_FWmemout_reg_20_ ( .D(i_data_Wmemout[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[20]) );
  DFC3 pipe_FWmemout_reg_18_ ( .D(i_data_Wmemout[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[18]) );
  DFC3 pipe_FWmemout_reg_17_ ( .D(i_data_Wmemout[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[17]) );
  DFC3 pipe_FWmemout_reg_16_ ( .D(i_data_Wmemout[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[16]) );
  DFC3 pipe_FWmemout_reg_15_ ( .D(i_data_Wmemout[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[15]) );
  DFC3 pipe_FWmemout_reg_14_ ( .D(i_data_Wmemout[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[14]) );
  DFC3 pipe_FWmemout_reg_13_ ( .D(i_data_Wmemout[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[13]) );
  DFC3 pipe_FWmemout_reg_11_ ( .D(i_data_Wmemout[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[11]) );
  DFC3 pipe_FWmemout_reg_10_ ( .D(i_data_Wmemout[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[10]) );
  DFC3 pipe_FWmemout_reg_9_ ( .D(i_data_Wmemout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[9]) );
  DFC3 pipe_FWmemout_reg_8_ ( .D(i_data_Wmemout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[8]) );
  DFC3 pipe_FWmemout_reg_6_ ( .D(i_data_Wmemout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[6]) );
  DFC3 pipe_FWmemout_reg_4_ ( .D(i_data_Wmemout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[4]) );
  DFC3 pipe_FWmemout_reg_2_ ( .D(i_data_Wmemout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[2]) );
  DFC3 pipe_FWmemout_reg_1_ ( .D(i_data_Wmemout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[1]) );
  DFC3 pipe_FWmemout_reg_0_ ( .D(i_data_Wmemout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[0]) );
  DFC3 pipe_addr_branch_reg_31_ ( .D(pcadd_o_addr_pcbranchE[31]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[31]) );
  DFC3 pipe_addr_branch_reg_30_ ( .D(pcadd_o_addr_pcbranchE[30]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[30]) );
  DFC3 pipe_addr_branch_reg_29_ ( .D(pcadd_o_addr_pcbranchE[29]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[29]) );
  DFC3 pipe_addr_branch_reg_28_ ( .D(pcadd_o_addr_pcbranchE[28]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[28]) );
  DFC3 pipe_addr_branch_reg_27_ ( .D(pcadd_o_addr_pcbranchE[27]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[27]) );
  DFC3 pipe_addr_branch_reg_26_ ( .D(pcadd_o_addr_pcbranchE[26]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[26]) );
  DFC3 pipe_addr_branch_reg_25_ ( .D(pcadd_o_addr_pcbranchE[25]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[25]) );
  DFC3 pipe_addr_branch_reg_24_ ( .D(pcadd_o_addr_pcbranchE[24]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[24]) );
  DFC3 pipe_addr_branch_reg_23_ ( .D(pcadd_o_addr_pcbranchE[23]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[23]) );
  DFC3 pipe_addr_branch_reg_22_ ( .D(pcadd_o_addr_pcbranchE[22]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[22]) );
  DFC3 pipe_addr_branch_reg_21_ ( .D(pcadd_o_addr_pcbranchE[21]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[21]) );
  DFC3 pipe_addr_branch_reg_20_ ( .D(pcadd_o_addr_pcbranchE[20]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[20]) );
  DFC3 pipe_addr_branch_reg_19_ ( .D(pcadd_o_addr_pcbranchE[19]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[19]) );
  DFC3 pipe_addr_branch_reg_18_ ( .D(pcadd_o_addr_pcbranchE[18]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[18]) );
  DFC3 pipe_addr_branch_reg_17_ ( .D(pcadd_o_addr_pcbranchE[17]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[17]) );
  DFC3 pipe_addr_branch_reg_16_ ( .D(pcadd_o_addr_pcbranchE[16]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[16]) );
  DFC3 pipe_addr_branch_reg_15_ ( .D(pcadd_o_addr_pcbranchE[15]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[15]) );
  DFC3 pipe_addr_branch_reg_14_ ( .D(pcadd_o_addr_pcbranchE[14]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[14]) );
  DFC3 pipe_addr_branch_reg_13_ ( .D(pcadd_o_addr_pcbranchE[13]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[13]) );
  DFC3 pipe_addr_branch_reg_12_ ( .D(pcadd_o_addr_pcbranchE[12]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[12]) );
  DFC3 pipe_addr_branch_reg_11_ ( .D(pcadd_o_addr_pcbranchE[11]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[11]) );
  DFC3 pipe_addr_branch_reg_10_ ( .D(pcadd_o_addr_pcbranchE[10]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[10]) );
  DFC3 pipe_addr_branch_reg_9_ ( .D(pcadd_o_addr_pcbranchE[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[9]) );
  DFC3 pipe_addr_branch_reg_8_ ( .D(pcadd_o_addr_pcbranchE[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[8]) );
  DFC3 pipe_addr_branch_reg_7_ ( .D(pcadd_o_addr_pcbranchE[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[7]) );
  DFC3 pipe_addr_branch_reg_6_ ( .D(pcadd_o_addr_pcbranchE[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[6]) );
  DFC3 pipe_addr_branch_reg_5_ ( .D(pcadd_o_addr_pcbranchE[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[5]) );
  DFC3 pipe_addr_branch_reg_4_ ( .D(pcadd_o_addr_pcbranchE[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[4]) );
  DFC3 pipe_addr_branch_reg_3_ ( .D(pcadd_o_addr_pcbranchE[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[3]) );
  DFC3 pipe_addr_branch_reg_2_ ( .D(pcadd_o_addr_pcbranchE[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[2]) );
  DFC3 pipe_addr_branch_reg_1_ ( .D(pcadd_o_addr_pcbranchE[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[1]) );
  DFC3 pipe_addr_branch_reg_0_ ( .D(pcadd_o_addr_pcbranchE[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[0]) );
  D_control u_control ( .o_con_regdst(control_o_con_regdst), .o_con_memread(
        control_o_con_memread), .o_con_memtoreg(control_o_con_memtoreg), 
        .o_con_memwrite(control_o_con_memwrite), .o_con_alusrc(
        control_o_con_alusrc), .o_con_regwrite(control_o_con_regwrite), 
        .o_con_ifsign(signext_i_con_signext), .o_con_aluop(control_o_con_aluop), .i_con_instru(i_data_instr[31:26]) );
  D_jb_control u_jb_control ( .o_con_jump(o_con_jump), .o_con_bop(
        jbcon_o_con_bop), .o_con_aluPC4(jbcon_o_con_aluPC4), .o_con_ifstall(
        o_con_ifstall), .i_con_instru(i_data_instr[31:26]), .i_con_func(
        i_data_instr[5:0]), .i_con_rt(i_data_instr[16]) );
  D_pcadd u_pcadd ( .i_addr_pcadd4E(i_addr_pc4), .i_data_immshiftl({
        pcadd_i_data_immshiftl, o_addr_jump[0], o_addr_jump[0]}), 
        .o_addr_pcbranchE(pcadd_o_addr_pcbranchE) );
  D_register_bank u_regbank ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_addr_Rs(
        i_data_instr[25:21]), .i_addr_Rt(i_data_instr[20:16]), .i_con_RegWr(
        i_con_Wregwrite), .i_addr_Rd(i_addr_Wregwrite), .i_data_Rd(
        i_data_Wregwrite), .o_data_Rs(o_data_jr), .o_data_Rt(regbank_o_data_Rt) );
  D_shiftleft u_sl ( .i_data_immE(i_data_instr[15:0]), .o_data_immshiftl({
        pcadd_i_data_immshiftl, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}) );
  D_sign_extend u_signext ( .i_data_immD(i_data_instr[15:0]), .i_con_signext(
        signext_i_con_signext), .o_data_immD(signext_o_data_immD) );
  D_jump_ext u_jump_ext ( .i_addr_j(i_data_instr[25:0]), .i_PC4_j(
        i_addr_pc4[31:28]), .o_addr_j({o_addr_jump[31:2], 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4}) );
  D_forward u_forward ( .i_addr_rs(i_data_instr[25:21]), .i_addr_rt(
        i_data_instr[20:16]), .i_addr_rdE(i_addr_Erd), .i_addr_rdM(i_addr_Mrd), 
        .i_addr_rtM(i_addr_rtM), .i_addr_rtW(i_addr_rtW), .i_con_regwriteE(
        i_con_Eregwrite), .i_con_regwriteM(i_con_Mregwrite), .i_con_memreadM(
        i_con_memreadM), .i_con_memreadW(i_con_memreadW), .o_con_fa(
        for_o_con_fa), .o_con_fb(for_o_con_fb) );
  DFC1 pipe_FWmemout_reg_3_ ( .D(i_data_Wmemout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[3]) );
  DFC1 pipe_FWmemout_reg_19_ ( .D(i_data_Wmemout[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[19]) );
  DFC1 pipe_FWmemout_reg_5_ ( .D(i_data_Wmemout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[5]) );
  DFC1 pipe_FWmemout_reg_12_ ( .D(i_data_Wmemout[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[12]) );
  DFC3 pipe_FWmemout_reg_7_ ( .D(i_data_Wmemout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[7]) );
  LOGIC0 U3 ( .Q(o_addr_jump[0]) );
endmodule


module E_alu_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392;

  NAND23 U2 ( .A(n220), .B(n197), .Q(n215) );
  CLKIN6 U3 ( .A(B[13]), .Q(n336) );
  NAND22 U4 ( .A(B[2]), .B(A[2]), .Q(n381) );
  XOR22 U5 ( .A(n99), .B(n100), .Q(SUM[28]) );
  NOR20 U6 ( .A(B[24]), .B(A[24]), .Q(n105) );
  INV1 U7 ( .A(B[24]), .Q(n113) );
  NOR22 U8 ( .A(n307), .B(n308), .Q(n306) );
  NAND26 U9 ( .A(n134), .B(n135), .Q(n102) );
  NOR32 U10 ( .A(n289), .B(n180), .C(n290), .Q(n288) );
  NAND23 U11 ( .A(n350), .B(n351), .Q(n289) );
  NAND23 U12 ( .A(n160), .B(n161), .Q(n299) );
  NAND33 U13 ( .A(n102), .B(n103), .C(n104), .Q(n78) );
  AOI220 U14 ( .A(B[27]), .B(A[27]), .C(n114), .D(n102), .Q(n107) );
  AOI312 U15 ( .A(n89), .B(n90), .C(n91), .D(n72), .Q(n88) );
  NOR21 U16 ( .A(n380), .B(n381), .Q(n293) );
  NOR22 U17 ( .A(n292), .B(n293), .Q(n379) );
  NOR23 U18 ( .A(n2), .B(n7), .Q(n8) );
  INV3 U19 ( .A(n1), .Q(n2) );
  NAND22 U20 ( .A(B[9]), .B(A[9]), .Q(n19) );
  INV3 U21 ( .A(n190), .Q(n196) );
  INV2 U22 ( .A(A[22]), .Q(n217) );
  OAI2112 U23 ( .A(n202), .B(n206), .C(n207), .D(n199), .Q(n205) );
  XOR21 U24 ( .A(n136), .B(n137), .Q(SUM[25]) );
  AOI212 U25 ( .A(n133), .B(n91), .C(n138), .Q(n137) );
  NOR21 U26 ( .A(A[3]), .B(B[3]), .Q(n389) );
  NOR23 U27 ( .A(A[1]), .B(B[1]), .Q(n86) );
  INV0 U28 ( .A(A[23]), .Q(n201) );
  NOR21 U29 ( .A(B[15]), .B(A[15]), .Q(n314) );
  NAND22 U30 ( .A(n386), .B(n387), .Q(n177) );
  NAND23 U31 ( .A(n336), .B(n337), .Q(n304) );
  INV3 U32 ( .A(n5), .Q(n6) );
  NAND22 U33 ( .A(n375), .B(n376), .Q(n290) );
  INV6 U34 ( .A(n322), .Q(n39) );
  NAND22 U35 ( .A(n261), .B(n4), .Q(n253) );
  NOR21 U36 ( .A(n310), .B(n267), .Q(n261) );
  AOI211 U37 ( .A(n236), .B(n237), .C(n266), .Q(n284) );
  XOR21 U38 ( .A(n268), .B(n269), .Q(SUM[18]) );
  AOI211 U39 ( .A(n12), .B(n117), .C(n118), .Q(n116) );
  NAND31 U40 ( .A(n178), .B(n162), .C(n179), .Q(n151) );
  AOI221 U41 ( .A(B[23]), .B(A[23]), .C(n194), .D(n195), .Q(n184) );
  INV3 U42 ( .A(n125), .Q(n77) );
  NAND24 U43 ( .A(n379), .B(n6), .Q(n322) );
  NAND22 U44 ( .A(n287), .B(n288), .Q(n260) );
  NAND22 U45 ( .A(n224), .B(n225), .Q(n190) );
  NOR21 U46 ( .A(n241), .B(n242), .Q(n148) );
  AOI211 U47 ( .A(n112), .B(n113), .C(n138), .Q(n142) );
  AOI211 U48 ( .A(n253), .B(n254), .C(n235), .Q(n252) );
  NOR21 U49 ( .A(n256), .B(n257), .Q(n254) );
  NAND22 U50 ( .A(n304), .B(n301), .Q(n331) );
  XOR21 U51 ( .A(n364), .B(n365), .Q(SUM[10]) );
  INV3 U52 ( .A(n289), .Q(n179) );
  NOR22 U53 ( .A(n8), .B(n129), .Q(n128) );
  NAND22 U54 ( .A(n120), .B(n123), .Q(n129) );
  NAND22 U55 ( .A(n15), .B(n16), .Q(n362) );
  NOR22 U56 ( .A(A[5]), .B(B[5]), .Q(n35) );
  NAND43 U57 ( .A(n181), .B(n183), .C(n286), .D(n260), .Q(n56) );
  INV3 U58 ( .A(n371), .Q(n374) );
  INV3 U59 ( .A(n265), .Q(n276) );
  INV3 U60 ( .A(n19), .Q(n349) );
  INV3 U61 ( .A(B[25]), .Q(n140) );
  NAND21 U62 ( .A(B[2]), .B(A[2]), .Q(n48) );
  NAND21 U63 ( .A(B[22]), .B(A[22]), .Q(n199) );
  NOR21 U64 ( .A(n125), .B(n132), .Q(n1) );
  INV3 U65 ( .A(n12), .Q(n7) );
  NAND22 U66 ( .A(n291), .B(n6), .Q(n287) );
  NAND31 U67 ( .A(n262), .B(n260), .C(n263), .Q(n3) );
  INV3 U68 ( .A(n3), .Q(n4) );
  INV0 U69 ( .A(n264), .Q(n263) );
  INV3 U70 ( .A(n16), .Q(n22) );
  INV0 U71 ( .A(n348), .Q(n391) );
  NOR20 U72 ( .A(n347), .B(n348), .Q(n358) );
  NOR21 U73 ( .A(n347), .B(n348), .Q(n351) );
  XOR22 U74 ( .A(n25), .B(n26), .Q(SUM[7]) );
  XOR22 U75 ( .A(n87), .B(n88), .Q(SUM[29]) );
  INV1 U76 ( .A(A[16]), .Q(n236) );
  NOR21 U77 ( .A(B[23]), .B(A[23]), .Q(n193) );
  XNR20 U78 ( .A(B[30]), .B(A[30]), .Q(n65) );
  INV0 U79 ( .A(n78), .Q(n90) );
  NOR22 U80 ( .A(A[6]), .B(B[6]), .Q(n371) );
  NAND33 U81 ( .A(n189), .B(n190), .C(n191), .Q(n150) );
  NOR22 U82 ( .A(n192), .B(n193), .Q(n191) );
  NAND31 U83 ( .A(n175), .B(n176), .C(n177), .Q(n172) );
  NAND21 U84 ( .A(n206), .B(n198), .Q(n214) );
  NAND21 U85 ( .A(n215), .B(n190), .Q(n206) );
  NOR22 U86 ( .A(A[10]), .B(B[10]), .Q(n348) );
  NAND21 U87 ( .A(n130), .B(n103), .Q(n123) );
  NOR32 U88 ( .A(n289), .B(n180), .C(n311), .Q(n310) );
  INV2 U89 ( .A(n180), .Q(n162) );
  NAND20 U90 ( .A(B[24]), .B(A[24]), .Q(n131) );
  INV1 U91 ( .A(A[24]), .Q(n112) );
  NAND23 U92 ( .A(n305), .B(n306), .Q(n183) );
  XNR22 U93 ( .A(n9), .B(n203), .Q(SUM[23]) );
  NOR20 U94 ( .A(B[12]), .B(A[12]), .Q(n354) );
  NOR20 U95 ( .A(A[12]), .B(B[12]), .Q(n335) );
  NAND34 U96 ( .A(n303), .B(n304), .C(n312), .Q(n180) );
  NOR22 U97 ( .A(A[3]), .B(B[3]), .Q(n380) );
  NAND24 U98 ( .A(n148), .B(n149), .Q(n125) );
  NAND21 U99 ( .A(n148), .B(n223), .Q(n210) );
  NAND20 U100 ( .A(B[1]), .B(A[1]), .Q(n82) );
  CLKIN0 U101 ( .A(A[1]), .Q(n384) );
  NOR21 U102 ( .A(n35), .B(n371), .Q(n376) );
  NAND32 U103 ( .A(n181), .B(n182), .C(n183), .Q(n146) );
  INV3 U104 ( .A(B[22]), .Q(n216) );
  NOR22 U105 ( .A(A[9]), .B(B[9]), .Q(n347) );
  NAND21 U106 ( .A(B[7]), .B(A[7]), .Q(n311) );
  NAND24 U107 ( .A(n144), .B(n145), .Q(n91) );
  NAND22 U108 ( .A(n177), .B(n174), .Q(n5) );
  NAND20 U109 ( .A(B[3]), .B(A[3]), .Q(n174) );
  AOI211 U110 ( .A(n178), .B(n322), .C(n323), .Q(n319) );
  NAND20 U111 ( .A(B[16]), .B(A[16]), .Q(n277) );
  INV1 U112 ( .A(B[16]), .Q(n237) );
  NAND21 U113 ( .A(B[21]), .B(A[21]), .Q(n198) );
  NAND20 U114 ( .A(B[0]), .B(A[0]), .Q(n250) );
  IMUX20 U115 ( .A(n392), .B(B[0]), .S(A[0]), .Q(SUM[0]) );
  BUF15 U116 ( .A(n56), .Q(n12) );
  NAND21 U117 ( .A(n298), .B(n19), .Q(n296) );
  AOI312 U118 ( .A(n294), .B(n169), .C(n295), .D(n180), .Q(n264) );
  NOR22 U119 ( .A(n52), .B(n380), .Q(n383) );
  NOR22 U120 ( .A(n389), .B(n52), .Q(n386) );
  NOR23 U121 ( .A(A[2]), .B(B[2]), .Q(n52) );
  XOR22 U122 ( .A(n127), .B(n128), .Q(SUM[26]) );
  NAND22 U123 ( .A(B[6]), .B(A[6]), .Q(n36) );
  INV0 U124 ( .A(n308), .Q(n367) );
  INV2 U125 ( .A(A[14]), .Q(n330) );
  NOR21 U126 ( .A(n188), .B(n222), .Q(n221) );
  NAND22 U127 ( .A(n221), .B(n187), .Q(n220) );
  CLKIN6 U128 ( .A(B[14]), .Q(n329) );
  OAI2111 U129 ( .A(n119), .B(n120), .C(n121), .D(n111), .Q(n118) );
  INV1 U130 ( .A(n174), .Q(n173) );
  NAND20 U131 ( .A(n122), .B(n102), .Q(n121) );
  CLKIN0 U132 ( .A(n233), .Q(n257) );
  CLKIN3 U133 ( .A(B[18]), .Q(n279) );
  NAND22 U134 ( .A(n184), .B(n185), .Q(n76) );
  NOR31 U135 ( .A(n35), .B(n372), .C(n373), .Q(n370) );
  NAND20 U136 ( .A(n171), .B(n19), .Q(n170) );
  INV2 U137 ( .A(n132), .Q(n126) );
  AOI211 U138 ( .A(n283), .B(n12), .C(n266), .Q(n282) );
  NAND20 U139 ( .A(n179), .B(n334), .Q(n320) );
  NOR20 U140 ( .A(n244), .B(n274), .Q(n259) );
  CLKIN1 U141 ( .A(n74), .Q(n73) );
  NAND20 U142 ( .A(n160), .B(n161), .Q(n158) );
  INV2 U143 ( .A(A[13]), .Q(n337) );
  NOR21 U144 ( .A(n258), .B(n259), .Q(n256) );
  XNR21 U145 ( .A(n331), .B(n327), .Q(SUM[13]) );
  CLKIN0 U146 ( .A(n274), .Q(n283) );
  NOR21 U147 ( .A(n97), .B(n79), .Q(n96) );
  NOR20 U148 ( .A(n81), .B(n52), .Q(n80) );
  CLKIN1 U149 ( .A(n157), .Q(n156) );
  NAND22 U150 ( .A(n158), .B(n159), .Q(n155) );
  INV0 U151 ( .A(n131), .Q(n138) );
  AOI312 U152 ( .A(n303), .B(n304), .C(n317), .D(n318), .Q(n316) );
  NOR22 U153 ( .A(n342), .B(n343), .Q(n168) );
  AOI221 U154 ( .A(n98), .B(n101), .C(n90), .D(n91), .Q(n100) );
  NOR20 U155 ( .A(n354), .B(n332), .Q(n338) );
  CLKIN3 U156 ( .A(B[4]), .Q(n373) );
  INV2 U157 ( .A(n139), .Q(n133) );
  NOR21 U158 ( .A(n377), .B(n378), .Q(n375) );
  CLKIN0 U159 ( .A(n79), .Q(n89) );
  NAND20 U160 ( .A(n303), .B(n159), .Q(n325) );
  NAND20 U161 ( .A(n189), .B(n199), .Q(n211) );
  NAND20 U162 ( .A(n190), .B(n198), .Q(n218) );
  CLKIN3 U163 ( .A(n165), .Q(n297) );
  NAND20 U164 ( .A(n208), .B(n189), .Q(n207) );
  NAND20 U165 ( .A(n276), .B(n277), .Q(n275) );
  NAND20 U166 ( .A(n190), .B(n189), .Q(n209) );
  NAND20 U167 ( .A(n233), .B(n255), .Q(n268) );
  NAND20 U168 ( .A(n131), .B(n115), .Q(n130) );
  XOR20 U169 ( .A(n50), .B(n80), .Q(SUM[2]) );
  NAND20 U170 ( .A(n103), .B(n115), .Q(n136) );
  XOR20 U171 ( .A(n33), .B(n37), .Q(SUM[5]) );
  NAND20 U172 ( .A(n133), .B(n103), .Q(n132) );
  NAND20 U173 ( .A(n102), .B(n111), .Q(n127) );
  NAND20 U174 ( .A(n126), .B(n102), .Q(n124) );
  NAND21 U175 ( .A(n24), .B(n362), .Q(n366) );
  NAND21 U176 ( .A(n162), .B(n163), .Q(n153) );
  INV0 U177 ( .A(n97), .Q(n101) );
  CLKIN1 U178 ( .A(n63), .Q(n70) );
  INV0 U179 ( .A(n197), .Q(n247) );
  NOR20 U180 ( .A(n188), .B(n230), .Q(n229) );
  XOR20 U181 ( .A(B[23]), .B(A[23]), .Q(n9) );
  XNR21 U182 ( .A(n10), .B(n116), .Q(SUM[27]) );
  XOR20 U183 ( .A(B[27]), .B(A[27]), .Q(n10) );
  NOR22 U184 ( .A(n86), .B(n388), .Q(n387) );
  NAND20 U185 ( .A(B[12]), .B(A[12]), .Q(n300) );
  AOI212 U186 ( .A(n27), .B(n374), .C(n28), .Q(n26) );
  NAND22 U187 ( .A(n368), .B(n369), .Q(n309) );
  NAND20 U188 ( .A(B[8]), .B(A[8]), .Q(n298) );
  INV2 U189 ( .A(n96), .Q(n93) );
  INV0 U190 ( .A(A[28]), .Q(n94) );
  INV0 U191 ( .A(B[28]), .Q(n95) );
  OAI2110 U192 ( .A(n341), .B(n165), .C(n169), .D(n294), .Q(n333) );
  AOI210 U193 ( .A(n15), .B(n16), .C(n17), .Q(n14) );
  NAND20 U194 ( .A(n18), .B(n19), .Q(n13) );
  IMUX20 U195 ( .A(n20), .B(n21), .S(n22), .Q(SUM[8]) );
  NOR20 U196 ( .A(B[20]), .B(A[20]), .Q(n192) );
  NOR20 U197 ( .A(A[20]), .B(B[20]), .Q(n222) );
  NAND20 U198 ( .A(B[15]), .B(A[15]), .Q(n182) );
  NAND20 U199 ( .A(B[17]), .B(A[17]), .Q(n278) );
  IMUX20 U200 ( .A(n143), .B(n142), .S(n91), .Q(SUM[24]) );
  IMUX20 U201 ( .A(n42), .B(n43), .S(n39), .Q(SUM[4]) );
  AOI210 U202 ( .A(n179), .B(n16), .C(n333), .Q(n340) );
  NAND20 U203 ( .A(B[8]), .B(A[8]), .Q(n171) );
  NAND20 U204 ( .A(B[12]), .B(A[12]), .Q(n355) );
  NAND20 U205 ( .A(A[30]), .B(B[30]), .Q(n61) );
  INV0 U206 ( .A(A[17]), .Q(n240) );
  INV0 U207 ( .A(A[20]), .Q(n245) );
  NOR21 U208 ( .A(n310), .B(n267), .Q(n272) );
  AOI211 U209 ( .A(n67), .B(n12), .C(n68), .Q(n66) );
  NAND22 U210 ( .A(n62), .B(n69), .Q(n68) );
  NOR21 U211 ( .A(n70), .B(n71), .Q(n69) );
  NAND22 U212 ( .A(n77), .B(n75), .Q(n64) );
  NOR21 U213 ( .A(n265), .B(n264), .Q(n286) );
  NOR21 U214 ( .A(n362), .B(n363), .Q(n360) );
  INV3 U215 ( .A(n358), .Q(n363) );
  INV3 U216 ( .A(n259), .Q(n273) );
  NAND22 U217 ( .A(n311), .B(n324), .Q(n323) );
  NAND22 U218 ( .A(n296), .B(n297), .Q(n295) );
  INV3 U219 ( .A(n168), .Q(n294) );
  OAI2111 U220 ( .A(n196), .B(n197), .C(n198), .D(n199), .Q(n195) );
  NOR31 U221 ( .A(n78), .B(n79), .C(n74), .Q(n75) );
  XOR21 U222 ( .A(n211), .B(n212), .Q(SUM[22]) );
  AOI2111 U223 ( .A(n55), .B(n12), .C(n57), .D(n58), .Q(n54) );
  NOR21 U224 ( .A(n64), .B(n59), .Q(n55) );
  OAI2111 U225 ( .A(n151), .B(n152), .C(n153), .D(n154), .Q(n147) );
  NOR21 U226 ( .A(n292), .B(n293), .Q(n291) );
  NAND22 U227 ( .A(n367), .B(n309), .Q(n324) );
  NAND22 U228 ( .A(n391), .B(n343), .Q(n364) );
  AOI211 U229 ( .A(n366), .B(n18), .C(n349), .Q(n365) );
  XOR21 U230 ( .A(n281), .B(n282), .Q(SUM[17]) );
  NAND22 U231 ( .A(n243), .B(n278), .Q(n281) );
  XOR21 U232 ( .A(n29), .B(n30), .Q(SUM[6]) );
  NAND22 U233 ( .A(n374), .B(n36), .Q(n29) );
  INV3 U234 ( .A(n222), .Q(n223) );
  NAND22 U235 ( .A(n126), .B(n76), .Q(n120) );
  XOR21 U236 ( .A(n325), .B(n326), .Q(SUM[14]) );
  XOR21 U237 ( .A(n218), .B(n219), .Q(SUM[21]) );
  NAND22 U238 ( .A(n72), .B(n73), .Q(n60) );
  NAND22 U239 ( .A(n75), .B(n76), .Q(n62) );
  NAND22 U240 ( .A(n303), .B(n304), .Q(n302) );
  NOR21 U241 ( .A(n180), .B(n289), .Q(n305) );
  INV3 U242 ( .A(n309), .Q(n307) );
  NOR22 U243 ( .A(n258), .B(n270), .Q(n269) );
  INV3 U244 ( .A(n310), .Q(n181) );
  NAND22 U245 ( .A(n31), .B(n32), .Q(n27) );
  NAND22 U246 ( .A(n33), .B(n34), .Q(n32) );
  INV3 U247 ( .A(n35), .Q(n34) );
  NOR21 U248 ( .A(n35), .B(n38), .Q(n37) );
  INV3 U249 ( .A(n31), .Q(n38) );
  XOR21 U250 ( .A(n65), .B(n66), .Q(SUM[30]) );
  NAND22 U251 ( .A(n155), .B(n156), .Q(n154) );
  NOR21 U252 ( .A(n236), .B(n237), .Q(n234) );
  INV3 U253 ( .A(n170), .Q(n164) );
  NOR21 U254 ( .A(n167), .B(n168), .Q(n166) );
  NOR21 U255 ( .A(n209), .B(n210), .Q(n204) );
  INV3 U256 ( .A(n293), .Q(n175) );
  INV3 U257 ( .A(n98), .Q(n92) );
  XOR21 U258 ( .A(n84), .B(n248), .Q(SUM[1]) );
  NOR21 U259 ( .A(n249), .B(n86), .Q(n248) );
  NAND22 U260 ( .A(n24), .B(n19), .Q(n359) );
  INV3 U261 ( .A(n347), .Q(n18) );
  NAND22 U262 ( .A(n82), .B(n83), .Q(n50) );
  NAND22 U263 ( .A(n84), .B(n85), .Q(n83) );
  INV3 U264 ( .A(n86), .Q(n85) );
  INV3 U265 ( .A(n52), .Q(n51) );
  XOR21 U266 ( .A(n13), .B(n14), .Q(SUM[9]) );
  XOR21 U267 ( .A(n315), .B(n316), .Q(SUM[15]) );
  NOR22 U268 ( .A(n313), .B(n314), .Q(n312) );
  NOR21 U269 ( .A(B[12]), .B(A[12]), .Q(n313) );
  INV3 U270 ( .A(A[21]), .Q(n225) );
  INV3 U271 ( .A(B[21]), .Q(n224) );
  NAND22 U272 ( .A(n140), .B(n141), .Q(n103) );
  NOR21 U273 ( .A(A[17]), .B(B[17]), .Q(n244) );
  NAND22 U274 ( .A(n233), .B(n243), .Q(n241) );
  INV3 U275 ( .A(n244), .Q(n243) );
  NAND22 U276 ( .A(n216), .B(n217), .Q(n189) );
  NOR21 U277 ( .A(n352), .B(n353), .Q(n350) );
  NOR21 U278 ( .A(B[11]), .B(A[11]), .Q(n352) );
  NAND22 U279 ( .A(n279), .B(n280), .Q(n233) );
  NOR21 U280 ( .A(n105), .B(n106), .Q(n104) );
  INV3 U281 ( .A(B[26]), .Q(n134) );
  NAND22 U282 ( .A(n231), .B(n232), .Q(n187) );
  AOI311 U283 ( .A(n243), .B(n233), .C(n234), .D(n235), .Q(n232) );
  NOR21 U284 ( .A(n239), .B(n240), .Q(n238) );
  NAND22 U285 ( .A(n370), .B(n374), .Q(n369) );
  NAND22 U286 ( .A(n344), .B(n345), .Q(n165) );
  INV3 U287 ( .A(n346), .Q(n345) );
  NOR22 U288 ( .A(n347), .B(n348), .Q(n344) );
  NAND24 U289 ( .A(n329), .B(n330), .Q(n303) );
  NAND22 U290 ( .A(n300), .B(n301), .Q(n161) );
  XOR21 U291 ( .A(n53), .B(n54), .Q(SUM[31]) );
  NAND22 U292 ( .A(n382), .B(n383), .Q(n176) );
  NOR21 U293 ( .A(n384), .B(n385), .Q(n382) );
  IMUX21 U294 ( .A(n226), .B(n227), .S(n228), .Q(SUM[20]) );
  AOI211 U295 ( .A(n245), .B(n246), .C(n247), .Q(n226) );
  AOI211 U296 ( .A(n148), .B(n12), .C(n229), .Q(n228) );
  AOI211 U297 ( .A(n200), .B(n201), .C(n202), .Q(n194) );
  INV3 U298 ( .A(B[23]), .Q(n200) );
  NAND22 U299 ( .A(n107), .B(n108), .Q(n98) );
  AOI311 U300 ( .A(n102), .B(n103), .C(n109), .D(n110), .Q(n108) );
  NOR21 U301 ( .A(n112), .B(n113), .Q(n109) );
  NOR21 U302 ( .A(n44), .B(n45), .Q(n42) );
  IMUX21 U303 ( .A(n285), .B(n284), .S(n12), .Q(SUM[16]) );
  NOR21 U304 ( .A(n23), .B(n17), .Q(n20) );
  IMUX21 U305 ( .A(n338), .B(n339), .S(n340), .Q(SUM[12]) );
  NOR21 U306 ( .A(n124), .B(n125), .Q(n117) );
  XOR21 U307 ( .A(n251), .B(n252), .Q(SUM[19]) );
  XOR21 U308 ( .A(n356), .B(n357), .Q(SUM[11]) );
  AOI2111 U309 ( .A(n358), .B(n359), .C(n360), .D(n361), .Q(n357) );
  INV3 U310 ( .A(n343), .Q(n361) );
  NAND22 U311 ( .A(n186), .B(n187), .Q(n185) );
  NOR21 U312 ( .A(n188), .B(n150), .Q(n186) );
  INV3 U313 ( .A(n390), .Q(n15) );
  INV3 U314 ( .A(n335), .Q(n334) );
  INV3 U315 ( .A(B[17]), .Q(n239) );
  INV3 U316 ( .A(B[1]), .Q(n385) );
  XOR21 U317 ( .A(n46), .B(n47), .Q(SUM[3]) );
  NAND22 U318 ( .A(n48), .B(n49), .Q(n46) );
  NAND22 U319 ( .A(n50), .B(n51), .Q(n49) );
  INV3 U320 ( .A(n250), .Q(n84) );
  INV3 U321 ( .A(B[0]), .Q(n392) );
  AOI211 U322 ( .A(n327), .B(n304), .C(n328), .Q(n326) );
  AOI221 U323 ( .A(B[19]), .B(A[19]), .C(n238), .D(n233), .Q(n231) );
  XNR21 U324 ( .A(B[28]), .B(A[28]), .Q(n99) );
  NOR21 U325 ( .A(A[28]), .B(B[28]), .Q(n79) );
  NAND22 U326 ( .A(B[0]), .B(A[0]), .Q(n388) );
  NAND22 U327 ( .A(B[18]), .B(A[18]), .Q(n255) );
  INV3 U328 ( .A(A[18]), .Q(n280) );
  NOR21 U329 ( .A(n172), .B(n173), .Q(n152) );
  NOR21 U330 ( .A(A[27]), .B(B[27]), .Q(n97) );
  NOR21 U331 ( .A(B[27]), .B(A[27]), .Q(n106) );
  INV3 U332 ( .A(A[26]), .Q(n135) );
  NOR20 U333 ( .A(A[16]), .B(B[16]), .Q(n274) );
  XNR20 U334 ( .A(B[16]), .B(A[16]), .Q(n285) );
  OAI220 U335 ( .A(B[19]), .B(A[19]), .C(B[16]), .D(A[16]), .Q(n242) );
  XNR21 U336 ( .A(B[29]), .B(A[29]), .Q(n87) );
  NAND22 U337 ( .A(B[29]), .B(A[29]), .Q(n63) );
  NOR21 U338 ( .A(A[29]), .B(B[29]), .Q(n74) );
  NAND22 U339 ( .A(B[10]), .B(A[10]), .Q(n343) );
  NAND22 U340 ( .A(B[26]), .B(A[26]), .Q(n111) );
  NOR21 U341 ( .A(A[11]), .B(B[11]), .Q(n342) );
  NAND21 U342 ( .A(B[11]), .B(A[11]), .Q(n169) );
  NOR21 U343 ( .A(A[11]), .B(B[11]), .Q(n346) );
  XNR20 U344 ( .A(B[11]), .B(A[11]), .Q(n356) );
  NAND22 U345 ( .A(B[5]), .B(A[5]), .Q(n31) );
  AOI312 U346 ( .A(A[5]), .B(B[5]), .C(n374), .D(n28), .Q(n368) );
  XNR20 U347 ( .A(B[19]), .B(A[19]), .Q(n251) );
  NOR21 U348 ( .A(A[19]), .B(B[19]), .Q(n188) );
  XNR20 U349 ( .A(B[12]), .B(A[12]), .Q(n339) );
  OAI2111 U350 ( .A(n319), .B(n320), .C(n321), .D(n301), .Q(n317) );
  NOR21 U351 ( .A(n264), .B(n275), .Q(n271) );
  XOR20 U352 ( .A(B[3]), .B(A[3]), .Q(n47) );
  XNR20 U353 ( .A(B[15]), .B(A[15]), .Q(n315) );
  NOR21 U354 ( .A(A[15]), .B(B[15]), .Q(n157) );
  INV0 U355 ( .A(A[25]), .Q(n141) );
  NAND22 U356 ( .A(B[25]), .B(A[25]), .Q(n115) );
  NOR21 U357 ( .A(B[4]), .B(A[4]), .Q(n377) );
  INV3 U358 ( .A(A[4]), .Q(n372) );
  NOR20 U359 ( .A(B[4]), .B(A[4]), .Q(n44) );
  NAND20 U360 ( .A(B[4]), .B(A[4]), .Q(n41) );
  XNR20 U361 ( .A(B[4]), .B(A[4]), .Q(n43) );
  NOR20 U362 ( .A(A[4]), .B(B[4]), .Q(n40) );
  XNR20 U363 ( .A(B[31]), .B(A[31]), .Q(n53) );
  NAND22 U364 ( .A(B[14]), .B(A[14]), .Q(n159) );
  NOR20 U365 ( .A(A[24]), .B(B[24]), .Q(n139) );
  NOR20 U366 ( .A(B[8]), .B(A[8]), .Q(n23) );
  NAND22 U367 ( .A(B[8]), .B(A[8]), .Q(n24) );
  NOR20 U368 ( .A(A[8]), .B(B[8]), .Q(n390) );
  NOR21 U369 ( .A(B[8]), .B(A[8]), .Q(n353) );
  XNR20 U370 ( .A(B[7]), .B(A[7]), .Q(n25) );
  NOR21 U371 ( .A(A[7]), .B(B[7]), .Q(n308) );
  NOR21 U372 ( .A(B[7]), .B(A[7]), .Q(n378) );
  NOR30 U373 ( .A(n265), .B(n258), .C(n266), .Q(n262) );
  NOR20 U374 ( .A(A[30]), .B(B[30]), .Q(n59) );
  NAND22 U375 ( .A(B[13]), .B(A[13]), .Q(n301) );
  XNR20 U376 ( .A(B[24]), .B(A[24]), .Q(n143) );
  CLKIN0 U377 ( .A(B[20]), .Q(n246) );
  NAND22 U378 ( .A(B[20]), .B(A[20]), .Q(n197) );
  XNR20 U379 ( .A(B[20]), .B(A[20]), .Q(n227) );
  XNR20 U380 ( .A(B[8]), .B(A[8]), .Q(n21) );
  AOI210 U381 ( .A(B[8]), .B(A[8]), .C(n349), .Q(n341) );
  CLKIN3 U382 ( .A(n24), .Q(n17) );
  CLKIN3 U383 ( .A(n27), .Q(n30) );
  OAI212 U384 ( .A(n39), .B(n40), .C(n41), .Q(n33) );
  CLKIN3 U385 ( .A(n41), .Q(n45) );
  OAI212 U386 ( .A(n59), .B(n60), .C(n61), .Q(n58) );
  OAI222 U387 ( .A(n59), .B(n62), .C(n59), .D(n63), .Q(n57) );
  CLKIN3 U388 ( .A(n60), .Q(n71) );
  CLKIN3 U389 ( .A(n64), .Q(n67) );
  CLKIN3 U390 ( .A(n48), .Q(n81) );
  OAI222 U391 ( .A(n92), .B(n93), .C(n94), .D(n95), .Q(n72) );
  CLKIN3 U392 ( .A(n111), .Q(n110) );
  CLKIN3 U393 ( .A(n115), .Q(n114) );
  CLKIN3 U394 ( .A(n123), .Q(n122) );
  CLKIN3 U395 ( .A(n102), .Q(n119) );
  OAI212 U396 ( .A(n146), .B(n147), .C(n77), .Q(n145) );
  CLKIN3 U397 ( .A(n150), .Q(n149) );
  OAI212 U398 ( .A(n164), .B(n165), .C(n166), .Q(n163) );
  CLKIN3 U399 ( .A(n169), .Q(n167) );
  CLKIN3 U400 ( .A(n76), .Q(n144) );
  AOI212 U401 ( .A(n12), .B(n204), .C(n205), .Q(n203) );
  CLKIN3 U402 ( .A(n198), .Q(n208) );
  CLKIN3 U403 ( .A(n189), .Q(n202) );
  AOI312 U404 ( .A(n190), .B(n213), .C(n12), .D(n214), .Q(n212) );
  AOI212 U405 ( .A(n213), .B(n12), .C(n215), .Q(n219) );
  CLKIN3 U406 ( .A(n210), .Q(n213) );
  CLKIN3 U407 ( .A(n187), .Q(n230) );
  CLKIN3 U408 ( .A(n82), .Q(n249) );
  CLKIN3 U409 ( .A(n255), .Q(n235) );
  AOI312 U410 ( .A(n271), .B(n260), .C(n272), .D(n273), .Q(n270) );
  CLKIN3 U411 ( .A(n183), .Q(n267) );
  CLKIN3 U412 ( .A(n278), .Q(n258) );
  CLKIN3 U413 ( .A(n176), .Q(n292) );
  AOI312 U414 ( .A(n182), .B(n159), .C(n299), .D(n157), .Q(n265) );
  CLKIN3 U415 ( .A(n302), .Q(n160) );
  CLKIN3 U416 ( .A(n277), .Q(n266) );
  CLKIN3 U417 ( .A(n159), .Q(n318) );
  CLKIN3 U418 ( .A(n290), .Q(n178) );
  CLKIN3 U419 ( .A(n301), .Q(n328) );
  OAI212 U420 ( .A(n22), .B(n320), .C(n321), .Q(n327) );
  OAI212 U421 ( .A(n332), .B(n333), .C(n334), .Q(n321) );
  CLKIN3 U422 ( .A(n355), .Q(n332) );
  OAI2112 U423 ( .A(n39), .B(n290), .C(n311), .D(n324), .Q(n16) );
  CLKIN3 U424 ( .A(n36), .Q(n28) );
endmodule


module E_alu_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393;

  NAND23 U3 ( .A(n293), .B(n359), .Q(n39) );
  NAND42 U4 ( .A(n294), .B(n295), .C(n296), .D(n297), .Q(n359) );
  NOR23 U5 ( .A(n288), .B(n289), .Q(n287) );
  NAND42 U6 ( .A(n298), .B(n299), .C(n300), .D(n301), .Q(n282) );
  NAND23 U7 ( .A(n71), .B(n381), .Q(n298) );
  NAND34 U8 ( .A(n276), .B(n277), .C(n287), .Q(n269) );
  NAND23 U9 ( .A(n310), .B(n275), .Q(n308) );
  NOR21 U10 ( .A(A[5]), .B(n360), .Q(n364) );
  NAND23 U11 ( .A(n375), .B(n16), .Q(n301) );
  NAND34 U12 ( .A(n385), .B(n58), .C(n386), .Q(n40) );
  NAND21 U13 ( .A(n294), .B(n295), .Q(n292) );
  INV1 U14 ( .A(B[24]), .Q(n135) );
  NAND24 U15 ( .A(n112), .B(n111), .Q(n265) );
  NAND22 U16 ( .A(n266), .B(n267), .Q(n111) );
  NAND33 U17 ( .A(n298), .B(n300), .C(n301), .Q(n367) );
  NAND22 U18 ( .A(n10), .B(n11), .Q(n12) );
  NAND22 U19 ( .A(n276), .B(n277), .Q(n274) );
  INV6 U20 ( .A(B[12]), .Q(n290) );
  INV3 U21 ( .A(n220), .Q(n166) );
  NAND23 U22 ( .A(B[1]), .B(n378), .Q(n100) );
  INV3 U23 ( .A(B[6]), .Q(n55) );
  NAND24 U24 ( .A(n108), .B(n109), .Q(n88) );
  NOR21 U25 ( .A(n358), .B(n342), .Q(n357) );
  NOR23 U26 ( .A(n243), .B(n244), .Q(n242) );
  CLKIN3 U27 ( .A(n242), .Q(n3) );
  NAND22 U28 ( .A(B[10]), .B(n392), .Q(n340) );
  NAND22 U29 ( .A(n8), .B(n9), .Q(DIFF[27]) );
  NAND22 U30 ( .A(n6), .B(n7), .Q(n9) );
  NAND22 U31 ( .A(A[9]), .B(n339), .Q(n34) );
  NAND22 U32 ( .A(A[10]), .B(n391), .Q(n338) );
  NAND34 U33 ( .A(n221), .B(n230), .C(n231), .Q(n211) );
  INV6 U34 ( .A(B[23]), .Q(n169) );
  XOR22 U35 ( .A(n195), .B(n196), .Q(DIFF[22]) );
  CLKIN6 U36 ( .A(n315), .Q(n311) );
  INV6 U37 ( .A(B[9]), .Q(n339) );
  AOI2112 U38 ( .A(n356), .B(n38), .C(n42), .D(n357), .Q(n32) );
  INV6 U39 ( .A(n324), .Q(n38) );
  OAI2111 U40 ( .A(n172), .B(n173), .C(n174), .D(n175), .Q(n171) );
  INV3 U41 ( .A(A[10]), .Q(n392) );
  INV3 U42 ( .A(n273), .Q(n10) );
  INV3 U43 ( .A(n274), .Q(n11) );
  NOR23 U44 ( .A(n278), .B(n279), .Q(n273) );
  INV3 U45 ( .A(A[0]), .Q(n240) );
  NOR22 U46 ( .A(n376), .B(n377), .Q(n375) );
  INV3 U47 ( .A(n15), .Q(n16) );
  NOR23 U48 ( .A(n345), .B(n343), .Q(n13) );
  NOR21 U49 ( .A(A[11]), .B(n334), .Q(n343) );
  INV3 U50 ( .A(B[17]), .Q(n228) );
  NOR22 U51 ( .A(n285), .B(n321), .Q(n26) );
  NAND22 U52 ( .A(n59), .B(n60), .Q(n54) );
  NAND22 U53 ( .A(A[14]), .B(n316), .Q(n275) );
  AOI211 U54 ( .A(B[23]), .B(n177), .C(n178), .Q(n170) );
  INV3 U55 ( .A(n32), .Q(n353) );
  INV3 U56 ( .A(n136), .Q(n6) );
  AOI211 U57 ( .A(n189), .B(n179), .C(n190), .Q(n188) );
  NOR21 U58 ( .A(A[17]), .B(n228), .Q(n227) );
  NAND22 U59 ( .A(n296), .B(n297), .Q(n291) );
  NOR23 U60 ( .A(n269), .B(n285), .Q(n284) );
  NAND22 U61 ( .A(n70), .B(n100), .Q(n371) );
  NOR21 U62 ( .A(A[9]), .B(n339), .Q(n346) );
  INV6 U63 ( .A(B[4]), .Q(n61) );
  NAND23 U64 ( .A(n12), .B(n275), .Q(n271) );
  NAND22 U65 ( .A(n166), .B(n218), .Q(n212) );
  NAND22 U66 ( .A(n17), .B(n18), .Q(n19) );
  INV3 U67 ( .A(n323), .Q(n279) );
  INV3 U68 ( .A(n137), .Q(n7) );
  INV3 U69 ( .A(n212), .Q(n200) );
  INV3 U70 ( .A(n26), .Q(n325) );
  NAND22 U71 ( .A(B[22]), .B(n206), .Q(n179) );
  INV3 U72 ( .A(B[22]), .Q(n205) );
  AOI211 U73 ( .A(n350), .B(n340), .C(n351), .Q(n349) );
  AOI211 U74 ( .A(n155), .B(n156), .C(n125), .Q(n154) );
  AOI311 U75 ( .A(n74), .B(n75), .C(n76), .D(n77), .Q(n73) );
  NOR21 U76 ( .A(A[6]), .B(n55), .Q(n365) );
  AOI211 U77 ( .A(n209), .B(n210), .C(n199), .Q(n208) );
  OAI211 U78 ( .A(n82), .B(n211), .C(n212), .Q(n209) );
  NAND21 U79 ( .A(n234), .B(A[16]), .Q(n20) );
  INV3 U80 ( .A(B[27]), .Q(n124) );
  INV3 U81 ( .A(n374), .Q(n393) );
  INV3 U82 ( .A(n39), .Q(n342) );
  INV3 U83 ( .A(n70), .Q(n379) );
  NAND23 U84 ( .A(B[2]), .B(n383), .Q(n70) );
  NAND22 U85 ( .A(n145), .B(n146), .Q(n144) );
  OAI2111 U86 ( .A(n278), .B(n311), .C(n276), .D(n277), .Q(n310) );
  NOR23 U87 ( .A(n361), .B(n387), .Q(n386) );
  NAND22 U88 ( .A(n156), .B(n126), .Q(n147) );
  NAND21 U89 ( .A(A[24]), .B(n135), .Q(n187) );
  INV2 U90 ( .A(n264), .Q(n1) );
  NAND22 U91 ( .A(n241), .B(n242), .Q(n4) );
  NAND24 U92 ( .A(n2), .B(n3), .Q(n5) );
  NAND24 U93 ( .A(n4), .B(n5), .Q(DIFF[19]) );
  INV3 U94 ( .A(n241), .Q(n2) );
  NAND22 U95 ( .A(n136), .B(n137), .Q(n8) );
  NOR24 U96 ( .A(n14), .B(n24), .Q(n286) );
  INV6 U97 ( .A(n13), .Q(n14) );
  INV12 U98 ( .A(n23), .Q(n24) );
  NOR24 U99 ( .A(A[8]), .B(n43), .Q(n345) );
  AOI211 U100 ( .A(n286), .B(n331), .C(n332), .Q(n330) );
  NAND22 U101 ( .A(n70), .B(n100), .Q(n15) );
  NAND22 U102 ( .A(n19), .B(n342), .Q(n331) );
  INV2 U103 ( .A(n64), .Q(n17) );
  INV0 U104 ( .A(n40), .Q(n18) );
  NAND22 U105 ( .A(n20), .B(n229), .Q(n222) );
  NAND22 U106 ( .A(n131), .B(n126), .Q(n21) );
  NAND22 U107 ( .A(n132), .B(n22), .Q(n130) );
  INV3 U108 ( .A(n21), .Q(n22) );
  CLKIN6 U109 ( .A(n286), .Q(n285) );
  OAI210 U110 ( .A(n82), .B(n148), .C(n157), .Q(n155) );
  NOR20 U111 ( .A(A[16]), .B(n234), .Q(n306) );
  NOR20 U112 ( .A(A[16]), .B(n234), .Q(n259) );
  NAND20 U113 ( .A(A[16]), .B(n234), .Q(n307) );
  INV2 U114 ( .A(A[13]), .Q(n327) );
  INV0 U115 ( .A(n59), .Q(n66) );
  NAND23 U116 ( .A(A[4]), .B(n61), .Q(n59) );
  NOR23 U117 ( .A(n183), .B(n184), .Q(n182) );
  NOR22 U118 ( .A(A[20]), .B(n185), .Q(n183) );
  NAND24 U119 ( .A(n380), .B(n381), .Q(n300) );
  AOI312 U120 ( .A(n111), .B(n112), .C(n1), .D(n83), .Q(n110) );
  NAND23 U121 ( .A(n113), .B(n114), .Q(n83) );
  NOR22 U122 ( .A(A[15]), .B(n272), .Q(n289) );
  CLKIN4 U123 ( .A(n110), .Q(n109) );
  NOR20 U124 ( .A(A[24]), .B(n135), .Q(n152) );
  NOR20 U125 ( .A(A[24]), .B(n135), .Q(n133) );
  NAND24 U126 ( .A(n248), .B(n146), .Q(n246) );
  NAND33 U127 ( .A(n53), .B(n48), .C(n59), .Q(n297) );
  NOR21 U128 ( .A(n268), .B(n269), .Q(n266) );
  INV2 U129 ( .A(A[3]), .Q(n370) );
  OAI2112 U130 ( .A(n291), .B(n292), .C(n293), .D(n40), .Q(n283) );
  NOR23 U131 ( .A(A[3]), .B(n373), .Q(n377) );
  INV2 U132 ( .A(A[5]), .Q(n388) );
  NAND22 U133 ( .A(A[1]), .B(n382), .Q(n97) );
  INV2 U134 ( .A(A[1]), .Q(n378) );
  NAND24 U135 ( .A(A[17]), .B(n228), .Q(n229) );
  NAND21 U136 ( .A(A[12]), .B(n290), .Q(n323) );
  NOR23 U137 ( .A(n341), .B(n42), .Q(n335) );
  NAND21 U138 ( .A(A[20]), .B(n185), .Q(n173) );
  NOR24 U139 ( .A(n344), .B(n346), .Q(n23) );
  XOR22 U140 ( .A(n312), .B(n313), .Q(DIFF[14]) );
  NAND20 U141 ( .A(n340), .B(n338), .Q(n354) );
  AOI211 U142 ( .A(n114), .B(n146), .C(n129), .Q(n162) );
  INV2 U143 ( .A(n340), .Q(n344) );
  AOI212 U144 ( .A(n104), .B(n88), .C(n92), .Q(n102) );
  NOR22 U145 ( .A(A[7]), .B(n362), .Q(n361) );
  AOI312 U146 ( .A(n245), .B(n229), .C(n246), .D(n247), .Q(n244) );
  NAND20 U147 ( .A(A[13]), .B(n326), .Q(n25) );
  NAND22 U148 ( .A(A[13]), .B(n326), .Q(n314) );
  INV2 U149 ( .A(B[13]), .Q(n326) );
  NOR24 U150 ( .A(n367), .B(n368), .Q(n324) );
  NOR21 U151 ( .A(A[0]), .B(n239), .Q(n238) );
  NOR23 U152 ( .A(A[0]), .B(n239), .Q(n376) );
  NOR21 U153 ( .A(A[12]), .B(n290), .Q(n288) );
  NOR20 U154 ( .A(A[12]), .B(n290), .Q(n321) );
  NAND22 U155 ( .A(A[5]), .B(n360), .Q(n53) );
  INV6 U156 ( .A(B[15]), .Q(n272) );
  OAI2112 U157 ( .A(n281), .B(n282), .C(n283), .D(n284), .Q(n27) );
  NAND42 U158 ( .A(n48), .B(n59), .C(n53), .D(n304), .Q(n281) );
  NAND22 U159 ( .A(A[6]), .B(n55), .Q(n48) );
  XOR22 U160 ( .A(n102), .B(n103), .Q(DIFF[29]) );
  INV3 U161 ( .A(n53), .Q(n57) );
  INV3 U162 ( .A(A[21]), .Q(n214) );
  OAI222 U163 ( .A(n270), .B(n271), .C(A[15]), .D(n272), .Q(n112) );
  INV6 U164 ( .A(n27), .Q(n264) );
  CLKIN0 U165 ( .A(A[17]), .Q(n260) );
  NOR21 U166 ( .A(A[23]), .B(n169), .Q(n184) );
  CLKIN1 U167 ( .A(n147), .Q(n149) );
  INV0 U168 ( .A(n69), .Q(n96) );
  CLKIN0 U169 ( .A(n152), .Q(n156) );
  CLKIN0 U170 ( .A(n268), .Q(n333) );
  CLKIN3 U171 ( .A(n101), .Q(n71) );
  INV0 U172 ( .A(A[14]), .Q(n317) );
  CLKIN0 U173 ( .A(B[26]), .Q(n142) );
  INV2 U174 ( .A(B[7]), .Q(n362) );
  NAND22 U175 ( .A(B[21]), .B(n214), .Q(n176) );
  INV0 U176 ( .A(B[25]), .Q(n158) );
  INV2 U177 ( .A(n119), .Q(n118) );
  INV12 U178 ( .A(n82), .Q(n146) );
  INV0 U179 ( .A(n204), .Q(n210) );
  NAND22 U180 ( .A(n33), .B(n353), .Q(n352) );
  CLKIN0 U181 ( .A(n122), .Q(n139) );
  NOR21 U182 ( .A(n302), .B(n303), .Q(n299) );
  OAI2112 U183 ( .A(n335), .B(n336), .C(n337), .D(n338), .Q(n267) );
  AOI221 U184 ( .A(A[23]), .B(n169), .C(n170), .D(n171), .Q(n163) );
  NAND24 U185 ( .A(n163), .B(n164), .Q(n129) );
  AOI211 U186 ( .A(n46), .B(n294), .C(n47), .Q(n45) );
  INV3 U187 ( .A(B[14]), .Q(n316) );
  CLKIN0 U188 ( .A(B[30]), .Q(n86) );
  CLKIN2 U189 ( .A(n92), .Q(n90) );
  INV0 U190 ( .A(A[29]), .Q(n91) );
  AOI212 U191 ( .A(n194), .B(n146), .C(n197), .Q(n196) );
  NOR20 U192 ( .A(n139), .B(n120), .Q(n140) );
  NOR20 U193 ( .A(n147), .B(n148), .Q(n145) );
  INV2 U194 ( .A(n369), .Q(n368) );
  NOR22 U195 ( .A(n305), .B(n302), .Q(n369) );
  INV1 U196 ( .A(n81), .Q(n75) );
  AOI2112 U197 ( .A(n26), .B(n39), .C(n319), .D(n320), .Q(n315) );
  NAND20 U198 ( .A(n245), .B(n229), .Q(n251) );
  INV0 U199 ( .A(n93), .Q(n104) );
  INV1 U200 ( .A(n54), .Q(n52) );
  NAND20 U201 ( .A(n276), .B(n275), .Q(n312) );
  AOI212 U202 ( .A(n311), .B(n277), .C(n278), .Q(n313) );
  INV6 U203 ( .A(n211), .Q(n180) );
  NOR22 U204 ( .A(n379), .B(n97), .Q(n380) );
  AOI312 U205 ( .A(n221), .B(n222), .C(n223), .D(n224), .Q(n220) );
  NAND20 U206 ( .A(n277), .B(n25), .Q(n318) );
  AOI210 U207 ( .A(n69), .B(n70), .C(n71), .Q(n68) );
  XOR20 U208 ( .A(n31), .B(n32), .Q(DIFF[9]) );
  NAND20 U209 ( .A(n252), .B(n230), .Q(n245) );
  INV0 U210 ( .A(n167), .Q(n218) );
  NAND20 U211 ( .A(n230), .B(n229), .Q(n257) );
  NAND20 U212 ( .A(n179), .B(n175), .Q(n195) );
  NAND20 U213 ( .A(n176), .B(n174), .Q(n207) );
  NAND20 U214 ( .A(n221), .B(n226), .Q(n249) );
  NAND20 U215 ( .A(n70), .B(n101), .Q(n95) );
  NAND20 U216 ( .A(n125), .B(n126), .Q(n151) );
  NAND20 U217 ( .A(n254), .B(n230), .Q(n253) );
  INV0 U218 ( .A(n99), .Q(n237) );
  NOR22 U219 ( .A(B[0]), .B(n240), .Q(n374) );
  NOR22 U220 ( .A(n232), .B(n233), .Q(n231) );
  INV0 U221 ( .A(n175), .Q(n190) );
  NOR23 U222 ( .A(n371), .B(n372), .Q(n305) );
  AOI210 U223 ( .A(B[24]), .B(n186), .C(n125), .Q(n160) );
  XNR20 U224 ( .A(B[30]), .B(A[30]), .Q(n28) );
  INV0 U225 ( .A(A[6]), .Q(n363) );
  NOR20 U226 ( .A(B[28]), .B(n105), .Q(n92) );
  INV0 U227 ( .A(A[28]), .Q(n105) );
  NOR20 U228 ( .A(A[20]), .B(n185), .Q(n204) );
  INV0 U229 ( .A(B[29]), .Q(n94) );
  INV0 U230 ( .A(B[28]), .Q(n106) );
  NOR20 U231 ( .A(n40), .B(n358), .Q(n356) );
  AOI210 U232 ( .A(B[12]), .B(n347), .C(n279), .Q(n328) );
  NAND21 U233 ( .A(B[26]), .B(n141), .Q(n131) );
  INV0 U234 ( .A(A[26]), .Q(n141) );
  INV0 U235 ( .A(A[9]), .Q(n390) );
  AOI210 U236 ( .A(n18), .B(n38), .C(n39), .Q(n37) );
  NOR20 U237 ( .A(n41), .B(n42), .Q(n35) );
  XOR20 U238 ( .A(n107), .B(n88), .Q(DIFF[28]) );
  NOR20 U239 ( .A(A[27]), .B(n124), .Q(n119) );
  INV0 U240 ( .A(n338), .Q(n351) );
  INV0 U241 ( .A(A[15]), .Q(n280) );
  NOR20 U242 ( .A(B[15]), .B(n280), .Q(n270) );
  INV0 U243 ( .A(A[23]), .Q(n177) );
  NAND20 U244 ( .A(A[30]), .B(n86), .Q(n79) );
  INV0 U245 ( .A(A[24]), .Q(n186) );
  INV0 U246 ( .A(A[12]), .Q(n347) );
  INV0 U247 ( .A(A[20]), .Q(n235) );
  NAND22 U248 ( .A(n194), .B(n146), .Q(n192) );
  NAND22 U249 ( .A(n193), .B(n191), .Q(n197) );
  NAND22 U250 ( .A(n201), .B(n180), .Q(n202) );
  INV3 U251 ( .A(n46), .Q(n50) );
  INV3 U252 ( .A(n148), .Q(n114) );
  NOR31 U253 ( .A(n324), .B(n325), .C(n40), .Q(n319) );
  NAND22 U254 ( .A(n78), .B(n79), .Q(n77) );
  AOI211 U255 ( .A(n254), .B(n146), .C(n252), .Q(n258) );
  AOI211 U256 ( .A(n248), .B(n146), .C(n251), .Q(n250) );
  XOR21 U257 ( .A(n354), .B(n355), .Q(DIFF[10]) );
  AOI211 U258 ( .A(n33), .B(n353), .C(n341), .Q(n355) );
  NOR21 U259 ( .A(n167), .B(n168), .Q(n165) );
  NOR21 U260 ( .A(n93), .B(n89), .Q(n74) );
  NOR22 U261 ( .A(n115), .B(n116), .Q(n108) );
  XOR21 U262 ( .A(n153), .B(n154), .Q(DIFF[25]) );
  XOR21 U263 ( .A(n49), .B(n50), .Q(DIFF[6]) );
  AOI211 U264 ( .A(n125), .B(n126), .C(n127), .Q(n121) );
  NAND24 U265 ( .A(n180), .B(n181), .Q(n148) );
  NAND22 U266 ( .A(n267), .B(n333), .Q(n322) );
  NAND22 U267 ( .A(n33), .B(n34), .Q(n31) );
  NAND22 U268 ( .A(n210), .B(n176), .Q(n203) );
  NAND22 U269 ( .A(n97), .B(n98), .Q(n69) );
  NAND22 U270 ( .A(n99), .B(n100), .Q(n98) );
  NAND22 U271 ( .A(n113), .B(n129), .Q(n85) );
  NAND22 U272 ( .A(n143), .B(n144), .Q(n138) );
  AOI211 U273 ( .A(n149), .B(n129), .C(n150), .Q(n143) );
  NAND22 U274 ( .A(n80), .B(n75), .Q(n78) );
  INV3 U275 ( .A(n227), .Q(n223) );
  NAND22 U276 ( .A(n225), .B(n226), .Q(n224) );
  INV3 U277 ( .A(n293), .Q(n303) );
  INV3 U278 ( .A(n305), .Q(n304) );
  NOR21 U279 ( .A(n57), .B(n51), .Q(n56) );
  NAND22 U280 ( .A(n294), .B(n48), .Q(n49) );
  NAND22 U281 ( .A(n100), .B(n97), .Q(n236) );
  NOR21 U282 ( .A(A[4]), .B(n61), .Q(n389) );
  NAND22 U283 ( .A(B[25]), .B(n159), .Q(n126) );
  NAND22 U284 ( .A(B[18]), .B(n256), .Q(n221) );
  INV3 U285 ( .A(B[1]), .Q(n382) );
  NAND22 U286 ( .A(B[17]), .B(n260), .Q(n230) );
  NAND22 U287 ( .A(A[21]), .B(n213), .Q(n174) );
  INV3 U288 ( .A(B[21]), .Q(n213) );
  NAND22 U289 ( .A(A[18]), .B(n255), .Q(n226) );
  INV3 U290 ( .A(B[18]), .Q(n255) );
  NOR21 U291 ( .A(A[6]), .B(n55), .Q(n387) );
  NAND22 U292 ( .A(B[13]), .B(n327), .Q(n277) );
  INV3 U293 ( .A(A[2]), .Q(n383) );
  NAND22 U294 ( .A(n192), .B(n30), .Q(n189) );
  XOR21 U295 ( .A(n236), .B(n237), .Q(DIFF[1]) );
  XNR21 U296 ( .A(n67), .B(n68), .Q(DIFF[3]) );
  IMUX21 U297 ( .A(n62), .B(n63), .S(n64), .Q(DIFF[4]) );
  XOR21 U298 ( .A(n54), .B(n56), .Q(DIFF[5]) );
  XOR21 U299 ( .A(n95), .B(n96), .Q(DIFF[2]) );
  NAND22 U300 ( .A(B[5]), .B(n388), .Q(n58) );
  XNR21 U301 ( .A(n87), .B(n28), .Q(DIFF[30]) );
  IMUX21 U302 ( .A(n261), .B(n262), .S(n263), .Q(DIFF[16]) );
  XOR21 U303 ( .A(n257), .B(n258), .Q(DIFF[17]) );
  XOR21 U304 ( .A(n249), .B(n250), .Q(DIFF[18]) );
  XOR21 U305 ( .A(n207), .B(n208), .Q(DIFF[21]) );
  XOR21 U306 ( .A(n72), .B(n73), .Q(DIFF[31]) );
  NOR21 U307 ( .A(B[3]), .B(n370), .Q(n302) );
  NOR21 U308 ( .A(n65), .B(n66), .Q(n62) );
  IMUX21 U309 ( .A(n215), .B(n216), .S(n217), .Q(DIFF[20]) );
  AOI211 U310 ( .A(n180), .B(n146), .C(n200), .Q(n217) );
  IMUX21 U311 ( .A(n160), .B(n161), .S(n162), .Q(DIFF[24]) );
  IMUX21 U312 ( .A(n35), .B(n36), .S(n37), .Q(DIFF[8]) );
  NAND22 U313 ( .A(A[2]), .B(n384), .Q(n101) );
  INV3 U314 ( .A(B[2]), .Q(n384) );
  NOR21 U315 ( .A(n133), .B(n134), .Q(n132) );
  NAND22 U316 ( .A(n393), .B(n238), .Q(n99) );
  XNR21 U317 ( .A(n44), .B(n45), .Q(DIFF[7]) );
  XOR21 U318 ( .A(n308), .B(n309), .Q(DIFF[15]) );
  NAND22 U319 ( .A(n165), .B(n166), .Q(n164) );
  INV3 U320 ( .A(B[8]), .Q(n43) );
  IMUX21 U321 ( .A(n328), .B(n329), .S(n330), .Q(DIFF[12]) );
  INV3 U322 ( .A(n361), .Q(n296) );
  INV3 U323 ( .A(n377), .Q(n381) );
  INV3 U324 ( .A(B[3]), .Q(n373) );
  INV3 U325 ( .A(B[5]), .Q(n360) );
  INV3 U326 ( .A(n365), .Q(n294) );
  XNR21 U327 ( .A(n348), .B(n349), .Q(DIFF[11]) );
  INV3 U328 ( .A(n259), .Q(n254) );
  INV6 U329 ( .A(B[20]), .Q(n185) );
  INV3 U330 ( .A(B[0]), .Q(n239) );
  INV3 U331 ( .A(B[16]), .Q(n234) );
  INV3 U332 ( .A(B[11]), .Q(n334) );
  INV3 U333 ( .A(B[19]), .Q(n219) );
  NAND22 U334 ( .A(B[9]), .B(n390), .Q(n33) );
  NOR21 U335 ( .A(n306), .B(n252), .Q(n261) );
  NAND22 U336 ( .A(A[22]), .B(n205), .Q(n175) );
  INV3 U337 ( .A(A[22]), .Q(n206) );
  NAND22 U338 ( .A(A[19]), .B(n219), .Q(n225) );
  XNR21 U339 ( .A(B[28]), .B(A[28]), .Q(n107) );
  NOR21 U340 ( .A(A[28]), .B(n106), .Q(n93) );
  OAI210 U341 ( .A(A[0]), .B(n239), .C(n393), .Q(DIFF[0]) );
  INV3 U342 ( .A(A[18]), .Q(n256) );
  XNR21 U343 ( .A(B[27]), .B(A[27]), .Q(n136) );
  NOR21 U344 ( .A(A[27]), .B(n124), .Q(n134) );
  NAND21 U345 ( .A(A[27]), .B(n124), .Q(n123) );
  INV3 U346 ( .A(n389), .Q(n385) );
  XOR20 U347 ( .A(B[16]), .B(A[16]), .Q(n262) );
  NOR21 U348 ( .A(A[16]), .B(n234), .Q(n232) );
  NAND22 U349 ( .A(n117), .B(n118), .Q(n84) );
  OAI2111 U350 ( .A(n120), .B(n121), .C(n122), .D(n123), .Q(n117) );
  INV3 U351 ( .A(n128), .Q(n127) );
  NAND22 U352 ( .A(n126), .B(n128), .Q(n153) );
  NAND22 U353 ( .A(n151), .B(n128), .Q(n150) );
  NAND22 U354 ( .A(A[25]), .B(n158), .Q(n128) );
  XOR21 U355 ( .A(B[29]), .B(A[29]), .Q(n103) );
  NOR21 U356 ( .A(A[29]), .B(n94), .Q(n89) );
  INV1 U357 ( .A(B[10]), .Q(n391) );
  NAND22 U358 ( .A(A[26]), .B(n142), .Q(n122) );
  NOR21 U359 ( .A(A[11]), .B(n334), .Q(n268) );
  NAND20 U360 ( .A(A[11]), .B(n334), .Q(n337) );
  XNR20 U361 ( .A(B[11]), .B(A[11]), .Q(n348) );
  OAI210 U362 ( .A(A[9]), .B(n339), .C(n340), .Q(n336) );
  XOR21 U363 ( .A(n138), .B(n140), .Q(DIFF[26]) );
  XNR20 U364 ( .A(B[19]), .B(A[19]), .Q(n241) );
  NOR21 U365 ( .A(A[19]), .B(n219), .Q(n167) );
  NOR21 U366 ( .A(A[19]), .B(n219), .Q(n233) );
  OAI211 U367 ( .A(B[6]), .B(n363), .C(n364), .Q(n295) );
  XOR20 U368 ( .A(B[12]), .B(A[12]), .Q(n329) );
  NAND22 U369 ( .A(n193), .B(n191), .Q(n29) );
  INV3 U370 ( .A(n29), .Q(n30) );
  OAI210 U371 ( .A(n198), .B(n199), .C(n176), .Q(n191) );
  NAND22 U372 ( .A(n200), .B(n201), .Q(n193) );
  XNR20 U373 ( .A(B[3]), .B(A[3]), .Q(n67) );
  XNR20 U374 ( .A(B[15]), .B(A[15]), .Q(n309) );
  OAI212 U375 ( .A(A[4]), .B(n61), .C(n38), .Q(n60) );
  INV0 U376 ( .A(A[25]), .Q(n159) );
  INV2 U377 ( .A(n226), .Q(n243) );
  NOR20 U378 ( .A(A[4]), .B(n61), .Q(n65) );
  XOR20 U379 ( .A(B[4]), .B(A[4]), .Q(n63) );
  XOR20 U380 ( .A(B[31]), .B(A[31]), .Q(n72) );
  NAND22 U381 ( .A(B[14]), .B(n317), .Q(n276) );
  INV2 U382 ( .A(n146), .Q(n263) );
  NAND22 U383 ( .A(n352), .B(n34), .Q(n350) );
  NOR20 U384 ( .A(A[8]), .B(n43), .Q(n41) );
  NOR20 U385 ( .A(A[8]), .B(n43), .Q(n358) );
  NAND22 U386 ( .A(A[8]), .B(n43), .Q(n366) );
  CLKIN3 U387 ( .A(n129), .Q(n157) );
  XNR20 U388 ( .A(B[7]), .B(A[7]), .Q(n44) );
  NAND22 U389 ( .A(A[7]), .B(n362), .Q(n293) );
  NOR20 U390 ( .A(A[30]), .B(n86), .Q(n81) );
  INV3 U391 ( .A(n168), .Q(n181) );
  XOR20 U392 ( .A(B[24]), .B(A[24]), .Q(n161) );
  AOI210 U393 ( .A(B[20]), .B(n235), .C(n199), .Q(n215) );
  XOR20 U394 ( .A(B[20]), .B(A[20]), .Q(n216) );
  XOR20 U395 ( .A(B[8]), .B(A[8]), .Q(n36) );
  XOR20 U396 ( .A(n318), .B(n315), .Q(DIFF[13]) );
  OAI2111 U397 ( .A(n82), .B(n83), .C(n84), .D(n85), .Q(n76) );
  CLKIN3 U398 ( .A(n48), .Q(n47) );
  OAI212 U399 ( .A(n51), .B(n52), .C(n53), .Q(n46) );
  CLKIN3 U400 ( .A(n58), .Q(n51) );
  AOI212 U401 ( .A(n74), .B(n88), .C(n80), .Q(n87) );
  OAI222 U402 ( .A(n89), .B(n90), .C(B[29]), .D(n91), .Q(n80) );
  CLKIN3 U403 ( .A(n84), .Q(n116) );
  CLKIN3 U404 ( .A(n85), .Q(n115) );
  CLKIN3 U405 ( .A(n130), .Q(n113) );
  AOI212 U406 ( .A(n138), .B(n131), .C(n139), .Q(n137) );
  CLKIN3 U407 ( .A(n131), .Q(n120) );
  CLKIN3 U408 ( .A(n176), .Q(n172) );
  CLKIN3 U409 ( .A(n179), .Q(n178) );
  NAND33 U410 ( .A(n179), .B(n176), .C(n182), .Q(n168) );
  CLKIN3 U411 ( .A(n187), .Q(n125) );
  XOR31 U412 ( .A(B[23]), .B(A[23]), .C(n188), .Q(DIFF[23]) );
  CLKIN3 U413 ( .A(n174), .Q(n198) );
  CLKIN3 U414 ( .A(n202), .Q(n194) );
  CLKIN3 U415 ( .A(n203), .Q(n201) );
  CLKIN3 U416 ( .A(n173), .Q(n199) );
  CLKIN3 U417 ( .A(n221), .Q(n247) );
  CLKIN3 U418 ( .A(n253), .Q(n248) );
  NOR24 U419 ( .A(n264), .B(n265), .Q(n82) );
  CLKIN3 U420 ( .A(n307), .Q(n252) );
  CLKIN3 U421 ( .A(n314), .Q(n278) );
  OAI212 U422 ( .A(n321), .B(n322), .C(n323), .Q(n320) );
  CLKIN3 U423 ( .A(n322), .Q(n332) );
  CLKIN3 U424 ( .A(n38), .Q(n64) );
  CLKIN3 U425 ( .A(n34), .Q(n341) );
  CLKIN3 U426 ( .A(n366), .Q(n42) );
  OAI212 U427 ( .A(A[3]), .B(n373), .C(n374), .Q(n372) );
endmodule


module E_alu_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265;

  NAND21 U1 ( .A(n209), .B(n136), .Q(n208) );
  NOR20 U2 ( .A(B[13]), .B(n148), .Q(n227) );
  NOR21 U3 ( .A(n158), .B(n159), .Q(n12) );
  INV1 U4 ( .A(A[23]), .Q(n262) );
  NAND22 U5 ( .A(n147), .B(n149), .Q(n225) );
  INV3 U6 ( .A(n224), .Q(n102) );
  INV0 U7 ( .A(A[3]), .Q(n78) );
  NOR20 U8 ( .A(B[2]), .B(n79), .Q(n76) );
  NAND30 U9 ( .A(n37), .B(n100), .C(n8), .Q(n34) );
  NOR31 U10 ( .A(n101), .B(n102), .C(n57), .Q(n100) );
  NOR21 U11 ( .A(n91), .B(n192), .Q(n218) );
  NAND42 U12 ( .A(n221), .B(n89), .C(n86), .D(n222), .Q(n215) );
  NAND22 U13 ( .A(n86), .B(n89), .Q(n1) );
  NAND31 U14 ( .A(n218), .B(n217), .C(n2), .Q(n216) );
  INV3 U15 ( .A(n1), .Q(n2) );
  NOR22 U16 ( .A(n111), .B(n110), .Q(n3) );
  NOR21 U17 ( .A(n4), .B(n109), .Q(n108) );
  INV3 U18 ( .A(n3), .Q(n4) );
  INV6 U19 ( .A(n89), .Q(n110) );
  NAND31 U20 ( .A(n48), .B(n112), .C(n50), .Q(n111) );
  NAND30 U21 ( .A(n10), .B(n87), .C(B[8]), .Q(n5) );
  NAND22 U22 ( .A(n86), .B(n6), .Q(n174) );
  INV3 U23 ( .A(n5), .Q(n6) );
  NOR20 U24 ( .A(A[16]), .B(n120), .Q(n214) );
  OAI2112 U25 ( .A(n175), .B(n199), .C(n200), .D(n201), .Q(n198) );
  AOI311 U26 ( .A(n36), .B(n37), .C(n38), .D(n25), .Q(n35) );
  NOR20 U27 ( .A(A[24]), .B(n205), .Q(n204) );
  OAI211 U28 ( .A(A[24]), .B(n205), .C(A[22]), .Q(n259) );
  AOI311 U29 ( .A(n178), .B(n179), .C(n37), .D(n180), .Q(n177) );
  NAND21 U30 ( .A(n50), .B(n48), .Q(n104) );
  NAND22 U31 ( .A(A[17]), .B(n153), .Q(n50) );
  NAND20 U32 ( .A(n147), .B(n148), .Q(n146) );
  NAND22 U33 ( .A(A[14]), .B(n230), .Q(n147) );
  NAND21 U34 ( .A(n108), .B(n37), .Q(n33) );
  NAND21 U35 ( .A(A[10]), .B(n191), .Q(n54) );
  NAND22 U36 ( .A(A[15]), .B(n229), .Q(n149) );
  NOR20 U37 ( .A(A[1]), .B(n82), .Q(n81) );
  INV0 U38 ( .A(A[1]), .Q(n74) );
  INV0 U39 ( .A(B[22]), .Q(n211) );
  CLKIN0 U40 ( .A(B[10]), .Q(n191) );
  OAI221 U41 ( .A(B[27]), .B(n241), .C(B[26]), .D(n242), .Q(n236) );
  INV1 U42 ( .A(A[26]), .Q(n242) );
  NAND21 U43 ( .A(n89), .B(n99), .Q(n7) );
  NOR31 U44 ( .A(n104), .B(n105), .C(n106), .Q(n99) );
  CLKIN0 U45 ( .A(B[16]), .Q(n232) );
  NOR42 U46 ( .A(n234), .B(n235), .C(n236), .D(n237), .Q(n233) );
  NAND22 U47 ( .A(n132), .B(n243), .Q(n234) );
  NAND21 U48 ( .A(n113), .B(n37), .Q(n32) );
  INV12 U49 ( .A(n175), .Q(n37) );
  NAND30 U50 ( .A(n131), .B(n132), .C(n133), .Q(n130) );
  NAND22 U51 ( .A(A[25]), .B(n157), .Q(n131) );
  INV1 U52 ( .A(A[0]), .Q(n75) );
  NAND21 U53 ( .A(B[23]), .B(n262), .Q(n261) );
  NAND42 U54 ( .A(n32), .B(n34), .C(n33), .D(n35), .Q(n31) );
  INV4 U55 ( .A(n233), .Q(n175) );
  NOR22 U56 ( .A(n30), .B(n31), .Q(n13) );
  INV1 U57 ( .A(A[27]), .Q(n241) );
  CLKIN3 U58 ( .A(n49), .Q(n105) );
  NAND21 U59 ( .A(n87), .B(n9), .Q(n101) );
  INV2 U60 ( .A(B[21]), .Q(n138) );
  INV3 U61 ( .A(n7), .Q(n8) );
  NAND22 U62 ( .A(A[21]), .B(n138), .Q(n243) );
  CLKIN3 U63 ( .A(n129), .Q(n136) );
  NAND42 U64 ( .A(n121), .B(n122), .C(n123), .D(n124), .Q(n30) );
  INV3 U65 ( .A(B[6]), .Q(n58) );
  NOR21 U66 ( .A(n119), .B(n120), .Q(n170) );
  NOR21 U67 ( .A(n90), .B(n91), .Q(n88) );
  INV6 U68 ( .A(n257), .Q(n89) );
  INV2 U69 ( .A(n260), .Q(n258) );
  INV3 U70 ( .A(B[25]), .Q(n157) );
  CLKIN0 U71 ( .A(A[13]), .Q(n148) );
  NAND22 U72 ( .A(B[6]), .B(n96), .Q(n67) );
  CLKIN0 U73 ( .A(A[6]), .Q(n96) );
  INV3 U74 ( .A(B[29]), .Q(n29) );
  BUF6 U75 ( .A(n103), .Q(n10) );
  NOR20 U76 ( .A(n120), .B(n219), .Q(n217) );
  NAND20 U77 ( .A(n48), .B(n220), .Q(n219) );
  NAND40 U78 ( .A(n132), .B(n10), .C(n135), .D(n136), .Q(n127) );
  NOR20 U79 ( .A(n120), .B(n231), .Q(n221) );
  NOR20 U80 ( .A(n91), .B(n223), .Q(n222) );
  NAND20 U81 ( .A(n48), .B(n228), .Q(n231) );
  NOR20 U82 ( .A(n129), .B(n181), .Q(n180) );
  NOR20 U83 ( .A(n110), .B(n185), .Q(n178) );
  OAI310 U84 ( .A(n245), .B(n110), .C(n246), .D(n247), .Q(n195) );
  NAND20 U85 ( .A(n10), .B(n140), .Q(n139) );
  NOR20 U86 ( .A(n102), .B(n91), .Q(n167) );
  NOR20 U87 ( .A(n110), .B(n169), .Q(n168) );
  INV2 U88 ( .A(n206), .Q(n200) );
  INV2 U89 ( .A(n254), .Q(n253) );
  NAND40 U90 ( .A(n50), .B(n48), .C(n188), .D(n89), .Q(n176) );
  NOR20 U91 ( .A(n105), .B(n189), .Q(n188) );
  INV0 U92 ( .A(A[8]), .Q(n190) );
  NAND40 U93 ( .A(B[19]), .B(n132), .C(n131), .D(n136), .Q(n245) );
  NAND40 U94 ( .A(B[16]), .B(n9), .C(n214), .D(n89), .Q(n199) );
  INV0 U95 ( .A(B[20]), .Q(n244) );
  NOR20 U96 ( .A(A[20]), .B(n251), .Q(n248) );
  NAND40 U97 ( .A(n9), .B(n248), .C(n89), .D(n249), .Q(n247) );
  NOR20 U98 ( .A(n129), .B(n250), .Q(n249) );
  INV0 U99 ( .A(B[27]), .Q(n165) );
  NAND20 U100 ( .A(B[28]), .B(n166), .Q(n162) );
  INV0 U101 ( .A(B[26]), .Q(n183) );
  INV2 U102 ( .A(n182), .Q(n181) );
  NOR20 U103 ( .A(A[14]), .B(n118), .Q(n117) );
  NAND21 U104 ( .A(n67), .B(n68), .Q(n59) );
  NAND20 U105 ( .A(n54), .B(n173), .Q(n172) );
  INV0 U106 ( .A(A[9]), .Q(n173) );
  INV0 U107 ( .A(A[5]), .Q(n97) );
  INV0 U108 ( .A(B[15]), .Q(n229) );
  NAND20 U109 ( .A(A[7]), .B(n57), .Q(n56) );
  INV0 U110 ( .A(B[28]), .Q(n27) );
  NOR20 U111 ( .A(n25), .B(n26), .Q(n24) );
  NOR20 U112 ( .A(n25), .B(n28), .Q(n23) );
  INV0 U113 ( .A(A[12]), .Q(n228) );
  NOR20 U114 ( .A(n210), .B(n211), .Q(n209) );
  NAND20 U115 ( .A(n10), .B(B[14]), .Q(n115) );
  INV0 U116 ( .A(A[7]), .Q(n107) );
  INV0 U117 ( .A(A[28]), .Q(n166) );
  NAND20 U118 ( .A(n10), .B(n252), .Q(n246) );
  NAND20 U119 ( .A(A[6]), .B(n58), .Q(n55) );
  NAND20 U120 ( .A(B[15]), .B(n9), .Q(n109) );
  INV0 U121 ( .A(A[11]), .Q(n220) );
  NAND20 U122 ( .A(n89), .B(n134), .Q(n128) );
  INV0 U123 ( .A(A[21]), .Q(n134) );
  CLKIN0 U124 ( .A(B[7]), .Q(n57) );
  INV0 U125 ( .A(A[15]), .Q(n112) );
  NAND20 U126 ( .A(A[30]), .B(n21), .Q(n20) );
  NOR20 U127 ( .A(A[10]), .B(n105), .Q(n187) );
  INV0 U128 ( .A(B[4]), .Q(n62) );
  NAND20 U129 ( .A(B[9]), .B(n37), .Q(n160) );
  NAND20 U130 ( .A(n202), .B(n136), .Q(n201) );
  NOR20 U131 ( .A(n137), .B(n203), .Q(n202) );
  NAND20 U132 ( .A(n152), .B(n37), .Q(n122) );
  NAND20 U133 ( .A(n10), .B(n155), .Q(n154) );
  INV0 U134 ( .A(A[17]), .Q(n155) );
  INV0 U135 ( .A(B[30]), .Q(n21) );
  NAND20 U136 ( .A(A[5]), .B(n98), .Q(n92) );
  NAND20 U137 ( .A(A[23]), .B(n256), .Q(n255) );
  INV0 U138 ( .A(B[12]), .Q(n223) );
  NOR21 U139 ( .A(n119), .B(n120), .Q(n116) );
  NOR21 U140 ( .A(n119), .B(n120), .Q(n144) );
  INV3 U141 ( .A(n10), .Q(n91) );
  NAND41 U142 ( .A(n48), .B(n49), .C(n50), .D(n51), .Q(n47) );
  NOR21 U143 ( .A(n52), .B(n53), .Q(n51) );
  NAND22 U144 ( .A(n55), .B(n56), .Q(n52) );
  NAND22 U145 ( .A(n54), .B(n107), .Q(n106) );
  NOR21 U146 ( .A(n137), .B(n138), .Q(n135) );
  AOI311 U147 ( .A(n44), .B(n45), .C(n46), .D(n47), .Q(n38) );
  NOR21 U148 ( .A(n84), .B(n85), .Q(n36) );
  NAND22 U149 ( .A(n69), .B(n70), .Q(n45) );
  AOI2111 U150 ( .A(n195), .B(n196), .C(n197), .D(n198), .Q(n11) );
  NOR21 U151 ( .A(n184), .B(n102), .Q(n179) );
  AOI311 U152 ( .A(n11), .B(n12), .C(n13), .D(n14), .Q(LT_LE) );
  NAND22 U153 ( .A(n86), .B(n87), .Q(n85) );
  NOR21 U154 ( .A(n118), .B(n146), .Q(n145) );
  NAND22 U155 ( .A(n141), .B(n37), .Q(n123) );
  NOR21 U156 ( .A(n142), .B(n143), .Q(n141) );
  NAND22 U157 ( .A(n89), .B(n150), .Q(n142) );
  NAND22 U158 ( .A(n144), .B(n145), .Q(n143) );
  NAND22 U159 ( .A(n156), .B(n136), .Q(n121) );
  NAND22 U160 ( .A(n167), .B(n168), .Q(n161) );
  NAND22 U161 ( .A(n170), .B(n171), .Q(n169) );
  BUF2 U162 ( .A(n103), .Q(n9) );
  NAND22 U163 ( .A(n15), .B(n16), .Q(n14) );
  NOR21 U164 ( .A(n17), .B(n18), .Q(n16) );
  NOR21 U165 ( .A(n23), .B(n24), .Q(n15) );
  NOR21 U166 ( .A(n40), .B(n20), .Q(n17) );
  NOR21 U167 ( .A(n207), .B(n208), .Q(n206) );
  NAND22 U168 ( .A(n212), .B(n131), .Q(n207) );
  NAND22 U169 ( .A(A[24]), .B(n205), .Q(n132) );
  NAND22 U170 ( .A(n54), .B(n190), .Q(n189) );
  INV3 U171 ( .A(B[19]), .Q(n240) );
  AOI311 U172 ( .A(B[18]), .B(n125), .C(n37), .D(n126), .Q(n124) );
  NOR21 U173 ( .A(n110), .B(n139), .Q(n125) );
  NAND22 U174 ( .A(n238), .B(n239), .Q(n237) );
  NAND22 U175 ( .A(n39), .B(n22), .Q(n25) );
  NOR21 U176 ( .A(n42), .B(n43), .Q(n39) );
  INV3 U177 ( .A(B[23]), .Q(n256) );
  AOI221 U178 ( .A(B[3]), .B(n78), .C(n80), .D(n81), .Q(n44) );
  NOR21 U179 ( .A(n63), .B(n83), .Q(n80) );
  INV3 U180 ( .A(B[1]), .Q(n83) );
  NAND22 U181 ( .A(B[5]), .B(n97), .Q(n68) );
  NOR21 U182 ( .A(n19), .B(n40), .Q(n18) );
  NOR21 U183 ( .A(n258), .B(n259), .Q(n257) );
  NOR31 U184 ( .A(n225), .B(n226), .C(n227), .Q(n224) );
  NOR21 U185 ( .A(B[12]), .B(n228), .Q(n226) );
  NOR21 U186 ( .A(n151), .B(n91), .Q(n150) );
  NOR21 U187 ( .A(B[3]), .B(n78), .Q(n63) );
  NOR21 U188 ( .A(n193), .B(n194), .Q(n87) );
  NOR21 U189 ( .A(B[9]), .B(n173), .Q(n194) );
  NOR31 U190 ( .A(n71), .B(n72), .C(n73), .Q(n70) );
  INV3 U191 ( .A(B[0]), .Q(n71) );
  NOR21 U192 ( .A(B[1]), .B(n74), .Q(n73) );
  NOR31 U193 ( .A(n59), .B(n60), .C(n61), .Q(n46) );
  NOR21 U194 ( .A(n63), .B(n64), .Q(n60) );
  NOR31 U195 ( .A(n76), .B(A[0]), .C(n77), .Q(n69) );
  NOR21 U196 ( .A(B[3]), .B(n78), .Q(n77) );
  NAND22 U197 ( .A(n88), .B(n89), .Q(n84) );
  AOI2111 U198 ( .A(n92), .B(n93), .C(n94), .D(n95), .Q(n90) );
  NOR21 U199 ( .A(n105), .B(n172), .Q(n171) );
  NOR31 U200 ( .A(n114), .B(n115), .C(n110), .Q(n113) );
  NAND22 U201 ( .A(n116), .B(n117), .Q(n114) );
  INV3 U202 ( .A(n263), .Q(n129) );
  NOR21 U203 ( .A(n264), .B(n265), .Q(n263) );
  NOR21 U204 ( .A(B[27]), .B(n241), .Q(n265) );
  NOR21 U205 ( .A(B[26]), .B(n242), .Q(n264) );
  NAND22 U206 ( .A(n186), .B(n187), .Q(n185) );
  NOR21 U207 ( .A(n119), .B(n120), .Q(n186) );
  INV3 U208 ( .A(B[24]), .Q(n205) );
  INV3 U209 ( .A(B[17]), .Q(n153) );
  INV3 U210 ( .A(n204), .Q(n203) );
  INV3 U211 ( .A(n40), .Q(n22) );
  INV3 U212 ( .A(B[31]), .Q(n41) );
  OAI2111 U213 ( .A(n160), .B(n161), .C(n162), .D(n163), .Q(n159) );
  NOR31 U214 ( .A(n153), .B(n110), .C(n154), .Q(n152) );
  NAND22 U215 ( .A(n210), .B(n253), .Q(n103) );
  INV3 U216 ( .A(B[11]), .Q(n192) );
  INV3 U217 ( .A(n164), .Q(n163) );
  INV3 U218 ( .A(B[5]), .Q(n98) );
  INV3 U219 ( .A(A[2]), .Q(n79) );
  INV3 U220 ( .A(n65), .Q(n64) );
  NOR21 U221 ( .A(A[2]), .B(n66), .Q(n65) );
  INV3 U222 ( .A(B[2]), .Q(n66) );
  NOR21 U223 ( .A(A[22]), .B(n213), .Q(n212) );
  NOR20 U224 ( .A(A[19]), .B(n251), .Q(n252) );
  NAND21 U225 ( .A(A[19]), .B(n240), .Q(n238) );
  NAND22 U226 ( .A(A[28]), .B(n27), .Q(n26) );
  INV3 U227 ( .A(A[18]), .Q(n140) );
  NOR21 U228 ( .A(A[24]), .B(n205), .Q(n254) );
  NOR21 U229 ( .A(A[27]), .B(n165), .Q(n164) );
  NAND22 U230 ( .A(A[29]), .B(n29), .Q(n28) );
  NOR21 U231 ( .A(A[29]), .B(n29), .Q(n42) );
  NAND20 U232 ( .A(B[10]), .B(n9), .Q(n184) );
  NOR21 U233 ( .A(A[26]), .B(n183), .Q(n182) );
  NAND22 U234 ( .A(A[11]), .B(n192), .Q(n49) );
  NOR21 U235 ( .A(B[2]), .B(n79), .Q(n82) );
  OAI212 U236 ( .A(B[18]), .B(n140), .C(n196), .Q(n235) );
  NAND21 U237 ( .A(A[20]), .B(n244), .Q(n196) );
  NAND22 U238 ( .A(A[16]), .B(n232), .Q(n48) );
  NOR20 U239 ( .A(A[25]), .B(n157), .Q(n156) );
  NAND21 U240 ( .A(A[25]), .B(n157), .Q(n239) );
  NAND22 U241 ( .A(A[4]), .B(n62), .Q(n93) );
  NOR21 U242 ( .A(A[4]), .B(n62), .Q(n61) );
  XNR20 U243 ( .A(B[31]), .B(A[31]), .Q(n19) );
  NOR21 U244 ( .A(A[31]), .B(n41), .Q(n40) );
  INV2 U245 ( .A(B[14]), .Q(n230) );
  NOR21 U246 ( .A(B[22]), .B(n133), .Q(n260) );
  NOR20 U247 ( .A(A[30]), .B(n21), .Q(n43) );
  CLKIN0 U248 ( .A(B[13]), .Q(n151) );
  NAND31 U249 ( .A(B[20]), .B(n132), .C(n131), .Q(n250) );
  NOR21 U250 ( .A(B[8]), .B(n190), .Q(n193) );
  NOR21 U251 ( .A(B[0]), .B(n75), .Q(n72) );
  CLKIN3 U252 ( .A(n54), .Q(n53) );
  CLKIN3 U253 ( .A(n67), .Q(n95) );
  CLKIN3 U254 ( .A(n68), .Q(n94) );
  OAI222 U255 ( .A(n127), .B(n128), .C(n129), .D(n130), .Q(n126) );
  CLKIN3 U256 ( .A(n149), .Q(n118) );
  OAI312 U257 ( .A(n174), .B(n175), .C(n176), .D(n177), .Q(n158) );
  CLKIN3 U258 ( .A(n48), .Q(n119) );
  CLKIN3 U259 ( .A(n131), .Q(n137) );
  CLKIN3 U260 ( .A(n132), .Q(n213) );
  OAI222 U261 ( .A(n175), .B(n215), .C(n175), .D(n216), .Q(n197) );
  CLKIN3 U262 ( .A(n102), .Q(n86) );
  CLKIN3 U263 ( .A(n50), .Q(n120) );
  CLKIN3 U264 ( .A(n243), .Q(n251) );
  CLKIN3 U265 ( .A(n255), .Q(n210) );
  CLKIN3 U266 ( .A(n261), .Q(n133) );
endmodule


module E_alu_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291;

  AOI221 U3 ( .A(A[30]), .B(n189), .C(A[31]), .D(n190), .Q(n270) );
  NAND20 U4 ( .A(A[31]), .B(n10), .Q(n240) );
  NAND21 U5 ( .A(A[31]), .B(n189), .Q(n158) );
  AOI221 U6 ( .A(A[28]), .B(n9), .C(A[29]), .D(n5), .Q(n271) );
  AOI220 U7 ( .A(A[16]), .B(n189), .C(A[17]), .D(n190), .Q(n257) );
  AOI220 U8 ( .A(A[16]), .B(n9), .C(n6), .D(A[17]), .Q(n277) );
  NAND21 U9 ( .A(n99), .B(n129), .Q(n128) );
  AOI220 U10 ( .A(n98), .B(n103), .C(n99), .D(n101), .Q(n131) );
  NAND21 U11 ( .A(n13), .B(n117), .Q(n127) );
  CLKIN2 U12 ( .A(n115), .Q(B[28]) );
  CLKIN2 U13 ( .A(n100), .Q(B[31]) );
  NAND20 U14 ( .A(n102), .B(n19), .Q(n100) );
  CLKIN3 U15 ( .A(n112), .Q(B[29]) );
  NOR20 U16 ( .A(n18), .B(n20), .Q(B[25]) );
  OAI211 U17 ( .A(n123), .B(n124), .C(n125), .Q(n122) );
  NAND21 U18 ( .A(n12), .B(n114), .Q(n125) );
  NAND22 U19 ( .A(n113), .B(n19), .Q(n112) );
  NAND20 U20 ( .A(n93), .B(n94), .Q(n89) );
  NAND20 U21 ( .A(n98), .B(n94), .Q(n170) );
  NAND41 U22 ( .A(n89), .B(n90), .C(n91), .D(n92), .Q(n88) );
  AOI220 U23 ( .A(A[30]), .B(n9), .C(A[31]), .D(n6), .Q(n245) );
  INV3 U24 ( .A(n140), .Q(n123) );
  NAND22 U25 ( .A(n40), .B(n121), .Q(n242) );
  NAND21 U26 ( .A(n97), .B(n94), .Q(n132) );
  NAND21 U27 ( .A(n33), .B(n44), .Q(n211) );
  NAND22 U28 ( .A(n40), .B(n41), .Q(n39) );
  NAND22 U29 ( .A(n40), .B(n63), .Q(n62) );
  INV2 U30 ( .A(n66), .Q(n60) );
  NAND21 U31 ( .A(n12), .B(n107), .Q(n243) );
  NAND22 U32 ( .A(n99), .B(n136), .Q(n244) );
  AOI220 U33 ( .A(n97), .B(n117), .C(n93), .D(n129), .Q(n269) );
  MUX22 U34 ( .A(n267), .B(n162), .S(n18), .Q(B[0]) );
  INV2 U35 ( .A(n181), .Q(n180) );
  INV3 U36 ( .A(n51), .Q(n130) );
  NAND20 U37 ( .A(n28), .B(n114), .Q(n183) );
  NAND20 U38 ( .A(n26), .B(n29), .Q(n182) );
  AOI220 U39 ( .A(n26), .B(n71), .C(n28), .D(n105), .Q(n250) );
  AOI220 U40 ( .A(n97), .B(n53), .C(n93), .D(n58), .Q(n96) );
  AOI220 U41 ( .A(n30), .B(n52), .C(n33), .D(n53), .Q(n49) );
  NAND20 U42 ( .A(n40), .B(n51), .Q(n50) );
  AOI220 U43 ( .A(n26), .B(n44), .C(n28), .D(n45), .Q(n37) );
  AOI220 U44 ( .A(n28), .B(n29), .C(n30), .D(n31), .Q(n24) );
  NAND20 U45 ( .A(n12), .B(n59), .Q(n91) );
  NAND20 U46 ( .A(n97), .B(n101), .Q(n92) );
  AOI220 U47 ( .A(n98), .B(n44), .C(n99), .D(n45), .Q(n268) );
  AOI220 U48 ( .A(n97), .B(n107), .C(n93), .D(n136), .Q(n153) );
  AOI220 U49 ( .A(n13), .B(n71), .C(n99), .D(n105), .Q(n152) );
  AOI220 U50 ( .A(n12), .B(n27), .C(n99), .D(n29), .Q(n155) );
  NAND30 U51 ( .A(n159), .B(n160), .C(n158), .Q(n157) );
  NAND20 U52 ( .A(n99), .B(n103), .Q(n90) );
  NAND20 U53 ( .A(n28), .B(n27), .Q(n77) );
  NAND20 U54 ( .A(n26), .B(n27), .Q(n25) );
  NAND20 U55 ( .A(n33), .B(n27), .Q(n198) );
  NAND21 U56 ( .A(n28), .B(n117), .Q(n213) );
  NAND20 U57 ( .A(n26), .B(n103), .Q(n168) );
  NAND20 U58 ( .A(n28), .B(n71), .Q(n68) );
  NAND20 U59 ( .A(n26), .B(n58), .Q(n57) );
  NAND20 U60 ( .A(n28), .B(n59), .Q(n56) );
  CLKIN3 U61 ( .A(n215), .Q(n116) );
  NAND20 U62 ( .A(n98), .B(n129), .Q(n215) );
  AOI220 U63 ( .A(n33), .B(n71), .C(n40), .D(n106), .Q(n172) );
  NAND20 U64 ( .A(n28), .B(n44), .Q(n84) );
  NAND20 U65 ( .A(n28), .B(n101), .Q(n167) );
  NAND20 U66 ( .A(n28), .B(n107), .Q(n176) );
  NAND20 U67 ( .A(n26), .B(n105), .Q(n177) );
  AOI220 U68 ( .A(n33), .B(n59), .C(n40), .D(n102), .Q(n163) );
  MUX22 U69 ( .A(n87), .B(n88), .S(n18), .Q(B[3]) );
  MUX21 U70 ( .A(n108), .B(n109), .S(n18), .Q(B[2]) );
  MUX21 U71 ( .A(n144), .B(n145), .S(n18), .Q(B[1]) );
  NAND20 U72 ( .A(n30), .B(n58), .Q(n169) );
  AOI220 U73 ( .A(A[15]), .B(n9), .C(A[16]), .D(n6), .Q(n225) );
  AOI220 U74 ( .A(A[24]), .B(n189), .C(A[25]), .D(n190), .Q(n251) );
  AOI220 U75 ( .A(A[15]), .B(n189), .C(A[16]), .D(n190), .Q(n185) );
  AOI220 U76 ( .A(A[11]), .B(n189), .C(A[12]), .D(n190), .Q(n201) );
  AOI220 U77 ( .A(A[14]), .B(n189), .C(A[15]), .D(n190), .Q(n280) );
  AOI220 U78 ( .A(A[11]), .B(n9), .C(A[12]), .D(n7), .Q(n223) );
  AOI220 U79 ( .A(A[3]), .B(n9), .C(A[4]), .D(n6), .Q(n235) );
  AOI220 U80 ( .A(A[29]), .B(n189), .C(A[30]), .D(n190), .Q(n238) );
  AOI220 U81 ( .A(A[27]), .B(n11), .C(A[28]), .D(n7), .Q(n239) );
  AOI220 U82 ( .A(A[25]), .B(n189), .C(A[26]), .D(n190), .Q(n230) );
  AOI220 U83 ( .A(A[24]), .B(n8), .C(A[25]), .D(n5), .Q(n273) );
  AOI220 U84 ( .A(A[26]), .B(n189), .C(A[27]), .D(n190), .Q(n272) );
  AOI220 U85 ( .A(A[28]), .B(n189), .C(A[29]), .D(n190), .Q(n246) );
  AOI220 U86 ( .A(A[26]), .B(n9), .C(A[27]), .D(n7), .Q(n247) );
  AOI220 U87 ( .A(A[27]), .B(n189), .C(A[28]), .D(n190), .Q(n191) );
  AOI220 U88 ( .A(A[25]), .B(n10), .C(A[26]), .D(n7), .Q(n192) );
  AOI220 U89 ( .A(A[14]), .B(n8), .C(A[15]), .D(n6), .Q(n258) );
  AOI220 U90 ( .A(A[3]), .B(n189), .C(A[4]), .D(n190), .Q(n195) );
  NAND20 U91 ( .A(A[29]), .B(n11), .Q(n160) );
  NAND20 U92 ( .A(A[30]), .B(n5), .Q(n159) );
  NAND20 U93 ( .A(n119), .B(n19), .Q(n118) );
  NAND20 U94 ( .A(n116), .B(n19), .Q(n115) );
  NOR21 U95 ( .A(n22), .B(n23), .Q(n21) );
  INV3 U96 ( .A(n32), .Q(n22) );
  NAND22 U97 ( .A(n24), .B(n25), .Q(n23) );
  NOR21 U98 ( .A(n74), .B(n75), .Q(n73) );
  NAND22 U99 ( .A(n78), .B(n79), .Q(n74) );
  NAND22 U100 ( .A(n76), .B(n77), .Q(n75) );
  AOI211 U101 ( .A(n40), .B(n113), .C(n197), .Q(n179) );
  INV3 U102 ( .A(n198), .Q(n197) );
  NAND22 U103 ( .A(n241), .B(n242), .Q(B[10]) );
  INV3 U104 ( .A(n248), .Q(n241) );
  NAND22 U105 ( .A(n249), .B(n250), .Q(n248) );
  NAND22 U106 ( .A(n207), .B(n208), .Q(B[12]) );
  NAND22 U107 ( .A(n40), .B(n116), .Q(n207) );
  NOR21 U108 ( .A(n209), .B(n210), .Q(n208) );
  NAND22 U109 ( .A(n211), .B(n212), .Q(n210) );
  NOR21 U110 ( .A(n123), .B(n205), .Q(n113) );
  INV3 U111 ( .A(n98), .Q(n205) );
  BUF2 U112 ( .A(n187), .Q(n10) );
  BUF2 U113 ( .A(n187), .Q(n11) );
  INV3 U114 ( .A(n19), .Q(n40) );
  NAND31 U115 ( .A(n159), .B(n160), .C(n158), .Q(n140) );
  NAND31 U116 ( .A(n182), .B(n183), .C(n184), .Q(n181) );
  NAND22 U117 ( .A(n30), .B(n34), .Q(n184) );
  AOI221 U118 ( .A(n30), .B(n65), .C(n33), .D(n70), .Q(n249) );
  NAND31 U119 ( .A(n38), .B(n39), .C(n37), .Q(B[8]) );
  AOI221 U120 ( .A(n30), .B(n42), .C(n33), .D(n43), .Q(n38) );
  NAND31 U121 ( .A(n60), .B(n61), .C(n62), .Q(B[6]) );
  AOI221 U122 ( .A(n30), .B(n64), .C(n33), .D(n65), .Q(n61) );
  NAND22 U123 ( .A(n138), .B(n139), .Q(n137) );
  NAND22 U124 ( .A(n97), .B(n140), .Q(n139) );
  AOI221 U125 ( .A(n12), .B(n29), .C(n99), .D(n114), .Q(n138) );
  NAND22 U126 ( .A(n142), .B(n143), .Q(n141) );
  NAND22 U127 ( .A(n97), .B(n129), .Q(n143) );
  AOI221 U128 ( .A(n98), .B(n45), .C(n99), .D(n117), .Q(n142) );
  AOI2111 U129 ( .A(n26), .B(n43), .C(n82), .D(n83), .Q(n81) );
  INV3 U130 ( .A(n86), .Q(n82) );
  NAND22 U131 ( .A(n84), .B(n85), .Q(n83) );
  NAND22 U132 ( .A(n236), .B(n237), .Q(n119) );
  NAND22 U133 ( .A(n99), .B(n94), .Q(n236) );
  NAND22 U134 ( .A(n13), .B(n101), .Q(n237) );
  NAND31 U135 ( .A(n48), .B(n49), .C(n50), .Q(B[7]) );
  INV3 U136 ( .A(n54), .Q(n48) );
  NAND22 U137 ( .A(n127), .B(n128), .Q(n41) );
  NAND22 U138 ( .A(n131), .B(n132), .Q(n51) );
  NAND22 U139 ( .A(n243), .B(n244), .Q(n121) );
  NAND22 U140 ( .A(n134), .B(n135), .Q(n63) );
  NAND22 U141 ( .A(n97), .B(n136), .Q(n135) );
  AOI221 U142 ( .A(n13), .B(n105), .C(n99), .D(n107), .Q(n134) );
  NAND22 U143 ( .A(n152), .B(n153), .Q(n109) );
  NAND22 U144 ( .A(n155), .B(n156), .Q(n145) );
  AOI221 U145 ( .A(n97), .B(n114), .C(n93), .D(n157), .Q(n156) );
  NAND22 U146 ( .A(n268), .B(n269), .Q(n162) );
  NAND22 U147 ( .A(n30), .B(n43), .Q(n212) );
  NAND22 U148 ( .A(n26), .B(n59), .Q(n227) );
  NAND22 U149 ( .A(n176), .B(n177), .Q(n175) );
  NAND22 U150 ( .A(n33), .B(n34), .Q(n32) );
  NAND22 U151 ( .A(n213), .B(n214), .Q(n209) );
  NAND22 U152 ( .A(n26), .B(n45), .Q(n214) );
  NAND22 U153 ( .A(n30), .B(n46), .Q(n85) );
  NAND22 U154 ( .A(n30), .B(n36), .Q(n79) );
  NOR21 U155 ( .A(n18), .B(n161), .Q(B[16]) );
  NAND22 U156 ( .A(n68), .B(n69), .Q(n66) );
  NAND22 U157 ( .A(n26), .B(n70), .Q(n69) );
  NAND22 U158 ( .A(n33), .B(n58), .Q(n220) );
  NAND22 U159 ( .A(n56), .B(n57), .Q(n54) );
  NOR21 U160 ( .A(n18), .B(n148), .Q(B[19]) );
  AOI2111 U161 ( .A(n93), .B(n94), .C(n149), .D(n150), .Q(n148) );
  INV3 U162 ( .A(n92), .Q(n150) );
  NAND22 U163 ( .A(n90), .B(n91), .Q(n149) );
  NAND22 U164 ( .A(n28), .B(n103), .Q(n226) );
  NOR21 U165 ( .A(n18), .B(n154), .Q(B[17]) );
  NOR21 U166 ( .A(n18), .B(n80), .Q(B[20]) );
  NOR21 U167 ( .A(n218), .B(n219), .Q(n217) );
  NAND22 U168 ( .A(n220), .B(n221), .Q(n219) );
  NAND22 U169 ( .A(n226), .B(n227), .Q(n218) );
  NAND22 U170 ( .A(n30), .B(n53), .Q(n221) );
  NOR21 U171 ( .A(n18), .B(n120), .Q(B[26]) );
  NOR21 U172 ( .A(n18), .B(n151), .Q(B[18]) );
  NOR21 U173 ( .A(n18), .B(n133), .Q(B[22]) );
  NAND22 U174 ( .A(n163), .B(n164), .Q(B[15]) );
  NOR21 U175 ( .A(n165), .B(n166), .Q(n164) );
  NAND22 U176 ( .A(n167), .B(n168), .Q(n166) );
  NAND22 U177 ( .A(n171), .B(n172), .Q(B[14]) );
  NOR21 U178 ( .A(n174), .B(n175), .Q(n171) );
  INV3 U179 ( .A(n178), .Q(n174) );
  NOR21 U180 ( .A(n40), .B(n72), .Q(B[21]) );
  INV3 U181 ( .A(n169), .Q(n165) );
  NAND22 U182 ( .A(n278), .B(n279), .Q(n267) );
  AOI221 U183 ( .A(n97), .B(n42), .C(n93), .D(n43), .Q(n279) );
  NAND22 U184 ( .A(n95), .B(n96), .Q(n87) );
  NAND22 U185 ( .A(n146), .B(n147), .Q(n144) );
  AOI221 U186 ( .A(n93), .B(n34), .C(n97), .D(n31), .Q(n147) );
  NAND22 U187 ( .A(n110), .B(n111), .Q(n108) );
  AOI221 U188 ( .A(n93), .B(n70), .C(n97), .D(n65), .Q(n111) );
  INV3 U189 ( .A(n206), .Q(n190) );
  NAND22 U190 ( .A(SH[1]), .B(SH[0]), .Q(n206) );
  BUF2 U191 ( .A(n188), .Q(n6) );
  NOR21 U192 ( .A(SH[1]), .B(SH[0]), .Q(n187) );
  NOR21 U193 ( .A(SH[1]), .B(SH[0]), .Q(n8) );
  NOR21 U194 ( .A(SH[1]), .B(SH[0]), .Q(n9) );
  NAND22 U195 ( .A(n33), .B(n42), .Q(n86) );
  NAND22 U196 ( .A(n30), .B(n70), .Q(n178) );
  BUF2 U197 ( .A(n188), .Q(n7) );
  BUF2 U198 ( .A(n188), .Q(n5) );
  NAND22 U199 ( .A(n26), .B(n34), .Q(n76) );
  NAND22 U200 ( .A(n33), .B(n31), .Q(n78) );
  NOR21 U201 ( .A(n18), .B(n126), .Q(B[24]) );
  INV3 U202 ( .A(n170), .Q(n102) );
  INV3 U203 ( .A(n173), .Q(n106) );
  NAND22 U204 ( .A(n13), .B(n136), .Q(n173) );
  NOR21 U205 ( .A(SH[3]), .B(SH[2]), .Q(n98) );
  NOR21 U206 ( .A(SH[3]), .B(SH[2]), .Q(n12) );
  NOR21 U207 ( .A(SH[3]), .B(SH[2]), .Q(n13) );
  INV3 U208 ( .A(n124), .Q(n99) );
  INV3 U209 ( .A(n282), .Q(n93) );
  NAND22 U210 ( .A(SH[3]), .B(SH[2]), .Q(n282) );
  NAND22 U211 ( .A(n203), .B(n204), .Q(n36) );
  NAND22 U212 ( .A(n263), .B(n264), .Q(n64) );
  NAND22 U213 ( .A(n199), .B(n200), .Q(n27) );
  NAND22 U214 ( .A(n185), .B(n186), .Q(n34) );
  NAND22 U215 ( .A(n238), .B(n239), .Q(n101) );
  NAND22 U216 ( .A(n270), .B(n271), .Q(n129) );
  NAND22 U217 ( .A(n228), .B(n229), .Q(n59) );
  NAND22 U218 ( .A(n224), .B(n225), .Q(n58) );
  NAND22 U219 ( .A(n230), .B(n231), .Q(n103) );
  AOI221 U220 ( .A(A[23]), .B(n8), .C(A[24]), .D(n6), .Q(n231) );
  NAND22 U221 ( .A(n280), .B(n281), .Q(n43) );
  NAND22 U222 ( .A(n193), .B(n194), .Q(n29) );
  AOI221 U223 ( .A(A[23]), .B(n189), .C(A[24]), .D(n190), .Q(n193) );
  NAND22 U224 ( .A(n251), .B(n252), .Q(n105) );
  NAND22 U225 ( .A(n254), .B(n255), .Q(n71) );
  NAND22 U226 ( .A(n246), .B(n247), .Q(n107) );
  NAND22 U227 ( .A(n191), .B(n192), .Q(n114) );
  NAND22 U228 ( .A(n272), .B(n273), .Q(n117) );
  NAND22 U229 ( .A(n276), .B(n277), .Q(n44) );
  NAND22 U230 ( .A(n274), .B(n275), .Q(n45) );
  NAND22 U231 ( .A(n201), .B(n202), .Q(n31) );
  NAND22 U232 ( .A(n283), .B(n284), .Q(n42) );
  NAND22 U233 ( .A(n260), .B(n261), .Q(n65) );
  NAND22 U234 ( .A(n222), .B(n223), .Q(n53) );
  NOR21 U235 ( .A(n18), .B(n130), .Q(B[23]) );
  INV3 U236 ( .A(n118), .Q(B[27]) );
  NAND22 U237 ( .A(n216), .B(n217), .Q(B[11]) );
  NAND22 U238 ( .A(n40), .B(n119), .Q(n216) );
  NAND22 U239 ( .A(n286), .B(n287), .Q(n46) );
  AOI221 U240 ( .A(n99), .B(n36), .C(n13), .D(n35), .Q(n146) );
  NAND22 U241 ( .A(n195), .B(n196), .Q(n35) );
  AOI221 U242 ( .A(n99), .B(n64), .C(n98), .D(n67), .Q(n110) );
  NAND22 U243 ( .A(n265), .B(n266), .Q(n67) );
  AOI221 U244 ( .A(n13), .B(n47), .C(n99), .D(n46), .Q(n278) );
  NAND22 U245 ( .A(n288), .B(n289), .Q(n47) );
  INV3 U246 ( .A(n245), .Q(n136) );
  INV3 U247 ( .A(n104), .Q(B[30]) );
  AOI221 U248 ( .A(n12), .B(n55), .C(n99), .D(n52), .Q(n95) );
  NAND22 U249 ( .A(n234), .B(n235), .Q(n55) );
  NAND22 U250 ( .A(n232), .B(n233), .Q(n52) );
  INV3 U251 ( .A(n291), .Q(n189) );
  NAND22 U252 ( .A(SH[1]), .B(n14), .Q(n291) );
  NAND22 U253 ( .A(n257), .B(n258), .Q(n70) );
  INV3 U254 ( .A(n240), .Q(n94) );
  INV3 U255 ( .A(n290), .Q(n188) );
  NAND22 U256 ( .A(SH[0]), .B(n15), .Q(n290) );
  NAND22 U257 ( .A(n106), .B(n19), .Q(n104) );
  INV3 U258 ( .A(n19), .Q(n18) );
  NAND22 U259 ( .A(SH[2]), .B(n17), .Q(n124) );
  INV3 U260 ( .A(n256), .Q(n26) );
  NAND22 U261 ( .A(n97), .B(n19), .Q(n256) );
  INV3 U262 ( .A(n262), .Q(n30) );
  NAND22 U263 ( .A(n12), .B(n19), .Q(n262) );
  INV3 U264 ( .A(n259), .Q(n33) );
  NAND22 U265 ( .A(n99), .B(n19), .Q(n259) );
  INV3 U266 ( .A(n253), .Q(n28) );
  NAND22 U267 ( .A(n93), .B(n19), .Q(n253) );
  INV3 U268 ( .A(n285), .Q(n97) );
  NAND22 U269 ( .A(SH[3]), .B(n16), .Q(n285) );
  INV3 U270 ( .A(SH[0]), .Q(n14) );
  INV3 U271 ( .A(SH[1]), .Q(n15) );
  INV3 U272 ( .A(SH[4]), .Q(n19) );
  INV3 U273 ( .A(SH[3]), .Q(n17) );
  INV3 U274 ( .A(SH[2]), .Q(n16) );
  OAI212 U275 ( .A(n72), .B(n19), .C(n73), .Q(B[5]) );
  AOI220 U276 ( .A(A[9]), .B(n189), .C(A[10]), .D(n190), .Q(n232) );
  AOI220 U277 ( .A(A[9]), .B(n11), .C(A[10]), .D(n7), .Q(n202) );
  AOI220 U278 ( .A(A[10]), .B(n189), .C(A[11]), .D(n190), .Q(n283) );
  AOI220 U279 ( .A(A[10]), .B(n187), .C(A[11]), .D(n7), .Q(n261) );
  AOI220 U280 ( .A(A[1]), .B(n11), .C(A[2]), .D(n7), .Q(n196) );
  AOI220 U281 ( .A(A[2]), .B(n10), .C(A[3]), .D(n5), .Q(n266) );
  AOI220 U282 ( .A(A[2]), .B(n189), .C(A[3]), .D(n190), .Q(n288) );
  AOI220 U283 ( .A(A[17]), .B(n10), .C(A[18]), .D(n6), .Q(n200) );
  AOI220 U284 ( .A(A[18]), .B(n10), .C(A[19]), .D(n7), .Q(n255) );
  AOI220 U285 ( .A(n189), .B(A[17]), .C(A[18]), .D(n190), .Q(n224) );
  AOI220 U286 ( .A(n189), .B(A[18]), .C(A[19]), .D(n190), .Q(n276) );
  AOI220 U287 ( .A(A[21]), .B(n189), .C(A[22]), .D(n190), .Q(n228) );
  AOI220 U288 ( .A(A[21]), .B(n10), .C(A[22]), .D(n6), .Q(n194) );
  AOI220 U289 ( .A(A[22]), .B(n9), .C(A[23]), .D(n6), .Q(n252) );
  AOI220 U290 ( .A(A[22]), .B(n189), .C(A[23]), .D(n190), .Q(n274) );
  AOI220 U291 ( .A(A[6]), .B(n189), .C(A[7]), .D(n190), .Q(n286) );
  AOI220 U292 ( .A(A[6]), .B(n11), .C(A[7]), .D(n5), .Q(n264) );
  AOI220 U293 ( .A(A[4]), .B(n189), .C(A[5]), .D(n190), .Q(n265) );
  AOI220 U294 ( .A(A[4]), .B(n8), .C(A[5]), .D(n5), .Q(n287) );
  AOI220 U295 ( .A(A[5]), .B(n189), .C(A[6]), .D(n190), .Q(n234) );
  AOI220 U296 ( .A(A[5]), .B(n9), .C(A[6]), .D(n6), .Q(n204) );
  AOI220 U297 ( .A(A[12]), .B(n8), .C(A[13]), .D(n5), .Q(n281) );
  AOI220 U298 ( .A(A[12]), .B(n189), .C(A[13]), .D(n190), .Q(n260) );
  AOI220 U299 ( .A(A[13]), .B(n189), .C(A[14]), .D(n190), .Q(n222) );
  AOI220 U300 ( .A(A[13]), .B(n10), .C(A[14]), .D(n6), .Q(n186) );
  AOI221 U301 ( .A(A[20]), .B(n9), .C(A[21]), .D(n5), .Q(n275) );
  AOI221 U302 ( .A(A[20]), .B(n189), .C(A[21]), .D(n190), .Q(n254) );
  AOI221 U303 ( .A(A[19]), .B(n8), .C(A[20]), .D(n7), .Q(n229) );
  AOI221 U304 ( .A(A[19]), .B(n189), .C(A[20]), .D(n190), .Q(n199) );
  AOI220 U305 ( .A(A[7]), .B(n10), .C(A[8]), .D(n7), .Q(n233) );
  AOI220 U306 ( .A(A[7]), .B(n189), .C(A[8]), .D(n190), .Q(n203) );
  AOI220 U307 ( .A(A[8]), .B(n189), .C(A[9]), .D(n190), .Q(n263) );
  AOI220 U308 ( .A(A[8]), .B(n10), .C(A[9]), .D(n5), .Q(n284) );
  AOI220 U309 ( .A(n11), .B(A[0]), .C(A[1]), .D(n5), .Q(n289) );
  OAI212 U310 ( .A(n20), .B(n19), .C(n21), .Q(B[9]) );
  OAI212 U311 ( .A(n80), .B(n19), .C(n81), .Q(B[4]) );
  CLKIN3 U312 ( .A(n121), .Q(n120) );
  CLKIN3 U313 ( .A(n122), .Q(n20) );
  CLKIN3 U314 ( .A(n41), .Q(n126) );
  CLKIN3 U315 ( .A(n63), .Q(n133) );
  CLKIN3 U316 ( .A(n137), .Q(n72) );
  CLKIN3 U317 ( .A(n141), .Q(n80) );
  CLKIN3 U318 ( .A(n109), .Q(n151) );
  CLKIN3 U319 ( .A(n145), .Q(n154) );
  CLKIN3 U320 ( .A(n162), .Q(n161) );
  NAND22 U321 ( .A(n179), .B(n180), .Q(B[13]) );
endmodule


module E_alu_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   ML_int_1__31_, ML_int_1__30_, ML_int_1__29_, ML_int_1__28_,
         ML_int_1__27_, ML_int_1__26_, ML_int_1__25_, ML_int_1__24_,
         ML_int_1__23_, ML_int_1__22_, ML_int_1__21_, ML_int_1__20_,
         ML_int_1__19_, ML_int_1__18_, ML_int_1__17_, ML_int_1__16_,
         ML_int_1__15_, ML_int_1__14_, ML_int_1__13_, ML_int_1__12_,
         ML_int_1__11_, ML_int_1__10_, ML_int_1__9_, ML_int_1__8_,
         ML_int_1__7_, ML_int_1__6_, ML_int_1__5_, ML_int_1__4_, ML_int_1__3_,
         ML_int_1__2_, ML_int_1__1_, ML_int_1__0_, ML_int_2__31_,
         ML_int_2__30_, ML_int_2__29_, ML_int_2__28_, ML_int_2__27_,
         ML_int_2__26_, ML_int_2__25_, ML_int_2__24_, ML_int_2__23_,
         ML_int_2__22_, ML_int_2__21_, ML_int_2__20_, ML_int_2__19_,
         ML_int_2__18_, ML_int_2__17_, ML_int_2__16_, ML_int_2__15_,
         ML_int_2__14_, ML_int_2__13_, ML_int_2__12_, ML_int_2__11_,
         ML_int_2__10_, ML_int_2__9_, ML_int_2__8_, ML_int_2__7_, ML_int_2__6_,
         ML_int_2__5_, ML_int_2__4_, ML_int_2__3_, ML_int_2__2_, ML_int_2__1_,
         ML_int_2__0_, ML_int_3__31_, ML_int_3__30_, ML_int_3__29_,
         ML_int_3__28_, ML_int_3__27_, ML_int_3__26_, ML_int_3__25_,
         ML_int_3__24_, ML_int_3__23_, ML_int_3__22_, ML_int_3__21_,
         ML_int_3__20_, ML_int_3__19_, ML_int_3__18_, ML_int_3__17_,
         ML_int_3__16_, ML_int_3__15_, ML_int_3__14_, ML_int_3__13_,
         ML_int_3__12_, ML_int_3__11_, ML_int_3__10_, ML_int_3__9_,
         ML_int_3__8_, ML_int_3__7_, ML_int_3__6_, ML_int_3__5_, ML_int_3__4_,
         ML_int_3__3_, ML_int_3__2_, ML_int_3__1_, ML_int_3__0_, ML_int_4__31_,
         ML_int_4__30_, ML_int_4__29_, ML_int_4__28_, ML_int_4__27_,
         ML_int_4__26_, ML_int_4__25_, ML_int_4__24_, ML_int_4__23_,
         ML_int_4__22_, ML_int_4__21_, ML_int_4__20_, ML_int_4__19_,
         ML_int_4__18_, ML_int_4__17_, ML_int_4__16_, ML_int_4__15_,
         ML_int_4__14_, ML_int_4__13_, ML_int_4__12_, ML_int_4__11_,
         ML_int_4__10_, ML_int_4__9_, ML_int_4__8_, ML_int_4__7_, ML_int_4__6_,
         ML_int_4__5_, ML_int_4__4_, ML_int_4__3_, ML_int_4__2_, ML_int_4__1_,
         ML_int_4__0_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56;

  MUX21 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n32), .Q(ML_int_1__1_) );
  MUX21 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n33), .Q(ML_int_1__8_) );
  MUX21 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n33), .Q(ML_int_1__9_) );
  MUX22 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n35), .Q(ML_int_1__20_) );
  MUX21 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n35), .Q(ML_int_1__21_) );
  MUX21 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n34), .Q(ML_int_1__13_) );
  MUX21 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n33), .Q(ML_int_1__5_) );
  MUX21 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n33), .Q(ML_int_1__6_) );
  MUX21 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n35), .Q(ML_int_1__22_) );
  MUX21 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n35), .Q(ML_int_1__23_) );
  MUX21 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n35), .Q(ML_int_1__18_) );
  MUX21 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n36), .Q(ML_int_1__19_) );
  MUX21 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n32), .Q(ML_int_1__3_) );
  MUX21 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n32), .Q(ML_int_1__2_) );
  MUX21 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n34), .Q(ML_int_1__11_) );
  MUX21 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n34), .Q(ML_int_1__10_) );
  MUX22 M1_3_23 ( .A(ML_int_3__23_), .B(ML_int_3__15_), .S(n54), .Q(
        ML_int_4__23_) );
  MUX22 M1_2_28 ( .A(ML_int_2__28_), .B(ML_int_2__24_), .S(n49), .Q(
        ML_int_3__28_) );
  MUX22 M1_3_28 ( .A(ML_int_3__28_), .B(ML_int_3__20_), .S(n55), .Q(
        ML_int_4__28_) );
  MUX22 M1_4_28 ( .A(ML_int_4__28_), .B(ML_int_4__12_), .S(SH[4]), .Q(B[28])
         );
  MUX22 M1_3_25 ( .A(ML_int_3__25_), .B(ML_int_3__17_), .S(n55), .Q(
        ML_int_4__25_) );
  MUX22 M1_4_25 ( .A(ML_int_4__25_), .B(ML_int_4__9_), .S(SH[4]), .Q(B[25]) );
  MUX22 M1_4_24 ( .A(ML_int_4__24_), .B(ML_int_4__8_), .S(SH[4]), .Q(B[24]) );
  MUX22 M1_4_20 ( .A(ML_int_4__20_), .B(ML_int_4__4_), .S(SH[4]), .Q(B[20]) );
  MUX22 M1_1_30 ( .A(ML_int_1__30_), .B(ML_int_1__28_), .S(n43), .Q(
        ML_int_2__30_) );
  MUX22 M1_2_30 ( .A(ML_int_2__30_), .B(ML_int_2__26_), .S(n49), .Q(
        ML_int_3__30_) );
  MUX22 M1_3_30 ( .A(ML_int_3__30_), .B(ML_int_3__22_), .S(n54), .Q(
        ML_int_4__30_) );
  MUX22 M1_4_30 ( .A(ML_int_4__30_), .B(ML_int_4__14_), .S(SH[4]), .Q(B[30])
         );
  MUX22 M1_1_31 ( .A(ML_int_1__31_), .B(ML_int_1__29_), .S(n43), .Q(
        ML_int_2__31_) );
  MUX22 M1_2_31 ( .A(ML_int_2__31_), .B(ML_int_2__27_), .S(n49), .Q(
        ML_int_3__31_) );
  MUX22 M1_3_31 ( .A(ML_int_3__31_), .B(ML_int_3__23_), .S(n50), .Q(
        ML_int_4__31_) );
  MUX22 M1_4_31 ( .A(ML_int_4__31_), .B(ML_int_4__15_), .S(SH[4]), .Q(B[31])
         );
  MUX22 M1_4_19 ( .A(ML_int_4__19_), .B(ML_int_4__3_), .S(SH[4]), .Q(B[19]) );
  MUX22 M1_1_29 ( .A(ML_int_1__29_), .B(ML_int_1__27_), .S(n42), .Q(
        ML_int_2__29_) );
  MUX22 M1_2_29 ( .A(ML_int_2__29_), .B(ML_int_2__25_), .S(n49), .Q(
        ML_int_3__29_) );
  MUX22 M1_3_29 ( .A(ML_int_3__29_), .B(ML_int_3__21_), .S(n55), .Q(
        ML_int_4__29_) );
  MUX22 M1_4_29 ( .A(ML_int_4__29_), .B(ML_int_4__13_), .S(SH[4]), .Q(B[29])
         );
  MUX22 M1_2_27 ( .A(ML_int_2__27_), .B(ML_int_2__23_), .S(n49), .Q(
        ML_int_3__27_) );
  MUX22 M1_1_3 ( .A(ML_int_1__3_), .B(ML_int_1__1_), .S(n38), .Q(ML_int_2__3_)
         );
  MUX22 M1_3_12 ( .A(ML_int_3__12_), .B(ML_int_3__4_), .S(n52), .Q(
        ML_int_4__12_) );
  MUX22 M1_3_14 ( .A(ML_int_3__14_), .B(ML_int_3__6_), .S(n52), .Q(
        ML_int_4__14_) );
  MUX22 M1_3_13 ( .A(ML_int_3__13_), .B(ML_int_3__5_), .S(n52), .Q(
        ML_int_4__13_) );
  MUX22 M1_3_10 ( .A(ML_int_3__10_), .B(ML_int_3__2_), .S(n52), .Q(
        ML_int_4__10_) );
  MUX22 M1_3_9 ( .A(ML_int_3__9_), .B(ML_int_3__1_), .S(n51), .Q(ML_int_4__9_)
         );
  MUX22 M1_3_8 ( .A(ML_int_3__8_), .B(ML_int_3__0_), .S(n51), .Q(ML_int_4__8_)
         );
  MUX22 M1_3_11 ( .A(ML_int_3__11_), .B(ML_int_3__3_), .S(n52), .Q(
        ML_int_4__11_) );
  MUX22 M1_2_5 ( .A(ML_int_2__5_), .B(ML_int_2__1_), .S(n45), .Q(ML_int_3__5_)
         );
  MUX22 M1_2_6 ( .A(ML_int_2__6_), .B(ML_int_2__2_), .S(n45), .Q(ML_int_3__6_)
         );
  MUX22 M1_2_16 ( .A(ML_int_2__16_), .B(ML_int_2__12_), .S(n47), .Q(
        ML_int_3__16_) );
  MUX22 M1_1_17 ( .A(ML_int_1__17_), .B(ML_int_1__15_), .S(n40), .Q(
        ML_int_2__17_) );
  MUX22 M1_2_14 ( .A(ML_int_2__14_), .B(ML_int_2__10_), .S(n46), .Q(
        ML_int_3__14_) );
  MUX22 M1_2_20 ( .A(ML_int_2__20_), .B(ML_int_2__16_), .S(n48), .Q(
        ML_int_3__20_) );
  MUX22 M1_2_12 ( .A(ML_int_2__12_), .B(ML_int_2__8_), .S(n46), .Q(
        ML_int_3__12_) );
  MUX22 M1_1_26 ( .A(ML_int_1__26_), .B(ML_int_1__24_), .S(n42), .Q(
        ML_int_2__26_) );
  MUX22 M1_2_21 ( .A(ML_int_2__21_), .B(ML_int_2__17_), .S(n48), .Q(
        ML_int_3__21_) );
  MUX22 M1_2_19 ( .A(ML_int_2__19_), .B(ML_int_2__15_), .S(n47), .Q(
        ML_int_3__19_) );
  MUX22 M1_2_18 ( .A(ML_int_2__18_), .B(ML_int_2__14_), .S(n47), .Q(
        ML_int_3__18_) );
  MUX22 M1_2_22 ( .A(ML_int_2__22_), .B(ML_int_2__18_), .S(n48), .Q(
        ML_int_3__22_) );
  MUX22 M1_2_13 ( .A(ML_int_2__13_), .B(ML_int_2__9_), .S(n46), .Q(
        ML_int_3__13_) );
  MUX22 M1_2_8 ( .A(ML_int_2__8_), .B(ML_int_2__4_), .S(n45), .Q(ML_int_3__8_)
         );
  MUX22 M1_2_11 ( .A(ML_int_2__11_), .B(ML_int_2__7_), .S(n46), .Q(
        ML_int_3__11_) );
  MUX22 M1_1_27 ( .A(ML_int_1__27_), .B(ML_int_1__25_), .S(n42), .Q(
        ML_int_2__27_) );
  MUX22 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n35), .Q(ML_int_1__24_) );
  MUX22 M1_1_14 ( .A(ML_int_1__14_), .B(ML_int_1__12_), .S(n42), .Q(
        ML_int_2__14_) );
  MUX22 M1_1_2 ( .A(ML_int_1__2_), .B(ML_int_1__0_), .S(n38), .Q(ML_int_2__2_)
         );
  MUX22 M1_1_25 ( .A(ML_int_1__25_), .B(ML_int_1__23_), .S(n42), .Q(
        ML_int_2__25_) );
  MUX22 M1_1_10 ( .A(ML_int_1__10_), .B(ML_int_1__8_), .S(n42), .Q(
        ML_int_2__10_) );
  MUX22 M1_1_11 ( .A(ML_int_1__11_), .B(ML_int_1__9_), .S(n43), .Q(
        ML_int_2__11_) );
  MUX22 M1_1_19 ( .A(ML_int_1__19_), .B(ML_int_1__17_), .S(n40), .Q(
        ML_int_2__19_) );
  MUX22 M1_1_21 ( .A(ML_int_1__21_), .B(ML_int_1__19_), .S(n41), .Q(
        ML_int_2__21_) );
  MUX22 M1_1_18 ( .A(ML_int_1__18_), .B(ML_int_1__16_), .S(n40), .Q(
        ML_int_2__18_) );
  MUX22 M1_1_22 ( .A(ML_int_1__22_), .B(ML_int_1__20_), .S(n41), .Q(
        ML_int_2__22_) );
  MUX22 M1_1_7 ( .A(ML_int_1__7_), .B(ML_int_1__5_), .S(n39), .Q(ML_int_2__7_)
         );
  MUX22 M1_1_6 ( .A(ML_int_1__6_), .B(ML_int_1__4_), .S(n39), .Q(ML_int_2__6_)
         );
  MUX22 M1_3_26 ( .A(ML_int_3__26_), .B(ML_int_3__18_), .S(n55), .Q(
        ML_int_4__26_) );
  MUX22 M1_4_26 ( .A(ML_int_4__26_), .B(ML_int_4__10_), .S(SH[4]), .Q(B[26])
         );
  MUX22 M1_4_22 ( .A(ML_int_4__22_), .B(ML_int_4__6_), .S(SH[4]), .Q(B[22]) );
  MUX22 M1_3_21 ( .A(ML_int_3__21_), .B(ML_int_3__13_), .S(n54), .Q(
        ML_int_4__21_) );
  MUX22 M1_4_21 ( .A(ML_int_4__21_), .B(ML_int_4__5_), .S(SH[4]), .Q(B[21]) );
  MUX22 M1_3_18 ( .A(ML_int_3__18_), .B(ML_int_3__10_), .S(n53), .Q(
        ML_int_4__18_) );
  MUX22 M1_4_18 ( .A(ML_int_4__18_), .B(ML_int_4__2_), .S(n56), .Q(B[18]) );
  MUX22 M1_3_17 ( .A(ML_int_3__17_), .B(ML_int_3__9_), .S(n53), .Q(
        ML_int_4__17_) );
  MUX22 M1_4_17 ( .A(ML_int_4__17_), .B(ML_int_4__1_), .S(n56), .Q(B[17]) );
  MUX22 M1_3_16 ( .A(ML_int_3__16_), .B(ML_int_3__8_), .S(n53), .Q(
        ML_int_4__16_) );
  MUX22 M1_4_16 ( .A(ML_int_4__16_), .B(ML_int_4__0_), .S(n56), .Q(B[16]) );
  MUX21 M1_4_27 ( .A(ML_int_4__27_), .B(ML_int_4__11_), .S(SH[4]), .Q(B[27])
         );
  MUX21 M1_2_25 ( .A(ML_int_2__25_), .B(ML_int_2__21_), .S(n49), .Q(
        ML_int_3__25_) );
  MUX21 M1_1_28 ( .A(ML_int_1__28_), .B(ML_int_1__26_), .S(n42), .Q(
        ML_int_2__28_) );
  MUX21 M1_3_20 ( .A(ML_int_3__20_), .B(ML_int_3__12_), .S(n54), .Q(
        ML_int_4__20_) );
  MUX21 M1_3_19 ( .A(ML_int_3__19_), .B(ML_int_3__11_), .S(n53), .Q(
        ML_int_4__19_) );
  MUX21 M1_2_26 ( .A(ML_int_2__26_), .B(ML_int_2__22_), .S(n49), .Q(
        ML_int_3__26_) );
  MUX21 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n37), .Q(ML_int_1__31_) );
  MUX21 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n37), .Q(ML_int_1__30_) );
  MUX21 M1_2_17 ( .A(ML_int_2__17_), .B(ML_int_2__13_), .S(n47), .Q(
        ML_int_3__17_) );
  MUX21 M1_1_16 ( .A(ML_int_1__16_), .B(ML_int_1__14_), .S(n40), .Q(
        ML_int_2__16_) );
  MUX21 M1_2_9 ( .A(ML_int_2__9_), .B(ML_int_2__5_), .S(n45), .Q(ML_int_3__9_)
         );
  MUX21 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n36), .Q(ML_int_1__16_) );
  MUX21 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n34), .Q(ML_int_1__12_) );
  MUX21 M1_1_12 ( .A(ML_int_1__12_), .B(ML_int_1__10_), .S(n41), .Q(
        ML_int_2__12_) );
  MUX21 M1_1_15 ( .A(ML_int_1__15_), .B(ML_int_1__13_), .S(n40), .Q(
        ML_int_2__15_) );
  MUX21 M1_1_24 ( .A(ML_int_1__24_), .B(ML_int_1__22_), .S(n41), .Q(
        ML_int_2__24_) );
  MUX21 M1_1_20 ( .A(ML_int_1__20_), .B(ML_int_1__18_), .S(n41), .Q(
        ML_int_2__20_) );
  MUX21 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n37), .Q(ML_int_1__15_) );
  MUX21 M1_1_13 ( .A(ML_int_1__13_), .B(ML_int_1__11_), .S(n41), .Q(
        ML_int_2__13_) );
  MUX21 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n32), .Q(ML_int_1__4_) );
  MUX21 M1_1_8 ( .A(ML_int_1__8_), .B(ML_int_1__6_), .S(n39), .Q(ML_int_2__8_)
         );
  MUX21 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n36), .Q(ML_int_1__25_) );
  MUX21 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n36), .Q(ML_int_1__26_) );
  MUX21 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n36), .Q(ML_int_1__27_) );
  MUX21 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n36), .Q(ML_int_1__29_) );
  MUX21 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n36), .Q(ML_int_1__28_) );
  MUX21 M1_2_7 ( .A(ML_int_2__7_), .B(ML_int_2__3_), .S(n45), .Q(ML_int_3__7_)
         );
  MUX21 M1_3_22 ( .A(ML_int_3__22_), .B(ML_int_3__14_), .S(n54), .Q(
        ML_int_4__22_) );
  MUX22 M1_2_24 ( .A(ML_int_2__24_), .B(ML_int_2__20_), .S(n48), .Q(
        ML_int_3__24_) );
  MUX22 M1_1_9 ( .A(ML_int_1__9_), .B(ML_int_1__7_), .S(n39), .Q(ML_int_2__9_)
         );
  MUX22 M1_2_15 ( .A(ML_int_2__15_), .B(ML_int_2__11_), .S(n47), .Q(
        ML_int_3__15_) );
  MUX22 M1_2_10 ( .A(ML_int_2__10_), .B(ML_int_2__6_), .S(n46), .Q(
        ML_int_3__10_) );
  MUX22 M1_4_23 ( .A(ML_int_4__23_), .B(ML_int_4__7_), .S(SH[4]), .Q(B[23]) );
  MUX22 M1_3_24 ( .A(ML_int_3__24_), .B(ML_int_3__16_), .S(n54), .Q(
        ML_int_4__24_) );
  MUX21 M1_1_5 ( .A(ML_int_1__5_), .B(ML_int_1__3_), .S(n39), .Q(ML_int_2__5_)
         );
  MUX22 M1_1_23 ( .A(ML_int_1__23_), .B(ML_int_1__21_), .S(n41), .Q(
        ML_int_2__23_) );
  MUX22 M1_2_23 ( .A(ML_int_2__23_), .B(ML_int_2__19_), .S(n48), .Q(
        ML_int_3__23_) );
  MUX21 M1_2_4 ( .A(ML_int_2__4_), .B(ML_int_2__0_), .S(n44), .Q(ML_int_3__4_)
         );
  MUX22 M1_3_27 ( .A(ML_int_3__27_), .B(ML_int_3__19_), .S(n55), .Q(
        ML_int_4__27_) );
  MUX22 M1_1_4 ( .A(ML_int_1__4_), .B(ML_int_1__2_), .S(n38), .Q(ML_int_2__4_)
         );
  MUX22 M1_3_15 ( .A(ML_int_3__15_), .B(ML_int_3__7_), .S(n53), .Q(
        ML_int_4__15_) );
  MUX21 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n35), .Q(ML_int_1__17_) );
  MUX21 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n34), .Q(ML_int_1__14_) );
  MUX21 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n33), .Q(ML_int_1__7_) );
  NOR21 U3 ( .A(n38), .B(n29), .Q(ML_int_2__1_) );
  INV2 U4 ( .A(ML_int_1__1_), .Q(n29) );
  CLKIN1 U5 ( .A(ML_int_3__6_), .Q(n18) );
  INV2 U6 ( .A(ML_int_2__0_), .Q(n28) );
  INV2 U7 ( .A(ML_int_3__0_), .Q(n24) );
  INV2 U8 ( .A(ML_int_1__0_), .Q(n30) );
  CLKIN0 U9 ( .A(ML_int_3__3_), .Q(n21) );
  INV2 U10 ( .A(ML_int_3__1_), .Q(n23) );
  CLKIN1 U11 ( .A(ML_int_4__6_), .Q(n10) );
  CLKIN1 U12 ( .A(ML_int_4__2_), .Q(n14) );
  INV1 U13 ( .A(ML_int_4__1_), .Q(n15) );
  INV1 U14 ( .A(ML_int_2__1_), .Q(n27) );
  INV2 U15 ( .A(ML_int_4__0_), .Q(n16) );
  CLKIN0 U16 ( .A(ML_int_3__5_), .Q(n19) );
  CLKIN1 U17 ( .A(ML_int_2__2_), .Q(n26) );
  CLKIN1 U18 ( .A(ML_int_3__2_), .Q(n22) );
  CLKIN0 U19 ( .A(ML_int_4__14_), .Q(n2) );
  CLKIN1 U20 ( .A(ML_int_4__3_), .Q(n13) );
  CLKIN2 U21 ( .A(ML_int_4__4_), .Q(n12) );
  CLKIN3 U22 ( .A(ML_int_4__7_), .Q(n9) );
  CLKIN2 U23 ( .A(ML_int_4__9_), .Q(n7) );
  CLKIN1 U24 ( .A(ML_int_4__5_), .Q(n11) );
  CLKIN2 U25 ( .A(ML_int_4__8_), .Q(n8) );
  INV3 U26 ( .A(ML_int_4__11_), .Q(n5) );
  INV3 U27 ( .A(ML_int_4__13_), .Q(n3) );
  NOR21 U28 ( .A(n56), .B(n5), .Q(B[11]) );
  NOR21 U29 ( .A(n32), .B(n31), .Q(ML_int_1__0_) );
  INV3 U30 ( .A(A[0]), .Q(n31) );
  NOR21 U31 ( .A(n38), .B(n30), .Q(ML_int_2__0_) );
  NOR21 U32 ( .A(n51), .B(n19), .Q(ML_int_4__5_) );
  NOR21 U33 ( .A(n51), .B(n18), .Q(ML_int_4__6_) );
  NOR21 U34 ( .A(n44), .B(n25), .Q(ML_int_3__3_) );
  INV3 U35 ( .A(ML_int_2__3_), .Q(n25) );
  NOR21 U36 ( .A(n44), .B(n27), .Q(ML_int_3__1_) );
  NOR21 U37 ( .A(n44), .B(n26), .Q(ML_int_3__2_) );
  NOR21 U38 ( .A(n50), .B(n23), .Q(ML_int_4__1_) );
  NOR21 U39 ( .A(n50), .B(n22), .Q(ML_int_4__2_) );
  NOR21 U40 ( .A(n50), .B(n21), .Q(ML_int_4__3_) );
  NOR21 U41 ( .A(n50), .B(n20), .Q(ML_int_4__4_) );
  INV3 U42 ( .A(ML_int_3__4_), .Q(n20) );
  NOR21 U43 ( .A(n56), .B(n3), .Q(B[13]) );
  NOR21 U44 ( .A(n56), .B(n9), .Q(B[7]) );
  NOR21 U45 ( .A(n56), .B(n8), .Q(B[8]) );
  NOR21 U46 ( .A(n56), .B(n7), .Q(B[9]) );
  NOR21 U47 ( .A(n56), .B(n6), .Q(B[10]) );
  INV3 U48 ( .A(ML_int_4__10_), .Q(n6) );
  NOR21 U49 ( .A(n56), .B(n4), .Q(B[12]) );
  INV3 U50 ( .A(ML_int_4__12_), .Q(n4) );
  NOR21 U51 ( .A(n56), .B(n2), .Q(B[14]) );
  NOR21 U52 ( .A(n56), .B(n1), .Q(B[15]) );
  INV3 U53 ( .A(ML_int_4__15_), .Q(n1) );
  NOR21 U54 ( .A(n56), .B(n10), .Q(B[6]) );
  NOR21 U55 ( .A(n51), .B(n17), .Q(ML_int_4__7_) );
  INV3 U56 ( .A(ML_int_3__7_), .Q(n17) );
  NOR21 U57 ( .A(n56), .B(n15), .Q(B[1]) );
  NOR21 U58 ( .A(n56), .B(n14), .Q(B[2]) );
  NOR21 U59 ( .A(n56), .B(n13), .Q(B[3]) );
  NOR21 U60 ( .A(n56), .B(n12), .Q(B[4]) );
  NOR21 U61 ( .A(n56), .B(n11), .Q(B[5]) );
  NOR21 U62 ( .A(n50), .B(n24), .Q(ML_int_4__0_) );
  NOR21 U63 ( .A(n56), .B(n16), .Q(B[0]) );
  NOR21 U64 ( .A(n44), .B(n28), .Q(ML_int_3__0_) );
  BUF2 U65 ( .A(SH[0]), .Q(n32) );
  BUF2 U66 ( .A(SH[0]), .Q(n34) );
  BUF2 U67 ( .A(SH[0]), .Q(n35) );
  BUF2 U68 ( .A(SH[0]), .Q(n33) );
  BUF2 U69 ( .A(SH[3]), .Q(n52) );
  BUF2 U70 ( .A(SH[3]), .Q(n53) );
  BUF2 U71 ( .A(SH[3]), .Q(n54) );
  BUF2 U72 ( .A(SH[3]), .Q(n55) );
  BUF2 U73 ( .A(SH[0]), .Q(n36) );
  BUF2 U74 ( .A(SH[1]), .Q(n41) );
  BUF2 U75 ( .A(SH[1]), .Q(n40) );
  BUF2 U76 ( .A(SH[1]), .Q(n42) );
  BUF2 U77 ( .A(SH[2]), .Q(n46) );
  BUF2 U78 ( .A(SH[2]), .Q(n47) );
  BUF2 U79 ( .A(SH[2]), .Q(n49) );
  BUF2 U80 ( .A(SH[2]), .Q(n48) );
  BUF2 U81 ( .A(SH[1]), .Q(n38) );
  BUF2 U82 ( .A(SH[3]), .Q(n51) );
  BUF2 U83 ( .A(SH[2]), .Q(n44) );
  BUF2 U84 ( .A(SH[3]), .Q(n50) );
  BUF2 U85 ( .A(SH[2]), .Q(n45) );
  BUF2 U86 ( .A(SH[1]), .Q(n39) );
  BUF2 U87 ( .A(SH[0]), .Q(n37) );
  BUF2 U88 ( .A(SH[1]), .Q(n43) );
  BUF2 U89 ( .A(SH[4]), .Q(n56) );
endmodule


module E_alu ( o_data_AluRes, i_data_A, i_data_B, i_con_AluCtrl, i_data_shamt
 );
  output [31:0] o_data_AluRes;
  input [31:0] i_data_A;
  input [31:0] i_data_B;
  input [3:0] i_con_AluCtrl;
  input [4:0] i_data_shamt;
  wire   N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159,
         N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N244, N245, N246,
         N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257,
         N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, N270, N271, N272, N273, N274, N275, N276, n13, n96, n97, n98,
         n99, n111, n118, n125, n129, n130, n131, n132, n136, n137, n138, n139,
         n143, n144, n145, n146, n153, n162, n166, n167, n168, n169, n176,
         n183, n190, n197, n204, n211, n218, n225, n232, n239, n243, n244,
         n245, n246, n253, n260, n267, n274, n281, n288, n295, n302, n309,
         n316, n328, n329, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n112,
         n113, n114, n115, n116, n117, n119, n120, n121, n122, n123, n124,
         n126, n127, n128, n133, n134, n135, n140, n141, n142, n147, n148,
         n149, n150, n151, n152, n154, n155, n156, n157, n158, n159, n160,
         n161, n163, n164, n165, n170, n171, n172, n173, n174, n175, n177,
         n178, n179, n180, n181, n182, n184, n185, n186, n187, n188, n189,
         n191, n192, n193, n194, n195, n196, n198, n199, n200, n201, n202,
         n203, n205, n206, n207, n208, n209, n210, n212, n213, n214, n215,
         n216, n217, n219, n220, n221, n222, n223, n224, n226, n227, n228,
         n229, n230, n231, n233, n234, n235, n236, n237, n238, n240, n241,
         n242, n247, n248, n249, n250, n251, n252, n254, n255, n256, n257,
         n258, n259, n261, n262, n263, n264, n265, n266, n268, n269, n270,
         n271, n272, n273, n275, n276, n277, n278, n279, n280, n282, n283,
         n284, n285, n286, n287, n289, n290, n291, n292, n293, n294, n296,
         n297, n298, n299, n300, n301, n303, n304, n305, n306, n307, n308,
         n310, n311, n312, n313, n314, n315, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n330, n331, n332, n333, n334,
         n335;

  OAI222 U88 ( .A(n34), .B(n333), .C(i_data_A[2]), .D(n99), .Q(n167) );
  E_alu_DW01_add_1 add_53 ( .A(i_data_A), .B({i_data_B[31:30], n18, 
        i_data_B[28:0]}), .CI(n13), .SUM({N147, N146, N145, N144, N143, N142, 
        N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, 
        N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, 
        N117, N116}) );
  E_alu_DW01_sub_1 sub_62 ( .A(i_data_A), .B({i_data_B[31:30], n18, 
        i_data_B[28:0]}), .CI(n13), .DIFF({N275, N274, N273, N272, N271, N270, 
        N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, 
        N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, 
        N245, N244}) );
  E_alu_DW01_cmp2_1 r65 ( .A(i_data_A), .B({i_data_B[31:30], n18, 
        i_data_B[28:7], n37, i_data_B[5:0]}), .LEQ(n13), .TC(n13), .LT_LE(N276) );
  E_alu_DW_rash_1 r63 ( .A({i_data_B[31:30], n18, i_data_B[28:7], n37, 
        i_data_B[5:0]}), .DATA_TC(n13), .SH(i_data_shamt), .SH_TC(n13), .B({
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, 
        N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, 
        N187, N186, N185, N184, N183, N182, N181, N180}) );
  E_alu_DW01_ash_1 sll_56 ( .A({i_data_B[31:30], n18, i_data_B[28:7], n37, 
        i_data_B[5:0]}), .DATA_TC(n13), .SH(i_data_shamt), .SH_TC(n13), .B({
        N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, 
        N155, N154, N153, N152, N151, N150, N149, N148}) );
  OAI2110 U2 ( .A(i_data_A[6]), .B(n34), .C(n125), .D(n43), .Q(n115) );
  NAND22 U3 ( .A(N154), .B(n1), .Q(n119) );
  INV0 U4 ( .A(i_data_B[7]), .Q(n249) );
  AOI222 U5 ( .A(N273), .B(n2), .C(N145), .D(n21), .Q(n299) );
  INV6 U6 ( .A(n55), .Q(n34) );
  INV6 U7 ( .A(n96), .Q(n55) );
  AOI222 U8 ( .A(N123), .B(n21), .C(N155), .D(n1), .Q(n133) );
  BUF6 U9 ( .A(n98), .Q(n3) );
  NAND22 U10 ( .A(i_con_AluCtrl[0]), .B(n58), .Q(n96) );
  NAND22 U11 ( .A(N207), .B(n40), .Q(n283) );
  IMUX30 U12 ( .A(n305), .B(n51), .C(n203), .S0(i_data_A[17]), .S1(
        i_data_B[17]), .Q(n205) );
  IMUX30 U13 ( .A(n305), .B(n51), .C(n264), .S0(i_data_A[25]), .S1(
        i_data_B[25]), .Q(n265) );
  IMUX30 U14 ( .A(n99), .B(n34), .C(n76), .S0(i_data_A[0]), .S1(i_data_B[0]), 
        .Q(n77) );
  IMUX30 U15 ( .A(n305), .B(n51), .C(n224), .S0(i_data_A[20]), .S1(
        i_data_B[20]), .Q(n226) );
  INV6 U16 ( .A(n71), .Q(n21) );
  BUF8 U17 ( .A(n319), .Q(n2) );
  BUF8 U18 ( .A(n20), .Q(n1) );
  AOI211 U19 ( .A(i_data_A[19]), .B(n47), .C(n219), .Q(n221) );
  NOR21 U20 ( .A(n329), .B(i_con_AluCtrl[1]), .Q(n98) );
  INV3 U21 ( .A(i_con_AluCtrl[0]), .Q(n17) );
  NAND21 U22 ( .A(n72), .B(i_con_AluCtrl[0]), .Q(n61) );
  NAND42 U23 ( .A(n236), .B(n235), .C(n234), .D(n233), .Q(o_data_AluRes[21])
         );
  BUF6 U24 ( .A(n318), .Q(n40) );
  AOI221 U25 ( .A(N170), .B(n1), .C(N266), .D(n2), .Q(n241) );
  INV3 U26 ( .A(n67), .Q(n20) );
  INV3 U27 ( .A(n73), .Q(n319) );
  INV6 U28 ( .A(n19), .Q(n4) );
  INV6 U29 ( .A(n19), .Q(n5) );
  NAND23 U30 ( .A(n58), .B(n17), .Q(n99) );
  INV3 U31 ( .A(i_con_AluCtrl[2]), .Q(n56) );
  NAND22 U32 ( .A(N187), .B(n41), .Q(n128) );
  AOI211 U33 ( .A(n53), .B(n122), .C(n121), .Q(n123) );
  NAND22 U34 ( .A(n205), .B(n208), .Q(n8) );
  AOI221 U35 ( .A(i_data_A[15]), .B(n48), .C(N131), .D(n21), .Q(n193) );
  NAND31 U36 ( .A(n271), .B(n270), .C(n269), .Q(o_data_AluRes[25]) );
  AOI221 U37 ( .A(N141), .B(n21), .C(N269), .D(n2), .Q(n271) );
  INV3 U38 ( .A(i_con_AluCtrl[3]), .Q(n196) );
  IMUX30 U39 ( .A(n305), .B(n51), .C(n256), .S0(i_data_A[24]), .S1(
        i_data_B[24]), .Q(n257) );
  AOI221 U40 ( .A(i_data_A[9]), .B(n48), .C(N125), .D(n21), .Q(n149) );
  NAND42 U41 ( .A(n303), .B(n301), .C(n300), .D(n299), .Q(o_data_AluRes[29])
         );
  INV3 U42 ( .A(n15), .Q(n16) );
  INV3 U43 ( .A(n6), .Q(n7) );
  NAND41 U44 ( .A(n202), .B(n201), .C(n200), .D(n199), .Q(o_data_AluRes[16])
         );
  NAND31 U45 ( .A(n206), .B(n207), .C(n9), .Q(o_data_AluRes[17]) );
  INV3 U46 ( .A(n8), .Q(n9) );
  AOI221 U47 ( .A(i_data_A[18]), .B(n47), .C(N134), .D(n21), .Q(n212) );
  NAND22 U48 ( .A(N271), .B(n2), .Q(n287) );
  INV3 U49 ( .A(n11), .Q(n12) );
  NAND31 U50 ( .A(n294), .B(n296), .C(n33), .Q(o_data_AluRes[28]) );
  NAND41 U51 ( .A(n142), .B(n141), .C(n140), .D(n135), .Q(o_data_AluRes[8]) );
  AOI221 U52 ( .A(i_data_A[23]), .B(n47), .C(N139), .D(n21), .Q(n255) );
  NAND41 U53 ( .A(n174), .B(n173), .C(n172), .D(n171), .Q(o_data_AluRes[12])
         );
  NAND22 U54 ( .A(N256), .B(n2), .Q(n173) );
  NAND23 U55 ( .A(n241), .B(n242), .Q(n15) );
  INV0 U56 ( .A(i_data_A[3]), .Q(n94) );
  NAND33 U57 ( .A(i_con_AluCtrl[0]), .B(n70), .C(n68), .Q(n335) );
  INV6 U58 ( .A(n99), .Q(n305) );
  NAND31 U59 ( .A(i_con_AluCtrl[1]), .B(i_con_AluCtrl[0]), .C(n70), .Q(n67) );
  NAND31 U60 ( .A(i_con_AluCtrl[1]), .B(n70), .C(n17), .Q(n71) );
  INV3 U61 ( .A(n98), .Q(n19) );
  CLKIN3 U62 ( .A(n55), .Q(n35) );
  OAI2111 U63 ( .A(i_data_A[30]), .B(n50), .C(n162), .D(n43), .Q(n304) );
  IMUX30 U64 ( .A(n305), .B(n51), .C(n304), .S0(i_data_A[30]), .S1(
        i_data_B[30]), .Q(n306) );
  CLKIN3 U65 ( .A(i_data_B[2]), .Q(n332) );
  AOI211 U66 ( .A(i_data_A[7]), .B(n48), .C(n124), .Q(n127) );
  NAND20 U67 ( .A(i_data_A[22]), .B(n5), .Q(n225) );
  NAND21 U68 ( .A(i_data_A[20]), .B(n4), .Q(n239) );
  BUF6 U69 ( .A(n55), .Q(n51) );
  AOI221 U70 ( .A(N135), .B(n21), .C(N167), .D(n1), .Q(n223) );
  AOI211 U71 ( .A(N120), .B(n21), .C(n105), .Q(n106) );
  NAND33 U72 ( .A(n127), .B(n133), .C(n128), .Q(n6) );
  NAND22 U73 ( .A(n126), .B(n7), .Q(o_data_AluRes[7]) );
  AOI221 U74 ( .A(i_data_B[1]), .B(n42), .C(N197), .D(n40), .Q(n208) );
  MUX22 U75 ( .A(n305), .B(n51), .S(i_data_A[27]), .Q(n10) );
  IMUX21 U76 ( .A(n10), .B(n282), .S(i_data_B[27]), .Q(n290) );
  NAND22 U77 ( .A(n290), .B(n289), .Q(n11) );
  NAND33 U78 ( .A(n291), .B(n287), .C(n12), .Q(o_data_AluRes[27]) );
  AOI211 U79 ( .A(N175), .B(n1), .C(n286), .Q(n289) );
  MUX22 U80 ( .A(n305), .B(n52), .S(i_data_A[6]), .Q(n14) );
  IMUX21 U81 ( .A(n14), .B(n115), .S(n37), .Q(n116) );
  CLKIN12 U82 ( .A(n36), .Q(n37) );
  NAND33 U83 ( .A(n240), .B(n238), .C(n16), .Q(o_data_AluRes[22]) );
  AOI220 U84 ( .A(i_data_A[22]), .B(n47), .C(N138), .D(n21), .Q(n240) );
  IMUX31 U85 ( .A(n305), .B(n51), .C(n215), .S0(i_data_A[19]), .S1(
        i_data_B[19]), .Q(n216) );
  OAI2111 U86 ( .A(i_data_A[24]), .B(n50), .C(n211), .D(n43), .Q(n256) );
  INV6 U87 ( .A(n49), .Q(n43) );
  NAND31 U89 ( .A(n117), .B(n116), .C(n119), .Q(n30) );
  NAND20 U90 ( .A(i_data_A[16]), .B(n4), .Q(n274) );
  NAND21 U91 ( .A(i_con_AluCtrl[2]), .B(n196), .Q(n60) );
  INV0 U92 ( .A(i_data_A[30]), .Q(n307) );
  AOI221 U93 ( .A(i_data_A[10]), .B(n48), .C(N126), .D(n21), .Q(n155) );
  NAND22 U94 ( .A(n288), .B(n44), .Q(n181) );
  CLKIN6 U95 ( .A(n49), .Q(n44) );
  OAI2111 U96 ( .A(i_data_A[26]), .B(n50), .C(n197), .D(n43), .Q(n272) );
  AOI211 U97 ( .A(i_data_A[24]), .B(n47), .C(n259), .Q(n261) );
  NAND22 U98 ( .A(N153), .B(n1), .Q(n113) );
  INV10 U99 ( .A(i_con_AluCtrl[1]), .Q(n68) );
  OAI2110 U100 ( .A(i_data_A[1]), .B(n35), .C(n45), .D(n246), .Q(n245) );
  OAI220 U101 ( .A(n34), .B(n83), .C(i_data_A[1]), .D(n99), .Q(n244) );
  NAND20 U102 ( .A(i_data_A[1]), .B(n4), .Q(n246) );
  BUF12 U103 ( .A(i_data_B[29]), .Q(n18) );
  AOI221 U104 ( .A(N186), .B(n41), .C(i_data_A[6]), .D(n46), .Q(n117) );
  AOI221 U105 ( .A(i_data_A[27]), .B(n46), .C(N143), .D(n21), .Q(n291) );
  AOI221 U106 ( .A(i_data_A[28]), .B(n46), .C(N144), .D(n21), .Q(n294) );
  AOI222 U107 ( .A(N258), .B(n2), .C(N162), .D(n1), .Q(n189) );
  NAND20 U108 ( .A(n3), .B(i_data_A[31]), .Q(n153) );
  NAND20 U109 ( .A(i_data_A[3]), .B(n5), .Q(n146) );
  NAND20 U110 ( .A(i_data_A[4]), .B(n3), .Q(n139) );
  NAND20 U111 ( .A(i_data_A[27]), .B(n4), .Q(n190) );
  NAND20 U112 ( .A(i_data_A[28]), .B(n3), .Q(n183) );
  NAND20 U113 ( .A(i_data_A[26]), .B(n5), .Q(n197) );
  NAND20 U114 ( .A(i_data_A[24]), .B(n5), .Q(n211) );
  NAND20 U115 ( .A(i_data_A[30]), .B(n3), .Q(n162) );
  CLKIN4 U116 ( .A(i_data_B[6]), .Q(n36) );
  OAI2111 U117 ( .A(i_data_A[11]), .B(n50), .C(n309), .D(n43), .Q(n158) );
  NAND22 U118 ( .A(n79), .B(n80), .Q(n22) );
  NAND32 U119 ( .A(n81), .B(n78), .C(n23), .Q(o_data_AluRes[0]) );
  INV3 U120 ( .A(n22), .Q(n23) );
  AOI212 U121 ( .A(N276), .B(n66), .C(n65), .Q(n81) );
  NAND31 U122 ( .A(n129), .B(n113), .C(n114), .Q(n24) );
  NAND22 U123 ( .A(n112), .B(n25), .Q(o_data_AluRes[5]) );
  INV3 U124 ( .A(n24), .Q(n25) );
  NOR21 U125 ( .A(n26), .B(n71), .Q(n27) );
  NOR21 U126 ( .A(n27), .B(n110), .Q(n112) );
  INV3 U127 ( .A(N121), .Q(n26) );
  OAI211 U128 ( .A(n335), .B(n330), .C(n109), .Q(n110) );
  NAND31 U129 ( .A(n322), .B(n324), .C(n325), .Q(n28) );
  NAND22 U130 ( .A(n323), .B(n29), .Q(o_data_AluRes[31]) );
  INV3 U131 ( .A(n28), .Q(n29) );
  AOI210 U132 ( .A(n326), .B(i_data_B[31]), .C(n321), .Q(n322) );
  NOR20 U133 ( .A(i_data_B[31]), .B(i_data_A[31]), .Q(n320) );
  NAND22 U134 ( .A(n120), .B(n31), .Q(o_data_AluRes[6]) );
  CLKIN3 U135 ( .A(n30), .Q(n31) );
  INV0 U136 ( .A(i_data_A[0]), .Q(n75) );
  NAND42 U137 ( .A(n195), .B(n194), .C(n193), .D(n192), .Q(o_data_AluRes[15])
         );
  NAND22 U138 ( .A(n293), .B(n297), .Q(n32) );
  INV3 U139 ( .A(n32), .Q(n33) );
  CLKIN3 U140 ( .A(n55), .Q(n50) );
  AOI222 U141 ( .A(N142), .B(n21), .C(N174), .D(n1), .Q(n280) );
  OAI2111 U142 ( .A(n44), .B(n161), .C(n160), .D(n159), .Q(n163) );
  OAI211 U143 ( .A(n44), .B(n307), .C(n306), .Q(n312) );
  OAI210 U144 ( .A(n44), .B(n104), .C(n103), .Q(n105) );
  OAI210 U145 ( .A(n44), .B(n83), .C(n82), .Q(n84) );
  OAI210 U146 ( .A(n44), .B(n333), .C(n88), .Q(n89) );
  OAI210 U147 ( .A(n44), .B(n94), .C(n93), .Q(n95) );
  CLKIN2 U148 ( .A(n329), .Q(n70) );
  AOI221 U149 ( .A(i_data_A[17]), .B(n47), .C(N133), .D(n21), .Q(n206) );
  AOI220 U150 ( .A(N173), .B(n1), .C(N205), .D(n41), .Q(n270) );
  AOI220 U151 ( .A(i_data_B[14]), .B(n42), .C(N210), .D(n40), .Q(n310) );
  CLKIN3 U152 ( .A(n63), .Q(n315) );
  AOI210 U153 ( .A(N117), .B(n21), .C(n84), .Q(n85) );
  AOI210 U154 ( .A(N119), .B(n21), .C(n95), .Q(n100) );
  IMUX30 U155 ( .A(n305), .B(n52), .C(n158), .S0(i_data_A[11]), .S1(
        i_data_B[11]), .Q(n160) );
  IMUX30 U156 ( .A(n305), .B(n53), .C(n247), .S0(i_data_A[23]), .S1(
        i_data_B[23]), .Q(n254) );
  NAND20 U157 ( .A(N178), .B(n1), .Q(n308) );
  NAND22 U158 ( .A(N255), .B(n2), .Q(n165) );
  AOI211 U159 ( .A(n53), .B(n75), .C(n74), .Q(n76) );
  OAI2110 U160 ( .A(i_data_A[19]), .B(n50), .C(n253), .D(n44), .Q(n215) );
  AOI220 U161 ( .A(i_data_A[16]), .B(n48), .C(N132), .D(n21), .Q(n200) );
  AOI221 U162 ( .A(n137), .B(n331), .C(i_data_B[4]), .D(n138), .Q(n136) );
  CLKIN3 U163 ( .A(n69), .Q(n318) );
  AOI210 U164 ( .A(N118), .B(n21), .C(n89), .Q(n90) );
  INV0 U165 ( .A(i_data_B[4]), .Q(n331) );
  AOI220 U166 ( .A(N188), .B(n40), .C(N156), .D(n1), .Q(n142) );
  AOI220 U167 ( .A(N189), .B(n41), .C(N157), .D(n1), .Q(n151) );
  AOI220 U168 ( .A(N195), .B(n40), .C(N163), .D(n1), .Q(n195) );
  AOI220 U169 ( .A(N176), .B(n1), .C(N272), .D(n2), .Q(n296) );
  AOI220 U170 ( .A(i_data_B[12]), .B(n42), .C(N208), .D(n40), .Q(n297) );
  NAND20 U171 ( .A(i_data_A[21]), .B(n5), .Q(n232) );
  NAND20 U172 ( .A(i_data_A[8]), .B(n4), .Q(n111) );
  NAND20 U173 ( .A(i_data_A[15]), .B(n5), .Q(n281) );
  NAND20 U174 ( .A(i_data_A[12]), .B(n4), .Q(n302) );
  NAND20 U175 ( .A(i_data_A[11]), .B(n3), .Q(n309) );
  AOI220 U176 ( .A(N177), .B(n1), .C(N209), .D(n41), .Q(n303) );
  AOI220 U177 ( .A(N148), .B(n1), .C(N180), .D(n40), .Q(n80) );
  AOI220 U178 ( .A(N116), .B(n21), .C(N244), .D(n2), .Q(n79) );
  AOI220 U179 ( .A(i_data_B[15]), .B(n42), .C(n315), .D(n52), .Q(n325) );
  AOI220 U180 ( .A(N211), .B(n41), .C(N179), .D(n1), .Q(n324) );
  OAI2110 U181 ( .A(i_data_A[23]), .B(n34), .C(n218), .D(n44), .Q(n247) );
  NAND20 U182 ( .A(i_data_A[23]), .B(n4), .Q(n218) );
  NAND20 U183 ( .A(i_data_A[13]), .B(n5), .Q(n295) );
  NAND20 U184 ( .A(i_data_A[6]), .B(n3), .Q(n125) );
  AOI220 U185 ( .A(N190), .B(n40), .C(N158), .D(n1), .Q(n157) );
  AOI220 U186 ( .A(N192), .B(n41), .C(N160), .D(n1), .Q(n174) );
  AOI210 U187 ( .A(N171), .B(n1), .C(n250), .Q(n252) );
  AOI220 U188 ( .A(N172), .B(n1), .C(N204), .D(n40), .Q(n262) );
  NAND20 U189 ( .A(i_data_A[0]), .B(n3), .Q(n328) );
  NAND20 U190 ( .A(i_data_A[14]), .B(n3), .Q(n288) );
  NAND20 U191 ( .A(i_data_A[7]), .B(n3), .Q(n118) );
  OAI2110 U192 ( .A(i_data_A[20]), .B(n50), .C(n239), .D(n335), .Q(n224) );
  AOI220 U193 ( .A(N129), .B(n21), .C(N193), .D(n40), .Q(n180) );
  NAND20 U194 ( .A(n5), .B(i_data_A[9]), .Q(n97) );
  BUF6 U195 ( .A(n317), .Q(n42) );
  OAI2110 U196 ( .A(i_data_A[17]), .B(n35), .C(n267), .D(n44), .Q(n203) );
  NAND20 U197 ( .A(i_data_A[17]), .B(n3), .Q(n267) );
  OAI2110 U198 ( .A(i_data_A[2]), .B(n35), .C(n45), .D(n169), .Q(n168) );
  OAI2110 U199 ( .A(i_data_A[10]), .B(n34), .C(n316), .D(n43), .Q(n152) );
  NAND20 U200 ( .A(i_data_A[10]), .B(n3), .Q(n316) );
  INV2 U201 ( .A(n153), .Q(n326) );
  NAND20 U202 ( .A(i_data_A[2]), .B(n4), .Q(n169) );
  NAND20 U203 ( .A(i_data_A[5]), .B(n4), .Q(n132) );
  IMUX20 U204 ( .A(n43), .B(n99), .S(n320), .Q(n321) );
  INV0 U205 ( .A(i_data_A[5]), .Q(n330) );
  BUF2 U206 ( .A(n318), .Q(n41) );
  INV3 U207 ( .A(n49), .Q(n45) );
  BUF2 U208 ( .A(n49), .Q(n47) );
  BUF2 U209 ( .A(n49), .Q(n46) );
  BUF2 U210 ( .A(n49), .Q(n48) );
  BUF2 U211 ( .A(n54), .Q(n52) );
  BUF2 U212 ( .A(n54), .Q(n53) );
  NAND31 U213 ( .A(i_con_AluCtrl[1]), .B(n72), .C(n17), .Q(n73) );
  NAND41 U214 ( .A(n166), .B(n92), .C(n91), .D(n90), .Q(o_data_AluRes[2]) );
  NAND41 U215 ( .A(n143), .B(n102), .C(n101), .D(n100), .Q(o_data_AluRes[3])
         );
  NAND41 U216 ( .A(n136), .B(n108), .C(n107), .D(n106), .Q(o_data_AluRes[4])
         );
  NAND41 U217 ( .A(n243), .B(n87), .C(n86), .D(n85), .Q(o_data_AluRes[1]) );
  AOI221 U218 ( .A(N250), .B(n2), .C(N122), .D(n21), .Q(n120) );
  NOR31 U219 ( .A(n64), .B(n63), .C(n62), .Q(n65) );
  INV3 U220 ( .A(n57), .Q(n58) );
  NAND31 U221 ( .A(i_con_AluCtrl[2]), .B(i_con_AluCtrl[3]), .C(n68), .Q(n57)
         );
  NAND22 U222 ( .A(n196), .B(n56), .Q(n329) );
  AOI2111 U223 ( .A(N274), .B(n2), .C(n312), .D(n311), .Q(n314) );
  INV3 U224 ( .A(n335), .Q(n49) );
  INV3 U225 ( .A(n96), .Q(n54) );
  INV3 U226 ( .A(i_data_B[5]), .Q(n327) );
  IMUX30 U227 ( .A(n99), .B(n34), .C(n184), .S0(i_data_A[14]), .S1(
        i_data_B[14]), .Q(n185) );
  AOI211 U228 ( .A(n53), .B(n182), .C(n181), .Q(n184) );
  NAND41 U229 ( .A(n212), .B(n213), .C(n214), .D(n210), .Q(o_data_AluRes[18])
         );
  AOI211 U230 ( .A(i_data_A[14]), .B(n48), .C(n185), .Q(n187) );
  NAND41 U231 ( .A(n151), .B(n150), .C(n149), .D(n148), .Q(o_data_AluRes[9])
         );
  AOI221 U232 ( .A(n144), .B(n217), .C(i_data_B[3]), .D(n145), .Q(n143) );
  AOI221 U233 ( .A(n244), .B(n334), .C(i_data_B[1]), .D(n245), .Q(n243) );
  INV3 U234 ( .A(i_data_B[1]), .Q(n334) );
  AOI221 U235 ( .A(N159), .B(n1), .C(N191), .D(n40), .Q(n159) );
  AOI221 U236 ( .A(N164), .B(n1), .C(N260), .D(n2), .Q(n201) );
  AOI221 U237 ( .A(N165), .B(n1), .C(N261), .D(n2), .Q(n207) );
  AOI221 U238 ( .A(N166), .B(n1), .C(N262), .D(n2), .Q(n213) );
  AOI221 U239 ( .A(N169), .B(n1), .C(N265), .D(n2), .Q(n235) );
  AOI221 U240 ( .A(N275), .B(n2), .C(N147), .D(n21), .Q(n323) );
  IMUX30 U241 ( .A(n305), .B(n51), .C(n272), .S0(i_data_A[26]), .S1(
        i_data_B[26]), .Q(n273) );
  NAND31 U242 ( .A(n230), .B(n229), .C(n228), .Q(o_data_AluRes[20]) );
  AOI221 U243 ( .A(N168), .B(n1), .C(N200), .D(n40), .Q(n229) );
  AOI211 U244 ( .A(i_data_A[20]), .B(n47), .C(n227), .Q(n228) );
  AOI221 U245 ( .A(N264), .B(n2), .C(N136), .D(n21), .Q(n230) );
  NAND31 U246 ( .A(n263), .B(n262), .C(n261), .Q(o_data_AluRes[24]) );
  AOI221 U247 ( .A(N268), .B(n2), .C(N140), .D(n21), .Q(n263) );
  NAND31 U248 ( .A(n180), .B(n178), .C(n39), .Q(o_data_AluRes[13]) );
  INV3 U249 ( .A(i_data_A[2]), .Q(n333) );
  LOGIC0 U250 ( .Q(n13) );
  NOR40 U251 ( .A(i_con_AluCtrl[2]), .B(n17), .C(i_con_AluCtrl[1]), .D(n196), 
        .Q(n59) );
  NOR40 U252 ( .A(i_con_AluCtrl[1]), .B(i_con_AluCtrl[0]), .C(i_con_AluCtrl[2]), .D(n196), .Q(n317) );
  OAI2111 U253 ( .A(i_data_A[13]), .B(n34), .C(n295), .D(n43), .Q(n175) );
  OAI2110 U254 ( .A(i_data_A[22]), .B(n35), .C(n225), .D(n44), .Q(n237) );
  INV0 U255 ( .A(i_data_A[1]), .Q(n83) );
  NAND20 U256 ( .A(i_data_A[19]), .B(n4), .Q(n253) );
  IMUX30 U257 ( .A(n305), .B(n51), .C(n292), .S0(i_data_A[28]), .S1(
        i_data_B[28]), .Q(n293) );
  OAI2111 U258 ( .A(i_data_A[28]), .B(n34), .C(n183), .D(n43), .Q(n292) );
  AOI210 U259 ( .A(i_data_A[0]), .B(n46), .C(n77), .Q(n78) );
  OAI2110 U260 ( .A(i_data_A[18]), .B(n34), .C(n260), .D(n44), .Q(n209) );
  NAND22 U261 ( .A(i_data_A[18]), .B(n5), .Q(n260) );
  OAI2111 U262 ( .A(i_data_A[27]), .B(n35), .C(n190), .D(n43), .Q(n282) );
  IMUX30 U263 ( .A(n305), .B(n51), .C(n198), .S0(i_data_A[16]), .S1(
        i_data_B[16]), .Q(n199) );
  OAI2110 U264 ( .A(i_data_A[16]), .B(n50), .C(n274), .D(n44), .Q(n198) );
  AOI221 U265 ( .A(i_data_A[21]), .B(n47), .C(N137), .D(n21), .Q(n234) );
  OAI2110 U266 ( .A(i_data_A[21]), .B(n34), .C(n232), .D(n44), .Q(n231) );
  IMUX30 U267 ( .A(n305), .B(n51), .C(n231), .S0(i_data_A[21]), .S1(
        i_data_B[21]), .Q(n233) );
  OAI2110 U268 ( .A(i_data_A[29]), .B(n35), .C(n176), .D(n43), .Q(n298) );
  NAND20 U269 ( .A(i_data_A[29]), .B(n4), .Q(n176) );
  IMUX30 U270 ( .A(n305), .B(n51), .C(n298), .S0(i_data_A[29]), .S1(n18), .Q(
        n301) );
  IMUX30 U271 ( .A(n305), .B(n52), .C(n152), .S0(i_data_A[10]), .S1(
        i_data_B[10]), .Q(n154) );
  INV0 U272 ( .A(i_data_B[10]), .Q(n275) );
  AOI211 U273 ( .A(i_data_A[26]), .B(n46), .C(n276), .Q(n278) );
  CLKIN2 U274 ( .A(i_data_A[11]), .Q(n161) );
  OAI2110 U275 ( .A(i_data_A[5]), .B(n35), .C(n45), .D(n132), .Q(n131) );
  OAI220 U276 ( .A(n50), .B(n330), .C(i_data_A[5]), .D(n99), .Q(n130) );
  AOI220 U277 ( .A(n37), .B(n42), .C(N202), .D(n40), .Q(n242) );
  OAI2110 U278 ( .A(i_data_A[9]), .B(n50), .C(n97), .D(n43), .Q(n147) );
  IMUX30 U279 ( .A(n305), .B(n52), .C(n147), .S0(i_data_A[9]), .S1(i_data_B[9]), .Q(n148) );
  AOI220 U280 ( .A(i_data_A[12]), .B(n48), .C(N128), .D(n21), .Q(n172) );
  OAI2110 U281 ( .A(i_data_A[12]), .B(n34), .C(n302), .D(n43), .Q(n170) );
  IMUX30 U282 ( .A(n305), .B(n52), .C(n170), .S0(i_data_A[12]), .S1(
        i_data_B[12]), .Q(n171) );
  AOI220 U283 ( .A(n167), .B(n332), .C(i_data_B[2]), .D(n168), .Q(n166) );
  AOI220 U284 ( .A(i_data_B[2]), .B(n42), .C(N198), .D(n40), .Q(n214) );
  OAI2110 U285 ( .A(i_data_A[3]), .B(n35), .C(n45), .D(n146), .Q(n145) );
  OAI220 U286 ( .A(n35), .B(n94), .C(i_data_A[3]), .D(n99), .Q(n144) );
  OAI2110 U287 ( .A(i_data_A[15]), .B(n35), .C(n281), .D(n43), .Q(n191) );
  IMUX30 U288 ( .A(n305), .B(n51), .C(n191), .S0(i_data_A[15]), .S1(
        i_data_B[15]), .Q(n192) );
  AOI211 U289 ( .A(i_data_A[25]), .B(n46), .C(n268), .Q(n269) );
  OAI2111 U290 ( .A(i_data_A[25]), .B(n34), .C(n204), .D(n43), .Q(n264) );
  NAND20 U291 ( .A(i_data_A[25]), .B(n5), .Q(n204) );
  IMUX30 U292 ( .A(n305), .B(n51), .C(n209), .S0(i_data_A[18]), .S1(
        i_data_B[18]), .Q(n210) );
  OAI2110 U293 ( .A(i_data_A[4]), .B(n35), .C(n45), .D(n139), .Q(n138) );
  OAI220 U294 ( .A(n35), .B(n104), .C(i_data_A[4]), .D(n99), .Q(n137) );
  CLKIN1 U295 ( .A(i_data_A[4]), .Q(n104) );
  INV2 U296 ( .A(i_data_A[31]), .Q(n62) );
  XNR20 U297 ( .A(i_data_B[31]), .B(i_data_A[31]), .Q(n63) );
  IMUX30 U298 ( .A(n305), .B(n51), .C(n237), .S0(i_data_A[22]), .S1(
        i_data_B[22]), .Q(n238) );
  AOI220 U299 ( .A(i_data_A[8]), .B(n48), .C(N124), .D(n21), .Q(n140) );
  OAI2110 U300 ( .A(i_data_A[8]), .B(n35), .C(n111), .D(n43), .Q(n134) );
  IMUX30 U301 ( .A(n99), .B(n35), .C(n123), .S0(i_data_A[7]), .S1(i_data_B[7]), 
        .Q(n124) );
  NAND22 U302 ( .A(n177), .B(n179), .Q(n38) );
  INV3 U303 ( .A(n38), .Q(n39) );
  AOI220 U304 ( .A(N257), .B(n2), .C(i_data_A[13]), .D(n46), .Q(n178) );
  AOI220 U305 ( .A(n130), .B(n327), .C(i_data_B[5]), .D(n131), .Q(n129) );
  AOI220 U306 ( .A(i_data_B[5]), .B(n42), .C(N201), .D(n40), .Q(n236) );
  AOI220 U307 ( .A(i_data_B[13]), .B(n42), .C(i_data_A[29]), .D(n46), .Q(n300)
         );
  IMUX30 U308 ( .A(n305), .B(n52), .C(n175), .S0(i_data_A[13]), .S1(
        i_data_B[13]), .Q(n177) );
  INV2 U309 ( .A(i_data_B[8]), .Q(n258) );
  IMUX30 U310 ( .A(n305), .B(n52), .C(n134), .S0(i_data_A[8]), .S1(i_data_B[8]), .Q(n135) );
  AOI220 U311 ( .A(i_data_B[0]), .B(n42), .C(N196), .D(n40), .Q(n202) );
  CLKIN3 U312 ( .A(n59), .Q(n64) );
  CLKIN3 U313 ( .A(n60), .Q(n72) );
  OAI222 U314 ( .A(n315), .B(n64), .C(n68), .D(n61), .Q(n66) );
  NAND22 U315 ( .A(n72), .B(n68), .Q(n69) );
  NAND22 U316 ( .A(n328), .B(n44), .Q(n74) );
  NAND22 U317 ( .A(N181), .B(n40), .Q(n87) );
  NAND22 U318 ( .A(N149), .B(n1), .Q(n86) );
  NAND22 U319 ( .A(N245), .B(n2), .Q(n82) );
  NAND22 U320 ( .A(N182), .B(n41), .Q(n92) );
  NAND22 U321 ( .A(N150), .B(n1), .Q(n91) );
  NAND22 U322 ( .A(N246), .B(n2), .Q(n88) );
  NAND22 U323 ( .A(N183), .B(n40), .Q(n102) );
  NAND22 U324 ( .A(N151), .B(n1), .Q(n101) );
  NAND22 U325 ( .A(N247), .B(n2), .Q(n93) );
  NAND22 U326 ( .A(N184), .B(n41), .Q(n108) );
  NAND22 U327 ( .A(N152), .B(n1), .Q(n107) );
  NAND22 U328 ( .A(N248), .B(n2), .Q(n103) );
  NAND22 U329 ( .A(N185), .B(n40), .Q(n114) );
  NAND22 U330 ( .A(N249), .B(n2), .Q(n109) );
  CLKIN3 U331 ( .A(i_data_A[7]), .Q(n122) );
  NAND22 U332 ( .A(n118), .B(n45), .Q(n121) );
  NAND22 U333 ( .A(N251), .B(n2), .Q(n126) );
  NAND22 U334 ( .A(N252), .B(n2), .Q(n141) );
  NAND22 U335 ( .A(N253), .B(n2), .Q(n150) );
  NAND22 U336 ( .A(N254), .B(n2), .Q(n156) );
  NAND42 U337 ( .A(n157), .B(n156), .C(n154), .D(n155), .Q(o_data_AluRes[10])
         );
  AOI212 U338 ( .A(N127), .B(n21), .C(n163), .Q(n164) );
  NAND22 U339 ( .A(n165), .B(n164), .Q(o_data_AluRes[11]) );
  NAND22 U340 ( .A(N161), .B(n1), .Q(n179) );
  NAND22 U341 ( .A(N194), .B(n40), .Q(n188) );
  CLKIN3 U342 ( .A(i_data_A[14]), .Q(n182) );
  NAND22 U343 ( .A(N130), .B(n21), .Q(n186) );
  NAND42 U344 ( .A(n189), .B(n188), .C(n187), .D(n186), .Q(o_data_AluRes[14])
         );
  NAND22 U345 ( .A(N259), .B(n2), .Q(n194) );
  NAND22 U346 ( .A(N199), .B(n41), .Q(n222) );
  CLKIN3 U347 ( .A(n42), .Q(n285) );
  CLKIN3 U348 ( .A(i_data_B[3]), .Q(n217) );
  OAI212 U349 ( .A(n285), .B(n217), .C(n216), .Q(n219) );
  NAND22 U350 ( .A(N263), .B(n2), .Q(n220) );
  NAND42 U351 ( .A(n220), .B(n222), .C(n221), .D(n223), .Q(o_data_AluRes[19])
         );
  OAI212 U352 ( .A(n285), .B(n331), .C(n226), .Q(n227) );
  NAND22 U353 ( .A(N203), .B(n40), .Q(n248) );
  OAI212 U354 ( .A(n285), .B(n249), .C(n248), .Q(n250) );
  NAND22 U355 ( .A(N267), .B(n2), .Q(n251) );
  NAND42 U356 ( .A(n255), .B(n254), .C(n252), .D(n251), .Q(o_data_AluRes[23])
         );
  OAI212 U357 ( .A(n285), .B(n258), .C(n257), .Q(n259) );
  CLKIN3 U358 ( .A(i_data_B[9]), .Q(n266) );
  OAI212 U359 ( .A(n285), .B(n266), .C(n265), .Q(n268) );
  NAND22 U360 ( .A(N206), .B(n41), .Q(n279) );
  OAI212 U361 ( .A(n285), .B(n275), .C(n273), .Q(n276) );
  NAND22 U362 ( .A(N270), .B(n2), .Q(n277) );
  NAND42 U363 ( .A(n277), .B(n279), .C(n278), .D(n280), .Q(o_data_AluRes[26])
         );
  CLKIN3 U364 ( .A(i_data_B[11]), .Q(n284) );
  OAI212 U365 ( .A(n285), .B(n284), .C(n283), .Q(n286) );
  NAND22 U366 ( .A(n310), .B(n308), .Q(n311) );
  NAND22 U367 ( .A(N146), .B(n21), .Q(n313) );
  NAND22 U368 ( .A(n314), .B(n313), .Q(o_data_AluRes[30]) );
endmodule


module E_alu_control ( o_con_AluCtrl, i_con_AluOp, i_con_FuncCode );
  output [3:0] o_con_AluCtrl;
  input [5:0] i_con_AluOp;
  input [5:0] i_con_FuncCode;
  wire   n59, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n54, n55, n56, n57,
         n58;

  OAI2112 U13 ( .A(n41), .B(n28), .C(n24), .D(n42), .Q(o_con_AluCtrl[0]) );
  OAI310 U3 ( .A(n32), .B(i_con_FuncCode[1]), .C(n58), .D(n52), .Q(n48) );
  NAND33 U4 ( .A(n49), .B(n32), .C(n33), .Q(n51) );
  CLKIN3 U5 ( .A(i_con_FuncCode[5]), .Q(n20) );
  BUF12 U6 ( .A(n59), .Q(o_con_AluCtrl[1]) );
  NAND31 U7 ( .A(i_con_FuncCode[5]), .B(n56), .C(i_con_FuncCode[2]), .Q(n32)
         );
  NAND41 U8 ( .A(n36), .B(n29), .C(n11), .D(n37), .Q(n59) );
  CLKIN3 U9 ( .A(i_con_FuncCode[3]), .Q(n56) );
  OAI2111 U10 ( .A(n15), .B(n22), .C(n23), .D(n24), .Q(o_con_AluCtrl[3]) );
  NOR21 U11 ( .A(n5), .B(n26), .Q(n27) );
  NOR31 U12 ( .A(i_con_FuncCode[2]), .B(i_con_FuncCode[3]), .C(n20), .Q(n35)
         );
  NOR21 U14 ( .A(i_con_AluOp[4]), .B(i_con_AluOp[3]), .Q(n1) );
  NOR31 U15 ( .A(n2), .B(n10), .C(n12), .Q(n44) );
  INV3 U16 ( .A(n1), .Q(n2) );
  AOI311 U17 ( .A(i_con_AluOp[3]), .B(i_con_AluOp[0]), .C(n43), .D(n8), .Q(n42) );
  NOR21 U18 ( .A(i_con_AluOp[5]), .B(i_con_AluOp[4]), .Q(n43) );
  NOR32 U19 ( .A(i_con_FuncCode[3]), .B(i_con_FuncCode[5]), .C(
        i_con_FuncCode[2]), .Q(n47) );
  OAI2112 U20 ( .A(n27), .B(n28), .C(n29), .D(n7), .Q(o_con_AluCtrl[2]) );
  OAI211 U21 ( .A(n35), .B(n40), .C(n14), .Q(n36) );
  NAND42 U22 ( .A(n49), .B(n18), .C(n16), .D(n55), .Q(n40) );
  INV6 U23 ( .A(i_con_FuncCode[1]), .Q(n57) );
  CLKIN0 U24 ( .A(n33), .Q(n21) );
  NAND22 U25 ( .A(n47), .B(i_con_FuncCode[1]), .Q(n33) );
  OAI211 U26 ( .A(n25), .B(n26), .C(n14), .Q(n23) );
  NOR41 U27 ( .A(n51), .B(n35), .C(n31), .D(n25), .Q(n50) );
  NOR22 U28 ( .A(n19), .B(i_con_FuncCode[0]), .Q(n25) );
  NOR31 U29 ( .A(n21), .B(n31), .C(n17), .Q(n4) );
  INV3 U30 ( .A(n4), .Q(n5) );
  NOR22 U31 ( .A(n58), .B(n19), .Q(n31) );
  OAI2112 U32 ( .A(n57), .B(n32), .C(n16), .D(n55), .Q(n26) );
  CLKIN0 U33 ( .A(i_con_AluOp[1]), .Q(n13) );
  INV1 U34 ( .A(n38), .Q(n6) );
  CLKIN1 U35 ( .A(n29), .Q(n8) );
  INV0 U36 ( .A(n31), .Q(n18) );
  NOR20 U37 ( .A(n13), .B(n6), .Q(n37) );
  NOR41 U38 ( .A(n20), .B(n56), .C(n57), .D(i_con_FuncCode[2]), .Q(n53) );
  CLKIN4 U39 ( .A(n53), .Q(n19) );
  CLKIN3 U40 ( .A(i_con_AluOp[2]), .Q(n12) );
  AOI2110 U41 ( .A(n47), .B(i_con_FuncCode[0]), .C(n48), .D(n40), .Q(n41) );
  NAND20 U42 ( .A(i_con_AluOp[1]), .B(n15), .Q(n28) );
  INV0 U43 ( .A(n32), .Q(n54) );
  AOI310 U44 ( .A(i_con_FuncCode[1]), .B(n58), .C(n54), .D(n25), .Q(n52) );
  NAND20 U45 ( .A(n44), .B(i_con_AluOp[0]), .Q(n29) );
  NOR30 U46 ( .A(i_con_AluOp[2]), .B(i_con_AluOp[3]), .C(n15), .Q(n39) );
  NAND40 U47 ( .A(n43), .B(i_con_AluOp[2]), .C(i_con_AluOp[3]), .D(
        i_con_AluOp[0]), .Q(n45) );
  CLKIN3 U48 ( .A(i_con_FuncCode[0]), .Q(n58) );
  CLKIN3 U49 ( .A(i_con_AluOp[5]), .Q(n10) );
  NAND20 U50 ( .A(i_con_FuncCode[1]), .B(n35), .Q(n34) );
  INV3 U51 ( .A(n39), .Q(n11) );
  INV3 U52 ( .A(n30), .Q(n7) );
  NAND31 U53 ( .A(n58), .B(n57), .C(n47), .Q(n49) );
  INV3 U54 ( .A(n22), .Q(n9) );
  INV3 U55 ( .A(n50), .Q(n16) );
  INV3 U56 ( .A(n28), .Q(n14) );
  AOI211 U57 ( .A(n13), .B(i_con_AluOp[0]), .C(n46), .Q(n38) );
  NOR40 U58 ( .A(n15), .B(n43), .C(n44), .D(n9), .Q(n46) );
  AOI311 U59 ( .A(n9), .B(n12), .C(i_con_AluOp[0]), .D(n30), .Q(n24) );
  NAND31 U60 ( .A(i_con_AluOp[3]), .B(n10), .C(i_con_AluOp[4]), .Q(n22) );
  INV3 U61 ( .A(i_con_AluOp[0]), .Q(n15) );
  NAND22 U62 ( .A(n38), .B(n45), .Q(n30) );
  INV3 U63 ( .A(n34), .Q(n17) );
  INV3 U64 ( .A(i_con_FuncCode[4]), .Q(n55) );
endmodule


module E_famux5 ( i_data_rs, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fa, o_data_alusra );
  input [31:0] i_data_rs;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fa;
  output [31:0] o_data_alusra;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128;

  NAND26 U1 ( .A(n32), .B(n4), .Q(o_data_alusra[1]) );
  NAND33 U2 ( .A(n74), .B(n73), .C(n72), .Q(o_data_alusra[14]) );
  NAND31 U3 ( .A(n122), .B(n121), .C(n120), .Q(o_data_alusra[30]) );
  AOI221 U4 ( .A(i_data_lwM[7]), .B(n125), .C(i_data_lwW[7]), .D(n20), .Q(n51)
         );
  AOI221 U5 ( .A(i_data_rs[7]), .B(n12), .C(i_data_writeres[7]), .D(n19), .Q(
        n53) );
  NAND22 U6 ( .A(i_data_alures[25]), .B(n13), .Q(n106) );
  NAND33 U7 ( .A(n77), .B(n76), .C(n75), .Q(o_data_alusra[15]) );
  AOI221 U8 ( .A(i_data_lwM[15]), .B(n125), .C(i_data_lwW[15]), .D(n20), .Q(
        n75) );
  NAND33 U9 ( .A(n101), .B(n100), .C(n99), .Q(o_data_alusra[23]) );
  AOI221 U10 ( .A(i_data_lwM[23]), .B(n125), .C(i_data_lwW[23]), .D(n20), .Q(
        n99) );
  AOI221 U11 ( .A(i_data_rs[23]), .B(n11), .C(i_data_writeres[23]), .D(n19), 
        .Q(n101) );
  AOI221 U12 ( .A(i_data_lwM[30]), .B(n125), .C(i_data_lwW[30]), .D(n20), .Q(
        n120) );
  AOI221 U13 ( .A(i_data_rs[30]), .B(n11), .C(i_data_writeres[30]), .D(n19), 
        .Q(n122) );
  AOI220 U14 ( .A(i_data_lwM[18]), .B(n125), .C(i_data_lwW[18]), .D(n20), .Q(
        n84) );
  NAND24 U15 ( .A(n93), .B(n10), .Q(o_data_alusra[21]) );
  INV3 U16 ( .A(n9), .Q(n10) );
  NAND22 U17 ( .A(n95), .B(n94), .Q(n9) );
  NAND31 U18 ( .A(n116), .B(n115), .C(n114), .Q(o_data_alusra[28]) );
  AOI221 U19 ( .A(i_data_lwM[8]), .B(n125), .C(i_data_lwW[8]), .D(n20), .Q(n54) );
  NAND33 U20 ( .A(n89), .B(n88), .C(n87), .Q(o_data_alusra[19]) );
  AOI221 U21 ( .A(i_data_lwM[10]), .B(n125), .C(i_data_lwW[10]), .D(n20), .Q(
        n60) );
  AOI221 U22 ( .A(i_data_rs[10]), .B(n12), .C(i_data_writeres[10]), .D(n19), 
        .Q(n62) );
  AOI221 U23 ( .A(i_data_lwM[11]), .B(n125), .C(i_data_lwW[11]), .D(n20), .Q(
        n63) );
  AOI221 U24 ( .A(i_data_rs[21]), .B(n12), .C(i_data_writeres[21]), .D(n19), 
        .Q(n95) );
  NAND22 U25 ( .A(i_data_alures[21]), .B(n13), .Q(n94) );
  NAND22 U26 ( .A(n34), .B(n33), .Q(n3) );
  AOI221 U27 ( .A(i_data_rs[4]), .B(n12), .C(i_data_writeres[4]), .D(n19), .Q(
        n44) );
  NAND33 U28 ( .A(n50), .B(n49), .C(n48), .Q(o_data_alusra[6]) );
  INV3 U29 ( .A(n28), .Q(n124) );
  INV12 U30 ( .A(n26), .Q(n125) );
  INV12 U31 ( .A(n24), .Q(n13) );
  INV3 U32 ( .A(n14), .Q(n15) );
  NAND31 U33 ( .A(n104), .B(n103), .C(n102), .Q(o_data_alusra[24]) );
  NAND33 U34 ( .A(n110), .B(n109), .C(n108), .Q(o_data_alusra[26]) );
  NAND26 U35 ( .A(n31), .B(n17), .Q(o_data_alusra[0]) );
  INV3 U36 ( .A(n16), .Q(n17) );
  AOI221 U37 ( .A(i_data_lwM[20]), .B(n125), .C(i_data_lwW[20]), .D(n20), .Q(
        n90) );
  AOI221 U38 ( .A(i_data_rs[20]), .B(n11), .C(i_data_writeres[20]), .D(n19), 
        .Q(n92) );
  AOI221 U39 ( .A(i_data_lwM[13]), .B(n125), .C(i_data_lwW[13]), .D(n20), .Q(
        n69) );
  AOI221 U40 ( .A(i_data_rs[13]), .B(n12), .C(i_data_writeres[13]), .D(n19), 
        .Q(n71) );
  AOI221 U41 ( .A(i_data_rs[2]), .B(n11), .C(i_data_writeres[2]), .D(n19), .Q(
        n38) );
  NAND22 U42 ( .A(n25), .B(n15), .Q(n24) );
  NAND33 U43 ( .A(n59), .B(n58), .C(n57), .Q(o_data_alusra[9]) );
  AOI221 U44 ( .A(i_data_lwM[26]), .B(n125), .C(i_data_lwW[26]), .D(n20), .Q(
        n108) );
  INV3 U45 ( .A(n21), .Q(n35) );
  NAND33 U46 ( .A(n41), .B(n40), .C(n39), .Q(o_data_alusra[3]) );
  NAND33 U47 ( .A(n119), .B(n118), .C(n117), .Q(o_data_alusra[29]) );
  AOI221 U48 ( .A(i_data_lwM[29]), .B(n125), .C(i_data_lwW[29]), .D(n20), .Q(
        n117) );
  NAND22 U49 ( .A(n23), .B(i_con_fa[0]), .Q(n1) );
  NAND22 U50 ( .A(n27), .B(n2), .Q(n22) );
  CLKIN3 U51 ( .A(n1), .Q(n2) );
  CLKIN6 U52 ( .A(i_con_fa[1]), .Q(n27) );
  INV3 U53 ( .A(n3), .Q(n4) );
  NAND24 U54 ( .A(n106), .B(n107), .Q(n5) );
  NAND24 U55 ( .A(n105), .B(n6), .Q(o_data_alusra[25]) );
  CLKIN6 U56 ( .A(n5), .Q(n6) );
  AOI222 U57 ( .A(i_data_rs[25]), .B(n11), .C(i_data_writeres[25]), .D(n19), 
        .Q(n107) );
  NAND22 U58 ( .A(i_con_fa[1]), .B(n21), .Q(n7) );
  NAND22 U59 ( .A(n27), .B(n35), .Q(n8) );
  NAND24 U60 ( .A(n7), .B(n8), .Q(n18) );
  BUF12 U61 ( .A(n18), .Q(n11) );
  BUF12 U62 ( .A(n18), .Q(n12) );
  AOI221 U63 ( .A(i_data_lwM[21]), .B(n125), .C(i_data_lwW[21]), .D(n20), .Q(
        n93) );
  AOI221 U64 ( .A(i_data_lwM[4]), .B(n125), .C(i_data_lwW[4]), .D(n20), .Q(n42) );
  NAND33 U65 ( .A(n68), .B(n67), .C(n66), .Q(o_data_alusra[12]) );
  NAND31 U66 ( .A(i_con_fa[2]), .B(i_con_fa[0]), .C(n27), .Q(n28) );
  NAND33 U67 ( .A(n47), .B(n46), .C(n45), .Q(o_data_alusra[5]) );
  AOI221 U68 ( .A(i_data_lwM[12]), .B(n125), .C(i_data_lwW[12]), .D(n20), .Q(
        n66) );
  BUF15 U69 ( .A(n124), .Q(n20) );
  NAND22 U70 ( .A(i_con_fa[1]), .B(n23), .Q(n14) );
  NAND34 U71 ( .A(n53), .B(n52), .C(n51), .Q(o_data_alusra[7]) );
  CLKBU15 U72 ( .A(n123), .Q(n19) );
  NAND22 U73 ( .A(n29), .B(n30), .Q(n16) );
  AOI221 U74 ( .A(i_data_rs[0]), .B(n12), .C(i_data_writeres[0]), .D(n19), .Q(
        n31) );
  AOI220 U75 ( .A(i_data_lwM[0]), .B(n125), .C(i_data_lwW[0]), .D(n20), .Q(n29) );
  AOI220 U76 ( .A(i_data_lwM[1]), .B(n125), .C(i_data_lwW[1]), .D(n20), .Q(n32) );
  NAND24 U77 ( .A(n23), .B(n25), .Q(n21) );
  AOI220 U78 ( .A(i_data_rs[28]), .B(n11), .C(i_data_writeres[28]), .D(n19), 
        .Q(n116) );
  AOI220 U79 ( .A(i_data_lwM[25]), .B(n125), .C(i_data_lwW[25]), .D(n20), .Q(
        n105) );
  CLKIN6 U80 ( .A(i_con_fa[0]), .Q(n25) );
  AOI220 U81 ( .A(i_data_rs[12]), .B(n11), .C(i_data_writeres[12]), .D(n19), 
        .Q(n68) );
  AOI221 U82 ( .A(i_data_lwM[27]), .B(n125), .C(i_data_lwW[27]), .D(n20), .Q(
        n111) );
  AOI221 U83 ( .A(i_data_rs[27]), .B(n12), .C(i_data_writeres[27]), .D(n19), 
        .Q(n113) );
  AOI220 U84 ( .A(i_data_lwM[28]), .B(n125), .C(i_data_lwW[28]), .D(n20), .Q(
        n114) );
  AOI221 U85 ( .A(i_data_lwM[19]), .B(n125), .C(i_data_lwW[19]), .D(n20), .Q(
        n87) );
  AOI221 U86 ( .A(i_data_rs[19]), .B(n11), .C(i_data_writeres[19]), .D(n19), 
        .Q(n89) );
  NAND34 U87 ( .A(n44), .B(n43), .C(n42), .Q(o_data_alusra[4]) );
  AOI220 U88 ( .A(i_data_rs[22]), .B(n11), .C(i_data_writeres[22]), .D(n19), 
        .Q(n98) );
  AOI220 U89 ( .A(i_data_lwM[22]), .B(n125), .C(i_data_lwW[22]), .D(n20), .Q(
        n96) );
  AOI220 U90 ( .A(i_data_rs[24]), .B(n11), .C(i_data_writeres[24]), .D(n19), 
        .Q(n104) );
  AOI221 U91 ( .A(i_data_lwM[24]), .B(n125), .C(i_data_lwW[24]), .D(n20), .Q(
        n102) );
  AOI221 U92 ( .A(i_data_lwM[16]), .B(n125), .C(i_data_lwW[16]), .D(n20), .Q(
        n78) );
  AOI221 U93 ( .A(i_data_rs[3]), .B(n12), .C(i_data_writeres[3]), .D(n19), .Q(
        n41) );
  AOI221 U94 ( .A(i_data_lwM[3]), .B(n125), .C(i_data_lwW[3]), .D(n20), .Q(n39) );
  AOI221 U95 ( .A(i_data_lwM[2]), .B(n125), .C(i_data_lwW[2]), .D(n20), .Q(n36) );
  NAND31 U96 ( .A(n38), .B(n37), .C(n36), .Q(o_data_alusra[2]) );
  INV3 U97 ( .A(n22), .Q(n123) );
  NAND33 U98 ( .A(n113), .B(n112), .C(n111), .Q(o_data_alusra[27]) );
  NAND22 U99 ( .A(i_data_alures[27]), .B(n13), .Q(n112) );
  NAND32 U100 ( .A(i_con_fa[2]), .B(n25), .C(n27), .Q(n26) );
  AOI220 U101 ( .A(i_data_rs[16]), .B(n12), .C(i_data_writeres[16]), .D(n19), 
        .Q(n80) );
  AOI221 U102 ( .A(i_data_rs[9]), .B(n11), .C(i_data_writeres[9]), .D(n19), 
        .Q(n59) );
  AOI221 U103 ( .A(i_data_rs[11]), .B(n12), .C(i_data_writeres[11]), .D(n19), 
        .Q(n65) );
  AOI221 U104 ( .A(i_data_rs[15]), .B(n12), .C(i_data_writeres[15]), .D(n19), 
        .Q(n77) );
  AOI220 U105 ( .A(i_data_rs[29]), .B(n11), .C(i_data_writeres[29]), .D(n19), 
        .Q(n119) );
  AOI220 U106 ( .A(i_data_rs[26]), .B(n12), .C(i_data_writeres[26]), .D(n19), 
        .Q(n110) );
  AOI221 U107 ( .A(i_data_rs[18]), .B(n11), .C(i_data_writeres[18]), .D(n19), 
        .Q(n86) );
  AOI221 U108 ( .A(i_data_rs[31]), .B(n11), .C(i_data_writeres[31]), .D(n19), 
        .Q(n128) );
  NAND34 U109 ( .A(n128), .B(n127), .C(n126), .Q(o_data_alusra[31]) );
  AOI221 U110 ( .A(i_data_lwM[31]), .B(n125), .C(i_data_lwW[31]), .D(n20), .Q(
        n126) );
  AOI221 U111 ( .A(i_data_rs[8]), .B(n12), .C(i_data_writeres[8]), .D(n19), 
        .Q(n56) );
  NAND34 U112 ( .A(n56), .B(n55), .C(n54), .Q(o_data_alusra[8]) );
  AOI221 U113 ( .A(i_data_rs[14]), .B(n12), .C(i_data_writeres[14]), .D(n19), 
        .Q(n74) );
  AOI221 U114 ( .A(i_data_lwM[14]), .B(n125), .C(i_data_lwW[14]), .D(n20), .Q(
        n72) );
  AOI221 U115 ( .A(i_data_rs[5]), .B(n12), .C(i_data_writeres[5]), .D(n19), 
        .Q(n47) );
  AOI221 U116 ( .A(i_data_lwM[5]), .B(n125), .C(i_data_lwW[5]), .D(n20), .Q(
        n45) );
  AOI221 U117 ( .A(i_data_rs[1]), .B(n11), .C(i_data_writeres[1]), .D(n19), 
        .Q(n34) );
  NAND34 U118 ( .A(n92), .B(n91), .C(n90), .Q(o_data_alusra[20]) );
  AOI221 U119 ( .A(i_data_lwM[9]), .B(n125), .C(i_data_lwW[9]), .D(n20), .Q(
        n57) );
  NAND34 U120 ( .A(n83), .B(n82), .C(n81), .Q(o_data_alusra[17]) );
  CLKIN6 U121 ( .A(i_con_fa[2]), .Q(n23) );
  NAND34 U122 ( .A(n65), .B(n64), .C(n63), .Q(o_data_alusra[11]) );
  NAND34 U123 ( .A(n80), .B(n79), .C(n78), .Q(o_data_alusra[16]) );
  NAND22 U124 ( .A(i_data_alures[0]), .B(n13), .Q(n30) );
  NAND22 U125 ( .A(i_data_alures[1]), .B(n13), .Q(n33) );
  NAND22 U126 ( .A(i_data_alures[2]), .B(n13), .Q(n37) );
  NAND22 U127 ( .A(i_data_alures[3]), .B(n13), .Q(n40) );
  NAND22 U128 ( .A(i_data_alures[4]), .B(n13), .Q(n43) );
  NAND22 U129 ( .A(i_data_alures[5]), .B(n13), .Q(n46) );
  AOI222 U130 ( .A(i_data_rs[6]), .B(n11), .C(i_data_writeres[6]), .D(n19), 
        .Q(n50) );
  NAND22 U131 ( .A(i_data_alures[6]), .B(n13), .Q(n49) );
  AOI222 U132 ( .A(i_data_lwM[6]), .B(n125), .C(i_data_lwW[6]), .D(n20), .Q(
        n48) );
  NAND22 U133 ( .A(i_data_alures[7]), .B(n13), .Q(n52) );
  NAND22 U134 ( .A(i_data_alures[8]), .B(n13), .Q(n55) );
  NAND22 U135 ( .A(i_data_alures[9]), .B(n13), .Q(n58) );
  NAND22 U136 ( .A(i_data_alures[10]), .B(n13), .Q(n61) );
  NAND33 U137 ( .A(n62), .B(n61), .C(n60), .Q(o_data_alusra[10]) );
  NAND22 U138 ( .A(i_data_alures[11]), .B(n13), .Q(n64) );
  NAND22 U139 ( .A(i_data_alures[12]), .B(n13), .Q(n67) );
  NAND22 U140 ( .A(i_data_alures[13]), .B(n13), .Q(n70) );
  NAND33 U141 ( .A(n71), .B(n70), .C(n69), .Q(o_data_alusra[13]) );
  NAND22 U142 ( .A(i_data_alures[14]), .B(n13), .Q(n73) );
  NAND22 U143 ( .A(i_data_alures[15]), .B(n13), .Q(n76) );
  NAND22 U144 ( .A(i_data_alures[16]), .B(n13), .Q(n79) );
  AOI222 U145 ( .A(i_data_rs[17]), .B(n12), .C(i_data_writeres[17]), .D(n19), 
        .Q(n83) );
  NAND22 U146 ( .A(i_data_alures[17]), .B(n13), .Q(n82) );
  AOI222 U147 ( .A(i_data_lwM[17]), .B(n125), .C(i_data_lwW[17]), .D(n20), .Q(
        n81) );
  NAND22 U148 ( .A(i_data_alures[18]), .B(n13), .Q(n85) );
  NAND33 U149 ( .A(n86), .B(n85), .C(n84), .Q(o_data_alusra[18]) );
  NAND22 U150 ( .A(i_data_alures[19]), .B(n13), .Q(n88) );
  NAND22 U151 ( .A(i_data_alures[20]), .B(n13), .Q(n91) );
  NAND22 U152 ( .A(i_data_alures[22]), .B(n13), .Q(n97) );
  NAND33 U153 ( .A(n98), .B(n97), .C(n96), .Q(o_data_alusra[22]) );
  NAND22 U154 ( .A(i_data_alures[23]), .B(n13), .Q(n100) );
  NAND22 U155 ( .A(i_data_alures[24]), .B(n13), .Q(n103) );
  NAND22 U156 ( .A(i_data_alures[26]), .B(n13), .Q(n109) );
  NAND22 U157 ( .A(i_data_alures[28]), .B(n13), .Q(n115) );
  NAND22 U158 ( .A(i_data_alures[29]), .B(n13), .Q(n118) );
  NAND22 U159 ( .A(i_data_alures[30]), .B(n13), .Q(n121) );
  NAND22 U160 ( .A(i_data_alures[31]), .B(n13), .Q(n127) );
endmodule


module E_fbmux5 ( i_data_rt, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fb, o_data_alusrb );
  input [31:0] i_data_rt;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fb;
  output [31:0] o_data_alusrb;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145;

  NAND34 U1 ( .A(n89), .B(n88), .C(n87), .Q(o_data_alusrb[15]) );
  CLKIN8 U2 ( .A(n140), .Q(n22) );
  INV3 U3 ( .A(n34), .Q(n141) );
  INV3 U4 ( .A(n31), .Q(n140) );
  INV12 U5 ( .A(n22), .Q(n23) );
  INV8 U6 ( .A(n29), .Q(n20) );
  INV12 U7 ( .A(n22), .Q(n24) );
  INV6 U8 ( .A(n68), .Q(n102) );
  NAND22 U9 ( .A(n8), .B(n9), .Q(n68) );
  NAND22 U10 ( .A(n112), .B(n113), .Q(n16) );
  NAND33 U11 ( .A(n45), .B(n44), .C(n43), .Q(o_data_alusrb[2]) );
  NAND33 U12 ( .A(n57), .B(n56), .C(n55), .Q(o_data_alusrb[5]) );
  NAND33 U13 ( .A(n63), .B(n62), .C(n61), .Q(o_data_alusrb[7]) );
  NAND22 U14 ( .A(n38), .B(n3), .Q(o_data_alusrb[0]) );
  NAND34 U15 ( .A(n60), .B(n59), .C(n58), .Q(o_data_alusrb[6]) );
  NAND33 U16 ( .A(n83), .B(n82), .C(n81), .Q(o_data_alusrb[13]) );
  AOI221 U17 ( .A(i_data_writeres[13]), .B(n138), .C(i_data_alures[13]), .D(
        n24), .Q(n83) );
  AOI222 U18 ( .A(i_data_lwM[19]), .B(n142), .C(i_data_lwW[19]), .D(n29), .Q(
        n99) );
  CLKIN15 U19 ( .A(n32), .Q(n142) );
  NAND24 U20 ( .A(n114), .B(n17), .Q(o_data_alusrb[23]) );
  AOI221 U21 ( .A(i_data_lwM[23]), .B(n142), .C(i_data_lwW[23]), .D(n29), .Q(
        n112) );
  CLKIN6 U22 ( .A(n36), .Q(n115) );
  NAND22 U23 ( .A(n40), .B(n15), .Q(o_data_alusrb[1]) );
  INV3 U24 ( .A(n14), .Q(n15) );
  INV3 U25 ( .A(n16), .Q(n17) );
  NAND33 U26 ( .A(n80), .B(n79), .C(n78), .Q(o_data_alusrb[12]) );
  AOI221 U27 ( .A(i_data_writeres[12]), .B(n138), .C(i_data_alures[12]), .D(
        n23), .Q(n80) );
  NAND33 U28 ( .A(n101), .B(n100), .C(n99), .Q(o_data_alusrb[19]) );
  NAND33 U29 ( .A(n116), .B(n117), .C(n118), .Q(o_data_alusrb[24]) );
  NAND31 U30 ( .A(n121), .B(n119), .C(n120), .Q(o_data_alusrb[25]) );
  AOI221 U31 ( .A(i_data_rt[1]), .B(n115), .C(i_data_writeres[1]), .D(n138), 
        .Q(n42) );
  NAND33 U32 ( .A(n54), .B(n53), .C(n52), .Q(o_data_alusrb[4]) );
  INV2 U33 ( .A(n32), .Q(n1) );
  AOI221 U34 ( .A(i_data_lwM[31]), .B(n1), .C(i_data_lwW[31]), .D(n21), .Q(
        n143) );
  NAND33 U35 ( .A(n71), .B(n70), .C(n69), .Q(o_data_alusrb[9]) );
  AOI221 U36 ( .A(i_data_writeres[11]), .B(n138), .C(i_data_alures[11]), .D(
        n24), .Q(n77) );
  NAND22 U37 ( .A(n39), .B(n37), .Q(n2) );
  INV3 U38 ( .A(n2), .Q(n3) );
  AOI221 U39 ( .A(i_data_writeres[0]), .B(n138), .C(i_data_alures[0]), .D(n23), 
        .Q(n39) );
  NAND21 U40 ( .A(i_data_rt[0]), .B(n115), .Q(n37) );
  NAND22 U41 ( .A(n134), .B(n133), .Q(n4) );
  NAND23 U42 ( .A(n132), .B(n5), .Q(o_data_alusrb[29]) );
  CLKIN3 U43 ( .A(n4), .Q(n5) );
  AOI220 U44 ( .A(i_data_rt[29]), .B(n139), .C(i_data_writeres[29]), .D(n138), 
        .Q(n134) );
  NAND21 U45 ( .A(n19), .B(n67), .Q(n8) );
  NAND22 U46 ( .A(n6), .B(n7), .Q(n9) );
  CLKIN0 U47 ( .A(n19), .Q(n6) );
  INV2 U48 ( .A(n67), .Q(n7) );
  NAND21 U49 ( .A(n19), .B(n67), .Q(n12) );
  NAND24 U50 ( .A(n10), .B(n11), .Q(n13) );
  NAND24 U51 ( .A(n12), .B(n13), .Q(n51) );
  INV1 U52 ( .A(n19), .Q(n10) );
  INV3 U53 ( .A(n67), .Q(n11) );
  CLKIN8 U54 ( .A(n51), .Q(n139) );
  CLKIN12 U55 ( .A(n51), .Q(n125) );
  NAND22 U56 ( .A(n42), .B(n41), .Q(n14) );
  NAND21 U57 ( .A(i_data_alures[1]), .B(n24), .Q(n41) );
  AOI221 U58 ( .A(i_data_rt[23]), .B(n115), .C(i_data_writeres[23]), .D(n138), 
        .Q(n114) );
  AOI222 U59 ( .A(i_data_writeres[5]), .B(n138), .C(i_data_alures[5]), .D(n23), 
        .Q(n57) );
  AOI221 U60 ( .A(i_data_rt[17]), .B(n102), .C(i_data_writeres[17]), .D(n138), 
        .Q(n95) );
  NAND22 U61 ( .A(i_data_rt[11]), .B(n125), .Q(n75) );
  AOI221 U62 ( .A(i_data_lwM[18]), .B(n142), .C(i_data_lwW[18]), .D(n29), .Q(
        n96) );
  NOR21 U63 ( .A(i_con_fb[2]), .B(n26), .Q(n25) );
  CLKIN6 U64 ( .A(i_con_fb[2]), .Q(n46) );
  INV15 U65 ( .A(n30), .Q(n138) );
  NAND24 U66 ( .A(n33), .B(n25), .Q(n30) );
  NAND32 U67 ( .A(i_con_fb[2]), .B(i_con_fb[0]), .C(n33), .Q(n34) );
  AOI221 U68 ( .A(i_data_writeres[8]), .B(n138), .C(i_data_alures[8]), .D(n23), 
        .Q(n66) );
  AOI221 U69 ( .A(i_data_lwM[26]), .B(n142), .C(i_data_lwW[26]), .D(n21), .Q(
        n122) );
  NAND22 U70 ( .A(n47), .B(i_con_fb[2]), .Q(n27) );
  AOI221 U71 ( .A(i_data_lwM[11]), .B(n142), .C(i_data_lwW[11]), .D(n29), .Q(
        n76) );
  NAND33 U72 ( .A(n128), .B(n127), .C(n126), .Q(o_data_alusrb[27]) );
  NAND34 U73 ( .A(n105), .B(n104), .C(n103), .Q(o_data_alusrb[20]) );
  AOI221 U74 ( .A(i_data_writeres[3]), .B(n138), .C(i_data_alures[3]), .D(n24), 
        .Q(n50) );
  AOI221 U75 ( .A(i_data_writeres[2]), .B(n138), .C(i_data_alures[2]), .D(n24), 
        .Q(n45) );
  NAND33 U76 ( .A(n66), .B(n65), .C(n64), .Q(o_data_alusrb[8]) );
  CLKIN15 U77 ( .A(n19), .Q(n33) );
  AOI222 U78 ( .A(i_data_rt[9]), .B(n102), .C(i_data_writeres[9]), .D(n138), 
        .Q(n71) );
  AOI222 U79 ( .A(i_data_lwM[9]), .B(n142), .C(i_data_lwW[9]), .D(n29), .Q(n69) );
  AOI221 U80 ( .A(i_data_lwM[13]), .B(n142), .C(i_data_lwW[13]), .D(n21), .Q(
        n82) );
  CLKIN12 U81 ( .A(n35), .Q(n67) );
  AOI222 U82 ( .A(i_data_lwM[5]), .B(n142), .C(i_data_lwW[5]), .D(n29), .Q(n56) );
  AOI221 U83 ( .A(i_data_lwM[12]), .B(n142), .C(i_data_lwW[12]), .D(n29), .Q(
        n79) );
  AOI221 U84 ( .A(i_data_lwM[3]), .B(n142), .C(i_data_lwW[3]), .D(n29), .Q(n49) );
  AOI221 U85 ( .A(i_data_writeres[10]), .B(n138), .C(i_data_alures[10]), .D(
        n23), .Q(n74) );
  AOI221 U86 ( .A(i_data_lwM[30]), .B(n1), .C(i_data_lwW[30]), .D(n21), .Q(
        n135) );
  AOI222 U87 ( .A(i_data_lwM[20]), .B(n142), .C(i_data_lwW[20]), .D(n21), .Q(
        n103) );
  CLKIN15 U88 ( .A(n20), .Q(n21) );
  AOI222 U89 ( .A(i_data_lwM[16]), .B(n1), .C(i_data_lwW[16]), .D(n21), .Q(n91) );
  AOI221 U90 ( .A(i_data_lwM[21]), .B(n1), .C(i_data_lwW[21]), .D(n21), .Q(
        n106) );
  AOI221 U91 ( .A(i_data_rt[18]), .B(n139), .C(i_data_writeres[18]), .D(n138), 
        .Q(n98) );
  NAND32 U92 ( .A(n111), .B(n110), .C(n109), .Q(o_data_alusrb[22]) );
  AOI221 U93 ( .A(i_data_rt[22]), .B(n139), .C(i_data_writeres[22]), .D(n138), 
        .Q(n111) );
  AOI221 U94 ( .A(i_data_lwM[8]), .B(n142), .C(i_data_lwW[8]), .D(n29), .Q(n65) );
  AOI221 U95 ( .A(i_data_lwM[10]), .B(n142), .C(i_data_lwW[10]), .D(n29), .Q(
        n73) );
  AOI221 U96 ( .A(i_data_writeres[7]), .B(n138), .C(i_data_alures[7]), .D(n24), 
        .Q(n63) );
  CLKIN6 U97 ( .A(i_con_fb[1]), .Q(n18) );
  INV12 U98 ( .A(n18), .Q(n19) );
  NAND22 U99 ( .A(i_data_rt[16]), .B(n139), .Q(n90) );
  NAND34 U100 ( .A(n92), .B(n91), .C(n90), .Q(o_data_alusrb[16]) );
  AOI221 U101 ( .A(i_data_lwM[7]), .B(n142), .C(i_data_lwW[7]), .D(n29), .Q(
        n62) );
  NAND22 U102 ( .A(i_data_rt[10]), .B(n125), .Q(n72) );
  AOI221 U103 ( .A(i_data_lwM[6]), .B(n142), .C(i_data_lwW[6]), .D(n21), .Q(
        n59) );
  NAND22 U104 ( .A(i_data_rt[3]), .B(n125), .Q(n48) );
  AOI221 U105 ( .A(i_data_lwM[2]), .B(n142), .C(i_data_lwW[2]), .D(n21), .Q(
        n44) );
  XNR22 U106 ( .A(n19), .B(n67), .Q(n36) );
  AOI221 U107 ( .A(i_data_lwM[4]), .B(n142), .C(i_data_lwW[4]), .D(n21), .Q(
        n53) );
  NAND21 U108 ( .A(i_data_rt[6]), .B(n125), .Q(n58) );
  AOI221 U109 ( .A(i_data_rt[15]), .B(n102), .C(i_data_writeres[15]), .D(n138), 
        .Q(n89) );
  AOI222 U110 ( .A(i_data_lwM[15]), .B(n142), .C(i_data_lwW[15]), .D(n21), .Q(
        n87) );
  NAND24 U111 ( .A(n47), .B(n46), .Q(n35) );
  NAND22 U112 ( .A(i_data_rt[5]), .B(n115), .Q(n55) );
  CLKIN3 U113 ( .A(i_con_fb[0]), .Q(n26) );
  AOI221 U114 ( .A(i_data_lwM[17]), .B(n142), .C(i_data_lwW[17]), .D(n21), .Q(
        n93) );
  AOI221 U115 ( .A(i_data_lwM[14]), .B(n1), .C(i_data_lwW[14]), .D(n21), .Q(
        n84) );
  AOI220 U116 ( .A(i_data_lwM[29]), .B(n1), .C(i_data_lwW[29]), .D(n21), .Q(
        n132) );
  AOI220 U117 ( .A(i_data_lwM[28]), .B(n142), .C(i_data_lwW[28]), .D(n21), .Q(
        n129) );
  AOI221 U118 ( .A(i_data_lwM[24]), .B(n142), .C(i_data_lwW[24]), .D(n21), .Q(
        n116) );
  NAND33 U119 ( .A(n145), .B(n144), .C(n143), .Q(o_data_alusrb[31]) );
  AOI221 U120 ( .A(i_data_lwM[25]), .B(n142), .C(i_data_lwW[25]), .D(n29), .Q(
        n119) );
  AOI221 U121 ( .A(i_data_rt[25]), .B(n125), .C(i_data_writeres[25]), .D(n138), 
        .Q(n121) );
  CLKBU15 U122 ( .A(n141), .Q(n29) );
  NAND24 U123 ( .A(i_data_rt[12]), .B(n139), .Q(n78) );
  INV2 U124 ( .A(n27), .Q(n28) );
  NAND24 U125 ( .A(n33), .B(n28), .Q(n32) );
  CLKIN6 U126 ( .A(i_con_fb[0]), .Q(n47) );
  AOI220 U127 ( .A(i_data_rt[21]), .B(n139), .C(i_data_writeres[21]), .D(n138), 
        .Q(n108) );
  AOI220 U128 ( .A(i_data_lwM[1]), .B(n142), .C(i_data_lwW[1]), .D(n29), .Q(
        n40) );
  NAND33 U129 ( .A(n50), .B(n49), .C(n48), .Q(o_data_alusrb[3]) );
  AOI220 U130 ( .A(i_data_rt[30]), .B(n139), .C(i_data_writeres[30]), .D(n138), 
        .Q(n137) );
  AOI220 U131 ( .A(i_data_writeres[4]), .B(n138), .C(i_data_alures[4]), .D(n23), .Q(n54) );
  AOI220 U132 ( .A(i_data_lwM[0]), .B(n142), .C(i_data_lwW[0]), .D(n29), .Q(
        n38) );
  AOI220 U133 ( .A(i_data_lwM[22]), .B(n142), .C(i_data_lwW[22]), .D(n29), .Q(
        n109) );
  AOI220 U134 ( .A(i_data_rt[14]), .B(n102), .C(i_data_writeres[14]), .D(n138), 
        .Q(n86) );
  NAND20 U135 ( .A(i_data_alures[14]), .B(n24), .Q(n85) );
  AOI220 U136 ( .A(i_data_lwM[27]), .B(n142), .C(i_data_lwW[27]), .D(n21), .Q(
        n126) );
  AOI220 U137 ( .A(i_data_rt[26]), .B(n139), .C(i_data_writeres[26]), .D(n138), 
        .Q(n124) );
  NAND31 U138 ( .A(n19), .B(n46), .C(n47), .Q(n31) );
  AOI221 U139 ( .A(i_data_rt[31]), .B(n139), .C(i_data_writeres[31]), .D(n138), 
        .Q(n145) );
  NAND31 U140 ( .A(n131), .B(n130), .C(n129), .Q(o_data_alusrb[28]) );
  AOI221 U141 ( .A(i_data_rt[28]), .B(n139), .C(i_data_writeres[28]), .D(n138), 
        .Q(n131) );
  NAND33 U142 ( .A(n86), .B(n85), .C(n84), .Q(o_data_alusrb[14]) );
  NAND33 U143 ( .A(n95), .B(n94), .C(n93), .Q(o_data_alusrb[17]) );
  NAND33 U144 ( .A(n77), .B(n76), .C(n75), .Q(o_data_alusrb[11]) );
  AOI221 U145 ( .A(i_data_writeres[6]), .B(n138), .C(i_data_alures[6]), .D(n24), .Q(n60) );
  AOI221 U146 ( .A(i_data_rt[19]), .B(n102), .C(i_data_writeres[19]), .D(n138), 
        .Q(n101) );
  AOI221 U147 ( .A(i_data_rt[20]), .B(n102), .C(i_data_writeres[20]), .D(n138), 
        .Q(n105) );
  NAND21 U148 ( .A(i_data_alures[20]), .B(n23), .Q(n104) );
  NAND21 U149 ( .A(i_data_alures[19]), .B(n24), .Q(n100) );
  AOI220 U150 ( .A(i_data_rt[27]), .B(n125), .C(i_data_writeres[27]), .D(n138), 
        .Q(n128) );
  NAND21 U151 ( .A(i_data_rt[13]), .B(n125), .Q(n81) );
  AOI221 U152 ( .A(i_data_writeres[16]), .B(n138), .C(i_data_alures[16]), .D(
        n24), .Q(n92) );
  AOI221 U153 ( .A(i_data_rt[24]), .B(n115), .C(i_data_writeres[24]), .D(n138), 
        .Q(n118) );
  NAND22 U154 ( .A(i_data_rt[2]), .B(n115), .Q(n43) );
  NAND22 U155 ( .A(i_data_rt[4]), .B(n139), .Q(n52) );
  NAND22 U156 ( .A(i_data_rt[7]), .B(n125), .Q(n61) );
  NAND22 U157 ( .A(i_data_rt[8]), .B(n125), .Q(n64) );
  NAND22 U158 ( .A(i_data_alures[9]), .B(n23), .Q(n70) );
  NAND33 U159 ( .A(n74), .B(n73), .C(n72), .Q(o_data_alusrb[10]) );
  NAND22 U160 ( .A(i_data_alures[15]), .B(n24), .Q(n88) );
  NAND22 U161 ( .A(i_data_alures[17]), .B(n23), .Q(n94) );
  NAND22 U162 ( .A(i_data_alures[18]), .B(n24), .Q(n97) );
  NAND33 U163 ( .A(n98), .B(n97), .C(n96), .Q(o_data_alusrb[18]) );
  NAND22 U164 ( .A(i_data_alures[21]), .B(n23), .Q(n107) );
  NAND33 U165 ( .A(n108), .B(n107), .C(n106), .Q(o_data_alusrb[21]) );
  NAND22 U166 ( .A(i_data_alures[22]), .B(n23), .Q(n110) );
  NAND22 U167 ( .A(i_data_alures[23]), .B(n23), .Q(n113) );
  NAND22 U168 ( .A(i_data_alures[24]), .B(n23), .Q(n117) );
  NAND22 U169 ( .A(i_data_alures[25]), .B(n24), .Q(n120) );
  NAND22 U170 ( .A(i_data_alures[26]), .B(n24), .Q(n123) );
  NAND33 U171 ( .A(n124), .B(n123), .C(n122), .Q(o_data_alusrb[26]) );
  NAND22 U172 ( .A(i_data_alures[27]), .B(n23), .Q(n127) );
  NAND22 U173 ( .A(i_data_alures[28]), .B(n24), .Q(n130) );
  NAND22 U174 ( .A(i_data_alures[29]), .B(n23), .Q(n133) );
  NAND22 U175 ( .A(i_data_alures[30]), .B(n24), .Q(n136) );
  NAND33 U176 ( .A(n137), .B(n136), .C(n135), .Q(o_data_alusrb[30]) );
  NAND22 U177 ( .A(i_data_alures[31]), .B(n23), .Q(n144) );
endmodule


module E_alubmux ( i_data_fb, i_data_imm, i_con_imm, o_data_alub );
  input [31:0] i_data_fb;
  input [31:0] i_data_imm;
  output [31:0] o_data_alub;
  input i_con_imm;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;

  INV12 U1 ( .A(n34), .Q(o_data_alub[15]) );
  CLKIN15 U2 ( .A(n36), .Q(o_data_alub[17]) );
  CLKIN12 U3 ( .A(n31), .Q(o_data_alub[12]) );
  CLKIN12 U4 ( .A(n33), .Q(o_data_alub[14]) );
  INV8 U5 ( .A(n18), .Q(o_data_alub[5]) );
  CLKIN12 U6 ( .A(n42), .Q(o_data_alub[23]) );
  INV6 U7 ( .A(n44), .Q(o_data_alub[26]) );
  AOI221 U8 ( .A(i_data_fb[26]), .B(n8), .C(i_data_imm[26]), .D(n4), .Q(n44)
         );
  NAND22 U9 ( .A(n2), .B(n3), .Q(o_data_alub[31]) );
  CLKIN6 U10 ( .A(n32), .Q(o_data_alub[13]) );
  AOI221 U11 ( .A(i_data_fb[18]), .B(n7), .C(i_data_imm[18]), .D(n4), .Q(n37)
         );
  INV8 U12 ( .A(n30), .Q(o_data_alub[11]) );
  BUF6 U13 ( .A(n5), .Q(n1) );
  INV6 U14 ( .A(n41), .Q(o_data_alub[22]) );
  CLKIN6 U15 ( .A(n38), .Q(o_data_alub[19]) );
  CLKIN6 U16 ( .A(n37), .Q(o_data_alub[18]) );
  INV6 U17 ( .A(n40), .Q(o_data_alub[21]) );
  INV6 U18 ( .A(n29), .Q(o_data_alub[10]) );
  CLKIN6 U19 ( .A(n24), .Q(o_data_alub[7]) );
  INV6 U20 ( .A(n28), .Q(o_data_alub[9]) );
  CLKIN15 U21 ( .A(n35), .Q(o_data_alub[16]) );
  INV8 U22 ( .A(n11), .Q(o_data_alub[0]) );
  BUF8 U23 ( .A(n10), .Q(n6) );
  INV6 U24 ( .A(n14), .Q(o_data_alub[3]) );
  INV6 U25 ( .A(n43), .Q(o_data_alub[24]) );
  CLKIN15 U26 ( .A(n39), .Q(o_data_alub[20]) );
  MUX21 U27 ( .A(i_data_fb[28]), .B(i_data_imm[28]), .S(n4), .Q(
        o_data_alub[28]) );
  MUX21 U28 ( .A(i_data_fb[29]), .B(i_data_imm[29]), .S(n4), .Q(
        o_data_alub[29]) );
  NAND20 U29 ( .A(i_data_fb[31]), .B(n9), .Q(n2) );
  NAND20 U30 ( .A(i_data_imm[31]), .B(n4), .Q(n3) );
  CLKIN3 U31 ( .A(n6), .Q(n4) );
  NAND20 U32 ( .A(i_data_imm[6]), .B(n5), .Q(n19) );
  INV6 U33 ( .A(n21), .Q(o_data_alub[6]) );
  INV3 U34 ( .A(n6), .Q(n5) );
  INV8 U35 ( .A(n12), .Q(o_data_alub[1]) );
  NAND20 U36 ( .A(i_data_imm[8]), .B(n5), .Q(n25) );
  INV8 U37 ( .A(n27), .Q(o_data_alub[8]) );
  INV8 U38 ( .A(n13), .Q(o_data_alub[2]) );
  AOI222 U39 ( .A(i_data_fb[22]), .B(n7), .C(i_data_imm[22]), .D(n4), .Q(n41)
         );
  AOI222 U40 ( .A(i_data_fb[21]), .B(n7), .C(i_data_imm[21]), .D(n4), .Q(n40)
         );
  AOI222 U41 ( .A(i_data_fb[13]), .B(n8), .C(i_data_imm[13]), .D(n1), .Q(n32)
         );
  CLKIN3 U42 ( .A(i_con_imm), .Q(n10) );
  BUF2 U43 ( .A(n10), .Q(n7) );
  BUF2 U44 ( .A(n6), .Q(n8) );
  BUF2 U45 ( .A(n6), .Q(n9) );
  INV8 U46 ( .A(n17), .Q(o_data_alub[4]) );
  AOI222 U47 ( .A(i_data_fb[0]), .B(n6), .C(i_data_imm[0]), .D(n4), .Q(n11) );
  AOI222 U48 ( .A(i_data_fb[1]), .B(n9), .C(i_data_imm[1]), .D(n1), .Q(n12) );
  AOI222 U49 ( .A(i_data_fb[2]), .B(n9), .C(i_data_imm[2]), .D(n1), .Q(n13) );
  AOI222 U50 ( .A(i_data_fb[3]), .B(n9), .C(i_data_imm[3]), .D(n1), .Q(n14) );
  NAND22 U51 ( .A(i_data_imm[4]), .B(n1), .Q(n15) );
  CLKIN3 U52 ( .A(n15), .Q(n16) );
  OAI222 U53 ( .A(i_data_fb[4]), .B(n16), .C(n16), .D(n9), .Q(n17) );
  AOI222 U54 ( .A(i_data_fb[5]), .B(n8), .C(i_data_imm[5]), .D(n1), .Q(n18) );
  CLKIN3 U55 ( .A(n19), .Q(n20) );
  OAI222 U56 ( .A(n20), .B(n9), .C(i_data_fb[6]), .D(n20), .Q(n21) );
  NAND22 U57 ( .A(i_data_imm[7]), .B(n1), .Q(n22) );
  CLKIN3 U58 ( .A(n22), .Q(n23) );
  OAI222 U59 ( .A(n23), .B(n8), .C(i_data_fb[7]), .D(n23), .Q(n24) );
  CLKIN3 U60 ( .A(n25), .Q(n26) );
  OAI222 U61 ( .A(n26), .B(n7), .C(i_data_fb[8]), .D(n26), .Q(n27) );
  AOI222 U62 ( .A(i_data_fb[9]), .B(n8), .C(i_data_imm[9]), .D(n1), .Q(n28) );
  AOI222 U63 ( .A(i_data_fb[10]), .B(n8), .C(i_data_imm[10]), .D(n1), .Q(n29)
         );
  AOI222 U64 ( .A(i_data_fb[11]), .B(n8), .C(i_data_imm[11]), .D(n1), .Q(n30)
         );
  AOI222 U65 ( .A(i_data_fb[12]), .B(n8), .C(i_data_imm[12]), .D(n1), .Q(n31)
         );
  AOI222 U66 ( .A(i_data_fb[14]), .B(n8), .C(i_data_imm[14]), .D(n1), .Q(n33)
         );
  AOI222 U67 ( .A(i_data_fb[15]), .B(n7), .C(i_data_imm[15]), .D(n1), .Q(n34)
         );
  AOI222 U68 ( .A(i_data_fb[16]), .B(n7), .C(i_data_imm[16]), .D(n1), .Q(n35)
         );
  AOI222 U69 ( .A(i_data_fb[17]), .B(n7), .C(i_data_imm[17]), .D(n4), .Q(n36)
         );
  AOI222 U70 ( .A(i_data_fb[19]), .B(n7), .C(i_data_imm[19]), .D(n4), .Q(n38)
         );
  AOI222 U71 ( .A(i_data_fb[20]), .B(n7), .C(i_data_imm[20]), .D(n4), .Q(n39)
         );
  AOI222 U72 ( .A(i_data_fb[23]), .B(n6), .C(i_data_imm[23]), .D(n4), .Q(n42)
         );
  AOI222 U73 ( .A(i_data_fb[24]), .B(n6), .C(i_data_imm[24]), .D(n4), .Q(n43)
         );
  MUX26 U74 ( .A(i_data_fb[25]), .B(i_data_imm[25]), .S(n4), .Q(
        o_data_alub[25]) );
  MUX26 U75 ( .A(i_data_fb[27]), .B(i_data_imm[27]), .S(n4), .Q(
        o_data_alub[27]) );
  MUX26 U76 ( .A(i_data_fb[30]), .B(i_data_imm[30]), .S(n4), .Q(
        o_data_alub[30]) );
endmodule


module E_rdmux ( i_data_rtE, i_data_rdE, i_con_regdst, i_con_aluPC4, 
        o_data_writeE );
  input [4:0] i_data_rtE;
  input [4:0] i_data_rdE;
  output [4:0] o_data_writeE;
  input i_con_regdst, i_con_aluPC4;
  wire   n7, n8, n9, n10, n11, n1, n2, n3, n4, n5, n6;

  OAI2111 U2 ( .A(i_con_regdst), .B(n5), .C(n6), .D(n11), .Q(o_data_writeE[0])
         );
  INV3 U3 ( .A(i_data_rtE[0]), .Q(n5) );
  NAND22 U4 ( .A(i_data_rdE[0]), .B(i_con_regdst), .Q(n11) );
  OAI2111 U5 ( .A(i_con_regdst), .B(n4), .C(n6), .D(n10), .Q(o_data_writeE[1])
         );
  INV3 U6 ( .A(i_data_rtE[1]), .Q(n4) );
  NAND22 U7 ( .A(i_data_rdE[1]), .B(i_con_regdst), .Q(n10) );
  OAI2111 U8 ( .A(i_con_regdst), .B(n3), .C(n6), .D(n9), .Q(o_data_writeE[2])
         );
  INV3 U9 ( .A(i_data_rtE[2]), .Q(n3) );
  NAND22 U10 ( .A(i_data_rdE[2]), .B(i_con_regdst), .Q(n9) );
  OAI2111 U11 ( .A(i_con_regdst), .B(n2), .C(n6), .D(n8), .Q(o_data_writeE[3])
         );
  INV3 U12 ( .A(i_data_rtE[3]), .Q(n2) );
  NAND22 U13 ( .A(i_data_rdE[3]), .B(i_con_regdst), .Q(n8) );
  OAI2111 U14 ( .A(i_con_regdst), .B(n1), .C(n6), .D(n7), .Q(o_data_writeE[4])
         );
  INV3 U15 ( .A(i_data_rtE[4]), .Q(n1) );
  NAND22 U16 ( .A(i_data_rdE[4]), .B(i_con_regdst), .Q(n7) );
  INV3 U17 ( .A(i_con_aluPC4), .Q(n6) );
endmodule


module D_compare_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166;

  NAND22 U1 ( .A(B[3]), .B(n55), .Q(n54) );
  CLKIN3 U2 ( .A(B[28]), .Q(n85) );
  INV1 U3 ( .A(B[15]), .Q(n40) );
  INV0 U4 ( .A(B[3]), .Q(n161) );
  NOR21 U5 ( .A(n51), .B(n52), .Q(n50) );
  INV3 U6 ( .A(A[6]), .Q(n56) );
  NOR22 U7 ( .A(n2), .B(n8), .Q(n4) );
  NAND20 U8 ( .A(B[20]), .B(n98), .Q(n97) );
  NAND23 U9 ( .A(n135), .B(n136), .Q(n129) );
  NAND22 U10 ( .A(A[25]), .B(n137), .Q(n136) );
  INV1 U11 ( .A(A[23]), .Q(n109) );
  INV3 U12 ( .A(B[25]), .Q(n137) );
  NAND22 U13 ( .A(n126), .B(n127), .Q(n7) );
  NAND22 U14 ( .A(n131), .B(n132), .Q(n130) );
  NAND22 U15 ( .A(A[22]), .B(n133), .Q(n132) );
  INV3 U16 ( .A(A[0]), .Q(n86) );
  NAND22 U17 ( .A(n152), .B(n153), .Q(n16) );
  INV3 U18 ( .A(A[2]), .Q(n59) );
  NOR21 U19 ( .A(n149), .B(n148), .Q(n124) );
  INV0 U20 ( .A(A[16]), .Q(n47) );
  CLKIN3 U21 ( .A(B[16]), .Q(n166) );
  NAND22 U22 ( .A(A[3]), .B(n161), .Q(n23) );
  NAND22 U23 ( .A(A[16]), .B(n166), .Q(n12) );
  INV3 U24 ( .A(A[5]), .Q(n69) );
  NAND22 U25 ( .A(A[8]), .B(n162), .Q(n22) );
  NOR21 U26 ( .A(n7), .B(n9), .Q(n1) );
  INV3 U27 ( .A(n1), .Q(n2) );
  NAND34 U28 ( .A(n3), .B(n4), .C(n5), .Q(NE) );
  XNR22 U29 ( .A(B[31]), .B(A[31]), .Q(n155) );
  INV3 U30 ( .A(A[19]), .Q(n99) );
  NAND21 U31 ( .A(A[23]), .B(n134), .Q(n131) );
  INV2 U32 ( .A(A[13]), .Q(n48) );
  XNR22 U33 ( .A(B[30]), .B(A[30]), .Q(n156) );
  NOR21 U34 ( .A(A[1]), .B(n80), .Q(n79) );
  NAND21 U35 ( .A(B[2]), .B(n59), .Q(n58) );
  NAND21 U36 ( .A(A[20]), .B(n143), .Q(n142) );
  NOR21 U37 ( .A(B[0]), .B(n86), .Q(n122) );
  INV1 U38 ( .A(B[22]), .Q(n133) );
  NAND21 U39 ( .A(A[13]), .B(n154), .Q(n152) );
  CLKIN1 U40 ( .A(A[24]), .Q(n108) );
  INV6 U41 ( .A(A[12]), .Q(n66) );
  INV2 U42 ( .A(A[3]), .Q(n55) );
  INV0 U43 ( .A(B[10]), .Q(n117) );
  AOI2110 U44 ( .A(B[10]), .B(n77), .C(n78), .D(n79), .Q(n76) );
  NOR21 U45 ( .A(A[14]), .B(n45), .Q(n44) );
  NAND22 U46 ( .A(A[14]), .B(n45), .Q(n21) );
  INV1 U47 ( .A(B[14]), .Q(n45) );
  NAND21 U48 ( .A(B[29]), .B(n87), .Q(n73) );
  INV2 U49 ( .A(B[29]), .Q(n144) );
  AOI2110 U50 ( .A(A[10]), .B(n117), .C(n118), .D(n119), .Q(n112) );
  AOI2110 U51 ( .A(A[1]), .B(n80), .C(n122), .D(n123), .Q(n121) );
  AOI2112 U52 ( .A(A[24]), .B(n128), .C(n129), .D(n130), .Q(n127) );
  CLKIN0 U53 ( .A(A[10]), .Q(n77) );
  NAND22 U54 ( .A(n112), .B(n113), .Q(n24) );
  NAND22 U55 ( .A(n13), .B(n12), .Q(n163) );
  NAND22 U56 ( .A(n11), .B(n10), .Q(n164) );
  CLKIN0 U57 ( .A(B[11]), .Q(n46) );
  NOR20 U58 ( .A(A[9]), .B(n81), .Q(n78) );
  NAND20 U59 ( .A(B[4]), .B(n60), .Q(n57) );
  CLKIN0 U60 ( .A(A[21]), .Q(n95) );
  CLKIN3 U61 ( .A(n121), .Q(n25) );
  NOR31 U62 ( .A(n114), .B(n115), .C(n116), .Q(n113) );
  INV0 U63 ( .A(A[25]), .Q(n105) );
  INV1 U64 ( .A(B[1]), .Q(n80) );
  CLKIN0 U65 ( .A(B[20]), .Q(n143) );
  NAND21 U66 ( .A(A[15]), .B(n40), .Q(n20) );
  NAND20 U67 ( .A(B[0]), .B(n86), .Q(n74) );
  NAND22 U68 ( .A(A[17]), .B(n41), .Q(n13) );
  INV3 U69 ( .A(A[7]), .Q(n65) );
  CLKIN0 U70 ( .A(B[21]), .Q(n138) );
  NAND22 U71 ( .A(B[8]), .B(n70), .Q(n67) );
  NAND21 U72 ( .A(B[19]), .B(n99), .Q(n96) );
  NAND22 U73 ( .A(B[24]), .B(n108), .Q(n107) );
  NAND22 U74 ( .A(n124), .B(n125), .Q(n27) );
  NAND40 U75 ( .A(n10), .B(n11), .C(n12), .D(n13), .Q(n9) );
  NOR23 U76 ( .A(n71), .B(n72), .Q(n29) );
  INV1 U77 ( .A(n7), .Q(n125) );
  NOR20 U78 ( .A(B[5]), .B(n69), .Q(n114) );
  CLKIN2 U79 ( .A(B[26]), .Q(n147) );
  NAND20 U80 ( .A(B[5]), .B(n69), .Q(n68) );
  NOR20 U81 ( .A(B[12]), .B(n66), .Q(n118) );
  NOR20 U82 ( .A(B[7]), .B(n65), .Q(n119) );
  INV0 U83 ( .A(B[8]), .Q(n162) );
  NAND20 U84 ( .A(A[9]), .B(n81), .Q(n26) );
  NOR20 U85 ( .A(B[6]), .B(n56), .Q(n115) );
  CLKIN3 U86 ( .A(B[13]), .Q(n154) );
  INV0 U87 ( .A(B[19]), .Q(n165) );
  NAND20 U88 ( .A(B[7]), .B(n65), .Q(n64) );
  NAND20 U89 ( .A(B[12]), .B(n66), .Q(n63) );
  INV0 U90 ( .A(B[9]), .Q(n81) );
  NAND20 U91 ( .A(B[23]), .B(n109), .Q(n106) );
  CLKIN0 U92 ( .A(B[23]), .Q(n134) );
  CLKIN0 U93 ( .A(B[24]), .Q(n128) );
  NAND42 U94 ( .A(n33), .B(n34), .C(n35), .D(n36), .Q(n32) );
  NAND22 U95 ( .A(B[13]), .B(n48), .Q(n33) );
  NOR31 U96 ( .A(n37), .B(n38), .C(n39), .Q(n36) );
  NAND22 U97 ( .A(n22), .B(n23), .Q(n18) );
  NAND22 U98 ( .A(n14), .B(n15), .Q(n8) );
  NOR21 U99 ( .A(n18), .B(n19), .Q(n14) );
  NOR21 U100 ( .A(n16), .B(n17), .Q(n15) );
  NAND22 U101 ( .A(n20), .B(n21), .Q(n19) );
  NAND22 U102 ( .A(n88), .B(n89), .Q(n71) );
  NOR21 U103 ( .A(n90), .B(n91), .Q(n89) );
  NOR21 U104 ( .A(n100), .B(n101), .Q(n88) );
  NAND22 U105 ( .A(n92), .B(n93), .Q(n91) );
  NAND22 U106 ( .A(n110), .B(n111), .Q(n28) );
  NOR21 U107 ( .A(n25), .B(n120), .Q(n110) );
  NAND22 U108 ( .A(n49), .B(n50), .Q(n31) );
  NOR21 U109 ( .A(n61), .B(n62), .Q(n49) );
  NAND22 U110 ( .A(n63), .B(n64), .Q(n62) );
  NOR21 U111 ( .A(n159), .B(n160), .Q(n158) );
  NAND22 U112 ( .A(n20), .B(n21), .Q(n160) );
  NAND22 U113 ( .A(n22), .B(n23), .Q(n159) );
  NOR21 U114 ( .A(n163), .B(n164), .Q(n157) );
  NAND22 U115 ( .A(n150), .B(n151), .Q(n149) );
  NAND22 U116 ( .A(n157), .B(n158), .Q(n148) );
  NOR21 U117 ( .A(A[17]), .B(n41), .Q(n38) );
  INV3 U118 ( .A(A[4]), .Q(n60) );
  NAND22 U119 ( .A(n155), .B(n156), .Q(n17) );
  AOI2111 U120 ( .A(A[21]), .B(n138), .C(n139), .D(n140), .Q(n126) );
  NAND22 U121 ( .A(n141), .B(n142), .Q(n140) );
  NAND22 U122 ( .A(n67), .B(n68), .Q(n61) );
  NAND22 U123 ( .A(n57), .B(n58), .Q(n51) );
  NAND22 U124 ( .A(n106), .B(n107), .Q(n100) );
  NAND22 U125 ( .A(n96), .B(n97), .Q(n90) );
  INV3 U126 ( .A(A[20]), .Q(n98) );
  NAND22 U127 ( .A(B[22]), .B(n94), .Q(n93) );
  NAND22 U128 ( .A(n102), .B(n103), .Q(n101) );
  NAND22 U129 ( .A(B[25]), .B(n105), .Q(n102) );
  NAND22 U130 ( .A(B[26]), .B(n104), .Q(n103) );
  NAND22 U131 ( .A(n53), .B(n54), .Q(n52) );
  NOR21 U132 ( .A(B[4]), .B(n60), .Q(n116) );
  NAND22 U133 ( .A(n145), .B(n146), .Q(n139) );
  NAND22 U134 ( .A(B[16]), .B(n47), .Q(n34) );
  NAND22 U135 ( .A(B[21]), .B(n95), .Q(n92) );
  INV3 U136 ( .A(B[18]), .Q(n42) );
  INV3 U137 ( .A(B[27]), .Q(n84) );
  NOR21 U138 ( .A(n43), .B(n44), .Q(n35) );
  NOR23 U139 ( .A(n31), .B(n32), .Q(n30) );
  INV6 U140 ( .A(n6), .Q(n5) );
  INV3 U141 ( .A(A[22]), .Q(n94) );
  NAND22 U142 ( .A(A[19]), .B(n165), .Q(n11) );
  NAND42 U143 ( .A(n73), .B(n74), .C(n75), .D(n76), .Q(n72) );
  NOR21 U144 ( .A(n82), .B(n83), .Q(n75) );
  NOR21 U145 ( .A(A[28]), .B(n85), .Q(n82) );
  NAND22 U146 ( .A(A[28]), .B(n85), .Q(n135) );
  NAND22 U147 ( .A(A[18]), .B(n42), .Q(n10) );
  NOR21 U148 ( .A(A[18]), .B(n42), .Q(n37) );
  NAND22 U149 ( .A(A[27]), .B(n84), .Q(n145) );
  NOR21 U150 ( .A(A[27]), .B(n84), .Q(n83) );
  INV3 U151 ( .A(A[26]), .Q(n104) );
  NAND22 U152 ( .A(A[29]), .B(n144), .Q(n141) );
  INV3 U153 ( .A(A[29]), .Q(n87) );
  NOR31 U154 ( .A(n24), .B(n25), .C(n120), .Q(n3) );
  NAND22 U155 ( .A(A[26]), .B(n147), .Q(n146) );
  NAND22 U156 ( .A(A[11]), .B(n46), .Q(n153) );
  NOR21 U157 ( .A(A[11]), .B(n46), .Q(n43) );
  INV3 U158 ( .A(A[8]), .Q(n70) );
  INV3 U159 ( .A(n24), .Q(n111) );
  NOR21 U160 ( .A(B[2]), .B(n59), .Q(n123) );
  NOR21 U161 ( .A(A[15]), .B(n40), .Q(n39) );
  INV3 U162 ( .A(n17), .Q(n150) );
  NAND21 U163 ( .A(B[6]), .B(n56), .Q(n53) );
  INV1 U164 ( .A(B[17]), .Q(n41) );
  NOR33 U165 ( .A(n27), .B(n28), .C(n6), .Q(EQ) );
  NAND24 U166 ( .A(n29), .B(n30), .Q(n6) );
  CLKIN3 U167 ( .A(n26), .Q(n120) );
  CLKIN3 U168 ( .A(n16), .Q(n151) );
endmodule


module D_compare ( o_con_ifbranch, i_data_rs, i_data_rt, i_con_bop );
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [2:0] i_con_bop;
  output o_con_ifbranch;
  wire   N32, N33, n4, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n1,
         n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  D_compare_DW01_cmp6_1 r49 ( .A(i_data_rs), .B(i_data_rt), .TC(n4), .EQ(N32), 
        .NE(N33) );
  CLKIN3 U2 ( .A(n1), .Q(n2) );
  NOR22 U3 ( .A(n18), .B(n17), .Q(n9) );
  NOR22 U4 ( .A(i_data_rs[25]), .B(i_data_rs[23]), .Q(n1) );
  NOR30 U5 ( .A(n2), .B(i_data_rs[24]), .C(i_data_rs[26]), .Q(n23) );
  INV1 U6 ( .A(i_data_rs[31]), .Q(n5) );
  IMUX24 U7 ( .A(N32), .B(i_data_rs[31]), .S(i_con_bop[2]), .Q(n10) );
  NOR30 U8 ( .A(i_data_rs[0]), .B(i_data_rs[11]), .C(i_data_rs[10]), .Q(n19)
         );
  NOR40 U9 ( .A(i_data_rs[19]), .B(i_data_rs[18]), .C(i_data_rs[17]), .D(
        i_data_rs[16]), .Q(n21) );
  NOR40 U10 ( .A(i_data_rs[9]), .B(i_data_rs[8]), .C(i_data_rs[7]), .D(
        i_data_rs[6]), .Q(n26) );
  NOR40 U11 ( .A(i_data_rs[5]), .B(i_data_rs[4]), .C(i_data_rs[3]), .D(
        i_data_rs[30]), .Q(n25) );
  NOR40 U12 ( .A(i_data_rs[15]), .B(i_data_rs[14]), .C(i_data_rs[13]), .D(
        i_data_rs[12]), .Q(n20) );
  NOR40 U13 ( .A(i_data_rs[22]), .B(i_data_rs[21]), .C(i_data_rs[20]), .D(
        i_data_rs[1]), .Q(n22) );
  NOR40 U14 ( .A(i_data_rs[2]), .B(i_data_rs[29]), .C(i_data_rs[28]), .D(
        i_data_rs[27]), .Q(n24) );
  IMUX22 U15 ( .A(n11), .B(n12), .S(n3), .Q(n13) );
  INV3 U16 ( .A(i_con_bop[0]), .Q(n3) );
  LOGIC0 U17 ( .Q(n4) );
  NAND42 U18 ( .A(n23), .B(n24), .C(n25), .D(n26), .Q(n17) );
  NAND42 U19 ( .A(n19), .B(n20), .C(n21), .D(n22), .Q(n18) );
  NOR24 U20 ( .A(i_con_bop[1]), .B(n10), .Q(n11) );
  CLKIN3 U21 ( .A(n9), .Q(n6) );
  NAND22 U22 ( .A(n6), .B(n5), .Q(n7) );
  IMUX23 U23 ( .A(N33), .B(n7), .S(i_con_bop[0]), .Q(n15) );
  CLKIN3 U24 ( .A(i_con_bop[1]), .Q(n14) );
  CLKIN3 U25 ( .A(i_con_bop[2]), .Q(n8) );
  AOI2112 U26 ( .A(n9), .B(n14), .C(i_data_rs[31]), .D(n8), .Q(n12) );
  OAI312 U27 ( .A(i_con_bop[2]), .B(n15), .C(n14), .D(n13), .Q(o_con_ifbranch)
         );
endmodule


module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Efamux, i_con_Efbmux, 
        i_con_Ealuop, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread, 
        i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_bop, o_data_pc4, o_data_alures, o_data_rt, o_addr_regdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_addr_Erd, o_addr_Mrt, o_con_ifbranch );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [5:0] i_con_Ealuop;
  input [2:0] i_con_bop;
  output [31:0] o_data_pc4;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [31:0] alu_o_data_AluRes;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;

  DFC3 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[0]) );
  DFC3 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC3 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  DFC3 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC3 pipe_rt_reg_25_ ( .D(compare_i_data_rt[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[25]) );
  DFC3 pipe_rt_reg_24_ ( .D(compare_i_data_rt[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[24]) );
  DFC3 pipe_rt_reg_22_ ( .D(compare_i_data_rt[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[22]) );
  DFC3 pipe_rt_reg_21_ ( .D(compare_i_data_rt[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[21]) );
  DFC3 pipe_rt_reg_19_ ( .D(compare_i_data_rt[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[19]) );
  DFC3 pipe_rt_reg_18_ ( .D(compare_i_data_rt[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[18]) );
  DFC3 pipe_rt_reg_17_ ( .D(compare_i_data_rt[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[17]) );
  DFC3 pipe_rt_reg_16_ ( .D(compare_i_data_rt[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[16]) );
  DFC3 pipe_rt_reg_15_ ( .D(compare_i_data_rt[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[15]) );
  DFC3 pipe_rt_reg_14_ ( .D(compare_i_data_rt[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[14]) );
  DFC3 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC3 pipe_rt_reg_11_ ( .D(compare_i_data_rt[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[11]) );
  DFC3 pipe_rt_reg_10_ ( .D(compare_i_data_rt[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[10]) );
  DFC3 pipe_rt_reg_9_ ( .D(compare_i_data_rt[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[9]) );
  DFC3 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC3 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC3 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC3 pipe_rt_reg_5_ ( .D(compare_i_data_rt[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[5]) );
  DFC3 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(compare_i_data_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[2]) );
  DFC3 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC3 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC3 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC3 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC3 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC3 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Malupc8_reg ( .D(i_con_Malupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Malupc8) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  E_alu u_alu ( .o_data_AluRes(alu_o_data_AluRes), .i_data_A({
        compare_i_data_rs[31], n1, compare_i_data_rs[29], n10, 
        compare_i_data_rs[27:26], n7, n3, compare_i_data_rs[23:13], n4, 
        compare_i_data_rs[11:6], n6, compare_i_data_rs[4:3], n11, 
        compare_i_data_rs[1:0]}), .i_data_B({alu_i_data_B[31:29], n8, 
        alu_i_data_B[27:0]}), .i_con_AluCtrl(alu_i_con_AluCtrl), 
        .i_data_shamt(i_data_immext[10:6]) );
  E_alu_control u_alu_control ( .o_con_AluCtrl(alu_i_con_AluCtrl), 
        .i_con_AluOp(i_con_Ealuop), .i_con_FuncCode(i_data_immext[5:0]) );
  E_famux5 u_famux5 ( .i_data_rs(i_data_rs), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fa(i_con_Efamux), .o_data_alusra(
        compare_i_data_rs) );
  E_fbmux5 u_fbmux ( .i_data_rt(i_data_rt), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fb(i_con_Efbmux), .o_data_alusrb(
        compare_i_data_rt) );
  E_alubmux u_alubmux ( .i_data_fb(compare_i_data_rt), .i_data_imm(
        i_data_immext), .i_con_imm(i_con_Ealusrc), .o_data_alub(alu_i_data_B)
         );
  E_rdmux u_rdmux ( .i_data_rtE(i_addr_rt), .i_data_rdE(i_addr_rd), 
        .i_con_regdst(i_con_Eregdst), .i_con_aluPC4(i_con_Malupc8), 
        .o_data_writeE(o_addr_Erd) );
  D_compare u_compare ( .o_con_ifbranch(o_con_ifbranch), .i_data_rs({
        compare_i_data_rs[31], n1, compare_i_data_rs[29], n10, 
        compare_i_data_rs[27:26], n7, n3, compare_i_data_rs[23:13], n4, 
        compare_i_data_rs[11:6], n6, compare_i_data_rs[4:3], n11, 
        compare_i_data_rs[1:0]}), .i_data_rt({compare_i_data_rt[31:14], n12, 
        compare_i_data_rt[12:0]}), .i_con_bop(i_con_bop) );
  DFC1 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC1 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC1 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC1 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC1 pipe_alures_reg_13_ ( .D(alu_o_data_AluRes[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[13]) );
  DFC1 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC1 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC1 pipe_rt_reg_28_ ( .D(compare_i_data_rt[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[28]) );
  DFC1 pipe_rt_reg_13_ ( .D(n12), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC1 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC1 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC1 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC1 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC1 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC1 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC1 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  DFC1 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC1 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC1 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC1 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC1 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC1 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC1 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC1 pipe_alures_reg_15_ ( .D(alu_o_data_AluRes[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[15]) );
  DFC1 pipe_alures_reg_14_ ( .D(alu_o_data_AluRes[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[14]) );
  DFC1 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC1 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC1 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC1 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC1 pipe_rt_reg_23_ ( .D(compare_i_data_rt[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[23]) );
  DFC1 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC1 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC1 pipe_rt_reg_0_ ( .D(compare_i_data_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[0]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC1 pipe_rt_reg_20_ ( .D(compare_i_data_rt[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[20]) );
  BUF6 U3 ( .A(compare_i_data_rs[2]), .Q(n11) );
  INV8 U4 ( .A(n2), .Q(n3) );
  BUF6 U5 ( .A(compare_i_data_rs[30]), .Q(n1) );
  INV6 U6 ( .A(n9), .Q(n10) );
  INV3 U7 ( .A(compare_i_data_rs[28]), .Q(n9) );
  INV3 U8 ( .A(compare_i_data_rs[5]), .Q(n5) );
  INV3 U9 ( .A(compare_i_data_rs[24]), .Q(n2) );
  BUF8 U10 ( .A(compare_i_data_rs[25]), .Q(n7) );
  INV6 U11 ( .A(n5), .Q(n6) );
  BUF15 U12 ( .A(compare_i_data_rs[12]), .Q(n4) );
  BUF12 U13 ( .A(alu_i_data_B[28]), .Q(n8) );
  BUF2 U14 ( .A(compare_i_data_rt[13]), .Q(n12) );
endmodule


module M_resmux ( i_data_alures, i_data_pc8, i_con_pc8, o_data_alu );
  input [31:0] i_data_alures;
  input [31:0] i_data_pc8;
  output [31:0] o_data_alu;
  input i_con_pc8;
  wire   n34, n35, n36, n37, n38, n39, n40, n43, n54, n60, n61, n62, n63, n64,
         n65, n1;

  INV3 U1 ( .A(n38), .Q(o_data_alu[5]) );
  INV3 U2 ( .A(n40), .Q(o_data_alu[3]) );
  INV3 U3 ( .A(n36), .Q(o_data_alu[7]) );
  INV3 U4 ( .A(n64), .Q(o_data_alu[10]) );
  INV3 U5 ( .A(n63), .Q(o_data_alu[11]) );
  INV3 U6 ( .A(n61), .Q(o_data_alu[13]) );
  INV3 U7 ( .A(n60), .Q(o_data_alu[14]) );
  MUX22 U8 ( .A(i_data_alures[30]), .B(i_data_pc8[30]), .S(i_con_pc8), .Q(
        o_data_alu[30]) );
  AOI220 U9 ( .A(i_data_alures[14]), .B(n1), .C(i_data_pc8[14]), .D(i_con_pc8), 
        .Q(n60) );
  AOI220 U10 ( .A(i_data_alures[12]), .B(n1), .C(i_data_pc8[12]), .D(i_con_pc8), .Q(n62) );
  AOI220 U11 ( .A(i_data_alures[7]), .B(n1), .C(i_data_pc8[7]), .D(i_con_pc8), 
        .Q(n36) );
  AOI221 U12 ( .A(i_data_alures[5]), .B(n1), .C(i_data_pc8[5]), .D(i_con_pc8), 
        .Q(n38) );
  AOI221 U13 ( .A(i_data_alures[10]), .B(n1), .C(i_data_pc8[10]), .D(i_con_pc8), .Q(n64) );
  AOI221 U14 ( .A(i_data_alures[11]), .B(n1), .C(i_data_pc8[11]), .D(i_con_pc8), .Q(n63) );
  AOI220 U15 ( .A(i_data_alures[13]), .B(n1), .C(i_data_pc8[13]), .D(i_con_pc8), .Q(n61) );
  AOI220 U16 ( .A(i_data_alures[2]), .B(n1), .C(i_data_pc8[2]), .D(i_con_pc8), 
        .Q(n43) );
  AOI220 U17 ( .A(i_data_alures[3]), .B(n1), .C(i_data_pc8[3]), .D(i_con_pc8), 
        .Q(n40) );
  MUX22 U18 ( .A(i_data_alures[23]), .B(i_data_pc8[23]), .S(i_con_pc8), .Q(
        o_data_alu[23]) );
  MUX22 U19 ( .A(i_data_alures[27]), .B(i_data_pc8[27]), .S(i_con_pc8), .Q(
        o_data_alu[27]) );
  MUX22 U20 ( .A(i_data_alures[17]), .B(i_data_pc8[17]), .S(i_con_pc8), .Q(
        o_data_alu[17]) );
  MUX22 U21 ( .A(i_data_alures[21]), .B(i_data_pc8[21]), .S(i_con_pc8), .Q(
        o_data_alu[21]) );
  MUX22 U22 ( .A(i_data_alures[25]), .B(i_data_pc8[25]), .S(i_con_pc8), .Q(
        o_data_alu[25]) );
  INV3 U23 ( .A(n34), .Q(o_data_alu[9]) );
  AOI221 U24 ( .A(i_data_alures[9]), .B(n1), .C(i_data_pc8[9]), .D(i_con_pc8), 
        .Q(n34) );
  INV3 U25 ( .A(n37), .Q(o_data_alu[6]) );
  AOI221 U26 ( .A(i_data_alures[6]), .B(n1), .C(i_data_pc8[6]), .D(i_con_pc8), 
        .Q(n37) );
  INV3 U27 ( .A(n62), .Q(o_data_alu[12]) );
  MUX22 U28 ( .A(i_data_alures[16]), .B(i_data_pc8[16]), .S(i_con_pc8), .Q(
        o_data_alu[16]) );
  MUX22 U29 ( .A(i_data_alures[26]), .B(i_data_pc8[26]), .S(i_con_pc8), .Q(
        o_data_alu[26]) );
  MUX22 U30 ( .A(i_data_alures[28]), .B(i_data_pc8[28]), .S(i_con_pc8), .Q(
        o_data_alu[28]) );
  MUX22 U31 ( .A(i_data_alures[15]), .B(i_data_pc8[15]), .S(i_con_pc8), .Q(
        o_data_alu[15]) );
  MUX22 U32 ( .A(i_data_alures[18]), .B(i_data_pc8[18]), .S(i_con_pc8), .Q(
        o_data_alu[18]) );
  MUX22 U33 ( .A(i_data_alures[20]), .B(i_data_pc8[20]), .S(i_con_pc8), .Q(
        o_data_alu[20]) );
  MUX22 U34 ( .A(i_data_alures[19]), .B(i_data_pc8[19]), .S(i_con_pc8), .Q(
        o_data_alu[19]) );
  MUX22 U35 ( .A(i_data_alures[22]), .B(i_data_pc8[22]), .S(i_con_pc8), .Q(
        o_data_alu[22]) );
  MUX22 U36 ( .A(i_data_alures[24]), .B(i_data_pc8[24]), .S(i_con_pc8), .Q(
        o_data_alu[24]) );
  MUX22 U37 ( .A(i_data_alures[29]), .B(i_data_pc8[29]), .S(i_con_pc8), .Q(
        o_data_alu[29]) );
  MUX22 U38 ( .A(i_data_alures[31]), .B(i_data_pc8[31]), .S(i_con_pc8), .Q(
        o_data_alu[31]) );
  INV3 U39 ( .A(i_con_pc8), .Q(n1) );
  INV3 U40 ( .A(n65), .Q(o_data_alu[0]) );
  AOI221 U41 ( .A(i_data_alures[0]), .B(n1), .C(i_data_pc8[0]), .D(i_con_pc8), 
        .Q(n65) );
  INV3 U42 ( .A(n43), .Q(o_data_alu[2]) );
  INV3 U43 ( .A(n39), .Q(o_data_alu[4]) );
  AOI221 U44 ( .A(i_data_alures[4]), .B(n1), .C(i_data_pc8[4]), .D(i_con_pc8), 
        .Q(n39) );
  INV3 U45 ( .A(n35), .Q(o_data_alu[8]) );
  AOI221 U46 ( .A(i_data_alures[8]), .B(n1), .C(i_data_pc8[8]), .D(i_con_pc8), 
        .Q(n35) );
  INV3 U47 ( .A(n54), .Q(o_data_alu[1]) );
  AOI221 U48 ( .A(i_data_alures[1]), .B(n1), .C(i_data_pc8[1]), .D(i_con_pc8), 
        .Q(n54) );
endmodule


module mem_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV3 U2 ( .A(n5), .Q(n7) );
  NOR21 U3 ( .A(n27), .B(n33), .Q(n31) );
  INV3 U4 ( .A(n48), .Q(n47) );
  NAND22 U5 ( .A(n38), .B(n22), .Q(n48) );
  INV3 U6 ( .A(n35), .Q(n34) );
  NAND22 U7 ( .A(n36), .B(n22), .Q(n35) );
  INV3 U8 ( .A(n58), .Q(n22) );
  NAND22 U9 ( .A(n59), .B(n60), .Q(n58) );
  NOR31 U10 ( .A(n61), .B(n62), .C(n63), .Q(n60) );
  NOR21 U11 ( .A(n65), .B(n66), .Q(n59) );
  INV3 U12 ( .A(n44), .Q(n43) );
  NAND22 U13 ( .A(n45), .B(A[21]), .Q(n44) );
  INV3 U14 ( .A(n64), .Q(n61) );
  INV3 U15 ( .A(n65), .Q(n3) );
  NOR21 U16 ( .A(n79), .B(n2), .Q(n78) );
  NOR21 U17 ( .A(n8), .B(n10), .Q(n5) );
  INV3 U18 ( .A(n20), .Q(n17) );
  NAND22 U19 ( .A(n21), .B(n22), .Q(n20) );
  NOR21 U20 ( .A(n23), .B(n24), .Q(n21) );
  NAND22 U21 ( .A(n78), .B(A[10]), .Q(n77) );
  NAND22 U22 ( .A(n5), .B(A[6]), .Q(n4) );
  INV3 U23 ( .A(n74), .Q(n73) );
  NAND22 U24 ( .A(n64), .B(n3), .Q(n74) );
  INV3 U25 ( .A(n70), .Q(n69) );
  NAND22 U26 ( .A(n71), .B(A[13]), .Q(n70) );
  INV3 U27 ( .A(n55), .Q(n54) );
  NAND22 U28 ( .A(n56), .B(A[17]), .Q(n55) );
  NOR31 U29 ( .A(n76), .B(n75), .C(n2), .Q(n64) );
  NAND22 U30 ( .A(A[11]), .B(A[8]), .Q(n75) );
  INV3 U31 ( .A(A[10]), .Q(n76) );
  NAND22 U32 ( .A(A[7]), .B(A[3]), .Q(n83) );
  XOR21 U33 ( .A(n42), .B(A[23]), .Q(SUM[23]) );
  NOR21 U34 ( .A(n41), .B(n44), .Q(n42) );
  NAND31 U35 ( .A(n80), .B(A[2]), .C(n81), .Q(n65) );
  NOR21 U36 ( .A(n6), .B(n8), .Q(n80) );
  NOR21 U37 ( .A(n82), .B(n83), .Q(n81) );
  INV3 U38 ( .A(A[4]), .Q(n82) );
  INV3 U39 ( .A(n46), .Q(n45) );
  NAND22 U40 ( .A(A[20]), .B(n47), .Q(n46) );
  INV3 U41 ( .A(n33), .Q(n32) );
  NAND22 U42 ( .A(A[24]), .B(n34), .Q(n33) );
  INV3 U43 ( .A(A[2]), .Q(SUM[2]) );
  XOR21 U44 ( .A(n29), .B(n30), .Q(SUM[27]) );
  INV3 U45 ( .A(A[27]), .Q(n29) );
  NAND22 U46 ( .A(n31), .B(A[26]), .Q(n30) );
  NOR31 U47 ( .A(n51), .B(n49), .C(n50), .Q(n38) );
  NAND22 U48 ( .A(A[19]), .B(A[16]), .Q(n49) );
  XOR21 U49 ( .A(n56), .B(A[17]), .Q(SUM[17]) );
  XOR21 U50 ( .A(n45), .B(A[21]), .Q(SUM[21]) );
  XOR21 U51 ( .A(n32), .B(A[25]), .Q(SUM[25]) );
  XOR21 U52 ( .A(A[30]), .B(n15), .Q(SUM[30]) );
  NAND22 U53 ( .A(n37), .B(n38), .Q(n23) );
  NOR31 U54 ( .A(n41), .B(n39), .C(n40), .Q(n37) );
  NAND22 U55 ( .A(A[23]), .B(A[20]), .Q(n39) );
  XNR21 U56 ( .A(n78), .B(n76), .Q(SUM[10]) );
  XNR21 U57 ( .A(n71), .B(n62), .Q(SUM[13]) );
  XNR21 U58 ( .A(n69), .B(n63), .Q(SUM[14]) );
  XOR21 U59 ( .A(n1), .B(A[9]), .Q(SUM[9]) );
  XNR21 U60 ( .A(A[7]), .B(n4), .Q(SUM[7]) );
  XNR21 U61 ( .A(A[11]), .B(n77), .Q(SUM[11]) );
  INV3 U62 ( .A(A[22]), .Q(n41) );
  INV3 U63 ( .A(A[25]), .Q(n27) );
  INV3 U64 ( .A(A[9]), .Q(n2) );
  INV3 U65 ( .A(A[18]), .Q(n51) );
  INV3 U66 ( .A(A[26]), .Q(n28) );
  INV3 U67 ( .A(A[13]), .Q(n62) );
  INV3 U68 ( .A(A[17]), .Q(n50) );
  INV3 U69 ( .A(A[21]), .Q(n40) );
  INV3 U70 ( .A(A[14]), .Q(n63) );
  INV3 U71 ( .A(A[5]), .Q(n8) );
  NOR21 U72 ( .A(n16), .B(n18), .Q(n15) );
  NAND22 U73 ( .A(A[28]), .B(n17), .Q(n16) );
  INV3 U74 ( .A(A[6]), .Q(n6) );
  NAND22 U75 ( .A(A[15]), .B(A[12]), .Q(n66) );
  NOR31 U76 ( .A(n28), .B(n26), .C(n27), .Q(n25) );
  NAND22 U77 ( .A(A[27]), .B(A[24]), .Q(n26) );
  INV3 U78 ( .A(n12), .Q(n11) );
  NAND22 U79 ( .A(A[3]), .B(A[2]), .Q(n12) );
  INV3 U80 ( .A(n57), .Q(n56) );
  NAND22 U81 ( .A(A[16]), .B(n22), .Q(n57) );
  INV3 U82 ( .A(n72), .Q(n71) );
  NAND22 U83 ( .A(A[12]), .B(n73), .Q(n72) );
  INV3 U84 ( .A(n79), .Q(n1) );
  NAND22 U85 ( .A(A[8]), .B(n3), .Q(n79) );
  INV3 U86 ( .A(n10), .Q(n9) );
  NAND22 U87 ( .A(A[4]), .B(n11), .Q(n10) );
  XNR21 U88 ( .A(n7), .B(A[6]), .Q(SUM[6]) );
  XOR21 U89 ( .A(n73), .B(A[12]), .Q(SUM[12]) );
  XOR21 U90 ( .A(n22), .B(A[16]), .Q(SUM[16]) );
  XOR21 U91 ( .A(n31), .B(A[26]), .Q(SUM[26]) );
  XOR21 U92 ( .A(n17), .B(A[28]), .Q(SUM[28]) );
  XOR21 U93 ( .A(n67), .B(n68), .Q(SUM[15]) );
  INV3 U94 ( .A(A[15]), .Q(n67) );
  NAND22 U95 ( .A(n69), .B(A[14]), .Q(n68) );
  XOR21 U96 ( .A(n54), .B(A[18]), .Q(SUM[18]) );
  XOR21 U97 ( .A(n47), .B(A[20]), .Q(SUM[20]) );
  XOR21 U98 ( .A(n52), .B(n53), .Q(SUM[19]) );
  INV3 U99 ( .A(A[19]), .Q(n52) );
  NAND22 U100 ( .A(n54), .B(A[18]), .Q(n53) );
  XOR21 U101 ( .A(n43), .B(A[22]), .Q(SUM[22]) );
  XOR21 U102 ( .A(n34), .B(A[24]), .Q(SUM[24]) );
  XOR21 U103 ( .A(n18), .B(n19), .Q(SUM[29]) );
  INV3 U104 ( .A(A[29]), .Q(n18) );
  NAND22 U105 ( .A(A[28]), .B(n17), .Q(n19) );
  XOR21 U106 ( .A(n13), .B(n14), .Q(SUM[31]) );
  INV3 U107 ( .A(A[31]), .Q(n13) );
  NAND22 U108 ( .A(A[30]), .B(n15), .Q(n14) );
  XNR21 U109 ( .A(n9), .B(n8), .Q(SUM[5]) );
  XNR21 U110 ( .A(A[3]), .B(SUM[2]), .Q(SUM[3]) );
  XOR21 U111 ( .A(n11), .B(A[4]), .Q(SUM[4]) );
  XOR21 U112 ( .A(n3), .B(A[8]), .Q(SUM[8]) );
  CLKIN3 U113 ( .A(n25), .Q(n24) );
  CLKIN3 U114 ( .A(n23), .Q(n36) );
endmodule


module mem ( i_clk, i_nrst, i_data_pc4, i_data_alures, i_data_memout, 
        i_addr_regdst, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_FWmemread, i_addr_Mrt, o_data_alures, o_data_memout, 
        o_addr_regdst, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread, 
        o_addr_Wrt );
  input [31:0] i_data_pc4;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [4:0] i_addr_regdst;
  input [4:0] i_addr_Mrt;
  output [31:0] o_data_alures;
  output [31:0] o_data_memout;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Wrt;
  input i_clk, i_nrst, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite,
         i_con_FWmemread;
  output o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread;
  wire   n_Logic1_, n_Logic0_;
  wire   [31:0] pc8;
  wire   [31:0] resmux_o_data_alu;

  DFC3 pipe_rt_reg_4_ ( .D(i_addr_Mrt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(i_addr_Mrt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(i_addr_Mrt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[2]) );
  DFC3 pipe_rt_reg_1_ ( .D(i_addr_Mrt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[1]) );
  DFC3 pipe_rt_reg_0_ ( .D(i_addr_Mrt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[0]) );
  DFC3 pipe_data_alures_reg_31_ ( .D(resmux_o_data_alu[31]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[31]) );
  DFC3 pipe_data_alures_reg_30_ ( .D(resmux_o_data_alu[30]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[30]) );
  DFC3 pipe_data_alures_reg_29_ ( .D(resmux_o_data_alu[29]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[29]) );
  DFC3 pipe_data_alures_reg_28_ ( .D(resmux_o_data_alu[28]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[28]) );
  DFC3 pipe_data_alures_reg_27_ ( .D(resmux_o_data_alu[27]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[27]) );
  DFC3 pipe_data_alures_reg_26_ ( .D(resmux_o_data_alu[26]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[26]) );
  DFC3 pipe_data_alures_reg_25_ ( .D(resmux_o_data_alu[25]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[25]) );
  DFC3 pipe_data_alures_reg_24_ ( .D(resmux_o_data_alu[24]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[24]) );
  DFC3 pipe_data_alures_reg_23_ ( .D(resmux_o_data_alu[23]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[23]) );
  DFC3 pipe_data_alures_reg_22_ ( .D(resmux_o_data_alu[22]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[22]) );
  DFC3 pipe_data_alures_reg_21_ ( .D(resmux_o_data_alu[21]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[21]) );
  DFC3 pipe_data_alures_reg_20_ ( .D(resmux_o_data_alu[20]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[20]) );
  DFC3 pipe_data_alures_reg_19_ ( .D(resmux_o_data_alu[19]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[19]) );
  DFC3 pipe_data_alures_reg_18_ ( .D(resmux_o_data_alu[18]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[18]) );
  DFC3 pipe_data_alures_reg_17_ ( .D(resmux_o_data_alu[17]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[17]) );
  DFC3 pipe_data_alures_reg_16_ ( .D(resmux_o_data_alu[16]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[16]) );
  DFC3 pipe_data_alures_reg_15_ ( .D(resmux_o_data_alu[15]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[15]) );
  DFC3 pipe_data_alures_reg_14_ ( .D(resmux_o_data_alu[14]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[14]) );
  DFC3 pipe_data_alures_reg_13_ ( .D(resmux_o_data_alu[13]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[13]) );
  DFC3 pipe_data_alures_reg_12_ ( .D(resmux_o_data_alu[12]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[12]) );
  DFC3 pipe_data_alures_reg_11_ ( .D(resmux_o_data_alu[11]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[11]) );
  DFC3 pipe_data_alures_reg_10_ ( .D(resmux_o_data_alu[10]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[10]) );
  DFC3 pipe_data_alures_reg_9_ ( .D(resmux_o_data_alu[9]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[9]) );
  DFC3 pipe_data_alures_reg_8_ ( .D(resmux_o_data_alu[8]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[8]) );
  DFC3 pipe_data_alures_reg_7_ ( .D(resmux_o_data_alu[7]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[7]) );
  DFC3 pipe_data_alures_reg_6_ ( .D(resmux_o_data_alu[6]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[6]) );
  DFC3 pipe_data_alures_reg_5_ ( .D(resmux_o_data_alu[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[5]) );
  DFC3 pipe_data_alures_reg_4_ ( .D(resmux_o_data_alu[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[4]) );
  DFC3 pipe_data_alures_reg_3_ ( .D(resmux_o_data_alu[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[3]) );
  DFC3 pipe_data_alures_reg_2_ ( .D(resmux_o_data_alu[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[2]) );
  DFC3 pipe_data_alures_reg_1_ ( .D(resmux_o_data_alu[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[1]) );
  DFC3 pipe_data_alures_reg_0_ ( .D(resmux_o_data_alu[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[0]) );
  DFC3 pipe_data_memout_reg_31_ ( .D(i_data_memout[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[31]) );
  DFC3 pipe_data_memout_reg_30_ ( .D(i_data_memout[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[30]) );
  DFC3 pipe_data_memout_reg_29_ ( .D(i_data_memout[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[29]) );
  DFC3 pipe_data_memout_reg_28_ ( .D(i_data_memout[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[28]) );
  DFC3 pipe_data_memout_reg_27_ ( .D(i_data_memout[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[27]) );
  DFC3 pipe_data_memout_reg_26_ ( .D(i_data_memout[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[26]) );
  DFC3 pipe_data_memout_reg_25_ ( .D(i_data_memout[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[25]) );
  DFC3 pipe_data_memout_reg_24_ ( .D(i_data_memout[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[24]) );
  DFC3 pipe_data_memout_reg_23_ ( .D(i_data_memout[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[23]) );
  DFC3 pipe_data_memout_reg_22_ ( .D(i_data_memout[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[22]) );
  DFC3 pipe_data_memout_reg_21_ ( .D(i_data_memout[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[21]) );
  DFC3 pipe_data_memout_reg_20_ ( .D(i_data_memout[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[20]) );
  DFC3 pipe_data_memout_reg_19_ ( .D(i_data_memout[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[19]) );
  DFC3 pipe_data_memout_reg_18_ ( .D(i_data_memout[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[18]) );
  DFC3 pipe_data_memout_reg_17_ ( .D(i_data_memout[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[17]) );
  DFC3 pipe_data_memout_reg_16_ ( .D(i_data_memout[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[16]) );
  DFC3 pipe_data_memout_reg_15_ ( .D(i_data_memout[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[15]) );
  DFC3 pipe_data_memout_reg_14_ ( .D(i_data_memout[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[14]) );
  DFC3 pipe_data_memout_reg_13_ ( .D(i_data_memout[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[13]) );
  DFC3 pipe_data_memout_reg_12_ ( .D(i_data_memout[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[12]) );
  DFC3 pipe_data_memout_reg_11_ ( .D(i_data_memout[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[11]) );
  DFC3 pipe_data_memout_reg_10_ ( .D(i_data_memout[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[10]) );
  DFC3 pipe_data_memout_reg_9_ ( .D(i_data_memout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[9]) );
  DFC3 pipe_data_memout_reg_8_ ( .D(i_data_memout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[8]) );
  DFC3 pipe_data_memout_reg_7_ ( .D(i_data_memout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[7]) );
  DFC3 pipe_data_memout_reg_6_ ( .D(i_data_memout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[6]) );
  DFC3 pipe_data_memout_reg_5_ ( .D(i_data_memout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[5]) );
  DFC3 pipe_data_memout_reg_4_ ( .D(i_data_memout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[4]) );
  DFC3 pipe_data_memout_reg_3_ ( .D(i_data_memout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[3]) );
  DFC3 pipe_data_memout_reg_2_ ( .D(i_data_memout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[2]) );
  DFC3 pipe_data_memout_reg_1_ ( .D(i_data_memout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[1]) );
  DFC3 pipe_data_memout_reg_0_ ( .D(i_data_memout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[0]) );
  DFC3 pipe_addr_regdst_reg_4_ ( .D(i_addr_regdst[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[4]) );
  DFC3 pipe_addr_regdst_reg_3_ ( .D(i_addr_regdst[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[3]) );
  DFC3 pipe_addr_regdst_reg_2_ ( .D(i_addr_regdst[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[2]) );
  DFC3 pipe_addr_regdst_reg_1_ ( .D(i_addr_regdst[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[1]) );
  DFC3 pipe_addr_regdst_reg_0_ ( .D(i_addr_regdst[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[0]) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_con_FWmemread_reg ( .D(i_con_FWmemread), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_FWmemread) );
  M_resmux u_resmux ( .i_data_alures(i_data_alures), .i_data_pc8(pc8), 
        .i_con_pc8(i_con_Malupc8), .o_data_alu(resmux_o_data_alu) );
  mem_DW01_add_1 add_27 ( .A(i_data_pc4), .B({n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic1_, n_Logic0_, n_Logic0_}), .CI(n_Logic0_), .SUM(pc8) );
  LOGIC0 U3 ( .Q(n_Logic0_) );
  LOGIC1 U4 ( .Q(n_Logic1_) );
endmodule


module W_datamux ( i_data_alu, i_data_load, i_con_memtoreg, o_data_toreg );
  input [31:0] i_data_alu;
  input [31:0] i_data_load;
  output [31:0] o_data_toreg;
  input i_con_memtoreg;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n1;

  AOI220 U1 ( .A(i_data_alu[19]), .B(n1), .C(i_data_load[19]), .D(
        i_con_memtoreg), .Q(n55) );
  AOI220 U2 ( .A(i_data_alu[21]), .B(n1), .C(i_data_load[21]), .D(
        i_con_memtoreg), .Q(n52) );
  AOI220 U3 ( .A(i_data_alu[5]), .B(n1), .C(i_data_load[5]), .D(i_con_memtoreg), .Q(n38) );
  AOI220 U4 ( .A(i_data_alu[7]), .B(n1), .C(i_data_load[7]), .D(i_con_memtoreg), .Q(n36) );
  AOI220 U5 ( .A(i_data_alu[12]), .B(n1), .C(i_data_load[12]), .D(
        i_con_memtoreg), .Q(n62) );
  AOI220 U6 ( .A(i_data_alu[1]), .B(n1), .C(i_data_load[1]), .D(i_con_memtoreg), .Q(n54) );
  AOI220 U7 ( .A(i_data_alu[2]), .B(n1), .C(i_data_load[2]), .D(i_con_memtoreg), .Q(n43) );
  AOI220 U8 ( .A(i_data_alu[3]), .B(n1), .C(i_data_load[3]), .D(i_con_memtoreg), .Q(n40) );
  AOI220 U9 ( .A(i_data_alu[9]), .B(n1), .C(i_data_load[9]), .D(i_con_memtoreg), .Q(n34) );
  AOI220 U10 ( .A(i_data_alu[10]), .B(n1), .C(i_data_load[10]), .D(
        i_con_memtoreg), .Q(n64) );
  AOI220 U11 ( .A(i_data_alu[11]), .B(n1), .C(i_data_load[11]), .D(
        i_con_memtoreg), .Q(n63) );
  AOI220 U12 ( .A(i_data_alu[13]), .B(n1), .C(i_data_load[13]), .D(
        i_con_memtoreg), .Q(n61) );
  INV3 U13 ( .A(n57), .Q(o_data_toreg[17]) );
  AOI221 U14 ( .A(i_data_alu[17]), .B(n1), .C(i_data_load[17]), .D(
        i_con_memtoreg), .Q(n57) );
  INV3 U15 ( .A(n51), .Q(o_data_toreg[22]) );
  AOI221 U16 ( .A(i_data_alu[22]), .B(n1), .C(i_data_load[22]), .D(
        i_con_memtoreg), .Q(n51) );
  INV3 U17 ( .A(n45), .Q(o_data_toreg[28]) );
  AOI221 U18 ( .A(i_data_alu[28]), .B(n1), .C(i_data_load[28]), .D(
        i_con_memtoreg), .Q(n45) );
  INV3 U19 ( .A(n42), .Q(o_data_toreg[30]) );
  AOI221 U20 ( .A(i_data_alu[30]), .B(n1), .C(i_data_load[30]), .D(
        i_con_memtoreg), .Q(n42) );
  INV3 U21 ( .A(n65), .Q(o_data_toreg[0]) );
  AOI221 U22 ( .A(i_data_alu[0]), .B(n1), .C(i_data_load[0]), .D(
        i_con_memtoreg), .Q(n65) );
  INV3 U23 ( .A(n43), .Q(o_data_toreg[2]) );
  INV3 U24 ( .A(n40), .Q(o_data_toreg[3]) );
  INV3 U25 ( .A(n39), .Q(o_data_toreg[4]) );
  AOI221 U26 ( .A(i_data_alu[4]), .B(n1), .C(i_data_load[4]), .D(
        i_con_memtoreg), .Q(n39) );
  INV3 U27 ( .A(n36), .Q(o_data_toreg[7]) );
  INV3 U28 ( .A(n64), .Q(o_data_toreg[10]) );
  INV3 U29 ( .A(n62), .Q(o_data_toreg[12]) );
  INV3 U30 ( .A(n61), .Q(o_data_toreg[13]) );
  INV3 U31 ( .A(n34), .Q(o_data_toreg[9]) );
  INV3 U32 ( .A(n60), .Q(o_data_toreg[14]) );
  AOI221 U33 ( .A(i_data_alu[14]), .B(n1), .C(i_data_load[14]), .D(
        i_con_memtoreg), .Q(n60) );
  INV3 U34 ( .A(n59), .Q(o_data_toreg[15]) );
  AOI221 U35 ( .A(i_data_alu[15]), .B(n1), .C(i_data_load[15]), .D(
        i_con_memtoreg), .Q(n59) );
  INV3 U36 ( .A(n56), .Q(o_data_toreg[18]) );
  AOI221 U37 ( .A(i_data_alu[18]), .B(n1), .C(i_data_load[18]), .D(
        i_con_memtoreg), .Q(n56) );
  INV3 U38 ( .A(n53), .Q(o_data_toreg[20]) );
  AOI221 U39 ( .A(i_data_alu[20]), .B(n1), .C(i_data_load[20]), .D(
        i_con_memtoreg), .Q(n53) );
  INV3 U40 ( .A(n52), .Q(o_data_toreg[21]) );
  INV3 U41 ( .A(n49), .Q(o_data_toreg[24]) );
  AOI221 U42 ( .A(i_data_alu[24]), .B(n1), .C(i_data_load[24]), .D(
        i_con_memtoreg), .Q(n49) );
  INV3 U43 ( .A(n41), .Q(o_data_toreg[31]) );
  AOI221 U44 ( .A(i_data_alu[31]), .B(n1), .C(i_data_load[31]), .D(
        i_con_memtoreg), .Q(n41) );
  INV3 U45 ( .A(n37), .Q(o_data_toreg[6]) );
  AOI221 U46 ( .A(i_data_alu[6]), .B(n1), .C(i_data_load[6]), .D(
        i_con_memtoreg), .Q(n37) );
  INV3 U47 ( .A(n38), .Q(o_data_toreg[5]) );
  INV3 U48 ( .A(n35), .Q(o_data_toreg[8]) );
  AOI221 U49 ( .A(i_data_alu[8]), .B(n1), .C(i_data_load[8]), .D(
        i_con_memtoreg), .Q(n35) );
  INV3 U50 ( .A(n63), .Q(o_data_toreg[11]) );
  INV3 U51 ( .A(n50), .Q(o_data_toreg[23]) );
  AOI221 U52 ( .A(i_data_alu[23]), .B(n1), .C(i_data_load[23]), .D(
        i_con_memtoreg), .Q(n50) );
  INV3 U53 ( .A(n48), .Q(o_data_toreg[25]) );
  AOI221 U54 ( .A(i_data_alu[25]), .B(n1), .C(i_data_load[25]), .D(
        i_con_memtoreg), .Q(n48) );
  INV3 U55 ( .A(n47), .Q(o_data_toreg[26]) );
  AOI221 U56 ( .A(i_data_alu[26]), .B(n1), .C(i_data_load[26]), .D(
        i_con_memtoreg), .Q(n47) );
  INV3 U57 ( .A(n46), .Q(o_data_toreg[27]) );
  AOI221 U58 ( .A(i_data_alu[27]), .B(n1), .C(i_data_load[27]), .D(
        i_con_memtoreg), .Q(n46) );
  INV3 U59 ( .A(n44), .Q(o_data_toreg[29]) );
  AOI221 U60 ( .A(i_data_alu[29]), .B(n1), .C(i_data_load[29]), .D(
        i_con_memtoreg), .Q(n44) );
  INV3 U61 ( .A(n54), .Q(o_data_toreg[1]) );
  INV3 U62 ( .A(n55), .Q(o_data_toreg[19]) );
  INV3 U63 ( .A(n58), .Q(o_data_toreg[16]) );
  AOI221 U64 ( .A(i_data_alu[16]), .B(n1), .C(i_data_load[16]), .D(
        i_con_memtoreg), .Q(n58) );
  INV3 U65 ( .A(i_con_memtoreg), .Q(n1) );
endmodule


module writeback ( i_data_alures, i_data_memout, i_con_Wmemtoreg, 
        o_data_regwrite );
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  output [31:0] o_data_regwrite;
  input i_con_Wmemtoreg;


  W_datamux u_datamux ( .i_data_alu(i_data_alures), .i_data_load(i_data_memout), .i_con_memtoreg(i_con_Wmemtoreg), .o_data_toreg(o_data_regwrite) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Mmemread, ex_con_Mmemwrite, ex_con_Malupc8, ex_con_Wmemtoreg,
         mem_con_Malupc8, mem_con_Wmemtoreg, wb_con_Wmemtoreg, n1,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2;
  wire   [31:0] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [31:0] id_addr_pc4;
  wire   [31:0] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] wb_data_memout;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] mem_data_alures;
  wire   [31:0] mem_data_pc4;

  fetch u_fetch ( .i_clk(clk), .i_nrst(rst_n), .i_addr_b(if_addr_b), 
        .i_addr_j({if_addr_j, n1, n1}), .i_addr_jr(id_data_jr), .i_con_b(
        if_con_b), .i_con_j(if_con_j), .i_data_instr(read_instruction), 
        .i_con_ifstall(if_con_ifstall), .o_addr_pc(instruction_address), 
        .o_addr_pc4(id_addr_pc4), .o_data_instr(id_data_instr) );
  decode u_decode ( .i_clk(clk), .i_nrst(rst_n), .i_addr_pc4(id_addr_pc4), 
        .i_data_instr(id_data_instr), .i_con_Wregwrite(id_con_Wregwrite), 
        .i_data_Wregwrite(id_data_Wregwrite), .i_addr_Wregwrite(
        id_addr_Wregwrite), .i_addr_Erd(for_o_addr_Erd), .i_addr_Mrd(
        mem_addr_regdst), .i_con_Eregwrite(ex_con_Wregwrite), 
        .i_con_Mregwrite(mem_con_Wregwrite), .i_addr_rtM(for_addr_rtM), 
        .i_addr_rtW(for_addr_rtW), .i_con_memreadM(mem_read), .i_con_memreadW(
        for_FWmemread), .i_data_Wmemout(wb_data_memout), .o_data_rs(id_data_rs), .o_data_rt(ex_data_rt), .o_addr_rd(ex_addr_rd), .o_addr_rt(ex_addr_rt), 
        .o_data_jr(id_data_jr), .o_con_jump(if_con_j), .o_addr_pc4(ex_data_pc4), .o_addr_branch(if_addr_b), .o_addr_jump({if_addr_j, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .o_con_Ealuop(ex_con_Ealuop), 
        .o_con_Ealusrc(ex_con_Ealusrc), .o_con_Eregdst(ex_con_Eregdst), 
        .o_con_Mmemread(ex_con_Mmemread), .o_con_Mmemwrite(ex_con_Mmemwrite), 
        .o_con_Malupc8(ex_con_Malupc8), .o_con_Wmemtoreg(ex_con_Wmemtoreg), 
        .o_con_Wregwrite(ex_con_Wregwrite), .o_con_ifstall(if_con_ifstall), 
        .o_con_Ebop(ex_con_bop), .o_data_signext(ex_data_immext), 
        .o_con_Efamux(for_o_con_Efamux), .o_con_Efbmux(for_o_con_Efbmux), 
        .o_data_Fmemout(for_memout) );
  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext(
        ex_data_immext), .i_addr_rt(ex_addr_rt), .i_addr_rd(ex_addr_rd), 
        .i_data_FEalures(data_address), .i_data_FMalures(mem_data_alures), 
        .i_data_FMmemout(wb_data_memout), .i_data_FWmemout(for_memout), 
        .i_con_Efamux(for_o_con_Efamux), .i_con_Efbmux(for_o_con_Efbmux), 
        .i_con_Ealuop(ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), 
        .i_con_Mmemwrite(ex_con_Mmemwrite), .i_con_Malupc8(ex_con_Malupc8), 
        .i_con_Wmemtoreg(ex_con_Wmemtoreg), .i_con_Wregwrite(ex_con_Wregwrite), 
        .i_con_bop(ex_con_bop), .o_data_pc4(mem_data_pc4), .o_data_alures(
        data_address), .o_data_rt(write_data), .o_addr_regdst(mem_addr_regdst), 
        .o_con_Mmemread(mem_read), .o_con_Mmemwrite(mem_write), 
        .o_con_Malupc8(mem_con_Malupc8), .o_con_Wmemtoreg(mem_con_Wmemtoreg), 
        .o_con_Wregwrite(mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), 
        .o_addr_Mrt(for_addr_rtM), .o_con_ifbranch(if_con_b) );
  mem u_mem ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(mem_data_pc4), 
        .i_data_alures(data_address), .i_data_memout(read_data), 
        .i_addr_regdst(mem_addr_regdst), .i_con_Malupc8(mem_con_Malupc8), 
        .i_con_Wmemtoreg(mem_con_Wmemtoreg), .i_con_Wregwrite(
        mem_con_Wregwrite), .i_con_FWmemread(ex_con_Mmemread), .i_addr_Mrt(
        for_addr_rtM), .o_data_alures(mem_data_alures), .o_data_memout(
        wb_data_memout), .o_addr_regdst(id_addr_Wregwrite), .o_con_Wmemtoreg(
        wb_con_Wmemtoreg), .o_con_Wregwrite(id_con_Wregwrite), 
        .o_con_FWmemread(for_FWmemread), .o_addr_Wrt(for_addr_rtW) );
  writeback u_writeback ( .i_data_alures(mem_data_alures), .i_data_memout(
        wb_data_memout), .i_con_Wmemtoreg(wb_con_Wmemtoreg), .o_data_regwrite(
        id_data_Wregwrite) );
  LOGIC0 U1 ( .Q(n1) );
endmodule

