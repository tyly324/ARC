
module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Efamux, i_con_Efbmux, 
        i_con_Ealuop, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread, 
        i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_bop, o_data_alures, o_data_rt, o_addr_regdst, o_con_Mmemread, 
        o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, o_con_Wregwrite, 
        o_addr_Erd, o_addr_Mrt, o_con_ifbranch, o_data_pc4_31_, o_data_pc4_30_, 
        o_data_pc4_29_, o_data_pc4_28_, o_data_pc4_27_, o_data_pc4_26_, 
        o_data_pc4_25_, o_data_pc4_24_, o_data_pc4_23_, o_data_pc4_22_, 
        o_data_pc4_21_, o_data_pc4_20_, o_data_pc4_19_, o_data_pc4_18_, 
        o_data_pc4_17_, o_data_pc4_16__BAR, o_data_pc4_15_, o_data_pc4_14_, 
        o_data_pc4_13_, o_data_pc4_12_, o_data_pc4_11_, o_data_pc4_10_, 
        o_data_pc4_9_, o_data_pc4_8_, o_data_pc4_7_, o_data_pc4_6_, 
        o_data_pc4_5_, o_data_pc4_4_, o_data_pc4_3_, o_data_pc4_2_, 
        o_data_pc4_1_, o_data_pc4_0_ );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [5:0] i_con_Ealuop;
  input [2:0] i_con_bop;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch, o_data_pc4_31_, o_data_pc4_30_,
         o_data_pc4_29_, o_data_pc4_28_, o_data_pc4_27_, o_data_pc4_26_,
         o_data_pc4_25_, o_data_pc4_24_, o_data_pc4_23_, o_data_pc4_22_,
         o_data_pc4_21_, o_data_pc4_20_, o_data_pc4_19_, o_data_pc4_18_,
         o_data_pc4_17_, o_data_pc4_16__BAR, o_data_pc4_15_, o_data_pc4_14_,
         o_data_pc4_13_, o_data_pc4_12_, o_data_pc4_11_, o_data_pc4_10_,
         o_data_pc4_9_, o_data_pc4_8_, o_data_pc4_7_, o_data_pc4_6_,
         o_data_pc4_5_, o_data_pc4_4_, o_data_pc4_3_, o_data_pc4_2_,
         o_data_pc4_1_, o_data_pc4_0_;
  wire   u_alu_N306, u_alu_N256, u_alu_N255, u_alu_N253, u_alu_N250,
         u_alu_N249, u_alu_N248, u_alu_N247, u_alu_N246, u_alu_N245,
         u_alu_N244, u_alu_N243, u_alu_N242, u_alu_N241, u_alu_N240,
         u_alu_N238, u_alu_N237, u_alu_N236, u_alu_N235, u_alu_N234,
         u_alu_N233, u_alu_N232, u_alu_N231, u_alu_N230, u_alu_N229,
         u_alu_N228, u_alu_N227, u_alu_N226, u_alu_N225, u_alu_N224,
         u_alu_N223, u_alu_N222, u_alu_N221, u_alu_N218, u_alu_N217,
         u_alu_N216, u_alu_N215, u_alu_N214, u_alu_N213, u_alu_N212,
         u_alu_N211, u_alu_N210, u_alu_N209, u_alu_N207, u_alu_N206,
         u_alu_N205, u_alu_N203, u_alu_N202, u_alu_N200, u_alu_N199,
         u_alu_N198, u_alu_N197, u_alu_N196, u_alu_N195, u_alu_N194,
         u_alu_N193, u_alu_N173, u_alu_N172, u_alu_N171, u_alu_N170,
         u_alu_N169, u_alu_N168, u_alu_N167, u_alu_N166, u_alu_N165,
         u_alu_half_sub_0_, u_alu_half_sub_1_, u_alu_half_sub_2_,
         u_alu_half_sub_3_, u_alu_half_sub_4_, u_alu_half_sub_5_,
         u_alu_half_sub_6_, u_alu_half_sub_7_, u_alu_half_sub_8_,
         u_alu_half_sub_9_, u_alu_half_sub_10_, u_alu_half_sub_11_,
         u_alu_half_sub_12_, u_alu_half_sub_13_, u_alu_half_sub_15_,
         u_alu_half_sub_16_, u_alu_sum_1_0_, u_alu_sum_1_1_, u_alu_sum_1_2_,
         u_alu_sum_1_3_, u_alu_sum_1_4_, u_alu_sum_1_5_, u_alu_sum_1_6_,
         u_alu_sum_1_7_, u_alu_sum_1_8_, u_alu_ashr_4_SH_3_,
         u_alu_ashr_4_SH_1_, u_alu_add_x_1_n51, u_alu_add_x_1_n50,
         u_alu_add_x_1_n49, u_alu_add_x_1_n48, u_alu_add_x_1_n47,
         u_alu_add_x_1_n46, u_alu_add_x_1_n45, u_alu_add_x_1_n44,
         u_alu_add_x_1_n43, u_alu_add_x_1_n42, u_alu_add_x_1_n41,
         u_alu_add_x_1_n40, u_alu_add_x_1_n39, u_alu_add_x_1_n38,
         u_alu_add_x_1_n37, u_alu_add_x_1_n36, u_alu_add_x_1_n35,
         u_alu_add_x_1_n34, u_alu_add_x_1_n33, u_alu_add_x_1_n32,
         u_alu_add_x_1_n31, u_alu_add_x_1_n30, u_alu_add_x_1_n29,
         u_alu_add_x_1_n28, u_alu_add_x_1_n27, u_alu_add_x_1_n26,
         u_alu_add_x_1_n24, u_alu_add_x_1_n23, u_alu_add_x_1_n22,
         u_alu_add_x_1_n21, u_alu_add_x_1_n20, u_alu_add_x_1_n19,
         u_alu_add_x_1_n18, u_alu_add_x_1_n17, u_alu_add_x_1_n16,
         u_alu_add_x_1_n15, u_alu_add_x_1_n14, u_alu_add_x_1_n13,
         u_alu_add_x_1_n12, u_alu_add_x_1_n11, u_alu_add_x_1_n10,
         u_alu_add_x_1_n8, u_alu_add_x_1_n7, u_alu_add_x_1_n6,
         u_alu_add_x_1_n5, u_alu_add_x_1_n4, u_alu_add_x_1_n3,
         u_alu_add_x_1_n2, u_alu_add_x_1_n1, u_alu_DP_OP_84J3_125_2615_n15,
         u_alu_DP_OP_84J3_125_2615_n14, u_alu_DP_OP_84J3_125_2615_n13,
         u_alu_DP_OP_84J3_125_2615_n12, u_alu_DP_OP_84J3_125_2615_n11,
         u_alu_DP_OP_84J3_125_2615_n10, u_alu_DP_OP_84J3_125_2615_n9,
         u_alu_DP_OP_84J3_125_2615_n6, u_alu_DP_OP_84J3_125_2615_n5,
         u_alu_DP_OP_84J3_125_2615_n4, u_alu_DP_OP_84J3_125_2615_n3,
         u_alu_DP_OP_84J3_125_2615_n2, u_alu_DP_OP_84J3_125_2615_n1,
         u_alu_lt_x_11_B_7_, u_alu_lt_x_11_B_2_, u_alu_sub_x_2_n107,
         u_alu_sub_x_2_n103, u_alu_sub_x_2_n99, u_alu_sub_x_2_n95,
         u_alu_sub_x_2_n94, u_alu_sub_x_2_n92, u_alu_sub_x_2_n91,
         u_alu_sub_x_2_n90, u_alu_sub_x_2_n89, u_alu_sub_x_2_n88,
         u_alu_sub_x_2_n87, u_alu_sub_x_2_n86, u_alu_sub_x_2_n85,
         u_alu_sub_x_2_n84, u_alu_sub_x_2_n83, u_alu_sub_x_2_n82,
         u_alu_sub_x_2_n81, u_alu_sub_x_2_n80, u_alu_sub_x_2_n79,
         u_alu_sub_x_2_n78, u_alu_sub_x_2_n76, u_alu_sub_x_2_n75,
         u_alu_sub_x_2_n74, u_alu_sub_x_2_n73, u_alu_sub_x_2_n72,
         u_alu_sub_x_2_n71, u_alu_sub_x_2_n70, u_alu_sub_x_2_n69,
         u_alu_sub_x_2_n64, u_alu_sub_x_2_n63, u_alu_sub_x_2_n62,
         u_alu_sub_x_2_n61, u_alu_sub_x_2_n60, u_alu_sub_x_2_n59,
         u_alu_sub_x_2_n58, u_alu_sub_x_2_n57, u_alu_sub_x_2_n56,
         u_alu_sub_x_2_n55, u_alu_sub_x_2_n54, u_alu_sub_x_2_n53,
         u_alu_sub_x_2_n52, u_alu_sub_x_2_n51, u_alu_sub_x_2_n50,
         u_alu_sub_x_2_n49, u_alu_sub_x_2_n48, u_alu_sub_x_2_n47,
         u_alu_sub_x_2_n46, u_alu_sub_x_2_n45, u_alu_sub_x_2_n44,
         u_alu_sub_x_2_n43, u_alu_sub_x_2_n42, u_alu_sub_x_2_n41,
         u_alu_sub_x_2_n40, u_alu_sub_x_2_n39, u_alu_sub_x_2_n38,
         u_alu_sub_x_2_n37, u_alu_sub_x_2_n36, u_alu_sub_x_2_n34,
         u_alu_sub_x_2_n33, u_alu_sub_x_2_n32, u_alu_sub_x_2_n31,
         u_alu_sub_x_2_n30, u_alu_sub_x_2_n29, u_alu_sub_x_2_n28,
         u_alu_sub_x_2_n27, u_alu_sub_x_2_n26, u_alu_sub_x_2_n25,
         u_alu_sub_x_2_n24, u_alu_sub_x_2_n23, u_alu_sub_x_2_n22,
         u_alu_sub_x_2_n21, u_alu_sub_x_2_n19, u_alu_sub_x_2_n18,
         u_alu_sub_x_2_n17, u_alu_sub_x_2_n16, u_alu_sub_x_2_n15,
         u_alu_sub_x_2_n12, u_alu_sub_x_2_n11, u_alu_sub_x_2_n9,
         u_alu_sub_x_2_n8, u_alu_sub_x_2_n7, u_alu_sub_x_2_n6,
         u_alu_sub_x_2_n5, u_alu_sub_x_2_n4, u_alu_sub_x_2_n3,
         u_alu_sub_x_2_n2, u_alu_sub_x_2_n1, u_alu_DP_OP_85J3_126_1427_n214,
         u_alu_DP_OP_85J3_126_1427_n203, u_alu_DP_OP_85J3_126_1427_n202,
         u_alu_DP_OP_85J3_126_1427_n201, u_alu_DP_OP_85J3_126_1427_n200,
         u_alu_DP_OP_85J3_126_1427_n199, u_alu_DP_OP_85J3_126_1427_n198,
         u_alu_DP_OP_85J3_126_1427_n197, u_alu_DP_OP_85J3_126_1427_n196,
         u_alu_DP_OP_85J3_126_1427_n195, u_alu_DP_OP_85J3_126_1427_n193,
         u_alu_DP_OP_85J3_126_1427_n192, u_alu_DP_OP_85J3_126_1427_n191,
         u_alu_DP_OP_85J3_126_1427_n187, u_alu_DP_OP_85J3_126_1427_n186,
         u_alu_DP_OP_85J3_126_1427_n179, u_alu_DP_OP_85J3_126_1427_n176,
         u_alu_DP_OP_85J3_126_1427_n175, u_alu_DP_OP_85J3_126_1427_n174,
         u_alu_DP_OP_85J3_126_1427_n173, u_alu_DP_OP_85J3_126_1427_n166,
         u_alu_DP_OP_85J3_126_1427_n164, u_alu_DP_OP_85J3_126_1427_n157,
         u_alu_DP_OP_85J3_126_1427_n156, u_alu_DP_OP_85J3_126_1427_n155,
         u_alu_DP_OP_85J3_126_1427_n152, u_alu_DP_OP_85J3_126_1427_n148,
         u_alu_DP_OP_85J3_126_1427_n145, u_alu_DP_OP_85J3_126_1427_n143,
         u_alu_DP_OP_85J3_126_1427_n140, u_alu_DP_OP_85J3_126_1427_n137,
         u_alu_DP_OP_85J3_126_1427_n135, u_alu_DP_OP_85J3_126_1427_n132,
         u_alu_DP_OP_85J3_126_1427_n129, u_alu_DP_OP_85J3_126_1427_n127,
         u_alu_DP_OP_85J3_126_1427_n124, u_alu_DP_OP_85J3_126_1427_n123,
         u_alu_DP_OP_85J3_126_1427_n122, u_alu_DP_OP_85J3_126_1427_n95,
         u_alu_DP_OP_85J3_126_1427_n94, u_alu_DP_OP_85J3_126_1427_n93,
         u_alu_DP_OP_85J3_126_1427_n92, u_alu_DP_OP_85J3_126_1427_n91,
         u_alu_DP_OP_85J3_126_1427_n90, u_alu_DP_OP_85J3_126_1427_n89,
         u_alu_DP_OP_85J3_126_1427_n88, u_alu_DP_OP_85J3_126_1427_n83,
         u_alu_DP_OP_85J3_126_1427_n81, u_alu_DP_OP_85J3_126_1427_n80,
         u_alu_DP_OP_85J3_126_1427_n79, u_alu_DP_OP_85J3_126_1427_n76,
         u_alu_DP_OP_85J3_126_1427_n75, u_alu_DP_OP_85J3_126_1427_n74,
         u_alu_DP_OP_85J3_126_1427_n73, u_alu_DP_OP_85J3_126_1427_n66,
         u_alu_DP_OP_85J3_126_1427_n65, u_alu_DP_OP_85J3_126_1427_n64,
         u_alu_DP_OP_85J3_126_1427_n57, u_alu_DP_OP_85J3_126_1427_n56,
         u_alu_DP_OP_85J3_126_1427_n55, u_alu_DP_OP_85J3_126_1427_n52,
         u_alu_DP_OP_85J3_126_1427_n51, u_alu_DP_OP_85J3_126_1427_n50,
         u_alu_DP_OP_85J3_126_1427_n49, u_alu_DP_OP_85J3_126_1427_n48,
         u_alu_DP_OP_85J3_126_1427_n45, u_alu_DP_OP_85J3_126_1427_n44,
         u_alu_DP_OP_85J3_126_1427_n42, u_alu_DP_OP_85J3_126_1427_n41,
         u_alu_DP_OP_85J3_126_1427_n40, u_alu_DP_OP_85J3_126_1427_n37,
         u_alu_DP_OP_85J3_126_1427_n36, u_alu_DP_OP_85J3_126_1427_n34,
         u_alu_DP_OP_85J3_126_1427_n33, u_alu_DP_OP_85J3_126_1427_n32,
         u_alu_DP_OP_85J3_126_1427_n29, u_alu_DP_OP_85J3_126_1427_n28,
         u_alu_DP_OP_85J3_126_1427_n27, u_alu_DP_OP_85J3_126_1427_n26,
         u_alu_DP_OP_85J3_126_1427_n25, u_alu_DP_OP_85J3_126_1427_n24,
         u_alu_DP_OP_85J3_126_1427_n23, u_alu_DP_OP_85J3_126_1427_n21,
         u_alu_DP_OP_85J3_126_1427_n20, u_alu_DP_OP_85J3_126_1427_n18,
         u_alu_DP_OP_85J3_126_1427_n17, u_alu_DP_OP_85J3_126_1427_n16,
         u_alu_DP_OP_85J3_126_1427_n15, u_alu_DP_OP_85J3_126_1427_n14,
         u_alu_DP_OP_85J3_126_1427_n13, u_alu_DP_OP_85J3_126_1427_n12,
         u_alu_DP_OP_85J3_126_1427_n11, u_alu_DP_OP_85J3_126_1427_n10,
         u_alu_DP_OP_85J3_126_1427_n9, u_alu_DP_OP_85J3_126_1427_n8,
         u_alu_DP_OP_85J3_126_1427_n7, u_alu_DP_OP_85J3_126_1427_n6,
         u_alu_DP_OP_85J3_126_1427_n5, u_alu_DP_OP_85J3_126_1427_n4,
         u_alu_DP_OP_85J3_126_1427_n3, u_alu_DP_OP_85J3_126_1427_n2,
         u_alu_DP_OP_85J3_126_1427_n1, u_alu_DP_OP_83J3_124_3384_n15,
         u_alu_DP_OP_83J3_124_3384_n14, u_alu_DP_OP_83J3_124_3384_n13,
         u_alu_DP_OP_83J3_124_3384_n12, u_alu_DP_OP_83J3_124_3384_n11,
         u_alu_DP_OP_83J3_124_3384_n10, u_alu_DP_OP_83J3_124_3384_n9,
         u_alu_DP_OP_83J3_124_3384_n7, u_alu_DP_OP_83J3_124_3384_n6,
         u_alu_DP_OP_83J3_124_3384_n5, u_alu_DP_OP_83J3_124_3384_n4,
         u_alu_DP_OP_83J3_124_3384_n3, u_alu_DP_OP_83J3_124_3384_n2,
         u_alu_DP_OP_83J3_124_3384_n1, DP_OP_77_130_260_n30,
         DP_OP_77_130_260_n29, DP_OP_77_130_260_n28, DP_OP_77_130_260_n27,
         DP_OP_77_130_260_n24, DP_OP_77_130_260_n23, DP_OP_77_130_260_n22,
         DP_OP_77_130_260_n20, DP_OP_77_130_260_n19, DP_OP_77_130_260_n18,
         DP_OP_77_130_260_n17, DP_OP_77_130_260_n16, DP_OP_77_130_260_n15,
         DP_OP_77_130_260_n14, DP_OP_77_130_260_n11, DP_OP_77_130_260_n10,
         DP_OP_77_130_260_n9, DP_OP_77_130_260_n8, DP_OP_77_130_260_n7,
         DP_OP_77_130_260_n6, DP_OP_77_130_260_n4, DP_OP_77_130_260_n3,
         DP_OP_77_130_260_n2, DP_OP_77_130_260_n1, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336;
  wire   [31:0] alu_o_data_AluRes;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;
  wire   [15:0] u_alu_pre_subb;
  wire   [15:1] u_alu_pre_suba;
  wire   [7:1] u_alu_pre_sum_4b;
  wire   [7:0] u_alu_pre_sum_4a;
  wire   [8:1] u_alu_pre_sum_3b;
  wire   [8:0] u_alu_pre_sum_3a;

  DFC1 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC1 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC1 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC1 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC1 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC1 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_31_) );
  DFC1 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_30_) );
  DFC1 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_29_) );
  DFC1 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_28_) );
  DFC1 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_27_) );
  DFC1 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_26_) );
  DFC1 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_25_) );
  DFC1 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_24_) );
  DFC1 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_23_) );
  DFC1 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_22_) );
  DFC1 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_21_) );
  DFC1 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_20_) );
  DFC1 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_19_) );
  DFC1 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_18_) );
  DFC1 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_17_) );
  DFC1 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_16__BAR) );
  DFC1 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_15_) );
  DFC1 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_14_) );
  DFC1 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_13_) );
  DFC1 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_12_) );
  DFC1 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_11_) );
  DFC1 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_10_) );
  DFC1 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_9_) );
  DFC1 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_8_) );
  DFC1 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_7_) );
  DFC1 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_6_) );
  DFC1 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_5_) );
  DFC1 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_4_) );
  DFC1 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_3_) );
  DFC1 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_2_) );
  DFC1 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_1_) );
  DFC1 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_0_) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  DFC1 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC1 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC1 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC1 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC1 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC1 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC1 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC1 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC1 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC1 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC1 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC1 pipe_alures_reg_15_ ( .D(alu_o_data_AluRes[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[15]) );
  DFC1 pipe_alures_reg_14_ ( .D(alu_o_data_AluRes[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[14]) );
  DFC1 pipe_alures_reg_13_ ( .D(alu_o_data_AluRes[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[13]) );
  DFC1 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC1 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC1 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC1 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC1 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC1 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC1 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC1 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC1 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC1 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC1 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC1 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC1 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC1 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC1 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC1 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC1 pipe_rt_reg_28_ ( .D(compare_i_data_rt[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[28]) );
  DFC1 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  DFC1 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC1 pipe_rt_reg_25_ ( .D(compare_i_data_rt[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[25]) );
  DFC1 pipe_rt_reg_24_ ( .D(compare_i_data_rt[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[24]) );
  DFC1 pipe_rt_reg_23_ ( .D(compare_i_data_rt[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[23]) );
  DFC1 pipe_rt_reg_22_ ( .D(compare_i_data_rt[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[22]) );
  DFC1 pipe_rt_reg_21_ ( .D(compare_i_data_rt[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[21]) );
  DFC1 pipe_rt_reg_20_ ( .D(compare_i_data_rt[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[20]) );
  DFC1 pipe_rt_reg_19_ ( .D(compare_i_data_rt[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[19]) );
  DFC1 pipe_rt_reg_18_ ( .D(compare_i_data_rt[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[18]) );
  DFC1 pipe_rt_reg_17_ ( .D(compare_i_data_rt[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[17]) );
  DFC1 pipe_rt_reg_16_ ( .D(compare_i_data_rt[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[16]) );
  DFC1 pipe_rt_reg_15_ ( .D(compare_i_data_rt[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[15]) );
  DFC1 pipe_rt_reg_14_ ( .D(compare_i_data_rt[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[14]) );
  DFC1 pipe_rt_reg_13_ ( .D(compare_i_data_rt[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[13]) );
  DFC1 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC1 pipe_rt_reg_11_ ( .D(compare_i_data_rt[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[11]) );
  DFC1 pipe_rt_reg_10_ ( .D(compare_i_data_rt[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[10]) );
  DFC1 pipe_rt_reg_9_ ( .D(compare_i_data_rt[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[9]) );
  DFC1 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC1 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC1 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC1 pipe_rt_reg_5_ ( .D(compare_i_data_rt[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[5]) );
  DFC1 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC1 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC1 pipe_rt_reg_2_ ( .D(compare_i_data_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[2]) );
  DFC1 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC1 pipe_rt_reg_0_ ( .D(compare_i_data_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[0]) );
  DFC1 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC1 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC1 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC1 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC1 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC1 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC1 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC1 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC1 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  XNR21 u_alu_add_x_1_U2 ( .A(u_alu_add_x_1_n1), .B(u_alu_add_x_1_n16), .Q(
        u_alu_sum_1_7_) );
  XNR21 u_alu_add_x_1_U34 ( .A(u_alu_add_x_1_n5), .B(u_alu_add_x_1_n35), .Q(
        u_alu_sum_1_3_) );
  XNR21 u_alu_add_x_1_U26 ( .A(u_alu_add_x_1_n4), .B(u_alu_add_x_1_n29), .Q(
        u_alu_sum_1_4_) );
  NAND22 u_alu_add_x_1_U60 ( .A(n81), .B(compare_i_data_rs[0]), .Q(
        u_alu_add_x_1_n43) );
  OAI212 u_alu_add_x_1_U51 ( .A(u_alu_add_x_1_n43), .B(u_alu_add_x_1_n40), .C(
        u_alu_add_x_1_n41), .Q(u_alu_add_x_1_n39) );
  OAI212 u_alu_add_x_1_U21 ( .A(u_alu_add_x_1_n28), .B(u_alu_add_x_1_n22), .C(
        u_alu_add_x_1_n23), .Q(u_alu_add_x_1_n21) );
  NAND22 u_alu_add_x_1_U17 ( .A(n112), .B(compare_i_data_rs[6]), .Q(
        u_alu_add_x_1_n18) );
  OAI212 u_alu_add_x_1_U3 ( .A(u_alu_add_x_1_n10), .B(u_alu_add_x_1_n30), .C(
        u_alu_add_x_1_n11), .Q(u_alu_sum_1_8_) );
  AOI211 u_alu_add_x_1_U27 ( .A(u_alu_add_x_1_n29), .B(u_alu_add_x_1_n47), .C(
        u_alu_add_x_1_n26), .Q(u_alu_add_x_1_n24) );
  XOR21 u_alu_add_x_1_U18 ( .A(u_alu_add_x_1_n3), .B(u_alu_add_x_1_n24), .Q(
        u_alu_sum_1_5_) );
  XOR21 u_alu_add_x_1_U43 ( .A(u_alu_add_x_1_n6), .B(u_alu_add_x_1_n38), .Q(
        u_alu_sum_1_2_) );
  NOR20 u_alu_add_x_1_U59 ( .A(compare_i_data_rs[0]), .B(n81), .Q(
        u_alu_add_x_1_n42) );
  OAI210 u_alu_add_x_1_U44 ( .A(u_alu_add_x_1_n36), .B(u_alu_add_x_1_n38), .C(
        u_alu_add_x_1_n37), .Q(u_alu_add_x_1_n35) );
  OAI212 u_alu_add_x_1_U38 ( .A(u_alu_add_x_1_n37), .B(u_alu_add_x_1_n33), .C(
        u_alu_add_x_1_n34), .Q(u_alu_add_x_1_n32) );
  NAND22 u_alu_add_x_1_U33 ( .A(alu_i_data_B[4]), .B(compare_i_data_rs[4]), 
        .Q(u_alu_add_x_1_n28) );
  OAI210 u_alu_add_x_1_U13 ( .A(u_alu_add_x_1_n17), .B(u_alu_add_x_1_n19), .C(
        u_alu_add_x_1_n18), .Q(u_alu_add_x_1_n16) );
  NAND22 u_alu_add_x_1_U48 ( .A(u_alu_lt_x_11_B_2_), .B(compare_i_data_rs[2]), 
        .Q(u_alu_add_x_1_n37) );
  NAND22 u_alu_add_x_1_U25 ( .A(alu_i_data_B[5]), .B(compare_i_data_rs[5]), 
        .Q(u_alu_add_x_1_n23) );
  NAND22 u_alu_add_x_1_U11 ( .A(alu_i_data_B[7]), .B(compare_i_data_rs[7]), 
        .Q(u_alu_add_x_1_n15) );
  AOI210 u_alu_add_x_1_U19 ( .A(u_alu_add_x_1_n29), .B(u_alu_add_x_1_n20), .C(
        u_alu_add_x_1_n21), .Q(u_alu_add_x_1_n19) );
  AOI212 u_alu_add_x_1_U36 ( .A(u_alu_add_x_1_n39), .B(u_alu_add_x_1_n31), .C(
        u_alu_add_x_1_n32), .Q(u_alu_add_x_1_n30) );
  XOR20 u_alu_add_x_1_U49 ( .A(u_alu_add_x_1_n43), .B(u_alu_add_x_1_n7), .Q(
        u_alu_sum_1_1_) );
  NOR22 u_alu_add_x_1_U41 ( .A(compare_i_data_rs[3]), .B(alu_i_data_B[3]), .Q(
        u_alu_add_x_1_n33) );
  OAI212 u_alu_add_x_1_U7 ( .A(u_alu_add_x_1_n18), .B(u_alu_add_x_1_n14), .C(
        u_alu_add_x_1_n15), .Q(u_alu_add_x_1_n13) );
  XOR20 u_alu_add_x_1_U12 ( .A(u_alu_add_x_1_n2), .B(u_alu_add_x_1_n19), .Q(
        u_alu_sum_1_6_) );
  NOR21 u_alu_add_x_1_U20 ( .A(u_alu_add_x_1_n27), .B(u_alu_add_x_1_n22), .Q(
        u_alu_add_x_1_n20) );
  NOR22 u_alu_add_x_1_U10 ( .A(compare_i_data_rs[7]), .B(alu_i_data_B[7]), .Q(
        u_alu_add_x_1_n14) );
  NOR22 u_alu_add_x_1_U6 ( .A(u_alu_add_x_1_n17), .B(u_alu_add_x_1_n14), .Q(
        u_alu_add_x_1_n12) );
  NOR21 u_alu_add_x_1_U37 ( .A(u_alu_add_x_1_n36), .B(u_alu_add_x_1_n33), .Q(
        u_alu_add_x_1_n31) );
  AOI211 u_alu_add_x_1_U5 ( .A(u_alu_add_x_1_n21), .B(u_alu_add_x_1_n12), .C(
        u_alu_add_x_1_n13), .Q(u_alu_add_x_1_n11) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U12 ( .A(compare_i_data_rs[29]), .B(
        alu_i_data_B[29]), .CI(u_alu_DP_OP_84J3_125_2615_n11), .CO(
        u_alu_DP_OP_84J3_125_2615_n10), .S(u_alu_pre_sum_4a[5]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U4 ( .A(u_alu_pre_sum_4a[4]), .B(
        u_alu_DP_OP_84J3_125_2615_n4), .CO(u_alu_DP_OP_84J3_125_2615_n3), .S(
        u_alu_pre_sum_4b[4]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U5 ( .A(u_alu_pre_sum_4a[3]), .B(
        u_alu_DP_OP_84J3_125_2615_n5), .CO(u_alu_DP_OP_84J3_125_2615_n4), .S(
        u_alu_pre_sum_4b[3]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U6 ( .A(u_alu_pre_sum_4a[2]), .B(
        u_alu_DP_OP_84J3_125_2615_n6), .CO(u_alu_DP_OP_84J3_125_2615_n5), .S(
        u_alu_pre_sum_4b[2]) );
  NAND22 u_alu_sub_x_2_U47 ( .A(u_alu_sub_x_2_n89), .B(u_alu_sub_x_2_n45), .Q(
        u_alu_sub_x_2_n6) );
  NAND22 u_alu_sub_x_2_U40 ( .A(u_alu_sub_x_2_n103), .B(compare_i_data_rs[10]), 
        .Q(u_alu_sub_x_2_n38) );
  NAND22 u_alu_sub_x_2_U50 ( .A(n116), .B(compare_i_data_rs[9]), .Q(
        u_alu_sub_x_2_n45) );
  NAND22 u_alu_sub_x_2_U81 ( .A(n232), .B(compare_i_data_rs[5]), .Q(
        u_alu_sub_x_2_n64) );
  NAND22 u_alu_sub_x_2_U104 ( .A(n111), .B(compare_i_data_rs[2]), .Q(
        u_alu_sub_x_2_n78) );
  NAND22 u_alu_sub_x_2_U89 ( .A(n115), .B(compare_i_data_rs[4]), .Q(
        u_alu_sub_x_2_n69) );
  XOR20 u_alu_sub_x_2_U17 ( .A(u_alu_sub_x_2_n3), .B(u_alu_sub_x_2_n27), .Q(
        u_alu_half_sub_12_) );
  NAND20 u_alu_sub_x_2_U19 ( .A(u_alu_sub_x_2_n86), .B(u_alu_sub_x_2_n26), .Q(
        u_alu_sub_x_2_n3) );
  NOR21 u_alu_sub_x_2_U80 ( .A(compare_i_data_rs[5]), .B(n232), .Q(
        u_alu_sub_x_2_n63) );
  XOR21 u_alu_sub_x_2_U68 ( .A(u_alu_sub_x_2_n9), .B(u_alu_sub_x_2_n60), .Q(
        u_alu_half_sub_6_) );
  AOI211 u_alu_sub_x_2_U75 ( .A(u_alu_sub_x_2_n70), .B(u_alu_sub_x_2_n61), .C(
        u_alu_sub_x_2_n62), .Q(u_alu_sub_x_2_n60) );
  NAND22 u_alu_sub_x_2_U70 ( .A(u_alu_sub_x_2_n92), .B(u_alu_sub_x_2_n59), .Q(
        u_alu_sub_x_2_n9) );
  OAI212 u_alu_sub_x_2_U42 ( .A(u_alu_sub_x_2_n40), .B(u_alu_sub_x_2_n49), .C(
        u_alu_sub_x_2_n41), .Q(u_alu_sub_x_2_n39) );
  XOR21 u_alu_sub_x_2_U51 ( .A(u_alu_sub_x_2_n7), .B(u_alu_sub_x_2_n49), .Q(
        u_alu_half_sub_8_) );
  OAI212 u_alu_sub_x_2_U4 ( .A(u_alu_sub_x_2_n17), .B(u_alu_sub_x_2_n19), .C(
        u_alu_sub_x_2_n18), .Q(u_alu_sub_x_2_n16) );
  NAND22 u_alu_sub_x_2_U8 ( .A(u_alu_sub_x_2_n99), .B(compare_i_data_rs[14]), 
        .Q(u_alu_sub_x_2_n18) );
  NAND22 u_alu_sub_x_2_U16 ( .A(n110), .B(compare_i_data_rs[13]), .Q(
        u_alu_sub_x_2_n23) );
  NOR21 u_alu_sub_x_2_U15 ( .A(compare_i_data_rs[13]), .B(n110), .Q(
        u_alu_sub_x_2_n22) );
  OAI212 u_alu_sub_x_2_U18 ( .A(u_alu_sub_x_2_n25), .B(u_alu_sub_x_2_n27), .C(
        u_alu_sub_x_2_n26), .Q(u_alu_sub_x_2_n24) );
  NAND22 u_alu_sub_x_2_U22 ( .A(n94), .B(compare_i_data_rs[12]), .Q(
        u_alu_sub_x_2_n26) );
  AOI211 u_alu_sub_x_2_U34 ( .A(u_alu_sub_x_2_n43), .B(u_alu_sub_x_2_n88), .C(
        u_alu_sub_x_2_n36), .Q(u_alu_sub_x_2_n34) );
  NAND22 u_alu_sub_x_2_U56 ( .A(n95), .B(compare_i_data_rs[8]), .Q(
        u_alu_sub_x_2_n48) );
  NOR21 u_alu_sub_x_2_U25 ( .A(u_alu_sub_x_2_n30), .B(u_alu_sub_x_2_n33), .Q(
        u_alu_sub_x_2_n28) );
  NAND22 u_alu_sub_x_2_U33 ( .A(u_alu_sub_x_2_n42), .B(u_alu_sub_x_2_n88), .Q(
        u_alu_sub_x_2_n33) );
  NOR21 u_alu_sub_x_2_U39 ( .A(compare_i_data_rs[10]), .B(u_alu_sub_x_2_n103), 
        .Q(u_alu_sub_x_2_n37) );
  NOR21 u_alu_sub_x_2_U45 ( .A(u_alu_sub_x_2_n47), .B(u_alu_sub_x_2_n44), .Q(
        u_alu_sub_x_2_n42) );
  NOR21 u_alu_sub_x_2_U49 ( .A(compare_i_data_rs[9]), .B(n116), .Q(
        u_alu_sub_x_2_n44) );
  NOR21 u_alu_sub_x_2_U55 ( .A(compare_i_data_rs[8]), .B(n95), .Q(
        u_alu_sub_x_2_n47) );
  NOR21 u_alu_sub_x_2_U29 ( .A(compare_i_data_rs[11]), .B(n96), .Q(
        u_alu_sub_x_2_n30) );
  OAI212 u_alu_sub_x_2_U59 ( .A(u_alu_sub_x_2_n51), .B(u_alu_sub_x_2_n71), .C(
        u_alu_sub_x_2_n52), .Q(u_alu_sub_x_2_n50) );
  AOI211 u_alu_sub_x_2_U61 ( .A(u_alu_sub_x_2_n62), .B(u_alu_sub_x_2_n53), .C(
        u_alu_sub_x_2_n54), .Q(u_alu_sub_x_2_n52) );
  NAND22 u_alu_sub_x_2_U73 ( .A(u_alu_sub_x_2_n107), .B(compare_i_data_rs[6]), 
        .Q(u_alu_sub_x_2_n59) );
  OAI212 u_alu_sub_x_2_U77 ( .A(u_alu_sub_x_2_n69), .B(u_alu_sub_x_2_n63), .C(
        u_alu_sub_x_2_n64), .Q(u_alu_sub_x_2_n62) );
  NOR21 u_alu_sub_x_2_U93 ( .A(n155), .B(u_alu_sub_x_2_n74), .Q(
        u_alu_sub_x_2_n72) );
  OAI212 u_alu_sub_x_2_U107 ( .A(u_alu_sub_x_2_n83), .B(u_alu_sub_x_2_n81), 
        .C(u_alu_sub_x_2_n82), .Q(u_alu_sub_x_2_n80) );
  NOR21 u_alu_sub_x_2_U113 ( .A(compare_i_data_rs[0]), .B(n114), .Q(
        u_alu_sub_x_2_n83) );
  NAND22 u_alu_sub_x_2_U60 ( .A(u_alu_sub_x_2_n61), .B(u_alu_sub_x_2_n53), .Q(
        u_alu_sub_x_2_n51) );
  NOR21 u_alu_sub_x_2_U62 ( .A(u_alu_sub_x_2_n58), .B(u_alu_sub_x_2_n55), .Q(
        u_alu_sub_x_2_n53) );
  NOR21 u_alu_sub_x_2_U66 ( .A(compare_i_data_rs[7]), .B(n233), .Q(
        u_alu_sub_x_2_n55) );
  NOR21 u_alu_sub_x_2_U72 ( .A(compare_i_data_rs[6]), .B(u_alu_sub_x_2_n107), 
        .Q(u_alu_sub_x_2_n58) );
  NOR21 u_alu_sub_x_2_U76 ( .A(n161), .B(u_alu_sub_x_2_n63), .Q(
        u_alu_sub_x_2_n61) );
  NOR21 u_alu_sub_x_2_U21 ( .A(compare_i_data_rs[12]), .B(n94), .Q(
        u_alu_sub_x_2_n25) );
  NOR21 u_alu_sub_x_2_U7 ( .A(compare_i_data_rs[14]), .B(u_alu_sub_x_2_n99), 
        .Q(u_alu_sub_x_2_n17) );
  XNR21 u_alu_sub_x_2_U112 ( .A(compare_i_data_rs[0]), .B(n114), .Q(
        u_alu_half_sub_0_) );
  XNR21 u_alu_sub_x_2_U82 ( .A(u_alu_sub_x_2_n11), .B(u_alu_sub_x_2_n70), .Q(
        u_alu_half_sub_4_) );
  XNR21 u_alu_sub_x_2_U90 ( .A(u_alu_sub_x_2_n12), .B(u_alu_sub_x_2_n76), .Q(
        u_alu_half_sub_3_) );
  XNR21 u_alu_sub_x_2_U9 ( .A(u_alu_sub_x_2_n2), .B(u_alu_sub_x_2_n24), .Q(
        u_alu_half_sub_13_) );
  XNR21 u_alu_sub_x_2_U57 ( .A(u_alu_sub_x_2_n8), .B(u_alu_sub_x_2_n57), .Q(
        u_alu_half_sub_7_) );
  XNR21 u_alu_sub_x_2_U41 ( .A(u_alu_sub_x_2_n6), .B(u_alu_sub_x_2_n46), .Q(
        u_alu_half_sub_9_) );
  XNR21 u_alu_sub_x_2_U31 ( .A(u_alu_sub_x_2_n5), .B(u_alu_sub_x_2_n39), .Q(
        u_alu_half_sub_10_) );
  XNR21 u_alu_sub_x_2_U23 ( .A(u_alu_sub_x_2_n4), .B(u_alu_sub_x_2_n32), .Q(
        u_alu_half_sub_11_) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U30 ( .A(u_alu_DP_OP_85J3_126_1427_n193), 
        .B(u_alu_DP_OP_85J3_126_1427_n33), .Q(u_alu_DP_OP_85J3_126_1427_n5) );
  AOI211 u_alu_DP_OP_85J3_126_1427_U73 ( .A(u_alu_DP_OP_85J3_126_1427_n75), 
        .B(u_alu_DP_OP_85J3_126_1427_n156), .C(u_alu_DP_OP_85J3_126_1427_n157), 
        .Q(u_alu_DP_OP_85J3_126_1427_n57) );
  AOI211 u_alu_DP_OP_85J3_126_1427_U181 ( .A(u_alu_DP_OP_85J3_126_1427_n173), 
        .B(u_alu_DP_OP_85J3_126_1427_n156), .C(u_alu_DP_OP_85J3_126_1427_n157), 
        .Q(u_alu_DP_OP_85J3_126_1427_n155) );
  NOR20 u_alu_DP_OP_85J3_126_1427_U4 ( .A(n91), .B(alu_i_data_B[31]), .Q(
        u_alu_DP_OP_85J3_126_1427_n16) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U25 ( .A(n113), .B(compare_i_data_rs[28]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n28) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U33 ( .A(n93), .B(compare_i_data_rs[27]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n33) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U39 ( .A(n85), .B(compare_i_data_rs[26]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n36) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U114 ( .A(n84), .B(compare_i_data_rs[18]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n83) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U127 ( .A(n90), .B(compare_i_data_rs[29]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n124), .CO(
        u_alu_DP_OP_85J3_126_1427_n123), .S(u_alu_pre_subb[13]) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U83 ( .A(n92), .B(compare_i_data_rs[21]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n65) );
  XOR20 u_alu_DP_OP_85J3_126_1427_U20 ( .A(u_alu_DP_OP_85J3_126_1427_n4), .B(
        u_alu_DP_OP_85J3_126_1427_n29), .Q(u_alu_pre_suba[12]) );
  XOR20 u_alu_DP_OP_85J3_126_1427_U142 ( .A(u_alu_DP_OP_85J3_126_1427_n6), .B(
        u_alu_DP_OP_85J3_126_1427_n135), .Q(u_alu_pre_subb[10]) );
  XOR20 u_alu_DP_OP_85J3_126_1427_U34 ( .A(u_alu_DP_OP_85J3_126_1427_n6), .B(
        u_alu_DP_OP_85J3_126_1427_n37), .Q(u_alu_pre_suba[10]) );
  XOR20 u_alu_DP_OP_85J3_126_1427_U156 ( .A(u_alu_DP_OP_85J3_126_1427_n8), .B(
        u_alu_DP_OP_85J3_126_1427_n143), .Q(u_alu_pre_subb[8]) );
  XOR20 u_alu_DP_OP_85J3_126_1427_U48 ( .A(u_alu_DP_OP_85J3_126_1427_n8), .B(
        u_alu_DP_OP_85J3_126_1427_n45), .Q(u_alu_pre_suba[8]) );
  XOR20 u_alu_DP_OP_85J3_126_1427_U128 ( .A(u_alu_DP_OP_85J3_126_1427_n4), .B(
        u_alu_DP_OP_85J3_126_1427_n127), .Q(u_alu_pre_subb[12]) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U117 ( .A(u_alu_DP_OP_85J3_126_1427_n92), 
        .B(u_alu_DP_OP_85J3_126_1427_n90), .C(u_alu_DP_OP_85J3_126_1427_n91), 
        .Q(u_alu_DP_OP_85J3_126_1427_n89) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U187 ( .A(u_alu_DP_OP_85J3_126_1427_n74), 
        .B(u_alu_DP_OP_85J3_126_1427_n64), .C(u_alu_DP_OP_85J3_126_1427_n65), 
        .Q(u_alu_DP_OP_85J3_126_1427_n157) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U208 ( .A(u_alu_DP_OP_85J3_126_1427_n83), 
        .B(u_alu_DP_OP_85J3_126_1427_n79), .C(u_alu_DP_OP_85J3_126_1427_n80), 
        .Q(u_alu_DP_OP_85J3_126_1427_n176) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U225 ( .A(u_alu_DP_OP_85J3_126_1427_n191), 
        .B(u_alu_DP_OP_85J3_126_1427_n90), .C(u_alu_DP_OP_85J3_126_1427_n91), 
        .Q(u_alu_DP_OP_85J3_126_1427_n187) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U36 ( .A(n219), .B(
        u_alu_DP_OP_85J3_126_1427_n36), .Q(u_alu_DP_OP_85J3_126_1427_n6) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U22 ( .A(u_alu_DP_OP_85J3_126_1427_n192), 
        .B(u_alu_DP_OP_85J3_126_1427_n28), .Q(u_alu_DP_OP_85J3_126_1427_n4) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U101 ( .A(u_alu_DP_OP_85J3_126_1427_n201), 
        .B(u_alu_DP_OP_85J3_126_1427_n80), .Q(u_alu_DP_OP_85J3_126_1427_n13)
         );
  NAND22 u_alu_DP_OP_85J3_126_1427_U92 ( .A(u_alu_DP_OP_85J3_126_1427_n200), 
        .B(u_alu_DP_OP_85J3_126_1427_n74), .Q(u_alu_DP_OP_85J3_126_1427_n12)
         );
  AOI211 u_alu_DP_OP_85J3_126_1427_U85 ( .A(u_alu_DP_OP_85J3_126_1427_n75), 
        .B(u_alu_DP_OP_85J3_126_1427_n200), .C(u_alu_DP_OP_85J3_126_1427_n166), 
        .Q(u_alu_DP_OP_85J3_126_1427_n66) );
  XOR21 u_alu_DP_OP_85J3_126_1427_U180 ( .A(u_alu_DP_OP_85J3_126_1427_n11), 
        .B(u_alu_DP_OP_85J3_126_1427_n164), .Q(u_alu_pre_subb[5]) );
  AOI211 u_alu_DP_OP_85J3_126_1427_U193 ( .A(u_alu_DP_OP_85J3_126_1427_n173), 
        .B(u_alu_DP_OP_85J3_126_1427_n200), .C(u_alu_DP_OP_85J3_126_1427_n166), 
        .Q(u_alu_DP_OP_85J3_126_1427_n164) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U80 ( .A(u_alu_DP_OP_85J3_126_1427_n199), 
        .B(u_alu_DP_OP_85J3_126_1427_n65), .Q(u_alu_DP_OP_85J3_126_1427_n11)
         );
  XOR21 u_alu_DP_OP_85J3_126_1427_U62 ( .A(u_alu_DP_OP_85J3_126_1427_n10), .B(
        u_alu_DP_OP_85J3_126_1427_n57), .Q(u_alu_pre_suba[6]) );
  XOR21 u_alu_DP_OP_85J3_126_1427_U170 ( .A(u_alu_DP_OP_85J3_126_1427_n10), 
        .B(u_alu_DP_OP_85J3_126_1427_n155), .Q(u_alu_pre_subb[6]) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U68 ( .A(u_alu_DP_OP_85J3_126_1427_n198), 
        .B(u_alu_DP_OP_85J3_126_1427_n56), .Q(u_alu_DP_OP_85J3_126_1427_n10)
         );
  NAND22 u_alu_DP_OP_85J3_126_1427_U44 ( .A(u_alu_DP_OP_85J3_126_1427_n195), 
        .B(u_alu_DP_OP_85J3_126_1427_n41), .Q(u_alu_DP_OP_85J3_126_1427_n7) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U7 ( .A(n145), .B(
        u_alu_DP_OP_85J3_126_1427_n21), .C(u_alu_DP_OP_85J3_126_1427_n20), .Q(
        u_alu_DP_OP_85J3_126_1427_n18) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U2 ( .A(u_alu_DP_OP_85J3_126_1427_n93), .B(
        u_alu_DP_OP_85J3_126_1427_n17), .Q(u_alu_DP_OP_85J3_126_1427_n1) );
  XOR21 u_alu_DP_OP_85J3_126_1427_U6 ( .A(u_alu_DP_OP_85J3_126_1427_n2), .B(
        u_alu_DP_OP_85J3_126_1427_n21), .Q(u_alu_pre_suba[14]) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U8 ( .A(u_alu_DP_OP_85J3_126_1427_n94), .B(
        u_alu_DP_OP_85J3_126_1427_n20), .Q(u_alu_DP_OP_85J3_126_1427_n2) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U50 ( .A(u_alu_DP_OP_85J3_126_1427_n196), 
        .B(u_alu_DP_OP_85J3_126_1427_n44), .Q(u_alu_DP_OP_85J3_126_1427_n8) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U129 ( .A(u_alu_DP_OP_85J3_126_1427_n27), 
        .B(u_alu_DP_OP_85J3_126_1427_n127), .C(u_alu_DP_OP_85J3_126_1427_n28), 
        .Q(u_alu_DP_OP_85J3_126_1427_n124) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U143 ( .A(n141), .B(
        u_alu_DP_OP_85J3_126_1427_n135), .C(u_alu_DP_OP_85J3_126_1427_n36), 
        .Q(u_alu_DP_OP_85J3_126_1427_n132) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U157 ( .A(n140), .B(
        u_alu_DP_OP_85J3_126_1427_n143), .C(u_alu_DP_OP_85J3_126_1427_n44), 
        .Q(u_alu_DP_OP_85J3_126_1427_n140) );
  AOI211 u_alu_DP_OP_85J3_126_1427_U163 ( .A(u_alu_DP_OP_85J3_126_1427_n148), 
        .B(u_alu_DP_OP_85J3_126_1427_n197), .C(u_alu_DP_OP_85J3_126_1427_n145), 
        .Q(u_alu_DP_OP_85J3_126_1427_n143) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U21 ( .A(u_alu_DP_OP_85J3_126_1427_n27), 
        .B(u_alu_DP_OP_85J3_126_1427_n29), .C(u_alu_DP_OP_85J3_126_1427_n28), 
        .Q(u_alu_DP_OP_85J3_126_1427_n26) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U35 ( .A(n141), .B(
        u_alu_DP_OP_85J3_126_1427_n37), .C(u_alu_DP_OP_85J3_126_1427_n36), .Q(
        u_alu_DP_OP_85J3_126_1427_n34) );
  AOI211 u_alu_DP_OP_85J3_126_1427_U41 ( .A(u_alu_DP_OP_85J3_126_1427_n42), 
        .B(u_alu_DP_OP_85J3_126_1427_n195), .C(u_alu_DP_OP_85J3_126_1427_n137), 
        .Q(u_alu_DP_OP_85J3_126_1427_n37) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U47 ( .A(u_alu_DP_OP_85J3_126_1427_n214), 
        .B(compare_i_data_rs[25]), .Q(u_alu_DP_OP_85J3_126_1427_n41) );
  NOR21 u_alu_DP_OP_85J3_126_1427_U46 ( .A(compare_i_data_rs[25]), .B(
        u_alu_DP_OP_85J3_126_1427_n214), .Q(u_alu_DP_OP_85J3_126_1427_n40) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U49 ( .A(n140), .B(
        u_alu_DP_OP_85J3_126_1427_n45), .C(u_alu_DP_OP_85J3_126_1427_n44), .Q(
        u_alu_DP_OP_85J3_126_1427_n42) );
  AOI211 u_alu_DP_OP_85J3_126_1427_U55 ( .A(u_alu_DP_OP_85J3_126_1427_n50), 
        .B(u_alu_DP_OP_85J3_126_1427_n197), .C(u_alu_DP_OP_85J3_126_1427_n145), 
        .Q(u_alu_DP_OP_85J3_126_1427_n45) );
  NOR21 u_alu_DP_OP_85J3_126_1427_U24 ( .A(compare_i_data_rs[28]), .B(n113), 
        .Q(u_alu_DP_OP_85J3_126_1427_n27) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U16 ( .A(u_alu_DP_OP_85J3_126_1427_n95), 
        .B(u_alu_DP_OP_85J3_126_1427_n25), .Q(u_alu_DP_OP_85J3_126_1427_n3) );
  XOR21 u_alu_DP_OP_85J3_126_1427_U105 ( .A(u_alu_DP_OP_85J3_126_1427_n14), 
        .B(u_alu_DP_OP_85J3_126_1427_n88), .Q(u_alu_pre_suba[2]) );
  XOR21 u_alu_DP_OP_85J3_126_1427_U213 ( .A(u_alu_DP_OP_85J3_126_1427_n14), 
        .B(u_alu_DP_OP_85J3_126_1427_n186), .Q(u_alu_pre_subb[2]) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U111 ( .A(u_alu_DP_OP_85J3_126_1427_n202), 
        .B(u_alu_DP_OP_85J3_126_1427_n83), .Q(u_alu_DP_OP_85J3_126_1427_n14)
         );
  OAI212 u_alu_DP_OP_85J3_126_1427_U63 ( .A(u_alu_DP_OP_85J3_126_1427_n51), 
        .B(u_alu_DP_OP_85J3_126_1427_n76), .C(u_alu_DP_OP_85J3_126_1427_n52), 
        .Q(u_alu_DP_OP_85J3_126_1427_n50) );
  AOI211 u_alu_DP_OP_85J3_126_1427_U98 ( .A(u_alu_DP_OP_85J3_126_1427_n89), 
        .B(u_alu_DP_OP_85J3_126_1427_n175), .C(u_alu_DP_OP_85J3_126_1427_n176), 
        .Q(u_alu_DP_OP_85J3_126_1427_n76) );
  OAI212 u_alu_DP_OP_85J3_126_1427_U171 ( .A(u_alu_DP_OP_85J3_126_1427_n51), 
        .B(u_alu_DP_OP_85J3_126_1427_n174), .C(u_alu_DP_OP_85J3_126_1427_n52), 
        .Q(u_alu_DP_OP_85J3_126_1427_n148) );
  AOI211 u_alu_DP_OP_85J3_126_1427_U65 ( .A(u_alu_DP_OP_85J3_126_1427_n157), 
        .B(u_alu_DP_OP_85J3_126_1427_n198), .C(u_alu_DP_OP_85J3_126_1427_n152), 
        .Q(u_alu_DP_OP_85J3_126_1427_n52) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U71 ( .A(n99), .B(compare_i_data_rs[22]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n56) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U95 ( .A(n82), .B(compare_i_data_rs[20]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n74) );
  AOI211 u_alu_DP_OP_85J3_126_1427_U206 ( .A(u_alu_DP_OP_85J3_126_1427_n187), 
        .B(u_alu_DP_OP_85J3_126_1427_n175), .C(u_alu_DP_OP_85J3_126_1427_n176), 
        .Q(u_alu_DP_OP_85J3_126_1427_n174) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U64 ( .A(u_alu_DP_OP_85J3_126_1427_n156), 
        .B(u_alu_DP_OP_85J3_126_1427_n198), .Q(u_alu_DP_OP_85J3_126_1427_n51)
         );
  NOR21 u_alu_DP_OP_85J3_126_1427_U70 ( .A(compare_i_data_rs[22]), .B(n99), 
        .Q(u_alu_DP_OP_85J3_126_1427_n55) );
  NOR21 u_alu_DP_OP_85J3_126_1427_U186 ( .A(u_alu_DP_OP_85J3_126_1427_n73), 
        .B(u_alu_DP_OP_85J3_126_1427_n64), .Q(u_alu_DP_OP_85J3_126_1427_n156)
         );
  NOR21 u_alu_DP_OP_85J3_126_1427_U94 ( .A(compare_i_data_rs[20]), .B(n82), 
        .Q(u_alu_DP_OP_85J3_126_1427_n73) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U58 ( .A(u_alu_DP_OP_85J3_126_1427_n197), 
        .B(u_alu_DP_OP_85J3_126_1427_n49), .Q(u_alu_DP_OP_85J3_126_1427_n9) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U61 ( .A(n109), .B(compare_i_data_rs[23]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n49) );
  NOR21 u_alu_DP_OP_85J3_126_1427_U60 ( .A(compare_i_data_rs[23]), .B(n109), 
        .Q(u_alu_DP_OP_85J3_126_1427_n48) );
  XOR21 u_alu_DP_OP_85J3_126_1427_U115 ( .A(u_alu_DP_OP_85J3_126_1427_n92), 
        .B(u_alu_DP_OP_85J3_126_1427_n15), .Q(u_alu_pre_suba[1]) );
  XOR21 u_alu_DP_OP_85J3_126_1427_U223 ( .A(u_alu_DP_OP_85J3_126_1427_n191), 
        .B(u_alu_DP_OP_85J3_126_1427_n15), .Q(u_alu_pre_subb[1]) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U118 ( .A(u_alu_DP_OP_85J3_126_1427_n203), 
        .B(u_alu_DP_OP_85J3_126_1427_n91), .Q(u_alu_DP_OP_85J3_126_1427_n15)
         );
  XNR21 u_alu_DP_OP_85J3_126_1427_U134 ( .A(u_alu_DP_OP_85J3_126_1427_n5), .B(
        u_alu_DP_OP_85J3_126_1427_n132), .Q(u_alu_pre_subb[11]) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U26 ( .A(u_alu_DP_OP_85J3_126_1427_n5), .B(
        u_alu_DP_OP_85J3_126_1427_n34), .Q(u_alu_pre_suba[11]) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U96 ( .A(u_alu_DP_OP_85J3_126_1427_n13), .B(
        u_alu_DP_OP_85J3_126_1427_n81), .Q(u_alu_pre_suba[3]) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U204 ( .A(u_alu_DP_OP_85J3_126_1427_n13), 
        .B(u_alu_DP_OP_85J3_126_1427_n179), .Q(u_alu_pre_subb[3]) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U192 ( .A(u_alu_DP_OP_85J3_126_1427_n12), 
        .B(u_alu_DP_OP_85J3_126_1427_n173), .Q(u_alu_pre_subb[4]) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U148 ( .A(u_alu_DP_OP_85J3_126_1427_n7), .B(
        u_alu_DP_OP_85J3_126_1427_n140), .Q(u_alu_pre_subb[9]) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U40 ( .A(u_alu_DP_OP_85J3_126_1427_n7), .B(
        u_alu_DP_OP_85J3_126_1427_n42), .Q(u_alu_pre_suba[9]) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U1 ( .A(u_alu_DP_OP_85J3_126_1427_n1), .B(
        u_alu_DP_OP_85J3_126_1427_n18), .Q(u_alu_pre_suba[15]) );
  NAND20 u_alu_DP_OP_85J3_126_1427_U5 ( .A(alu_i_data_B[31]), .B(n91), .Q(
        u_alu_DP_OP_85J3_126_1427_n17) );
  NAND20 u_alu_DP_OP_85J3_126_1427_U11 ( .A(n89), .B(compare_i_data_rs[30]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n20) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U12 ( .A(u_alu_DP_OP_85J3_126_1427_n3), .B(
        u_alu_DP_OP_85J3_126_1427_n26), .Q(u_alu_pre_suba[13]) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U54 ( .A(u_alu_DP_OP_85J3_126_1427_n9), .B(
        u_alu_DP_OP_85J3_126_1427_n50), .Q(u_alu_pre_suba[7]) );
  XNR21 u_alu_DP_OP_85J3_126_1427_U162 ( .A(u_alu_DP_OP_85J3_126_1427_n9), .B(
        u_alu_DP_OP_85J3_126_1427_n148), .Q(u_alu_pre_subb[7]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U7 ( .A(u_alu_pre_sum_3a[2]), .B(
        u_alu_DP_OP_83J3_124_3384_n7), .CO(u_alu_DP_OP_83J3_124_3384_n6), .S(
        u_alu_pre_sum_3b[2]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U2 ( .A(u_alu_pre_sum_3a[7]), .B(
        u_alu_DP_OP_83J3_124_3384_n2), .CO(u_alu_DP_OP_83J3_124_3384_n1), .S(
        u_alu_pre_sum_3b[7]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U8 ( .A(u_alu_pre_sum_3a[1]), .B(
        u_alu_pre_sum_3a[0]), .CO(u_alu_DP_OP_83J3_124_3384_n7), .S(
        u_alu_pre_sum_3b[1]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U16 ( .A(alu_i_data_B[17]), .B(
        compare_i_data_rs[17]), .CI(u_alu_DP_OP_83J3_124_3384_n15), .CO(
        u_alu_DP_OP_83J3_124_3384_n14), .S(u_alu_pre_sum_3a[1]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U11 ( .A(alu_i_data_B[22]), .B(
        compare_i_data_rs[22]), .CI(u_alu_DP_OP_83J3_124_3384_n10), .CO(
        u_alu_DP_OP_83J3_124_3384_n9), .S(u_alu_pre_sum_3a[6]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U10 ( .A(alu_i_data_B[23]), .B(
        compare_i_data_rs[23]), .CI(u_alu_DP_OP_83J3_124_3384_n9), .CO(
        u_alu_pre_sum_3a[8]), .S(u_alu_pre_sum_3a[7]) );
  NOR21 DP_OP_77_130_260_U32 ( .A(compare_i_data_rs[8]), .B(alu_i_data_B[8]), 
        .Q(DP_OP_77_130_260_n23) );
  AOI212 DP_OP_77_130_260_U27 ( .A(u_alu_sum_1_8_), .B(DP_OP_77_130_260_n30), 
        .C(DP_OP_77_130_260_n22), .Q(DP_OP_77_130_260_n20) );
  OAI212 DP_OP_77_130_260_U7 ( .A(DP_OP_77_130_260_n10), .B(n123), .C(
        DP_OP_77_130_260_n11), .Q(DP_OP_77_130_260_n9) );
  NAND22 DP_OP_77_130_260_U11 ( .A(alu_i_data_B[11]), .B(compare_i_data_rs[11]), .Q(DP_OP_77_130_260_n11) );
  NAND22 DP_OP_77_130_260_U19 ( .A(alu_i_data_B[10]), .B(compare_i_data_rs[10]), .Q(DP_OP_77_130_260_n16) );
  NOR21 DP_OP_77_130_260_U18 ( .A(compare_i_data_rs[10]), .B(alu_i_data_B[10]), 
        .Q(DP_OP_77_130_260_n15) );
  OAI212 DP_OP_77_130_260_U21 ( .A(DP_OP_77_130_260_n18), .B(
        DP_OP_77_130_260_n20), .C(DP_OP_77_130_260_n19), .Q(
        DP_OP_77_130_260_n17) );
  NAND22 DP_OP_77_130_260_U25 ( .A(alu_i_data_B[9]), .B(compare_i_data_rs[9]), 
        .Q(DP_OP_77_130_260_n19) );
  NAND22 DP_OP_77_130_260_U33 ( .A(alu_i_data_B[8]), .B(compare_i_data_rs[8]), 
        .Q(DP_OP_77_130_260_n24) );
  NOR21 DP_OP_77_130_260_U10 ( .A(compare_i_data_rs[11]), .B(alu_i_data_B[11]), 
        .Q(DP_OP_77_130_260_n10) );
  XNR21 DP_OP_77_130_260_U12 ( .A(DP_OP_77_130_260_n2), .B(
        DP_OP_77_130_260_n17), .Q(u_alu_N167) );
  NOR21 DP_OP_77_130_260_U24 ( .A(compare_i_data_rs[9]), .B(alu_i_data_B[9]), 
        .Q(DP_OP_77_130_260_n18) );
  NAND21 u_alu_sub_x_2_U30 ( .A(n96), .B(compare_i_data_rs[11]), .Q(
        u_alu_sub_x_2_n31) );
  OAI211 u_alu_sub_x_2_U46 ( .A(u_alu_sub_x_2_n48), .B(u_alu_sub_x_2_n44), .C(
        u_alu_sub_x_2_n45), .Q(u_alu_sub_x_2_n43) );
  NOR21 u_alu_DP_OP_85J3_126_1427_U32 ( .A(compare_i_data_rs[27]), .B(n93), 
        .Q(u_alu_DP_OP_85J3_126_1427_n32) );
  NAND22 u_alu_add_x_1_U45 ( .A(u_alu_add_x_1_n49), .B(u_alu_add_x_1_n37), .Q(
        u_alu_add_x_1_n6) );
  NOR21 u_alu_DP_OP_85J3_126_1427_U18 ( .A(compare_i_data_rs[29]), .B(n90), 
        .Q(u_alu_DP_OP_85J3_126_1427_n24) );
  NAND21 u_alu_DP_OP_85J3_126_1427_U19 ( .A(n90), .B(compare_i_data_rs[29]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n25) );
  NAND21 DP_OP_77_130_260_U16 ( .A(DP_OP_77_130_260_n28), .B(
        DP_OP_77_130_260_n16), .Q(DP_OP_77_130_260_n2) );
  NAND22 DP_OP_77_130_260_U30 ( .A(DP_OP_77_130_260_n30), .B(
        DP_OP_77_130_260_n24), .Q(DP_OP_77_130_260_n4) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U7 ( .A(u_alu_pre_sum_4a[1]), .B(
        u_alu_pre_sum_4a[0]), .CO(u_alu_DP_OP_84J3_125_2615_n6), .S(
        u_alu_pre_sum_4b[1]) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U15 ( .A(compare_i_data_rs[26]), .B(
        alu_i_data_B[26]), .CI(u_alu_DP_OP_84J3_125_2615_n14), .CO(
        u_alu_DP_OP_84J3_125_2615_n13), .S(u_alu_pre_sum_4a[2]) );
  NAND21 u_alu_add_x_1_U39 ( .A(u_alu_add_x_1_n48), .B(u_alu_add_x_1_n34), .Q(
        u_alu_add_x_1_n5) );
  NAND22 u_alu_add_x_1_U8 ( .A(u_alu_add_x_1_n44), .B(u_alu_add_x_1_n15), .Q(
        u_alu_add_x_1_n1) );
  NAND21 DP_OP_77_130_260_U8 ( .A(DP_OP_77_130_260_n27), .B(
        DP_OP_77_130_260_n11), .Q(DP_OP_77_130_260_n1) );
  NAND21 DP_OP_77_130_260_U22 ( .A(DP_OP_77_130_260_n29), .B(
        DP_OP_77_130_260_n19), .Q(DP_OP_77_130_260_n3) );
  NAND21 u_alu_sub_x_2_U13 ( .A(u_alu_sub_x_2_n85), .B(u_alu_sub_x_2_n23), .Q(
        u_alu_sub_x_2_n2) );
  NAND22 u_alu_sub_x_2_U37 ( .A(u_alu_sub_x_2_n88), .B(u_alu_sub_x_2_n38), .Q(
        u_alu_sub_x_2_n5) );
  NAND22 u_alu_sub_x_2_U27 ( .A(u_alu_sub_x_2_n87), .B(u_alu_sub_x_2_n31), .Q(
        u_alu_sub_x_2_n4) );
  NAND22 u_alu_sub_x_2_U53 ( .A(u_alu_sub_x_2_n90), .B(u_alu_sub_x_2_n48), .Q(
        u_alu_sub_x_2_n7) );
  OAI211 u_alu_sub_x_2_U63 ( .A(u_alu_sub_x_2_n59), .B(u_alu_sub_x_2_n55), .C(
        u_alu_sub_x_2_n56), .Q(u_alu_sub_x_2_n54) );
  OAI211 u_alu_sub_x_2_U26 ( .A(u_alu_sub_x_2_n30), .B(u_alu_sub_x_2_n34), .C(
        u_alu_sub_x_2_n31), .Q(u_alu_sub_x_2_n29) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U14 ( .A(compare_i_data_rs[27]), .B(
        alu_i_data_B[27]), .CI(u_alu_DP_OP_84J3_125_2615_n13), .CO(
        u_alu_DP_OP_84J3_125_2615_n12), .S(u_alu_pre_sum_4a[3]) );
  AOI211 u_alu_sub_x_2_U92 ( .A(u_alu_sub_x_2_n80), .B(u_alu_sub_x_2_n72), .C(
        u_alu_sub_x_2_n73), .Q(u_alu_sub_x_2_n71) );
  OAI211 u_alu_DP_OP_85J3_126_1427_U214 ( .A(n189), .B(
        u_alu_DP_OP_85J3_126_1427_n186), .C(u_alu_DP_OP_85J3_126_1427_n83), 
        .Q(u_alu_DP_OP_85J3_126_1427_n179) );
  OAI211 u_alu_DP_OP_85J3_126_1427_U106 ( .A(n189), .B(
        u_alu_DP_OP_85J3_126_1427_n88), .C(u_alu_DP_OP_85J3_126_1427_n83), .Q(
        u_alu_DP_OP_85J3_126_1427_n81) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U13 ( .A(compare_i_data_rs[28]), .B(
        alu_i_data_B[28]), .CI(u_alu_DP_OP_84J3_125_2615_n12), .CO(
        u_alu_DP_OP_84J3_125_2615_n11), .S(u_alu_pre_sum_4a[4]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U6 ( .A(u_alu_pre_sum_3a[3]), .B(
        u_alu_DP_OP_83J3_124_3384_n6), .CO(u_alu_DP_OP_83J3_124_3384_n5), .S(
        u_alu_pre_sum_3b[3]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U3 ( .A(u_alu_pre_sum_4a[5]), .B(
        u_alu_DP_OP_84J3_125_2615_n3), .CO(u_alu_DP_OP_84J3_125_2615_n2), .S(
        u_alu_pre_sum_4b[5]) );
  AOI211 u_alu_sub_x_2_U24 ( .A(u_alu_sub_x_2_n50), .B(u_alu_sub_x_2_n28), .C(
        u_alu_sub_x_2_n29), .Q(u_alu_sub_x_2_n27) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U11 ( .A(compare_i_data_rs[30]), .B(
        alu_i_data_B[30]), .CI(u_alu_DP_OP_84J3_125_2615_n10), .CO(
        u_alu_DP_OP_84J3_125_2615_n9), .S(u_alu_pre_sum_4a[6]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U2 ( .A(u_alu_pre_sum_4a[6]), .B(
        u_alu_DP_OP_84J3_125_2615_n2), .CO(u_alu_DP_OP_84J3_125_2615_n1), .S(
        u_alu_pre_sum_4b[6]) );
  OAI211 u_alu_sub_x_2_U69 ( .A(u_alu_sub_x_2_n58), .B(u_alu_sub_x_2_n60), .C(
        u_alu_sub_x_2_n59), .Q(u_alu_sub_x_2_n57) );
  OAI212 u_alu_sub_x_2_U52 ( .A(u_alu_sub_x_2_n47), .B(u_alu_sub_x_2_n49), .C(
        u_alu_sub_x_2_n48), .Q(u_alu_sub_x_2_n46) );
  OAI211 u_alu_sub_x_2_U32 ( .A(u_alu_sub_x_2_n33), .B(u_alu_sub_x_2_n49), .C(
        u_alu_sub_x_2_n34), .Q(u_alu_sub_x_2_n32) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U5 ( .A(u_alu_pre_sum_3a[4]), .B(
        u_alu_DP_OP_83J3_124_3384_n5), .CO(u_alu_DP_OP_83J3_124_3384_n4), .S(
        u_alu_pre_sum_3b[4]) );
  AOI211 u_alu_sub_x_2_U10 ( .A(u_alu_sub_x_2_n24), .B(u_alu_sub_x_2_n85), .C(
        u_alu_sub_x_2_n21), .Q(u_alu_sub_x_2_n19) );
  ADD32 u_alu_sub_x_2_U2 ( .A(n86), .B(n80), .CI(u_alu_sub_x_2_n16), .CO(
        u_alu_sub_x_2_n15), .S(u_alu_half_sub_15_) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U126 ( .A(n89), .B(compare_i_data_rs[30]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n123), .CO(
        u_alu_DP_OP_85J3_126_1427_n122), .S(u_alu_pre_subb[14]) );
  NAND22 u_alu_add_x_1_U52 ( .A(u_alu_add_x_1_n50), .B(u_alu_add_x_1_n41), .Q(
        u_alu_add_x_1_n7) );
  NAND22 u_alu_add_x_1_U30 ( .A(u_alu_add_x_1_n47), .B(u_alu_add_x_1_n28), .Q(
        u_alu_add_x_1_n4) );
  NAND22 u_alu_sub_x_2_U67 ( .A(n233), .B(compare_i_data_rs[7]), .Q(
        u_alu_sub_x_2_n56) );
  NAND21 u_alu_add_x_1_U57 ( .A(u_alu_add_x_1_n51), .B(u_alu_add_x_1_n43), .Q(
        u_alu_add_x_1_n8) );
  NAND21 u_alu_add_x_1_U22 ( .A(u_alu_add_x_1_n46), .B(u_alu_add_x_1_n23), .Q(
        u_alu_add_x_1_n3) );
  NAND21 u_alu_sub_x_2_U86 ( .A(u_alu_sub_x_2_n94), .B(u_alu_sub_x_2_n69), .Q(
        u_alu_sub_x_2_n11) );
  NAND22 u_alu_add_x_1_U14 ( .A(u_alu_add_x_1_n45), .B(u_alu_add_x_1_n18), .Q(
        u_alu_add_x_1_n2) );
  OAI210 u_alu_sub_x_2_U100 ( .A(n155), .B(u_alu_sub_x_2_n79), .C(
        u_alu_sub_x_2_n78), .Q(u_alu_sub_x_2_n76) );
  OAI211 u_alu_sub_x_2_U94 ( .A(u_alu_sub_x_2_n78), .B(u_alu_sub_x_2_n74), .C(
        u_alu_sub_x_2_n75), .Q(u_alu_sub_x_2_n73) );
  NAND22 u_alu_sub_x_2_U64 ( .A(u_alu_sub_x_2_n91), .B(u_alu_sub_x_2_n56), .Q(
        u_alu_sub_x_2_n8) );
  NOR21 u_alu_add_x_1_U24 ( .A(compare_i_data_rs[5]), .B(alu_i_data_B[5]), .Q(
        u_alu_add_x_1_n22) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U16 ( .A(compare_i_data_rs[25]), .B(
        alu_i_data_B[25]), .CI(u_alu_DP_OP_84J3_125_2615_n15), .CO(
        u_alu_DP_OP_84J3_125_2615_n14), .S(u_alu_pre_sum_4a[1]) );
  NAND22 u_alu_DP_OP_85J3_126_1427_U104 ( .A(n105), .B(compare_i_data_rs[19]), 
        .Q(u_alu_DP_OP_85J3_126_1427_n80) );
  NAND20 u_alu_sub_x_2_U5 ( .A(u_alu_sub_x_2_n84), .B(u_alu_sub_x_2_n18), .Q(
        u_alu_sub_x_2_n1) );
  NAND21 u_alu_sub_x_2_U95 ( .A(u_alu_sub_x_2_n95), .B(u_alu_sub_x_2_n75), .Q(
        u_alu_sub_x_2_n12) );
  DFC3 pipe_con_Malupc8_reg ( .D(i_con_Malupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Malupc8) );
  NAND22 U3 ( .A(u_alu_DP_OP_83J3_124_3384_n11), .B(compare_i_data_rs[21]), 
        .Q(n129) );
  XOR21 U4 ( .A(u_alu_DP_OP_83J3_124_3384_n13), .B(n135), .Q(
        u_alu_pre_sum_3a[3]) );
  INV3 U5 ( .A(n82), .Q(n83) );
  NAND41 U6 ( .A(n944), .B(n943), .C(n942), .D(n941), .Q(n945) );
  INV3 U7 ( .A(i_con_Efamux[2]), .Q(n531) );
  NAND23 U8 ( .A(n873), .B(n872), .Q(compare_i_data_rs[17]) );
  INV3 U9 ( .A(alu_i_data_B[18]), .Q(n84) );
  NAND24 U10 ( .A(n611), .B(n624), .Q(alu_i_data_B[19]) );
  MUX22 U11 ( .A(compare_i_data_rt[8]), .B(i_data_immext[8]), .S(n235), .Q(
        alu_i_data_B[8]) );
  INV3 U12 ( .A(alu_i_data_B[26]), .Q(n85) );
  MUX22 U13 ( .A(compare_i_data_rt[11]), .B(i_data_immext[11]), .S(n235), .Q(
        alu_i_data_B[11]) );
  INV3 U14 ( .A(n235), .Q(n623) );
  NOR21 U15 ( .A(compare_i_data_rs[2]), .B(u_alu_lt_x_11_B_2_), .Q(
        u_alu_add_x_1_n36) );
  INV3 U16 ( .A(n221), .Q(n112) );
  NAND23 U17 ( .A(n736), .B(n735), .Q(compare_i_data_rs[7]) );
  INV3 U18 ( .A(alu_i_data_B[16]), .Q(n87) );
  AOI2111 U19 ( .A(n121), .B(i_data_FEalures[16]), .C(n905), .D(n904), .Q(n907) );
  NAND22 U20 ( .A(u_alu_DP_OP_83J3_124_3384_n12), .B(compare_i_data_rs[20]), 
        .Q(n126) );
  NAND22 U21 ( .A(n818), .B(n817), .Q(compare_i_data_rs[26]) );
  INV3 U22 ( .A(n1263), .Q(n1247) );
  NAND23 U23 ( .A(n791), .B(n790), .Q(compare_i_data_rs[30]) );
  INV12 U24 ( .A(n522), .Q(n521) );
  NAND33 U25 ( .A(n537), .B(n536), .C(n535), .Q(compare_i_data_rs[5]) );
  NOR22 U26 ( .A(n545), .B(n1069), .Q(n1264) );
  NOR21 U27 ( .A(n1069), .B(n771), .Q(n1263) );
  NOR22 U28 ( .A(n764), .B(n763), .Q(n1250) );
  AOI211 U29 ( .A(n1169), .B(u_alu_pre_sum_3a[3]), .C(n1115), .Q(n1116) );
  INV3 U30 ( .A(n222), .Q(n1171) );
  INV12 U31 ( .A(n525), .Q(n121) );
  INV3 U32 ( .A(i_con_Efbmux[1]), .Q(n554) );
  BUF8 U33 ( .A(n900), .Q(n122) );
  NAND22 U34 ( .A(n230), .B(i_data_rt[16]), .Q(n622) );
  NAND22 U35 ( .A(n230), .B(i_data_rt[21]), .Q(n602) );
  NAND31 U36 ( .A(n1226), .B(n1225), .C(n1224), .Q(alu_o_data_AluRes[29]) );
  NOR23 U37 ( .A(n554), .B(n547), .Q(n670) );
  CLKIN0 U38 ( .A(compare_i_data_rs[27]), .Q(n1) );
  CLKIN0 U39 ( .A(alu_i_data_B[27]), .Q(n2) );
  IMAJ30 U40 ( .A(n1), .B(n1264), .C(n2), .Q(n3) );
  AOI310 U41 ( .A(n1247), .B(n1), .C(n2), .D(n3), .Q(n1198) );
  OAI2110 U42 ( .A(n86), .B(n1062), .C(n1061), .D(n1060), .Q(n4) );
  AOI210 U43 ( .A(u_alu_N172), .B(n1159), .C(n4), .Q(n5) );
  CLKIN0 U44 ( .A(i_data_immext[10]), .Q(n6) );
  NAND30 U45 ( .A(n1250), .B(n355), .C(n6), .Q(n7) );
  NAND20 U46 ( .A(u_alu_half_sub_15_), .B(n1064), .Q(n8) );
  NAND30 U47 ( .A(n8), .B(n7), .C(n5), .Q(alu_o_data_AluRes[15]) );
  INV3 U48 ( .A(n1068), .Q(n9) );
  NOR21 U49 ( .A(n1069), .B(n9), .Q(n1242) );
  IMAJ30 U50 ( .A(compare_i_data_rs[29]), .B(n138), .C(n90), .Q(n10) );
  MAJ31 U51 ( .A(n91), .B(alu_i_data_B[31]), .C(n145), .Q(n11) );
  AOI210 U52 ( .A(n146), .B(n10), .C(n11), .Q(n12) );
  NOR40 U53 ( .A(n186), .B(n193), .C(n185), .D(n184), .Q(n13) );
  OAI2110 U54 ( .A(n199), .B(n198), .C(n197), .D(n196), .Q(n14) );
  NOR40 U55 ( .A(n201), .B(n203), .C(n202), .D(n220), .Q(n15) );
  OAI210 U56 ( .A(n13), .B(n14), .C(n15), .Q(n16) );
  OAI2110 U57 ( .A(n201), .B(n144), .C(n12), .D(n16), .Q(u_alu_N306) );
  AOI210 U58 ( .A(n1058), .B(alu_i_data_B[14]), .C(n1057), .Q(n17) );
  AOI220 U59 ( .A(n1250), .B(u_alu_N207), .C(u_alu_N171), .D(n1159), .Q(n18)
         );
  CLKIN0 U60 ( .A(u_alu_sub_x_2_n19), .Q(n19) );
  IMUX20 U61 ( .A(n19), .B(u_alu_sub_x_2_n19), .S(u_alu_sub_x_2_n1), .Q(n20)
         );
  IMUX20 U62 ( .A(n420), .B(n468), .S(n378), .Q(n21) );
  AOI220 U63 ( .A(n1064), .B(n20), .C(n1251), .D(n21), .Q(n22) );
  NAND30 U64 ( .A(n17), .B(n18), .C(n22), .Q(alu_o_data_AluRes[14]) );
  NOR20 U65 ( .A(n879), .B(n886), .Q(n23) );
  AOI310 U66 ( .A(n1308), .B(n878), .C(n23), .D(i_data_immext[4]), .Q(n1262)
         );
  NAND22 U67 ( .A(i_data_rs[21]), .B(n118), .Q(n24) );
  OAI222 U68 ( .A(n120), .B(n840), .C(n842), .D(n119), .Q(n25) );
  AOI210 U69 ( .A(n121), .B(i_data_FEalures[21]), .C(n25), .Q(n26) );
  NAND33 U70 ( .A(n24), .B(n26), .C(n841), .Q(compare_i_data_rs[21]) );
  CLKIN0 U71 ( .A(i_data_immext[10]), .Q(n27) );
  XNR20 U72 ( .A(compare_i_data_rs[29]), .B(alu_i_data_B[29]), .Q(n28) );
  OAI2110 U73 ( .A(n1266), .B(n28), .C(n1219), .D(n1218), .Q(n29) );
  AOI310 U74 ( .A(n1251), .B(n458), .C(n27), .D(n29), .Q(n1221) );
  NOR20 U75 ( .A(alu_i_data_B[12]), .B(n1247), .Q(n30) );
  OAI210 U76 ( .A(n1266), .B(alu_i_data_B[12]), .C(n526), .Q(n31) );
  IMUX20 U77 ( .A(n30), .B(n31), .S(compare_i_data_rs[12]), .Q(n1039) );
  NOR20 U78 ( .A(i_data_immext[10]), .B(n372), .Q(n32) );
  NAND20 U79 ( .A(n1250), .B(n32), .Q(n33) );
  NAND40 U80 ( .A(n1009), .B(n1007), .C(n1008), .D(n33), .Q(
        alu_o_data_AluRes[8]) );
  IMUX20 U81 ( .A(n1252), .B(n1258), .S(u_alu_pre_subb[0]), .Q(n34) );
  AOI210 U82 ( .A(n1169), .B(u_alu_pre_sum_3a[0]), .C(n1078), .Q(n35) );
  NAND20 U83 ( .A(n34), .B(n35), .Q(alu_o_data_AluRes[16]) );
  NAND22 U84 ( .A(i_data_rs[29]), .B(n118), .Q(n36) );
  OAI222 U85 ( .A(n120), .B(n795), .C(n797), .D(n119), .Q(n37) );
  AOI210 U86 ( .A(n121), .B(i_data_FEalures[29]), .C(n37), .Q(n38) );
  NAND33 U87 ( .A(n36), .B(n38), .C(n796), .Q(compare_i_data_rs[29]) );
  CLKIN0 U88 ( .A(u_alu_sub_x_2_n78), .Q(n39) );
  NOR20 U89 ( .A(n155), .B(n39), .Q(n40) );
  XNR20 U90 ( .A(u_alu_sub_x_2_n79), .B(n40), .Q(u_alu_half_sub_2_) );
  NOR20 U91 ( .A(alu_i_data_B[13]), .B(n1247), .Q(n41) );
  OAI210 U92 ( .A(n1266), .B(alu_i_data_B[13]), .C(n526), .Q(n42) );
  IMUX20 U93 ( .A(n41), .B(n42), .S(compare_i_data_rs[13]), .Q(n1047) );
  CLKIN0 U94 ( .A(u_alu_DP_OP_85J3_126_1427_n191), .Q(n43) );
  NOR20 U95 ( .A(u_alu_DP_OP_85J3_126_1427_n92), .B(n43), .Q(u_alu_pre_subb[0]) );
  NAND20 U96 ( .A(u_alu_pre_sum_3b[5]), .B(n1150), .Q(n44) );
  AOI220 U97 ( .A(n1250), .B(u_alu_N214), .C(n1251), .D(u_alu_N246), .Q(n45)
         );
  AOI2110 U98 ( .A(n98), .B(compare_i_data_rs[21]), .C(n1130), .D(n1129), .Q(
        n46) );
  NAND30 U99 ( .A(n44), .B(n45), .C(n46), .Q(n1131) );
  IMUX20 U100 ( .A(n319), .B(n318), .S(i_data_immext[10]), .Q(n47) );
  CLKIN0 U101 ( .A(n1250), .Q(n48) );
  OAI310 U102 ( .A(compare_i_data_rs[26]), .B(n1247), .C(alu_i_data_B[26]), 
        .D(n1191), .Q(n49) );
  AOI2110 U103 ( .A(compare_i_data_rs[26]), .B(n98), .C(n1192), .D(n49), .Q(
        n50) );
  NOR20 U104 ( .A(i_data_immext[10]), .B(n510), .Q(n51) );
  NAND20 U105 ( .A(n1251), .B(n51), .Q(n52) );
  OAI2110 U106 ( .A(n47), .B(n48), .C(n50), .D(n52), .Q(n1193) );
  IMUX20 U107 ( .A(n325), .B(n324), .S(i_data_immext[10]), .Q(n53) );
  CLKIN0 U108 ( .A(n1250), .Q(n54) );
  AOI210 U109 ( .A(n98), .B(compare_i_data_rs[27]), .C(n1198), .Q(n55) );
  OAI310 U110 ( .A(n1267), .B(n93), .C(n1292), .D(n1197), .Q(n56) );
  NOR20 U111 ( .A(n378), .B(n519), .Q(n57) );
  AOI210 U112 ( .A(n57), .B(n1251), .C(n56), .Q(n58) );
  OAI2110 U113 ( .A(n53), .B(n54), .C(n55), .D(n58), .Q(n1199) );
  XNR20 U114 ( .A(u_alu_DP_OP_85J3_126_1427_n12), .B(
        u_alu_DP_OP_85J3_126_1427_n75), .Q(n59) );
  AOI210 U115 ( .A(n59), .B(n1252), .C(n1124), .Q(n60) );
  AOI220 U116 ( .A(u_alu_pre_sum_3a[4]), .B(n1169), .C(u_alu_pre_subb[4]), .D(
        n1258), .Q(n61) );
  NAND20 U117 ( .A(n60), .B(n61), .Q(alu_o_data_AluRes[20]) );
  CLKIN0 U118 ( .A(u_alu_sub_x_2_n82), .Q(n62) );
  NOR20 U119 ( .A(u_alu_sub_x_2_n81), .B(n62), .Q(n63) );
  XNR20 U120 ( .A(u_alu_sub_x_2_n83), .B(n63), .Q(u_alu_half_sub_1_) );
  CLKIN0 U121 ( .A(u_alu_sub_x_2_n69), .Q(n64) );
  AOI210 U122 ( .A(u_alu_sub_x_2_n70), .B(u_alu_sub_x_2_n94), .C(n64), .Q(n65)
         );
  CLKIN0 U123 ( .A(u_alu_sub_x_2_n64), .Q(n66) );
  NOR20 U124 ( .A(u_alu_sub_x_2_n63), .B(n66), .Q(n67) );
  XNR20 U125 ( .A(n65), .B(n67), .Q(u_alu_half_sub_5_) );
  OAI210 U126 ( .A(n1266), .B(alu_i_data_B[15]), .C(n526), .Q(n68) );
  NOR20 U127 ( .A(alu_i_data_B[15]), .B(n1247), .Q(n69) );
  IMUX20 U128 ( .A(n69), .B(n68), .S(n80), .Q(n1060) );
  AOI220 U129 ( .A(n1250), .B(u_alu_N213), .C(n1251), .D(u_alu_N245), .Q(n70)
         );
  AOI2110 U130 ( .A(n98), .B(compare_i_data_rs[20]), .C(n1123), .D(n1122), .Q(
        n71) );
  NAND20 U131 ( .A(u_alu_pre_sum_3b[4]), .B(n1150), .Q(n72) );
  NAND30 U132 ( .A(n72), .B(n70), .C(n71), .Q(n1124) );
  XOR30 U133 ( .A(alu_i_data_B[31]), .B(n91), .C(
        u_alu_DP_OP_85J3_126_1427_n122), .Q(u_alu_pre_subb[15]) );
  CLKIN0 U134 ( .A(n378), .Q(n73) );
  NAND30 U135 ( .A(n1250), .B(n324), .C(n73), .Q(n74) );
  NAND40 U136 ( .A(n1037), .B(n1035), .C(n1036), .D(n74), .Q(
        alu_o_data_AluRes[11]) );
  CLKIN0 U137 ( .A(u_alu_DP_OP_85J3_126_1427_n11), .Q(n75) );
  IMUX20 U138 ( .A(n75), .B(u_alu_DP_OP_85J3_126_1427_n11), .S(
        u_alu_DP_OP_85J3_126_1427_n66), .Q(n76) );
  AOI220 U139 ( .A(n1252), .B(n76), .C(n1258), .D(u_alu_pre_subb[5]), .Q(n77)
         );
  AOI210 U140 ( .A(u_alu_pre_sum_3a[5]), .B(n1169), .C(n1131), .Q(n78) );
  NAND20 U141 ( .A(n77), .B(n78), .Q(alu_o_data_AluRes[21]) );
  CLKIN4 U142 ( .A(n1170), .Q(n1150) );
  NAND22 U143 ( .A(n230), .B(i_data_rt[5]), .Q(n557) );
  NAND23 U144 ( .A(n225), .B(u_alu_pre_sum_3b[8]), .Q(n224) );
  NAND24 U145 ( .A(n859), .B(n858), .Q(compare_i_data_rs[19]) );
  AOI2110 U146 ( .A(n121), .B(i_data_FEalures[19]), .C(n857), .D(n856), .Q(
        n858) );
  NAND23 U147 ( .A(n235), .B(i_data_immext[16]), .Q(n624) );
  MUX26 U148 ( .A(compare_i_data_rt[5]), .B(i_data_immext[5]), .S(n235), .Q(
        alu_i_data_B[5]) );
  INV3 U149 ( .A(alu_i_data_B[17]), .Q(n108) );
  NAND23 U150 ( .A(n599), .B(n624), .Q(alu_i_data_B[22]) );
  NAND33 U151 ( .A(n602), .B(n601), .C(n600), .Q(compare_i_data_rt[21]) );
  NOR22 U152 ( .A(compare_i_data_rs[19]), .B(n105), .Q(
        u_alu_DP_OP_85J3_126_1427_n79) );
  NOR22 U153 ( .A(n189), .B(u_alu_DP_OP_85J3_126_1427_n79), .Q(
        u_alu_DP_OP_85J3_126_1427_n175) );
  NOR22 U154 ( .A(compare_i_data_rs[18]), .B(n84), .Q(n189) );
  NAND33 U155 ( .A(n618), .B(n617), .C(n616), .Q(compare_i_data_rt[17]) );
  NAND33 U156 ( .A(n622), .B(n621), .C(n620), .Q(compare_i_data_rt[16]) );
  AOI212 U157 ( .A(DP_OP_77_130_260_n17), .B(DP_OP_77_130_260_n28), .C(
        DP_OP_77_130_260_n14), .Q(n123) );
  NOR22 U158 ( .A(compare_i_data_rs[1]), .B(alu_i_data_B[1]), .Q(
        u_alu_add_x_1_n40) );
  BUF6 U159 ( .A(compare_i_data_rs[15]), .Q(n80) );
  OAI210 U160 ( .A(n119), .B(n1330), .C(n680), .Q(compare_i_data_rs[15]) );
  AOI2112 U161 ( .A(n1251), .B(u_alu_N249), .C(n1172), .D(n1171), .Q(n1173) );
  NAND24 U162 ( .A(n118), .B(i_data_rs[5]), .Q(n537) );
  NAND24 U163 ( .A(n543), .B(n542), .Q(n1267) );
  NOR20 U164 ( .A(n544), .B(alu_i_con_AluCtrl[2]), .Q(n542) );
  AOI221 U165 ( .A(n231), .B(i_data_FMmemout[1]), .C(n672), .D(
        i_data_FWmemout[1]), .Q(n667) );
  MUX26 U166 ( .A(compare_i_data_rt[4]), .B(i_data_immext[4]), .S(n235), .Q(
        alu_i_data_B[4]) );
  NAND33 U167 ( .A(n660), .B(n659), .C(n658), .Q(compare_i_data_rt[4]) );
  AOI221 U168 ( .A(n671), .B(i_data_FMalures[2]), .C(n521), .D(
        i_data_FEalures[2]), .Q(n665) );
  AOI2110 U169 ( .A(n121), .B(i_data_FEalures[30]), .C(n789), .D(n788), .Q(
        n790) );
  AOI221 U170 ( .A(n231), .B(i_data_FMmemout[5]), .C(n672), .D(
        i_data_FWmemout[5]), .Q(n555) );
  MUX26 U171 ( .A(compare_i_data_rt[3]), .B(i_data_immext[3]), .S(n235), .Q(
        alu_i_data_B[3]) );
  NAND33 U172 ( .A(n663), .B(n662), .C(n661), .Q(compare_i_data_rt[3]) );
  XOR20 U173 ( .A(compare_i_data_rs[19]), .B(alu_i_data_B[19]), .Q(n135) );
  NAND23 U174 ( .A(u_alu_DP_OP_83J3_124_3384_n13), .B(alu_i_data_B[19]), .Q(
        n133) );
  NAND33 U175 ( .A(n666), .B(n665), .C(n664), .Q(compare_i_data_rt[2]) );
  CLKBU15 U176 ( .A(alu_i_data_B[0]), .Q(n81) );
  NOR22 U177 ( .A(compare_i_data_rs[6]), .B(n112), .Q(u_alu_add_x_1_n17) );
  NAND24 U178 ( .A(n743), .B(n742), .Q(compare_i_data_rs[6]) );
  XOR20 U179 ( .A(alu_i_data_B[21]), .B(compare_i_data_rs[21]), .Q(n131) );
  NAND24 U180 ( .A(n603), .B(n624), .Q(alu_i_data_B[21]) );
  INV3 U181 ( .A(alu_i_data_B[20]), .Q(n82) );
  IMUX23 U182 ( .A(compare_i_data_rt[6]), .B(i_data_immext[6]), .S(n235), .Q(
        n221) );
  NAND33 U183 ( .A(n657), .B(n656), .C(n655), .Q(compare_i_data_rt[6]) );
  NAND34 U184 ( .A(n134), .B(n133), .C(n132), .Q(u_alu_DP_OP_83J3_124_3384_n12) );
  NAND21 U185 ( .A(u_alu_N206), .B(n1250), .Q(n1053) );
  NAND21 U186 ( .A(u_alu_N203), .B(n1250), .Q(n1025) );
  NAND21 U187 ( .A(u_alu_N200), .B(n1250), .Q(n999) );
  NAND21 U188 ( .A(u_alu_N202), .B(n1250), .Q(n1019) );
  NAND21 U189 ( .A(u_alu_N205), .B(n1250), .Q(n1045) );
  NAND20 U190 ( .A(u_alu_N216), .B(n1250), .Q(n1153) );
  NAND20 U191 ( .A(u_alu_N242), .B(n1251), .Q(n1086) );
  NAND20 U192 ( .A(u_alu_N243), .B(n1251), .Q(n1100) );
  NAND20 U193 ( .A(u_alu_N215), .B(n1250), .Q(n1139) );
  NAND21 U194 ( .A(u_alu_N199), .B(n1250), .Q(n989) );
  NAND20 U195 ( .A(u_alu_N244), .B(n1251), .Q(n1113) );
  NOR21 U196 ( .A(n378), .B(n516), .Q(u_alu_N246) );
  CLKIN3 U197 ( .A(n361), .Q(n371) );
  INV2 U198 ( .A(u_alu_sub_x_2_n71), .Q(u_alu_sub_x_2_n70) );
  INV2 U199 ( .A(n347), .Q(n377) );
  CLKIN3 U200 ( .A(n360), .Q(n370) );
  IMUX21 U201 ( .A(n490), .B(n449), .S(u_alu_ashr_4_SH_3_), .Q(n420) );
  IMUX20 U202 ( .A(n1263), .B(n1264), .S(u_alu_lt_x_11_B_2_), .Q(n1285) );
  IMUX20 U203 ( .A(n1263), .B(n1264), .S(alu_i_data_B[4]), .Q(n1273) );
  IMUX20 U204 ( .A(n1263), .B(n1264), .S(alu_i_data_B[1]), .Q(n1299) );
  IMUX20 U205 ( .A(n1263), .B(n1264), .S(alu_i_data_B[3]), .Q(n1278) );
  IMUX20 U206 ( .A(n1263), .B(n1264), .S(alu_i_data_B[5]), .Q(n1268) );
  CLKIN3 U207 ( .A(u_alu_add_x_1_n39), .Q(u_alu_add_x_1_n38) );
  INV3 U208 ( .A(u_alu_sub_x_2_n38), .Q(u_alu_sub_x_2_n36) );
  NOR20 U209 ( .A(alu_i_data_B[31]), .B(n91), .Q(n137) );
  IMUX20 U210 ( .A(n300), .B(n290), .S(u_alu_ashr_4_SH_1_), .Q(n315) );
  IMUX21 U211 ( .A(n389), .B(n392), .S(u_alu_ashr_4_SH_1_), .Q(n400) );
  NAND21 U212 ( .A(n95), .B(n1003), .Q(n1002) );
  INV1 U213 ( .A(u_alu_DP_OP_85J3_126_1427_n27), .Q(
        u_alu_DP_OP_85J3_126_1427_n192) );
  INV3 U214 ( .A(alu_i_data_B[15]), .Q(n86) );
  INV3 U215 ( .A(alu_i_data_B[29]), .Q(n90) );
  INV3 U216 ( .A(compare_i_data_rs[31]), .Q(n91) );
  NAND21 U217 ( .A(alu_i_data_B[21]), .B(compare_i_data_rs[21]), .Q(n128) );
  INV1 U218 ( .A(u_alu_add_x_1_n33), .Q(u_alu_add_x_1_n48) );
  INV3 U219 ( .A(alu_i_data_B[27]), .Q(n93) );
  INV3 U220 ( .A(alu_i_data_B[8]), .Q(n95) );
  INV3 U221 ( .A(alu_i_data_B[12]), .Q(n94) );
  NAND21 U222 ( .A(compare_i_data_rt[24]), .B(n623), .Q(n591) );
  MUX22 U223 ( .A(compare_i_data_rt[9]), .B(u_alu_ashr_4_SH_3_), .S(n235), .Q(
        alu_i_data_B[9]) );
  INV3 U224 ( .A(alu_i_data_B[11]), .Q(n96) );
  OAI211 U225 ( .A(n704), .B(n119), .C(n703), .Q(n705) );
  OAI211 U226 ( .A(n725), .B(n119), .C(n724), .Q(n726) );
  OAI211 U227 ( .A(n119), .B(n807), .C(n806), .Q(n808) );
  OAI212 U228 ( .A(n683), .B(n119), .C(n682), .Q(n684) );
  INV12 U229 ( .A(n524), .Q(n119) );
  INV2 U230 ( .A(n885), .Q(n887) );
  NAND21 U231 ( .A(n122), .B(i_data_FMmemout[8]), .Q(n724) );
  NAND21 U232 ( .A(n122), .B(i_data_FMmemout[11]), .Q(n703) );
  NAND22 U233 ( .A(n227), .B(n531), .Q(n528) );
  INV1 U234 ( .A(i_data_FMalures[14]), .Q(n681) );
  INV3 U235 ( .A(i_data_FEalures[31]), .Q(n780) );
  NAND21 U236 ( .A(i_con_bop[1]), .B(i_con_bop[2]), .Q(n955) );
  INV3 U237 ( .A(n1065), .Q(n1258) );
  INV3 U238 ( .A(u_alu_sub_x_2_n15), .Q(u_alu_half_sub_16_) );
  IMUX21 U239 ( .A(n97), .B(u_alu_pre_sum_4a[7]), .S(
        u_alu_DP_OP_84J3_125_2615_n1), .Q(u_alu_pre_sum_4b[7]) );
  NAND20 U240 ( .A(u_alu_N196), .B(n1250), .Q(n777) );
  NAND20 U241 ( .A(u_alu_N198), .B(n1250), .Q(n770) );
  NOR20 U242 ( .A(i_data_immext[10]), .B(n377), .Q(u_alu_N207) );
  AOI211 U243 ( .A(n971), .B(compare_i_data_rs[0]), .C(n970), .Q(n972) );
  INV3 U244 ( .A(n331), .Q(n375) );
  OAI211 U245 ( .A(n98), .B(n1302), .C(compare_i_data_rs[1]), .Q(n1301) );
  NAND20 U246 ( .A(u_alu_N197), .B(n1250), .Q(n774) );
  INV3 U247 ( .A(n338), .Q(n376) );
  OAI211 U248 ( .A(n98), .B(n1271), .C(compare_i_data_rs[5]), .Q(n1270) );
  NAND20 U249 ( .A(u_alu_N194), .B(n1250), .Q(n852) );
  OAI211 U250 ( .A(n98), .B(n1288), .C(compare_i_data_rs[2]), .Q(n1287) );
  NAND20 U251 ( .A(u_alu_N195), .B(n1250), .Q(n794) );
  OAI211 U252 ( .A(n98), .B(n1276), .C(compare_i_data_rs[4]), .Q(n1275) );
  OAI211 U253 ( .A(n98), .B(n1281), .C(compare_i_data_rs[3]), .Q(n1280) );
  MUX22 U254 ( .A(n503), .B(n502), .S(n378), .Q(u_alu_N233) );
  INV6 U255 ( .A(n526), .Q(n98) );
  OAI310 U256 ( .A(n108), .B(n1306), .C(n1267), .D(n1079), .Q(n1083) );
  OAI310 U257 ( .A(n84), .B(n1305), .C(n1267), .D(n1092), .Q(n1097) );
  OAI310 U258 ( .A(n109), .B(n1295), .C(n1267), .D(n1145), .Q(n1149) );
  IMUX21 U259 ( .A(n479), .B(n444), .S(u_alu_ashr_4_SH_3_), .Q(n404) );
  INV1 U260 ( .A(n191), .Q(n213) );
  CLKIN6 U261 ( .A(n1265), .Q(n526) );
  IMUX21 U262 ( .A(n421), .B(n424), .S(i_data_immext[8]), .Q(n434) );
  IMUX21 U263 ( .A(n247), .B(n246), .S(n381), .Q(n265) );
  MUX22 U264 ( .A(n403), .B(n402), .S(i_data_immext[8]), .Q(n444) );
  INV2 U265 ( .A(u_alu_DP_OP_85J3_126_1427_n25), .Q(
        u_alu_DP_OP_85J3_126_1427_n23) );
  IMUX21 U266 ( .A(n245), .B(n244), .S(n381), .Q(n266) );
  INV0 U267 ( .A(u_alu_sub_x_2_n17), .Q(u_alu_sub_x_2_n84) );
  XNR20 U268 ( .A(n1228), .B(alu_i_data_B[30]), .Q(n1229) );
  NAND21 U269 ( .A(alu_i_con_AluCtrl[2]), .B(n766), .Q(n767) );
  INV3 U270 ( .A(alu_i_data_B[19]), .Q(n105) );
  NAND21 U271 ( .A(compare_i_data_rs[19]), .B(alu_i_data_B[19]), .Q(n132) );
  NAND22 U272 ( .A(n962), .B(alu_i_con_AluCtrl[0]), .Q(n764) );
  NAND22 U273 ( .A(n715), .B(n714), .Q(compare_i_data_rs[10]) );
  INV3 U274 ( .A(alu_i_data_B[24]), .Q(n88) );
  INV3 U275 ( .A(alu_i_data_B[30]), .Q(n89) );
  INV6 U276 ( .A(alu_i_data_B[21]), .Q(n92) );
  NAND22 U277 ( .A(n722), .B(n721), .Q(compare_i_data_rs[9]) );
  NAND26 U278 ( .A(n615), .B(n624), .Q(alu_i_data_B[18]) );
  MUX22 U279 ( .A(compare_i_data_rt[10]), .B(i_data_immext[10]), .S(n235), .Q(
        alu_i_data_B[10]) );
  OAI211 U280 ( .A(n758), .B(n119), .C(n757), .Q(n759) );
  OAI211 U281 ( .A(n697), .B(n119), .C(n696), .Q(n698) );
  OAI211 U282 ( .A(n892), .B(n119), .C(n891), .Q(n893) );
  NAND31 U283 ( .A(n645), .B(n644), .C(n643), .Q(compare_i_data_rt[10]) );
  OAI211 U284 ( .A(n119), .B(n814), .C(n813), .Q(n815) );
  NAND32 U285 ( .A(n557), .B(n556), .C(n555), .Q(compare_i_data_rt[5]) );
  OAI211 U286 ( .A(n119), .B(n821), .C(n820), .Q(n822) );
  OAI211 U287 ( .A(n119), .B(n845), .C(n844), .Q(n846) );
  OAI211 U288 ( .A(n119), .B(n828), .C(n827), .Q(n829) );
  OAI211 U289 ( .A(n119), .B(n835), .C(n834), .Q(n836) );
  OAI211 U290 ( .A(n690), .B(n119), .C(n689), .Q(n691) );
  OAI211 U291 ( .A(n119), .B(n800), .C(n799), .Q(n801) );
  NAND31 U292 ( .A(n642), .B(n641), .C(n640), .Q(compare_i_data_rt[11]) );
  OAI211 U293 ( .A(n887), .B(n886), .C(n1325), .Q(n1323) );
  OAI221 U294 ( .A(n525), .B(n780), .C(n120), .D(n779), .Q(n781) );
  NAND22 U295 ( .A(n121), .B(i_data_FEalures[15]), .Q(n677) );
  BUF15 U296 ( .A(n228), .Q(n230) );
  INV3 U297 ( .A(n898), .Q(n523) );
  INV2 U298 ( .A(n528), .Q(n527) );
  AOI221 U299 ( .A(i_con_Ealuop[4]), .B(n1312), .C(i_con_Ealuop[5]), .D(n1309), 
        .Q(n1310) );
  INV1 U300 ( .A(i_data_FWmemout[0]), .Q(n758) );
  INV3 U301 ( .A(i_con_Efamux[0]), .Q(n227) );
  INV1 U302 ( .A(i_data_FMalures[31]), .Q(n779) );
  INV2 U303 ( .A(i_data_FWmemout[6]), .Q(n739) );
  INV2 U304 ( .A(i_data_FWmemout[9]), .Q(n718) );
  INV2 U305 ( .A(i_data_FWmemout[8]), .Q(n725) );
  INV2 U306 ( .A(i_data_FWmemout[7]), .Q(n732) );
  OAI2111 U307 ( .A(n1261), .B(n223), .C(n1174), .D(n1173), .Q(
        alu_o_data_AluRes[24]) );
  AOI211 U308 ( .A(n1252), .B(u_alu_pre_suba[13]), .C(n1223), .Q(n1225) );
  AOI211 U309 ( .A(n1169), .B(u_alu_pre_sum_3a[1]), .C(n1088), .Q(n1089) );
  NAND41 U310 ( .A(n1114), .B(n1113), .C(n1112), .D(n1111), .Q(n1115) );
  NAND41 U311 ( .A(n1087), .B(n1086), .C(n1085), .D(n1084), .Q(n1088) );
  NAND26 U312 ( .A(n226), .B(n224), .Q(n1241) );
  NAND41 U313 ( .A(n1140), .B(n1139), .C(n1138), .D(n1137), .Q(n1141) );
  NAND23 U314 ( .A(n1160), .B(n1159), .Q(n1261) );
  NAND42 U315 ( .A(n1256), .B(n1255), .C(n1254), .D(n1253), .Q(n1257) );
  AOI221 U316 ( .A(n1252), .B(u_alu_pre_suba[8]), .C(n1258), .D(
        u_alu_pre_subb[8]), .Q(n1174) );
  AOI221 U317 ( .A(n1252), .B(u_alu_pre_suba[10]), .C(n1258), .D(
        u_alu_pre_subb[10]), .Q(n1195) );
  AOI221 U318 ( .A(n1252), .B(u_alu_pre_suba[9]), .C(n1258), .D(
        u_alu_pre_subb[9]), .Q(n1186) );
  NAND23 U319 ( .A(n1169), .B(u_alu_pre_sum_3a[8]), .Q(n226) );
  OAI211 U320 ( .A(u_alu_pre_sum_3a[0]), .B(n1170), .C(n1077), .Q(n1078) );
  AOI221 U321 ( .A(n1252), .B(u_alu_pre_suba[11]), .C(n1258), .D(
        u_alu_pre_subb[11]), .Q(n1201) );
  NOR23 U322 ( .A(n1066), .B(u_alu_N173), .Q(n1169) );
  NAND23 U323 ( .A(u_alu_N173), .B(n1159), .Q(n1170) );
  NOR23 U324 ( .A(n1063), .B(u_alu_half_sub_16_), .Q(n1252) );
  OAI211 U325 ( .A(alu_i_data_B[31]), .B(n965), .C(n964), .Q(n967) );
  NAND21 U326 ( .A(u_alu_N170), .B(n1159), .Q(n1051) );
  INV2 U327 ( .A(u_alu_N306), .Q(n965) );
  NAND21 U328 ( .A(u_alu_N169), .B(n1159), .Q(n1043) );
  NAND21 U329 ( .A(u_alu_N168), .B(n1159), .Q(n1037) );
  NAND21 U330 ( .A(u_alu_half_sub_10_), .B(n1064), .Q(n1026) );
  AOI211 U331 ( .A(u_alu_DP_OP_85J3_126_1427_n34), .B(
        u_alu_DP_OP_85J3_126_1427_n193), .C(u_alu_DP_OP_85J3_126_1427_n129), 
        .Q(u_alu_DP_OP_85J3_126_1427_n29) );
  NAND31 U332 ( .A(n130), .B(n129), .C(n128), .Q(u_alu_DP_OP_83J3_124_3384_n10) );
  AOI211 U333 ( .A(u_alu_DP_OP_85J3_126_1427_n132), .B(
        u_alu_DP_OP_85J3_126_1427_n193), .C(u_alu_DP_OP_85J3_126_1427_n129), 
        .Q(u_alu_DP_OP_85J3_126_1427_n127) );
  XOR20 U334 ( .A(DP_OP_77_130_260_n1), .B(n123), .Q(u_alu_N168) );
  NAND21 U335 ( .A(u_alu_half_sub_8_), .B(n1064), .Q(n1007) );
  AOI211 U336 ( .A(u_alu_DP_OP_85J3_126_1427_n140), .B(
        u_alu_DP_OP_85J3_126_1427_n195), .C(u_alu_DP_OP_85J3_126_1427_n137), 
        .Q(u_alu_DP_OP_85J3_126_1427_n135) );
  INV3 U337 ( .A(u_alu_pre_sum_4a[7]), .Q(n97) );
  OAI311 U338 ( .A(n91), .B(n961), .C(n960), .D(n959), .Q(o_con_ifbranch) );
  NAND21 U339 ( .A(u_alu_N230), .B(n1251), .Q(n768) );
  NOR21 U340 ( .A(i_data_immext[10]), .B(n376), .Q(u_alu_N206) );
  NOR21 U341 ( .A(n958), .B(n957), .Q(n959) );
  NOR21 U342 ( .A(i_data_immext[10]), .B(n371), .Q(u_alu_N200) );
  NAND21 U343 ( .A(u_alu_N224), .B(n1250), .Q(n1255) );
  NAND21 U344 ( .A(u_alu_N222), .B(n1250), .Q(n1220) );
  NAND21 U345 ( .A(u_alu_N218), .B(n1250), .Q(n1181) );
  NAND21 U346 ( .A(u_alu_N210), .B(n1250), .Q(n1085) );
  NAND21 U347 ( .A(u_alu_N211), .B(n1250), .Q(n1099) );
  NAND21 U348 ( .A(u_alu_N233), .B(n1251), .Q(n1009) );
  NOR20 U349 ( .A(n378), .B(n514), .Q(u_alu_N250) );
  NAND21 U350 ( .A(u_alu_N226), .B(n1251), .Q(n850) );
  OAI311 U351 ( .A(alu_i_data_B[10]), .B(n1247), .C(compare_i_data_rs[10]), 
        .D(n1022), .Q(n1023) );
  NAND21 U352 ( .A(u_alu_N227), .B(n1251), .Q(n792) );
  OAI211 U353 ( .A(n1266), .B(compare_i_data_rs[10]), .C(n1020), .Q(n1024) );
  NAND21 U354 ( .A(u_alu_N247), .B(n1251), .Q(n1138) );
  INV2 U355 ( .A(u_alu_pre_sum_4a[5]), .Q(n1222) );
  NAND21 U356 ( .A(u_alu_N248), .B(n1251), .Q(n1152) );
  NAND21 U357 ( .A(u_alu_N212), .B(n1250), .Q(n1112) );
  NOR21 U358 ( .A(i_data_immext[10]), .B(n375), .Q(u_alu_N205) );
  NAND21 U359 ( .A(u_alu_N228), .B(n1251), .Q(n775) );
  OAI221 U360 ( .A(n1004), .B(n1003), .C(n1247), .D(n1002), .Q(n1005) );
  NAND21 U361 ( .A(u_alu_N236), .B(n1251), .Q(n1035) );
  INV2 U362 ( .A(n488), .Q(n516) );
  INV2 U363 ( .A(n440), .Q(n515) );
  INV2 U364 ( .A(n426), .Q(n513) );
  MUX22 U365 ( .A(n507), .B(n506), .S(i_data_immext[10]), .Q(u_alu_N234) );
  MUX22 U366 ( .A(n386), .B(n426), .S(n378), .Q(u_alu_N225) );
  INV2 U367 ( .A(u_alu_pre_sum_4a[4]), .Q(n1214) );
  NAND21 U368 ( .A(n1021), .B(compare_i_data_rs[10]), .Q(n1022) );
  INV2 U369 ( .A(n466), .Q(n509) );
  INV2 U370 ( .A(n477), .Q(n518) );
  AOI2111 U371 ( .A(n956), .B(n955), .C(i_con_bop[0]), .D(
        compare_i_data_rs[31]), .Q(n957) );
  IMUX21 U372 ( .A(n494), .B(n493), .S(n378), .Q(u_alu_N231) );
  INV1 U373 ( .A(n506), .Q(n514) );
  INV2 U374 ( .A(n359), .Q(n369) );
  AOI211 U375 ( .A(n992), .B(compare_i_data_rs[7]), .C(n991), .Q(n993) );
  IMUX21 U376 ( .A(n499), .B(n498), .S(i_data_immext[10]), .Q(u_alu_N232) );
  INV2 U377 ( .A(n502), .Q(n512) );
  IMUX21 U378 ( .A(n404), .B(n457), .S(i_data_immext[10]), .Q(u_alu_N237) );
  INV2 U379 ( .A(n357), .Q(n367) );
  NOR20 U380 ( .A(n378), .B(n498), .Q(u_alu_N248) );
  AOI211 U381 ( .A(n1012), .B(compare_i_data_rs[9]), .C(n1011), .Q(n1013) );
  IMUX21 U382 ( .A(n434), .B(n433), .S(u_alu_ashr_4_SH_3_), .Q(n477) );
  NOR20 U383 ( .A(n378), .B(n365), .Q(u_alu_N194) );
  IMUX21 U384 ( .A(n282), .B(n283), .S(u_alu_ashr_4_SH_3_), .Q(n331) );
  IMUX21 U385 ( .A(n444), .B(n443), .S(u_alu_ashr_4_SH_3_), .Q(n482) );
  IMUX21 U386 ( .A(n432), .B(n431), .S(u_alu_ashr_4_SH_3_), .Q(n466) );
  NOR20 U387 ( .A(n378), .B(n366), .Q(u_alu_N195) );
  IMUX21 U388 ( .A(n449), .B(n448), .S(u_alu_ashr_4_SH_3_), .Q(n493) );
  IMUX21 U389 ( .A(n452), .B(n451), .S(u_alu_ashr_4_SH_3_), .Q(n498) );
  NOR20 U390 ( .A(n378), .B(n368), .Q(u_alu_N197) );
  NOR31 U391 ( .A(u_alu_lt_x_11_B_7_), .B(compare_i_data_rs[7]), .C(n1247), 
        .Q(n991) );
  IMUX21 U392 ( .A(n312), .B(n311), .S(u_alu_ashr_4_SH_3_), .Q(n363) );
  INV1 U393 ( .A(u_alu_add_x_1_n30), .Q(u_alu_add_x_1_n29) );
  IMUX21 U394 ( .A(n297), .B(n298), .S(u_alu_ashr_4_SH_3_), .Q(n355) );
  INV2 U395 ( .A(n455), .Q(n510) );
  IMUX21 U396 ( .A(n271), .B(n272), .S(u_alu_ashr_4_SH_3_), .Q(n318) );
  INV2 U397 ( .A(u_alu_pre_sum_4a[3]), .Q(n1202) );
  INV2 U398 ( .A(n456), .Q(n519) );
  IMUX21 U399 ( .A(n500), .B(n453), .S(u_alu_ashr_4_SH_3_), .Q(n426) );
  IMUX21 U400 ( .A(n292), .B(n293), .S(u_alu_ashr_4_SH_3_), .Q(n347) );
  OAI211 U401 ( .A(n175), .B(n174), .C(n183), .Q(n176) );
  INV1 U402 ( .A(n193), .Q(n216) );
  IMUX21 U403 ( .A(n504), .B(n454), .S(u_alu_ashr_4_SH_3_), .Q(n440) );
  IMUX21 U404 ( .A(n287), .B(n288), .S(u_alu_ashr_4_SH_3_), .Q(n338) );
  OAI211 U405 ( .A(i_con_bop[1]), .B(i_con_bop[2]), .C(n954), .Q(n956) );
  AOI211 U406 ( .A(n954), .B(n952), .C(n951), .Q(n961) );
  IMUX21 U407 ( .A(n254), .B(n256), .S(i_data_immext[8]), .Q(n276) );
  IMUX21 U408 ( .A(n250), .B(n252), .S(i_data_immext[8]), .Q(n271) );
  NAND21 U409 ( .A(n1242), .B(alu_i_data_B[3]), .Q(n1106) );
  INV2 U410 ( .A(u_alu_add_x_1_n8), .Q(u_alu_sum_1_0_) );
  INV2 U411 ( .A(n279), .Q(n365) );
  NOR20 U412 ( .A(n378), .B(n469), .Q(u_alu_N256) );
  INV2 U413 ( .A(u_alu_sub_x_2_n55), .Q(u_alu_sub_x_2_n91) );
  IMUX21 U414 ( .A(n265), .B(n267), .S(i_data_immext[8]), .Q(n288) );
  IMUX21 U415 ( .A(n264), .B(n266), .S(i_data_immext[8]), .Q(n287) );
  IMUX21 U416 ( .A(n256), .B(n255), .S(i_data_immext[8]), .Q(n298) );
  INV2 U417 ( .A(u_alu_pre_sum_4a[2]), .Q(n1196) );
  IMUX21 U418 ( .A(n430), .B(n429), .S(i_data_immext[8]), .Q(n454) );
  IMUX21 U419 ( .A(n266), .B(n265), .S(i_data_immext[8]), .Q(n312) );
  NOR20 U420 ( .A(i_data_immext[8]), .B(n511), .Q(n443) );
  IMUX21 U421 ( .A(n258), .B(n260), .S(i_data_immext[8]), .Q(n282) );
  INV2 U422 ( .A(n340), .Q(n366) );
  INV1 U423 ( .A(n1242), .Q(n1176) );
  IMUX21 U424 ( .A(n505), .B(n504), .S(u_alu_ashr_4_SH_3_), .Q(n507) );
  INV3 U425 ( .A(n1066), .Q(n1159) );
  IMUX21 U426 ( .A(n260), .B(n259), .S(i_data_immext[8]), .Q(n305) );
  INV2 U427 ( .A(n358), .Q(n368) );
  IMUX21 U428 ( .A(n402), .B(n442), .S(i_data_immext[8]), .Q(n453) );
  INV3 U429 ( .A(n1063), .Q(n1064) );
  NOR20 U430 ( .A(i_data_immext[8]), .B(n517), .Q(n451) );
  IMUX21 U431 ( .A(n270), .B(n250), .S(i_data_immext[8]), .Q(n292) );
  MUX22 U432 ( .A(n419), .B(n418), .S(i_data_immext[8]), .Q(n449) );
  NOR20 U433 ( .A(i_data_immext[8]), .B(n508), .Q(n448) );
  OAI211 U434 ( .A(alu_i_data_B[16]), .B(n212), .C(n191), .Q(n185) );
  INV1 U435 ( .A(u_alu_sub_x_2_n74), .Q(u_alu_sub_x_2_n95) );
  NAND22 U436 ( .A(n950), .B(n949), .Q(n954) );
  IMUX20 U437 ( .A(n470), .B(n473), .S(u_alu_ashr_4_SH_1_), .Q(n485) );
  INV2 U438 ( .A(u_alu_DP_OP_85J3_126_1427_n90), .Q(
        u_alu_DP_OP_85J3_126_1427_n203) );
  IMUX21 U439 ( .A(n252), .B(n251), .S(i_data_immext[8]), .Q(n293) );
  IMUX21 U440 ( .A(n428), .B(n427), .S(i_data_immext[8]), .Q(n504) );
  INV2 U441 ( .A(n141), .Q(n219) );
  INV2 U442 ( .A(n447), .Q(n508) );
  NOR40 U443 ( .A(n928), .B(n927), .C(n926), .D(n925), .Q(n950) );
  INV2 U444 ( .A(u_alu_sub_x_2_n80), .Q(u_alu_sub_x_2_n79) );
  INV2 U445 ( .A(u_alu_sub_x_2_n42), .Q(u_alu_sub_x_2_n40) );
  INV2 U446 ( .A(n145), .Q(u_alu_DP_OP_85J3_126_1427_n94) );
  IMUX21 U447 ( .A(n423), .B(n450), .S(i_data_immext[8]), .Q(n433) );
  INV2 U448 ( .A(u_alu_DP_OP_85J3_126_1427_n64), .Q(
        u_alu_DP_OP_85J3_126_1427_n199) );
  INV2 U449 ( .A(u_alu_DP_OP_85J3_126_1427_n79), .Q(
        u_alu_DP_OP_85J3_126_1427_n201) );
  IMUX21 U450 ( .A(n418), .B(n447), .S(i_data_immext[8]), .Q(n431) );
  INV2 U451 ( .A(n450), .Q(n517) );
  INV2 U452 ( .A(n140), .Q(u_alu_DP_OP_85J3_126_1427_n196) );
  IMUX21 U453 ( .A(n275), .B(n254), .S(i_data_immext[8]), .Q(n297) );
  IMUX21 U454 ( .A(n393), .B(n396), .S(n381), .Q(n402) );
  INV2 U455 ( .A(u_alu_pre_sum_4a[1]), .Q(n1187) );
  IMUX21 U456 ( .A(n400), .B(n403), .S(i_data_immext[8]), .Q(n500) );
  INV2 U457 ( .A(n188), .Q(n214) );
  IMUX21 U458 ( .A(n484), .B(n438), .S(i_data_immext[8]), .Q(n505) );
  INV2 U459 ( .A(n189), .Q(u_alu_DP_OP_85J3_126_1427_n202) );
  INV1 U460 ( .A(n963), .Q(n763) );
  INV1 U461 ( .A(n198), .Q(n215) );
  INV2 U462 ( .A(u_alu_sub_x_2_n58), .Q(u_alu_sub_x_2_n92) );
  INV1 U463 ( .A(n442), .Q(n511) );
  IMUX21 U464 ( .A(n244), .B(n247), .S(u_alu_ashr_4_SH_1_), .Q(n256) );
  IMUX21 U465 ( .A(n238), .B(n237), .S(u_alu_ashr_4_SH_1_), .Q(n260) );
  INV2 U466 ( .A(n200), .Q(n220) );
  INV2 U467 ( .A(u_alu_DP_OP_85J3_126_1427_n56), .Q(
        u_alu_DP_OP_85J3_126_1427_n152) );
  INV1 U468 ( .A(n1069), .Q(n966) );
  IMUX20 U469 ( .A(n301), .B(n281), .S(i_data_immext[8]), .Q(n329) );
  IMUX21 U470 ( .A(n246), .B(n248), .S(n381), .Q(n255) );
  IMUX21 U471 ( .A(n480), .B(n401), .S(i_data_immext[8]), .Q(n501) );
  INV2 U472 ( .A(u_alu_sub_x_2_n43), .Q(u_alu_sub_x_2_n41) );
  IMUX21 U473 ( .A(n412), .B(n411), .S(u_alu_ashr_4_SH_1_), .Q(n430) );
  INV2 U474 ( .A(u_alu_DP_OP_85J3_126_1427_n16), .Q(
        u_alu_DP_OP_85J3_126_1427_n93) );
  NOR20 U475 ( .A(n378), .B(n364), .Q(u_alu_N193) );
  NOR40 U476 ( .A(n948), .B(n947), .C(n946), .D(n945), .Q(n949) );
  INV1 U477 ( .A(u_alu_sub_x_2_n47), .Q(u_alu_sub_x_2_n90) );
  IMUX21 U478 ( .A(n391), .B(n394), .S(u_alu_ashr_4_SH_1_), .Q(n403) );
  INV2 U479 ( .A(u_alu_sub_x_2_n44), .Q(u_alu_sub_x_2_n89) );
  INV2 U480 ( .A(n261), .Q(n364) );
  INV2 U481 ( .A(u_alu_add_x_1_n42), .Q(u_alu_add_x_1_n51) );
  IMUX21 U482 ( .A(n414), .B(n413), .S(n381), .Q(n429) );
  INV1 U483 ( .A(DP_OP_77_130_260_n10), .Q(DP_OP_77_130_260_n27) );
  INV1 U484 ( .A(DP_OP_77_130_260_n18), .Q(DP_OP_77_130_260_n29) );
  INV2 U485 ( .A(u_alu_add_x_1_n14), .Q(u_alu_add_x_1_n44) );
  NOR21 U486 ( .A(compare_i_data_rs[21]), .B(n92), .Q(
        u_alu_DP_OP_85J3_126_1427_n64) );
  INV1 U487 ( .A(u_alu_sub_x_2_n30), .Q(u_alu_sub_x_2_n87) );
  INV1 U488 ( .A(n161), .Q(u_alu_sub_x_2_n94) );
  IMUX21 U489 ( .A(n259), .B(n242), .S(i_data_immext[8]), .Q(n283) );
  XNR20 U490 ( .A(n1093), .B(alu_i_data_B[18]), .Q(n1094) );
  IMUX21 U491 ( .A(alu_i_data_B[8]), .B(u_alu_lt_x_11_B_7_), .S(
        i_data_immext[6]), .Q(n238) );
  IMUX21 U492 ( .A(n237), .B(n240), .S(n381), .Q(n252) );
  IMUX21 U493 ( .A(n263), .B(n253), .S(u_alu_ashr_4_SH_1_), .Q(n275) );
  XNR20 U494 ( .A(n1126), .B(alu_i_data_B[21]), .Q(n1127) );
  IMUX21 U495 ( .A(n396), .B(n395), .S(u_alu_ashr_4_SH_1_), .Q(n418) );
  IMUX21 U496 ( .A(alu_i_data_B[3]), .B(u_alu_lt_x_11_B_2_), .S(
        i_data_immext[6]), .Q(n246) );
  IMUX21 U497 ( .A(alu_i_data_B[5]), .B(alu_i_data_B[4]), .S(i_data_immext[6]), 
        .Q(n247) );
  NOR21 U498 ( .A(n766), .B(alu_i_con_AluCtrl[3]), .Q(n963) );
  NOR20 U499 ( .A(alu_i_data_B[25]), .B(n218), .Q(n202) );
  IMUX21 U500 ( .A(n249), .B(n236), .S(u_alu_ashr_4_SH_1_), .Q(n258) );
  INV1 U501 ( .A(u_alu_add_x_1_n22), .Q(u_alu_add_x_1_n46) );
  NOR20 U502 ( .A(n381), .B(n241), .Q(n242) );
  INV1 U503 ( .A(compare_i_data_rs[16]), .Q(n212) );
  INV1 U504 ( .A(u_alu_add_x_1_n36), .Q(u_alu_add_x_1_n49) );
  INV1 U505 ( .A(u_alu_add_x_1_n27), .Q(u_alu_add_x_1_n47) );
  INV2 U506 ( .A(u_alu_add_x_1_n28), .Q(u_alu_add_x_1_n26) );
  INV1 U507 ( .A(compare_i_data_rs[25]), .Q(n218) );
  INV2 U508 ( .A(alu_i_data_B[31]), .Q(n1244) );
  INV2 U509 ( .A(compare_i_data_rs[8]), .Q(n1003) );
  IMUX21 U510 ( .A(alu_i_data_B[30]), .B(alu_i_data_B[31]), .S(
        i_data_immext[6]), .Q(n397) );
  IMUX21 U511 ( .A(n240), .B(n239), .S(u_alu_ashr_4_SH_1_), .Q(n259) );
  XOR21 U512 ( .A(compare_i_data_rs[20]), .B(n83), .Q(n127) );
  INV1 U513 ( .A(u_alu_add_x_1_n40), .Q(u_alu_add_x_1_n50) );
  IMUX21 U514 ( .A(n243), .B(n245), .S(n381), .Q(n254) );
  NAND24 U515 ( .A(n908), .B(n907), .Q(compare_i_data_rs[16]) );
  INV3 U516 ( .A(alu_i_data_B[22]), .Q(n99) );
  INV1 U517 ( .A(compare_i_data_rs[22]), .Q(n100) );
  INV1 U518 ( .A(compare_i_data_rs[19]), .Q(n101) );
  NOR21 U519 ( .A(compare_i_data_rs[4]), .B(alu_i_data_B[4]), .Q(
        u_alu_add_x_1_n27) );
  INV2 U520 ( .A(compare_i_data_rs[11]), .Q(n102) );
  INV1 U521 ( .A(compare_i_data_rs[20]), .Q(n103) );
  IMUX21 U522 ( .A(alu_i_data_B[9]), .B(alu_i_data_B[8]), .S(i_data_immext[6]), 
        .Q(n245) );
  INV1 U523 ( .A(compare_i_data_rs[23]), .Q(n104) );
  IMUX21 U524 ( .A(alu_i_data_B[4]), .B(alu_i_data_B[3]), .S(i_data_immext[6]), 
        .Q(n240) );
  IMUX21 U525 ( .A(u_alu_lt_x_11_B_2_), .B(alu_i_data_B[1]), .S(
        i_data_immext[6]), .Q(n239) );
  INV1 U526 ( .A(compare_i_data_rs[28]), .Q(n106) );
  INV1 U527 ( .A(compare_i_data_rs[17]), .Q(n107) );
  NAND26 U528 ( .A(n625), .B(n624), .Q(alu_i_data_B[16]) );
  NAND41 U529 ( .A(n81), .B(n379), .C(n380), .D(n382), .Q(n304) );
  NAND22 U530 ( .A(compare_i_data_rt[16]), .B(n623), .Q(n625) );
  INV3 U531 ( .A(alu_i_data_B[23]), .Q(n109) );
  INV3 U532 ( .A(alu_i_data_B[13]), .Q(n110) );
  INV3 U533 ( .A(u_alu_lt_x_11_B_2_), .Q(n111) );
  NAND21 U534 ( .A(compare_i_data_rt[27]), .B(n623), .Q(n579) );
  NAND22 U535 ( .A(compare_i_data_rt[18]), .B(n623), .Q(n615) );
  INV3 U536 ( .A(alu_i_data_B[28]), .Q(n113) );
  INV3 U537 ( .A(n81), .Q(n114) );
  NAND21 U538 ( .A(compare_i_data_rt[31]), .B(n623), .Q(n563) );
  NAND21 U539 ( .A(compare_i_data_rt[29]), .B(n623), .Q(n571) );
  INV3 U540 ( .A(alu_i_data_B[4]), .Q(n115) );
  INV2 U541 ( .A(compare_i_data_rt[25]), .Q(n587) );
  NAND21 U542 ( .A(compare_i_data_rt[26]), .B(n623), .Q(n583) );
  NAND21 U543 ( .A(compare_i_data_rt[30]), .B(n623), .Q(n567) );
  INV2 U544 ( .A(alu_i_con_AluCtrl[2]), .Q(n962) );
  INV3 U545 ( .A(alu_i_data_B[9]), .Q(n116) );
  INV3 U546 ( .A(alu_i_data_B[1]), .Q(n117) );
  INV2 U547 ( .A(alu_i_con_AluCtrl[3]), .Q(n543) );
  NAND31 U548 ( .A(n648), .B(n647), .C(n646), .Q(compare_i_data_rt[9]) );
  INV2 U549 ( .A(n1324), .Q(n1317) );
  OAI2111 U550 ( .A(n1329), .B(n1328), .C(n1327), .D(n1326), .Q(
        alu_i_con_AluCtrl[3]) );
  NAND31 U551 ( .A(n1324), .B(n1327), .C(n1323), .Q(alu_i_con_AluCtrl[2]) );
  NAND21 U552 ( .A(compare_i_data_rt[28]), .B(n623), .Q(n575) );
  NAND31 U553 ( .A(n606), .B(n605), .C(n604), .Q(compare_i_data_rt[20]) );
  NAND21 U554 ( .A(n897), .B(i_data_rs[26]), .Q(n818) );
  NAND22 U555 ( .A(n229), .B(i_data_rt[27]), .Q(n578) );
  NAND22 U556 ( .A(n229), .B(i_data_rt[26]), .Q(n582) );
  NAND22 U557 ( .A(n229), .B(i_data_rt[25]), .Q(n586) );
  NAND22 U558 ( .A(n229), .B(i_data_rt[31]), .Q(n562) );
  AOI221 U559 ( .A(n1316), .B(n1325), .C(i_con_Ealuop[0]), .D(i_con_Ealuop[5]), 
        .Q(n1324) );
  NAND21 U560 ( .A(n897), .B(i_data_rs[28]), .Q(n804) );
  NAND22 U561 ( .A(n897), .B(i_data_rs[31]), .Q(n784) );
  OAI211 U562 ( .A(n889), .B(n888), .C(n1325), .Q(n1326) );
  INV2 U563 ( .A(n1262), .Q(n1316) );
  NAND22 U564 ( .A(n521), .B(i_data_FEalures[15]), .Q(n626) );
  BUF15 U565 ( .A(n897), .Q(n118) );
  NOR21 U566 ( .A(i_con_Efamux[1]), .B(n527), .Q(n529) );
  AOI2111 U567 ( .A(n1308), .B(i_data_immext[2]), .C(n882), .D(n881), .Q(n883)
         );
  INV15 U568 ( .A(n523), .Q(n120) );
  NOR21 U569 ( .A(n539), .B(n538), .Q(n879) );
  OAI211 U570 ( .A(i_con_Ealuop[5]), .B(n1313), .C(i_con_Ealuop[0]), .Q(n1314)
         );
  NOR22 U571 ( .A(n534), .B(n528), .Q(n906) );
  INV2 U572 ( .A(u_alu_ashr_4_SH_3_), .Q(n520) );
  NOR21 U573 ( .A(i_con_Ealuop[2]), .B(n1312), .Q(n1313) );
  NAND31 U574 ( .A(n540), .B(n874), .C(n877), .Q(n878) );
  NOR21 U575 ( .A(i_con_Ealuop[4]), .B(n1328), .Q(n1311) );
  INV2 U576 ( .A(i_data_FWmemout[20]), .Q(n845) );
  INV3 U577 ( .A(i_data_FWmemout[31]), .Q(n778) );
  INV3 U578 ( .A(i_data_FWmemout[15]), .Q(n1330) );
  INV2 U579 ( .A(i_data_FWmemout[22]), .Q(n835) );
  INV2 U580 ( .A(i_data_FWmemout[21]), .Q(n842) );
  INV2 U581 ( .A(i_data_FWmemout[27]), .Q(n807) );
  INV2 U582 ( .A(i_data_FWmemout[17]), .Q(n869) );
  INV2 U583 ( .A(i_data_FWmemout[14]), .Q(n683) );
  INV2 U584 ( .A(i_data_FWmemout[16]), .Q(n903) );
  INV2 U585 ( .A(i_con_bop[0]), .Q(n953) );
  AOI211 U586 ( .A(i_con_bop[0]), .B(i_con_bop[2]), .C(i_con_bop[1]), .Q(n960)
         );
  INV2 U587 ( .A(i_con_bop[1]), .Q(n951) );
  INV2 U588 ( .A(i_con_bop[2]), .Q(n952) );
  INV2 U589 ( .A(i_data_FWmemout[10]), .Q(n711) );
  INV2 U590 ( .A(i_data_FWmemout[12]), .Q(n697) );
  INV2 U591 ( .A(i_data_FWmemout[13]), .Q(n690) );
  INV2 U592 ( .A(i_data_FWmemout[11]), .Q(n704) );
  INV2 U593 ( .A(i_con_Ealuop[3]), .Q(n1312) );
  INV3 U594 ( .A(i_con_Efamux[1]), .Q(n534) );
  INV2 U595 ( .A(i_data_FWmemout[29]), .Q(n797) );
  INV1 U596 ( .A(i_con_Ealuop[2]), .Q(n1309) );
  NAND21 U597 ( .A(i_data_immext[1]), .B(i_data_immext[3]), .Q(n539) );
  INV2 U598 ( .A(i_data_FWmemout[24]), .Q(n892) );
  INV1 U599 ( .A(i_data_immext[0]), .Q(n881) );
  INV3 U600 ( .A(i_con_Ealuop[1]), .Q(n1318) );
  INV2 U601 ( .A(i_con_Ealuop[4]), .Q(n1329) );
  INV2 U602 ( .A(i_data_FWmemout[28]), .Q(n800) );
  INV2 U603 ( .A(i_data_FWmemout[30]), .Q(n787) );
  INV2 U604 ( .A(i_data_FWmemout[18]), .Q(n862) );
  INV2 U605 ( .A(i_data_FWmemout[26]), .Q(n814) );
  INV3 U606 ( .A(i_con_Malupc8), .Q(n1336) );
  BUF6 U607 ( .A(i_con_Ealusrc), .Q(n235) );
  INV2 U608 ( .A(i_data_FWmemout[19]), .Q(n855) );
  INV2 U609 ( .A(i_data_FWmemout[25]), .Q(n821) );
  INV2 U610 ( .A(i_data_FWmemout[23]), .Q(n828) );
  BUF6 U611 ( .A(i_data_immext[10]), .Q(n378) );
  XNR21 U612 ( .A(DP_OP_77_130_260_n4), .B(u_alu_sum_1_8_), .Q(u_alu_N165) );
  INV3 U613 ( .A(DP_OP_77_130_260_n23), .Q(DP_OP_77_130_260_n30) );
  INV3 U614 ( .A(DP_OP_77_130_260_n24), .Q(DP_OP_77_130_260_n22) );
  INV3 U615 ( .A(DP_OP_77_130_260_n15), .Q(DP_OP_77_130_260_n28) );
  INV3 U616 ( .A(DP_OP_77_130_260_n16), .Q(DP_OP_77_130_260_n14) );
  XOR20 U617 ( .A(DP_OP_77_130_260_n3), .B(DP_OP_77_130_260_n20), .Q(
        u_alu_N166) );
  ADD32 U618 ( .A(alu_i_data_B[12]), .B(compare_i_data_rs[12]), .CI(
        DP_OP_77_130_260_n9), .CO(DP_OP_77_130_260_n8), .S(u_alu_N169) );
  ADD32 U619 ( .A(alu_i_data_B[13]), .B(compare_i_data_rs[13]), .CI(
        DP_OP_77_130_260_n8), .CO(DP_OP_77_130_260_n7), .S(u_alu_N170) );
  ADD32 U620 ( .A(alu_i_data_B[14]), .B(compare_i_data_rs[14]), .CI(
        DP_OP_77_130_260_n7), .CO(DP_OP_77_130_260_n6), .S(u_alu_N171) );
  ADD32 U621 ( .A(alu_i_data_B[15]), .B(n80), .CI(DP_OP_77_130_260_n6), .CO(
        u_alu_N173), .S(u_alu_N172) );
  NAND22 U622 ( .A(compare_i_data_rs[16]), .B(alu_i_data_B[16]), .Q(n136) );
  INV3 U623 ( .A(n136), .Q(u_alu_DP_OP_83J3_124_3384_n15) );
  XOR21 U624 ( .A(compare_i_data_rs[16]), .B(alu_i_data_B[16]), .Q(
        u_alu_pre_sum_3a[0]) );
  NAND22 U625 ( .A(u_alu_DP_OP_83J3_124_3384_n11), .B(alu_i_data_B[21]), .Q(
        n130) );
  XOR21 U626 ( .A(u_alu_DP_OP_83J3_124_3384_n11), .B(n131), .Q(
        u_alu_pre_sum_3a[5]) );
  XOR21 U627 ( .A(u_alu_DP_OP_83J3_124_3384_n12), .B(n127), .Q(
        u_alu_pre_sum_3a[4]) );
  NAND22 U628 ( .A(u_alu_DP_OP_83J3_124_3384_n13), .B(compare_i_data_rs[19]), 
        .Q(n134) );
  NAND22 U629 ( .A(u_alu_DP_OP_83J3_124_3384_n12), .B(n83), .Q(n125) );
  NAND22 U630 ( .A(compare_i_data_rs[20]), .B(n83), .Q(n124) );
  NAND33 U631 ( .A(n126), .B(n125), .C(n124), .Q(u_alu_DP_OP_83J3_124_3384_n11) );
  XOR22 U632 ( .A(u_alu_DP_OP_83J3_124_3384_n1), .B(u_alu_pre_sum_3a[8]), .Q(
        u_alu_pre_sum_3b[8]) );
  ADD32 U633 ( .A(alu_i_data_B[18]), .B(compare_i_data_rs[18]), .CI(
        u_alu_DP_OP_83J3_124_3384_n14), .CO(u_alu_DP_OP_83J3_124_3384_n13), 
        .S(u_alu_pre_sum_3a[2]) );
  ADD22 U634 ( .A(u_alu_pre_sum_3a[5]), .B(u_alu_DP_OP_83J3_124_3384_n4), .CO(
        u_alu_DP_OP_83J3_124_3384_n3), .S(u_alu_pre_sum_3b[5]) );
  ADD22 U635 ( .A(u_alu_pre_sum_3a[6]), .B(u_alu_DP_OP_83J3_124_3384_n3), .CO(
        u_alu_DP_OP_83J3_124_3384_n2), .S(u_alu_pre_sum_3b[6]) );
  NAND22 U636 ( .A(n87), .B(compare_i_data_rs[16]), .Q(
        u_alu_DP_OP_85J3_126_1427_n191) );
  NOR21 U637 ( .A(compare_i_data_rs[17]), .B(n108), .Q(
        u_alu_DP_OP_85J3_126_1427_n90) );
  NAND22 U638 ( .A(n108), .B(compare_i_data_rs[17]), .Q(
        u_alu_DP_OP_85J3_126_1427_n91) );
  NOR21 U639 ( .A(compare_i_data_rs[16]), .B(n87), .Q(
        u_alu_DP_OP_85J3_126_1427_n92) );
  INV3 U640 ( .A(u_alu_DP_OP_85J3_126_1427_n48), .Q(
        u_alu_DP_OP_85J3_126_1427_n197) );
  INV3 U641 ( .A(u_alu_DP_OP_85J3_126_1427_n55), .Q(
        u_alu_DP_OP_85J3_126_1427_n198) );
  INV3 U642 ( .A(u_alu_DP_OP_85J3_126_1427_n187), .Q(
        u_alu_DP_OP_85J3_126_1427_n186) );
  INV3 U643 ( .A(u_alu_DP_OP_85J3_126_1427_n89), .Q(
        u_alu_DP_OP_85J3_126_1427_n88) );
  INV3 U644 ( .A(u_alu_DP_OP_85J3_126_1427_n24), .Q(
        u_alu_DP_OP_85J3_126_1427_n95) );
  INV3 U645 ( .A(u_alu_DP_OP_85J3_126_1427_n49), .Q(
        u_alu_DP_OP_85J3_126_1427_n145) );
  NAND22 U646 ( .A(n88), .B(compare_i_data_rs[24]), .Q(
        u_alu_DP_OP_85J3_126_1427_n44) );
  INV3 U647 ( .A(alu_i_data_B[25]), .Q(u_alu_DP_OP_85J3_126_1427_n214) );
  INV3 U648 ( .A(u_alu_DP_OP_85J3_126_1427_n40), .Q(
        u_alu_DP_OP_85J3_126_1427_n195) );
  INV3 U649 ( .A(u_alu_DP_OP_85J3_126_1427_n41), .Q(
        u_alu_DP_OP_85J3_126_1427_n137) );
  INV3 U650 ( .A(u_alu_DP_OP_85J3_126_1427_n32), .Q(
        u_alu_DP_OP_85J3_126_1427_n193) );
  INV3 U651 ( .A(u_alu_DP_OP_85J3_126_1427_n33), .Q(
        u_alu_DP_OP_85J3_126_1427_n129) );
  INV3 U652 ( .A(u_alu_DP_OP_85J3_126_1427_n174), .Q(
        u_alu_DP_OP_85J3_126_1427_n173) );
  INV3 U653 ( .A(u_alu_DP_OP_85J3_126_1427_n76), .Q(
        u_alu_DP_OP_85J3_126_1427_n75) );
  INV3 U654 ( .A(u_alu_DP_OP_85J3_126_1427_n73), .Q(
        u_alu_DP_OP_85J3_126_1427_n200) );
  INV3 U655 ( .A(u_alu_DP_OP_85J3_126_1427_n74), .Q(
        u_alu_DP_OP_85J3_126_1427_n166) );
  AOI212 U656 ( .A(u_alu_DP_OP_85J3_126_1427_n26), .B(
        u_alu_DP_OP_85J3_126_1427_n95), .C(u_alu_DP_OP_85J3_126_1427_n23), .Q(
        u_alu_DP_OP_85J3_126_1427_n21) );
  INV0 U657 ( .A(u_alu_sub_x_2_n25), .Q(u_alu_sub_x_2_n86) );
  INV3 U658 ( .A(alu_i_data_B[14]), .Q(u_alu_sub_x_2_n99) );
  INV3 U659 ( .A(n112), .Q(u_alu_sub_x_2_n107) );
  INV3 U660 ( .A(alu_i_data_B[10]), .Q(u_alu_sub_x_2_n103) );
  INV3 U661 ( .A(u_alu_sub_x_2_n37), .Q(u_alu_sub_x_2_n88) );
  INV3 U662 ( .A(u_alu_sub_x_2_n22), .Q(u_alu_sub_x_2_n85) );
  INV3 U663 ( .A(u_alu_sub_x_2_n23), .Q(u_alu_sub_x_2_n21) );
  INV3 U664 ( .A(u_alu_sub_x_2_n50), .Q(u_alu_sub_x_2_n49) );
  NOR21 U665 ( .A(compare_i_data_rs[3]), .B(n234), .Q(u_alu_sub_x_2_n74) );
  NOR21 U666 ( .A(compare_i_data_rs[1]), .B(n117), .Q(u_alu_sub_x_2_n81) );
  NAND22 U667 ( .A(n117), .B(compare_i_data_rs[1]), .Q(u_alu_sub_x_2_n82) );
  NAND22 U668 ( .A(n234), .B(compare_i_data_rs[3]), .Q(u_alu_sub_x_2_n75) );
  NAND20 U669 ( .A(n106), .B(alu_i_data_B[28]), .Q(n138) );
  NAND20 U670 ( .A(compare_i_data_rs[29]), .B(n90), .Q(n139) );
  AOI220 U671 ( .A(n93), .B(compare_i_data_rs[27]), .C(n85), .D(
        compare_i_data_rs[26]), .Q(n200) );
  NOR20 U672 ( .A(compare_i_data_rs[24]), .B(n88), .Q(n140) );
  MAJ31 U673 ( .A(alu_i_data_B[25]), .B(n218), .C(n140), .Q(n143) );
  NOR20 U674 ( .A(compare_i_data_rs[26]), .B(n85), .Q(n141) );
  IMAJ30 U675 ( .A(n93), .B(compare_i_data_rs[27]), .C(n219), .Q(n142) );
  NOR20 U676 ( .A(compare_i_data_rs[30]), .B(n89), .Q(n145) );
  NOR20 U677 ( .A(alu_i_data_B[17]), .B(n107), .Q(n186) );
  OAI220 U678 ( .A(n104), .B(alu_i_data_B[23]), .C(n100), .D(alu_i_data_B[22]), 
        .Q(n198) );
  NAND20 U679 ( .A(compare_i_data_rs[21]), .B(n92), .Q(n147) );
  NOR20 U680 ( .A(alu_i_data_B[19]), .B(n101), .Q(n148) );
  AOI210 U681 ( .A(compare_i_data_rs[18]), .B(n84), .C(n148), .Q(n191) );
  NOR20 U682 ( .A(alu_i_data_B[13]), .B(n210), .Q(n150) );
  NAND20 U683 ( .A(n80), .B(n86), .Q(n149) );
  NOR20 U684 ( .A(alu_i_data_B[9]), .B(n208), .Q(n151) );
  OAI220 U685 ( .A(alu_i_data_B[11]), .B(n102), .C(alu_i_data_B[10]), .D(n209), 
        .Q(n172) );
  OAI210 U686 ( .A(n112), .B(n207), .C(n152), .Q(n167) );
  AOI210 U687 ( .A(compare_i_data_rs[2]), .B(n111), .C(n153), .Q(n158) );
  OAI210 U688 ( .A(alu_i_data_B[1]), .B(n204), .C(n81), .Q(n154) );
  OAI220 U689 ( .A(compare_i_data_rs[0]), .B(n154), .C(compare_i_data_rs[1]), 
        .D(n117), .Q(n157) );
  NOR20 U690 ( .A(compare_i_data_rs[2]), .B(n111), .Q(n155) );
  MAJ31 U691 ( .A(alu_i_data_B[3]), .B(n205), .C(n155), .Q(n156) );
  AOI2110 U692 ( .A(compare_i_data_rs[4]), .B(n115), .C(n160), .D(n159), .Q(
        n163) );
  NOR20 U693 ( .A(compare_i_data_rs[4]), .B(n115), .Q(n161) );
  MAJ31 U694 ( .A(alu_i_data_B[5]), .B(n206), .C(n161), .Q(n162) );
  NAND20 U695 ( .A(n112), .B(n207), .Q(n164) );
  MAJ31 U696 ( .A(compare_i_data_rs[7]), .B(n233), .C(n164), .Q(n165) );
  NOR20 U697 ( .A(n94), .B(compare_i_data_rs[12]), .Q(n168) );
  IMAJ30 U698 ( .A(n210), .B(alu_i_data_B[13]), .C(n168), .Q(n179) );
  NAND20 U699 ( .A(alu_i_data_B[14]), .B(n211), .Q(n169) );
  MAJ31 U700 ( .A(n80), .B(n86), .C(n169), .Q(n177) );
  NAND20 U701 ( .A(n209), .B(alu_i_data_B[10]), .Q(n170) );
  IMAJ30 U702 ( .A(n96), .B(compare_i_data_rs[11]), .C(n170), .Q(n175) );
  IMAJ30 U703 ( .A(n208), .B(alu_i_data_B[9]), .C(n171), .Q(n173) );
  NAND20 U704 ( .A(n83), .B(n103), .Q(n187) );
  MAJ31 U705 ( .A(compare_i_data_rs[21]), .B(n92), .C(n187), .Q(n199) );
  NAND20 U706 ( .A(alu_i_data_B[22]), .B(n100), .Q(n188) );
  IMAJ30 U707 ( .A(n104), .B(alu_i_data_B[23]), .C(n214), .Q(n197) );
  MAJ31 U708 ( .A(alu_i_data_B[19]), .B(n101), .C(n189), .Q(n195) );
  NAND20 U709 ( .A(alu_i_data_B[16]), .B(n212), .Q(n190) );
  MAJ31 U710 ( .A(compare_i_data_rs[17]), .B(n108), .C(n190), .Q(n192) );
  NOR20 U711 ( .A(alu_i_data_B[24]), .B(n217), .Q(n203) );
  INV0 U712 ( .A(compare_i_data_rs[13]), .Q(n210) );
  INV0 U713 ( .A(compare_i_data_rs[14]), .Q(n211) );
  INV0 U714 ( .A(compare_i_data_rs[9]), .Q(n208) );
  INV0 U715 ( .A(compare_i_data_rs[10]), .Q(n209) );
  INV0 U716 ( .A(compare_i_data_rs[6]), .Q(n207) );
  INV0 U717 ( .A(compare_i_data_rs[5]), .Q(n206) );
  INV0 U718 ( .A(compare_i_data_rs[3]), .Q(n205) );
  INV0 U719 ( .A(compare_i_data_rs[1]), .Q(n204) );
  INV0 U720 ( .A(compare_i_data_rs[24]), .Q(n217) );
  AOI211 U721 ( .A(compare_i_data_rs[30]), .B(n89), .C(n137), .Q(n146) );
  OAI2111 U722 ( .A(alu_i_data_B[28]), .B(n106), .C(n146), .D(n139), .Q(n201)
         );
  AOI211 U723 ( .A(n200), .B(n143), .C(n142), .Q(n144) );
  AOI211 U724 ( .A(n158), .B(n157), .C(n156), .Q(n159) );
  NOR21 U725 ( .A(n163), .B(n162), .Q(n166) );
  OAI212 U726 ( .A(n167), .B(n166), .C(n165), .Q(n181) );
  NOR21 U727 ( .A(n173), .B(n172), .Q(n174) );
  OAI2111 U728 ( .A(n179), .B(n178), .C(n177), .D(n176), .Q(n180) );
  AOI311 U729 ( .A(n183), .B(n182), .C(n181), .D(n180), .Q(n184) );
  NOR21 U730 ( .A(n192), .B(n213), .Q(n194) );
  OAI212 U731 ( .A(n195), .B(n194), .C(n216), .Q(n196) );
  OAI2111 U732 ( .A(n83), .B(n103), .C(n215), .D(n147), .Q(n193) );
  AOI2110 U733 ( .A(compare_i_data_rs[8]), .B(n95), .C(n151), .D(n172), .Q(
        n182) );
  NAND20 U734 ( .A(compare_i_data_rs[7]), .B(n233), .Q(n152) );
  NOR20 U735 ( .A(n95), .B(compare_i_data_rs[8]), .Q(n171) );
  NOR20 U736 ( .A(alu_i_data_B[5]), .B(n206), .Q(n160) );
  NOR20 U737 ( .A(alu_i_data_B[3]), .B(n205), .Q(n153) );
  OAI210 U738 ( .A(alu_i_data_B[14]), .B(n211), .C(n149), .Q(n178) );
  AOI2110 U739 ( .A(compare_i_data_rs[12]), .B(n94), .C(n150), .D(n178), .Q(
        n183) );
  XOR31 U740 ( .A(alu_i_data_B[31]), .B(u_alu_DP_OP_84J3_125_2615_n9), .C(
        compare_i_data_rs[31]), .Q(u_alu_pre_sum_4a[7]) );
  ADD22 U741 ( .A(compare_i_data_rs[24]), .B(alu_i_data_B[24]), .CO(
        u_alu_DP_OP_84J3_125_2615_n15), .S(u_alu_pre_sum_4a[0]) );
  AOI221 U742 ( .A(n671), .B(i_data_FMalures[6]), .C(n521), .D(
        i_data_FEalures[6]), .Q(n656) );
  NAND33 U743 ( .A(n676), .B(n675), .C(n674), .Q(compare_i_data_rt[0]) );
  AOI221 U744 ( .A(n671), .B(i_data_FMalures[16]), .C(n521), .D(
        i_data_FEalures[16]), .Q(n621) );
  AOI220 U745 ( .A(n673), .B(i_data_FMmemout[11]), .C(n672), .D(
        i_data_FWmemout[11]), .Q(n640) );
  AOI220 U746 ( .A(n673), .B(i_data_FMmemout[10]), .C(n672), .D(
        i_data_FWmemout[10]), .Q(n643) );
  AOI220 U747 ( .A(n673), .B(i_data_FMmemout[9]), .C(n672), .D(
        i_data_FWmemout[9]), .Q(n646) );
  CLKBU15 U748 ( .A(n673), .Q(n231) );
  NAND24 U749 ( .A(n550), .B(n554), .Q(n558) );
  INV15 U750 ( .A(n558), .Q(n671) );
  MUX26 U751 ( .A(compare_i_data_rt[2]), .B(i_data_immext[2]), .S(n235), .Q(
        u_alu_lt_x_11_B_2_) );
  AOI221 U752 ( .A(n231), .B(i_data_FMmemout[21]), .C(n672), .D(
        i_data_FWmemout[21]), .Q(n600) );
  NAND22 U753 ( .A(n1252), .B(u_alu_pre_suba[14]), .Q(n1233) );
  NAND33 U754 ( .A(n669), .B(n668), .C(n667), .Q(compare_i_data_rt[1]) );
  MUX26 U755 ( .A(compare_i_data_rt[1]), .B(i_data_immext[1]), .S(n235), .Q(
        alu_i_data_B[1]) );
  OAI212 U756 ( .A(n903), .B(n119), .C(n901), .Q(n904) );
  IMUX21 U757 ( .A(u_alu_pre_sum_3a[8]), .B(u_alu_pre_sum_3b[8]), .S(
        u_alu_N173), .Q(n1160) );
  OAI210 U758 ( .A(n1244), .B(u_alu_N306), .C(compare_i_data_rs[31]), .Q(n964)
         );
  AOI211 U759 ( .A(u_alu_N306), .B(n963), .C(n962), .Q(n979) );
  IMUX20 U760 ( .A(n459), .B(n462), .S(n381), .Q(n481) );
  IMUX20 U761 ( .A(n473), .B(n472), .S(n381), .Q(n497) );
  NAND20 U762 ( .A(u_alu_sum_1_7_), .B(n1159), .Q(n994) );
  NAND22 U763 ( .A(u_alu_N234), .B(n1251), .Q(n1017) );
  NAND22 U764 ( .A(u_alu_N231), .B(n1251), .Q(n987) );
  NAND20 U765 ( .A(u_alu_sum_1_6_), .B(n1159), .Q(n983) );
  NAND20 U766 ( .A(u_alu_N221), .B(n1250), .Q(n1210) );
  NAND22 U767 ( .A(u_alu_pre_sum_4b[7]), .B(n1241), .Q(n1260) );
  NAND20 U768 ( .A(u_alu_N223), .B(n1250), .Q(n1235) );
  IMUX20 U769 ( .A(n315), .B(n291), .S(i_data_immext[8]), .Q(n345) );
  NAND22 U770 ( .A(u_alu_pre_sum_4b[6]), .B(n1241), .Q(n1239) );
  IMUX20 U771 ( .A(n491), .B(n417), .S(i_data_immext[8]), .Q(n464) );
  AOI211 U772 ( .A(alu_i_data_B[10]), .B(n1024), .C(n1023), .Q(n1028) );
  IMUX20 U773 ( .A(n496), .B(n422), .S(i_data_immext[8]), .Q(n475) );
  NAND20 U774 ( .A(u_alu_N217), .B(n1250), .Q(n1167) );
  IMUX20 U775 ( .A(n290), .B(n280), .S(n381), .Q(n301) );
  IMUX20 U776 ( .A(n461), .B(n388), .S(n381), .Q(n480) );
  IMUX20 U777 ( .A(n308), .B(n286), .S(i_data_immext[8]), .Q(n336) );
  NAND30 U778 ( .A(n1263), .B(n1217), .C(n90), .Q(n1218) );
  IMUX20 U779 ( .A(n291), .B(n270), .S(i_data_immext[8]), .Q(n316) );
  INV3 U780 ( .A(i_data_immext[6]), .Q(n382) );
  IMUX20 U781 ( .A(n281), .B(n258), .S(i_data_immext[8]), .Q(n302) );
  IMUX21 U782 ( .A(n269), .B(n257), .S(u_alu_ashr_4_SH_1_), .Q(n281) );
  NAND22 U783 ( .A(n122), .B(i_data_FMmemout[21]), .Q(n841) );
  AOI2111 U784 ( .A(i_data_FMmemout[31]), .B(n122), .C(n782), .D(n781), .Q(
        n783) );
  NAND22 U785 ( .A(n230), .B(i_data_rt[22]), .Q(n598) );
  AOI221 U786 ( .A(n231), .B(i_data_FMmemout[20]), .C(n672), .D(
        i_data_FWmemout[20]), .Q(n604) );
  NAND22 U787 ( .A(n229), .B(i_data_rt[20]), .Q(n606) );
  AOI2111 U788 ( .A(n98), .B(compare_i_data_rs[17]), .C(n1083), .D(n1082), .Q(
        n1087) );
  INV3 U789 ( .A(i_con_Ealuop[0]), .Q(n1328) );
  AOI211 U790 ( .A(n882), .B(n874), .C(n884), .Q(n541) );
  NAND22 U791 ( .A(n885), .B(n878), .Q(n884) );
  NAND22 U792 ( .A(n879), .B(i_data_immext[0]), .Q(n885) );
  INV3 U793 ( .A(n538), .Q(n882) );
  NOR21 U794 ( .A(n1318), .B(i_con_Ealuop[0]), .Q(n1325) );
  AOI221 U795 ( .A(n231), .B(i_data_FMmemout[13]), .C(n672), .D(
        i_data_FWmemout[13]), .Q(n634) );
  NAND31 U796 ( .A(n651), .B(n650), .C(n649), .Q(compare_i_data_rt[8]) );
  NAND22 U797 ( .A(n729), .B(n728), .Q(compare_i_data_rs[8]) );
  NAND22 U798 ( .A(n228), .B(i_data_rt[11]), .Q(n642) );
  AOI220 U799 ( .A(n231), .B(i_data_FMmemout[3]), .C(n672), .D(
        i_data_FWmemout[3]), .Q(n661) );
  AOI220 U800 ( .A(n671), .B(i_data_FMalures[3]), .C(n521), .D(
        i_data_FEalures[3]), .Q(n662) );
  AOI220 U801 ( .A(n671), .B(i_data_FMalures[1]), .C(n521), .D(
        i_data_FEalures[1]), .Q(n668) );
  NAND20 U802 ( .A(n230), .B(i_data_rt[0]), .Q(n676) );
  BUF6 U803 ( .A(i_data_immext[7]), .Q(u_alu_ashr_4_SH_1_) );
  AOI220 U804 ( .A(n671), .B(i_data_FMalures[7]), .C(n521), .D(
        i_data_FEalures[7]), .Q(n653) );
  NAND20 U805 ( .A(n122), .B(i_data_FMmemout[6]), .Q(n738) );
  AOI220 U806 ( .A(n671), .B(i_data_FMalures[4]), .C(n521), .D(
        i_data_FEalures[4]), .Q(n659) );
  NAND20 U807 ( .A(n230), .B(i_data_rt[4]), .Q(n660) );
  NAND22 U808 ( .A(n229), .B(i_data_rt[12]), .Q(n639) );
  NAND22 U809 ( .A(n229), .B(i_data_rt[14]), .Q(n633) );
  INV6 U810 ( .A(n902), .Q(n524) );
  NAND20 U811 ( .A(u_alu_N229), .B(n1251), .Q(n772) );
  AOI220 U812 ( .A(n1159), .B(u_alu_sum_1_5_), .C(u_alu_half_sub_5_), .D(n1064), .Q(n769) );
  IMUX21 U813 ( .A(n472), .B(n437), .S(u_alu_ashr_4_SH_1_), .Q(n484) );
  IMUX21 U814 ( .A(n462), .B(n461), .S(u_alu_ashr_4_SH_1_), .Q(n492) );
  OAI2111 U815 ( .A(n985), .B(n221), .C(n984), .D(n983), .Q(n986) );
  IMUX21 U816 ( .A(n388), .B(n387), .S(u_alu_ashr_4_SH_1_), .Q(n491) );
  IMUX21 U817 ( .A(n437), .B(n406), .S(u_alu_ashr_4_SH_1_), .Q(n496) );
  IMUX21 U818 ( .A(n387), .B(n390), .S(u_alu_ashr_4_SH_1_), .Q(n401) );
  IMUX21 U819 ( .A(n295), .B(n285), .S(u_alu_ashr_4_SH_1_), .Q(n308) );
  IMUX21 U820 ( .A(n239), .B(n241), .S(u_alu_ashr_4_SH_1_), .Q(n251) );
  IMUX21 U821 ( .A(n257), .B(n249), .S(u_alu_ashr_4_SH_1_), .Q(n270) );
  AOI2110 U822 ( .A(n98), .B(compare_i_data_rs[18]), .C(n1097), .D(n1096), .Q(
        n1101) );
  IMUX21 U823 ( .A(n321), .B(n296), .S(i_data_immext[8]), .Q(n353) );
  IMUX21 U824 ( .A(n285), .B(n274), .S(u_alu_ashr_4_SH_1_), .Q(n296) );
  IMUX21 U825 ( .A(n307), .B(n295), .S(u_alu_ashr_4_SH_1_), .Q(n321) );
  NAND22 U826 ( .A(n866), .B(n865), .Q(compare_i_data_rs[18]) );
  NOR31 U827 ( .A(n884), .B(n888), .C(n883), .Q(n1315) );
  AOI211 U828 ( .A(alu_i_data_B[3]), .B(n98), .C(n1282), .Q(n1279) );
  NAND22 U829 ( .A(n1252), .B(u_alu_pre_suba[15]), .Q(n1253) );
  AOI2111 U830 ( .A(u_alu_N165), .B(n1159), .C(n1006), .D(n1005), .Q(n1008) );
  NAND20 U831 ( .A(n122), .B(i_data_FMmemout[20]), .Q(n844) );
  NOR23 U832 ( .A(n767), .B(alu_i_con_AluCtrl[3]), .Q(n1251) );
  NAND24 U833 ( .A(n619), .B(n624), .Q(alu_i_data_B[17]) );
  AOI221 U834 ( .A(n231), .B(i_data_FMmemout[17]), .C(n672), .D(
        i_data_FWmemout[17]), .Q(n616) );
  NAND22 U835 ( .A(n122), .B(i_data_FMmemout[17]), .Q(n868) );
  AOI211 U836 ( .A(i_data_immext[2]), .B(n877), .C(n876), .Q(n886) );
  AOI220 U837 ( .A(n671), .B(i_data_FMalures[13]), .C(n521), .D(
        i_data_FEalures[13]), .Q(n635) );
  AOI221 U838 ( .A(n671), .B(i_data_FMalures[8]), .C(n521), .D(
        i_data_FEalures[8]), .Q(n650) );
  AOI221 U839 ( .A(n122), .B(i_data_FMmemout[3]), .C(n524), .D(
        i_data_FWmemout[3]), .Q(n747) );
  NAND22 U840 ( .A(n229), .B(i_data_rt[2]), .Q(n666) );
  AOI221 U841 ( .A(n122), .B(i_data_FMmemout[1]), .C(n524), .D(
        i_data_FWmemout[1]), .Q(n753) );
  AOI221 U842 ( .A(n523), .B(i_data_FMalures[1]), .C(n121), .D(
        i_data_FEalures[1]), .Q(n754) );
  AOI220 U843 ( .A(n673), .B(i_data_FMmemout[12]), .C(n672), .D(
        i_data_FWmemout[12]), .Q(n637) );
  AOI220 U844 ( .A(n671), .B(i_data_FMalures[12]), .C(n521), .D(
        i_data_FEalures[12]), .Q(n638) );
  NOR24 U845 ( .A(n548), .B(n670), .Q(n228) );
  AOI2111 U846 ( .A(n98), .B(compare_i_data_rs[23]), .C(n1149), .D(n1148), .Q(
        n1154) );
  OAI212 U847 ( .A(n119), .B(n787), .C(n786), .Q(n788) );
  NOR21 U848 ( .A(n785), .B(n120), .Q(n789) );
  NAND22 U849 ( .A(n122), .B(i_data_FMmemout[18]), .Q(n861) );
  NAND22 U850 ( .A(n122), .B(i_data_FMmemout[19]), .Q(n854) );
  NAND20 U851 ( .A(n230), .B(i_data_rt[30]), .Q(n566) );
  NAND20 U852 ( .A(n230), .B(i_data_rt[29]), .Q(n570) );
  NAND20 U853 ( .A(n230), .B(i_data_rt[24]), .Q(n590) );
  NAND22 U854 ( .A(alu_i_data_B[3]), .B(compare_i_data_rs[3]), .Q(
        u_alu_add_x_1_n34) );
  NAND22 U855 ( .A(alu_i_data_B[1]), .B(compare_i_data_rs[1]), .Q(
        u_alu_add_x_1_n41) );
  AOI221 U856 ( .A(n231), .B(i_data_FMmemout[16]), .C(n672), .D(
        i_data_FWmemout[16]), .Q(n620) );
  AOI311 U857 ( .A(i_con_Ealuop[3]), .B(i_con_Ealuop[2]), .C(n1311), .D(n1320), 
        .Q(n1327) );
  NOR40 U858 ( .A(n1320), .B(n1319), .C(n1318), .D(n1317), .Q(n1321) );
  MUX22 U859 ( .A(compare_i_data_rt[13]), .B(i_data_immext[13]), .S(n235), .Q(
        alu_i_data_B[13]) );
  NAND31 U860 ( .A(n636), .B(n635), .C(n634), .Q(compare_i_data_rt[13]) );
  NAND22 U861 ( .A(n122), .B(i_data_FMmemout[10]), .Q(n710) );
  NAND22 U862 ( .A(n122), .B(i_data_FMmemout[9]), .Q(n717) );
  NAND33 U863 ( .A(n749), .B(n748), .C(n747), .Q(compare_i_data_rs[3]) );
  AOI221 U864 ( .A(n231), .B(i_data_FMmemout[2]), .C(n672), .D(
        i_data_FWmemout[2]), .Q(n664) );
  NAND22 U865 ( .A(n118), .B(i_data_rs[2]), .Q(n752) );
  NAND33 U866 ( .A(n755), .B(n754), .C(n753), .Q(compare_i_data_rs[1]) );
  AOI221 U867 ( .A(n231), .B(i_data_FMmemout[0]), .C(n672), .D(
        i_data_FWmemout[0]), .Q(n674) );
  NAND22 U868 ( .A(n230), .B(i_data_rt[7]), .Q(n654) );
  NAND22 U869 ( .A(n230), .B(i_data_rt[6]), .Q(n657) );
  OAI212 U870 ( .A(n739), .B(n119), .C(n738), .Q(n740) );
  AOI221 U871 ( .A(n122), .B(i_data_FMmemout[4]), .C(n524), .D(
        i_data_FWmemout[4]), .Q(n744) );
  AOI220 U872 ( .A(n671), .B(i_data_FMalures[14]), .C(n521), .D(
        i_data_FEalures[14]), .Q(n632) );
  INV6 U873 ( .A(n670), .Q(n522) );
  NOR33 U874 ( .A(n551), .B(i_con_Efbmux[1]), .C(i_con_Efbmux[0]), .Q(n673) );
  NAND24 U875 ( .A(n549), .B(n551), .Q(n547) );
  INV6 U876 ( .A(i_con_Efbmux[0]), .Q(n549) );
  AOI220 U877 ( .A(n1252), .B(u_alu_pre_suba[12]), .C(n1258), .D(
        u_alu_pre_subb[12]), .Q(n1213) );
  IMUX20 U878 ( .A(n333), .B(n320), .S(n381), .Q(n351) );
  IMUX20 U879 ( .A(n326), .B(n314), .S(n381), .Q(n343) );
  AOI211 U880 ( .A(u_alu_N241), .B(n1251), .C(n1076), .Q(n1077) );
  NAND22 U881 ( .A(n784), .B(n783), .Q(compare_i_data_rs[31]) );
  INV3 U882 ( .A(n380), .Q(n381) );
  AOI221 U883 ( .A(n231), .B(i_data_FMmemout[19]), .C(n672), .D(
        i_data_FWmemout[19]), .Q(n608) );
  AOI221 U884 ( .A(n231), .B(i_data_FMmemout[18]), .C(n672), .D(
        i_data_FWmemout[18]), .Q(n612) );
  OAI212 U885 ( .A(n119), .B(n869), .C(n868), .Q(n870) );
  AOI221 U886 ( .A(n671), .B(i_data_FMalures[10]), .C(n521), .D(
        i_data_FEalures[10]), .Q(n644) );
  AOI221 U887 ( .A(n671), .B(i_data_FMalures[9]), .C(n521), .D(
        i_data_FEalures[9]), .Q(n647) );
  AOI221 U888 ( .A(n231), .B(i_data_FMmemout[8]), .C(n672), .D(
        i_data_FWmemout[8]), .Q(n649) );
  NAND33 U889 ( .A(n752), .B(n751), .C(n750), .Q(compare_i_data_rs[2]) );
  AOI2111 U890 ( .A(n121), .B(i_data_FEalures[0]), .C(n760), .D(n759), .Q(n761) );
  AOI221 U891 ( .A(n231), .B(i_data_FMmemout[7]), .C(n672), .D(
        i_data_FWmemout[7]), .Q(n652) );
  OAI212 U892 ( .A(n732), .B(n119), .C(n731), .Q(n733) );
  AOI221 U893 ( .A(n231), .B(i_data_FMmemout[6]), .C(n672), .D(
        i_data_FWmemout[6]), .Q(n655) );
  AOI221 U894 ( .A(n671), .B(i_data_FMalures[5]), .C(n521), .D(
        i_data_FEalures[5]), .Q(n556) );
  AOI221 U895 ( .A(n231), .B(i_data_FMmemout[4]), .C(n672), .D(
        i_data_FWmemout[4]), .Q(n658) );
  NAND33 U896 ( .A(n746), .B(n745), .C(n744), .Q(compare_i_data_rs[4]) );
  MUX22 U897 ( .A(compare_i_data_rt[14]), .B(i_data_immext[14]), .S(n235), .Q(
        alu_i_data_B[14]) );
  AOI220 U898 ( .A(n673), .B(i_data_FMmemout[14]), .C(n672), .D(
        i_data_FWmemout[14]), .Q(n631) );
  INV12 U899 ( .A(n630), .Q(n672) );
  NAND24 U900 ( .A(n554), .B(n553), .Q(n630) );
  INV0 U901 ( .A(u_alu_add_x_1_n17), .Q(u_alu_add_x_1_n45) );
  AOI2111 U902 ( .A(n121), .B(i_data_FEalures[27]), .C(n809), .D(n808), .Q(
        n810) );
  AOI2111 U903 ( .A(n121), .B(i_data_FEalures[25]), .C(n823), .D(n822), .Q(
        n824) );
  AOI2111 U904 ( .A(n121), .B(i_data_FEalures[24]), .C(n894), .D(n893), .Q(
        n895) );
  OAI212 U905 ( .A(n119), .B(n862), .C(n861), .Q(n863) );
  OAI212 U906 ( .A(n119), .B(n855), .C(n854), .Q(n856) );
  OAI212 U907 ( .A(n235), .B(n587), .C(n624), .Q(alu_i_data_B[25]) );
  NOR21 U908 ( .A(n978), .B(n1267), .Q(n1265) );
  OAI212 U909 ( .A(n711), .B(n119), .C(n710), .Q(n712) );
  NAND22 U910 ( .A(n229), .B(i_data_rt[9]), .Q(n648) );
  OAI212 U911 ( .A(n718), .B(n119), .C(n717), .Q(n719) );
  NAND22 U912 ( .A(n229), .B(i_data_rt[8]), .Q(n651) );
  AOI2111 U913 ( .A(n121), .B(i_data_FEalures[8]), .C(n727), .D(n726), .Q(n728) );
  AOI221 U914 ( .A(n671), .B(i_data_FMalures[11]), .C(n521), .D(
        i_data_FEalures[11]), .Q(n641) );
  NOR21 U915 ( .A(n756), .B(n120), .Q(n760) );
  AOI2111 U916 ( .A(n121), .B(i_data_FEalures[7]), .C(n734), .D(n733), .Q(n735) );
  NOR21 U917 ( .A(n730), .B(n120), .Q(n734) );
  MUX22 U918 ( .A(compare_i_data_rt[15]), .B(i_data_immext[15]), .S(n235), .Q(
        alu_i_data_B[15]) );
  NOR22 U919 ( .A(i_con_Efbmux[1]), .B(n546), .Q(n548) );
  INV6 U920 ( .A(i_con_Efbmux[2]), .Q(n551) );
  AOI210 U921 ( .A(n982), .B(compare_i_data_rs[6]), .C(n981), .Q(n984) );
  NAND20 U922 ( .A(n1242), .B(n112), .Q(n1132) );
  AOI220 U923 ( .A(u_alu_N235), .B(n1251), .C(u_alu_N167), .D(n1159), .Q(n1027) );
  NOR21 U924 ( .A(n378), .B(n513), .Q(u_alu_N241) );
  AOI2111 U925 ( .A(n121), .B(i_data_FEalures[26]), .C(n816), .D(n815), .Q(
        n817) );
  AOI2111 U926 ( .A(n121), .B(i_data_FEalures[28]), .C(n802), .D(n801), .Q(
        n803) );
  AOI2111 U927 ( .A(n121), .B(i_data_FEalures[20]), .C(n847), .D(n846), .Q(
        n848) );
  BUF6 U928 ( .A(i_data_immext[9]), .Q(u_alu_ashr_4_SH_3_) );
  AOI2111 U929 ( .A(n121), .B(i_data_FEalures[9]), .C(n720), .D(n719), .Q(n721) );
  AOI221 U930 ( .A(n122), .B(i_data_FMmemout[2]), .C(n524), .D(
        i_data_FWmemout[2]), .Q(n750) );
  NAND22 U931 ( .A(n118), .B(i_data_rs[0]), .Q(n762) );
  AOI2111 U932 ( .A(n121), .B(i_data_FEalures[6]), .C(n741), .D(n740), .Q(n742) );
  NOR32 U933 ( .A(n531), .B(i_con_Efamux[1]), .C(i_con_Efamux[0]), .Q(n900) );
  NOR24 U934 ( .A(n529), .B(n121), .Q(n897) );
  NOR21 U935 ( .A(n378), .B(n518), .Q(u_alu_N244) );
  IMUX21 U936 ( .A(n446), .B(n445), .S(u_alu_ashr_4_SH_3_), .Q(n488) );
  IMUX20 U937 ( .A(n1179), .B(n1178), .S(alu_i_data_B[25]), .Q(n1182) );
  AOI211 U938 ( .A(u_alu_half_sub_11_), .B(n1064), .C(n1034), .Q(n1036) );
  IMUX21 U939 ( .A(n276), .B(n277), .S(u_alu_ashr_4_SH_3_), .Q(n324) );
  NAND22 U940 ( .A(n1241), .B(n223), .Q(n222) );
  IMUX21 U941 ( .A(n305), .B(n304), .S(u_alu_ashr_4_SH_3_), .Q(n362) );
  NOR21 U942 ( .A(n378), .B(n509), .Q(u_alu_N243) );
  NAND20 U943 ( .A(n1242), .B(u_alu_lt_x_11_B_7_), .Q(n1145) );
  INV6 U944 ( .A(n1264), .Q(n1266) );
  IMUX21 U945 ( .A(n395), .B(n397), .S(u_alu_ashr_4_SH_1_), .Q(n442) );
  AOI2111 U946 ( .A(n121), .B(i_data_FEalures[18]), .C(n864), .D(n863), .Q(
        n865) );
  AOI2111 U947 ( .A(n121), .B(i_data_FEalures[23]), .C(n830), .D(n829), .Q(
        n831) );
  AOI2111 U948 ( .A(n121), .B(i_data_FEalures[22]), .C(n837), .D(n836), .Q(
        n838) );
  NOR21 U949 ( .A(n378), .B(n515), .Q(u_alu_N242) );
  AOI2110 U950 ( .A(n231), .B(i_data_FMmemout[31]), .C(n560), .D(n559), .Q(
        n561) );
  NAND22 U951 ( .A(compare_i_data_rt[23]), .B(n623), .Q(n595) );
  NAND22 U952 ( .A(compare_i_data_rt[22]), .B(n623), .Q(n599) );
  NAND22 U953 ( .A(compare_i_data_rt[21]), .B(n623), .Q(n603) );
  NAND22 U954 ( .A(compare_i_data_rt[20]), .B(n623), .Q(n607) );
  NAND22 U955 ( .A(compare_i_data_rt[19]), .B(n623), .Q(n611) );
  NAND22 U956 ( .A(alu_i_con_AluCtrl[0]), .B(alu_i_con_AluCtrl[2]), .Q(n545)
         );
  NAND22 U957 ( .A(compare_i_data_rt[17]), .B(n623), .Q(n619) );
  AOI2111 U958 ( .A(n121), .B(i_data_FEalures[17]), .C(n871), .D(n870), .Q(
        n872) );
  NOR21 U959 ( .A(i_data_immext[3]), .B(i_data_immext[1]), .Q(n1307) );
  NOR31 U960 ( .A(i_data_immext[2]), .B(i_data_immext[0]), .C(i_data_immext[1]), .Q(n540) );
  AOI2111 U961 ( .A(n121), .B(i_data_FEalures[13]), .C(n692), .D(n691), .Q(
        n693) );
  AOI2111 U962 ( .A(n121), .B(i_data_FEalures[10]), .C(n713), .D(n712), .Q(
        n714) );
  AOI2111 U963 ( .A(n121), .B(i_data_FEalures[11]), .C(n706), .D(n705), .Q(
        n707) );
  MUX22 U964 ( .A(compare_i_data_rt[7]), .B(u_alu_ashr_4_SH_1_), .S(n235), .Q(
        alu_i_data_B[7]) );
  AOI221 U965 ( .A(n122), .B(i_data_FMmemout[5]), .C(n524), .D(
        i_data_FWmemout[5]), .Q(n535) );
  AOI2111 U966 ( .A(n121), .B(i_data_FEalures[12]), .C(n699), .D(n698), .Q(
        n700) );
  INV6 U967 ( .A(n906), .Q(n525) );
  NAND22 U968 ( .A(n1336), .B(n1331), .Q(o_addr_Erd[0]) );
  NAND22 U969 ( .A(n1336), .B(n1333), .Q(o_addr_Erd[2]) );
  NAND22 U970 ( .A(n1336), .B(n1335), .Q(o_addr_Erd[4]) );
  NAND22 U971 ( .A(n1336), .B(n1334), .Q(o_addr_Erd[3]) );
  NAND22 U972 ( .A(n1336), .B(n1332), .Q(o_addr_Erd[1]) );
  OAI311 U973 ( .A(n979), .B(n978), .C(n977), .D(n976), .Q(
        alu_o_data_AluRes[0]) );
  AOI211 U974 ( .A(n1251), .B(u_alu_N225), .C(n975), .Q(n976) );
  OAI2111 U975 ( .A(n974), .B(n114), .C(n973), .D(n972), .Q(n975) );
  IMUX20 U976 ( .A(n81), .B(alu_i_data_B[1]), .S(i_data_immext[6]), .Q(n383)
         );
  AOI211 U977 ( .A(n967), .B(n966), .C(alu_i_con_AluCtrl[2]), .Q(n977) );
  OAI2111 U978 ( .A(n1261), .B(n1196), .C(n1195), .D(n1194), .Q(
        alu_o_data_AluRes[26]) );
  AOI211 U979 ( .A(n1241), .B(u_alu_pre_sum_4b[2]), .C(n1193), .Q(n1194) );
  OAI2111 U980 ( .A(compare_i_data_rs[4]), .B(n1273), .C(n1274), .D(n1275), 
        .Q(alu_o_data_AluRes[4]) );
  IMUX20 U981 ( .A(n1266), .B(n1267), .S(alu_i_data_B[4]), .Q(n1276) );
  AOI211 U982 ( .A(alu_i_data_B[4]), .B(n98), .C(n1277), .Q(n1274) );
  NAND31 U983 ( .A(n774), .B(n773), .C(n772), .Q(n1277) );
  OAI2111 U984 ( .A(compare_i_data_rs[2]), .B(n1285), .C(n1286), .D(n1287), 
        .Q(alu_o_data_AluRes[2]) );
  IMUX20 U985 ( .A(n1266), .B(n1267), .S(u_alu_lt_x_11_B_2_), .Q(n1288) );
  AOI211 U986 ( .A(u_alu_lt_x_11_B_2_), .B(n98), .C(n1289), .Q(n1286) );
  NAND31 U987 ( .A(n794), .B(n793), .C(n792), .Q(n1289) );
  IMUX20 U988 ( .A(alu_i_data_B[4]), .B(alu_i_data_B[5]), .S(i_data_immext[6]), 
        .Q(n459) );
  IMUX20 U989 ( .A(u_alu_lt_x_11_B_2_), .B(alu_i_data_B[3]), .S(
        i_data_immext[6]), .Q(n460) );
  OAI2111 U990 ( .A(compare_i_data_rs[5]), .B(n1268), .C(n1269), .D(n1270), 
        .Q(alu_o_data_AluRes[5]) );
  AOI211 U991 ( .A(alu_i_data_B[5]), .B(n98), .C(n1272), .Q(n1269) );
  NAND31 U992 ( .A(n770), .B(n769), .C(n768), .Q(n1272) );
  OAI2111 U993 ( .A(compare_i_data_rs[3]), .B(n1278), .C(n1279), .D(n1280), 
        .Q(alu_o_data_AluRes[3]) );
  NAND31 U994 ( .A(n777), .B(n776), .C(n775), .Q(n1282) );
  OAI2111 U995 ( .A(compare_i_data_rs[1]), .B(n1299), .C(n1300), .D(n1301), 
        .Q(alu_o_data_AluRes[1]) );
  IMUX20 U996 ( .A(n1266), .B(n1267), .S(alu_i_data_B[1]), .Q(n1302) );
  AOI211 U997 ( .A(alu_i_data_B[1]), .B(n98), .C(n1303), .Q(n1300) );
  NAND31 U998 ( .A(n852), .B(n851), .C(n850), .Q(n1303) );
  IMUX20 U999 ( .A(alu_i_data_B[5]), .B(n112), .S(i_data_immext[6]), .Q(n470)
         );
  IMUX20 U1000 ( .A(alu_i_data_B[3]), .B(alu_i_data_B[4]), .S(i_data_immext[6]), .Q(n471) );
  IMUX20 U1001 ( .A(alu_i_data_B[1]), .B(u_alu_lt_x_11_B_2_), .S(
        i_data_immext[6]), .Q(n435) );
  NAND31 U1002 ( .A(n1053), .B(n1052), .C(n1051), .Q(alu_o_data_AluRes[13]) );
  AOI211 U1003 ( .A(n1064), .B(u_alu_half_sub_13_), .C(n1050), .Q(n1052) );
  OAI2111 U1004 ( .A(n1049), .B(n110), .C(n1048), .D(n1047), .Q(n1050) );
  MUX21 U1005 ( .A(n415), .B(n458), .S(i_data_immext[10]), .Q(u_alu_N238) );
  NAND31 U1006 ( .A(n1045), .B(n1044), .C(n1043), .Q(alu_o_data_AluRes[12]) );
  AOI211 U1007 ( .A(u_alu_N237), .B(n1251), .C(n1042), .Q(n1044) );
  OAI2111 U1008 ( .A(n1041), .B(n94), .C(n1040), .D(n1039), .Q(n1042) );
  NAND31 U1009 ( .A(n999), .B(n998), .C(n997), .Q(alu_o_data_AluRes[7]) );
  NAND22 U1010 ( .A(u_alu_N232), .B(n1251), .Q(n997) );
  IMUX20 U1011 ( .A(u_alu_lt_x_11_B_7_), .B(alu_i_data_B[8]), .S(
        i_data_immext[6]), .Q(n473) );
  AOI211 U1012 ( .A(n1064), .B(u_alu_half_sub_7_), .C(n996), .Q(n998) );
  OAI2111 U1013 ( .A(n995), .B(n233), .C(n994), .D(n993), .Q(n996) );
  NAND31 U1014 ( .A(n1019), .B(n1018), .C(n1017), .Q(alu_o_data_AluRes[9]) );
  IMUX20 U1015 ( .A(alu_i_data_B[9]), .B(alu_i_data_B[10]), .S(
        i_data_immext[6]), .Q(n472) );
  AOI211 U1016 ( .A(n1064), .B(u_alu_half_sub_9_), .C(n1016), .Q(n1018) );
  OAI2111 U1017 ( .A(n1015), .B(n116), .C(n1014), .D(n1013), .Q(n1016) );
  NOR21 U1018 ( .A(n378), .B(n373), .Q(u_alu_N202) );
  INV3 U1019 ( .A(n363), .Q(n373) );
  NAND31 U1020 ( .A(n989), .B(n988), .C(n987), .Q(alu_o_data_AluRes[6]) );
  IMUX20 U1021 ( .A(n112), .B(u_alu_lt_x_11_B_7_), .S(i_data_immext[6]), .Q(
        n462) );
  AOI211 U1022 ( .A(n1064), .B(u_alu_half_sub_6_), .C(n986), .Q(n988) );
  NOR21 U1023 ( .A(n378), .B(n370), .Q(u_alu_N199) );
  IMUX20 U1024 ( .A(n425), .B(n469), .S(i_data_immext[10]), .Q(u_alu_N240) );
  OAI2111 U1025 ( .A(n1261), .B(n1202), .C(n1201), .D(n1200), .Q(
        alu_o_data_AluRes[27]) );
  AOI211 U1026 ( .A(n1241), .B(u_alu_pre_sum_4b[3]), .C(n1199), .Q(n1200) );
  OAI2111 U1027 ( .A(n1261), .B(n1214), .C(n1213), .D(n1212), .Q(
        alu_o_data_AluRes[28]) );
  AOI211 U1028 ( .A(n1241), .B(u_alu_pre_sum_4b[4]), .C(n1211), .Q(n1212) );
  NAND31 U1029 ( .A(n1210), .B(n1209), .C(n1208), .Q(n1211) );
  NAND31 U1030 ( .A(n520), .B(n379), .C(n442), .Q(n457) );
  MUX21 U1031 ( .A(n332), .B(n331), .S(i_data_immext[10]), .Q(u_alu_N221) );
  NAND31 U1032 ( .A(n1118), .B(n1117), .C(n1116), .Q(alu_o_data_AluRes[19]) );
  NAND22 U1033 ( .A(n1150), .B(u_alu_pre_sum_3b[3]), .Q(n1111) );
  NOR21 U1034 ( .A(u_alu_ashr_4_SH_3_), .B(n277), .Q(n357) );
  NAND22 U1035 ( .A(n1252), .B(u_alu_pre_suba[3]), .Q(n1117) );
  NAND22 U1036 ( .A(n1258), .B(u_alu_pre_subb[3]), .Q(n1118) );
  NOR21 U1037 ( .A(u_alu_ashr_4_SH_3_), .B(n283), .Q(n358) );
  MUX21 U1038 ( .A(n289), .B(n359), .S(i_data_immext[10]), .Q(u_alu_N214) );
  NOR21 U1039 ( .A(u_alu_ashr_4_SH_3_), .B(n288), .Q(n359) );
  NAND31 U1040 ( .A(n1144), .B(n1143), .C(n1142), .Q(alu_o_data_AluRes[22]) );
  AOI211 U1041 ( .A(n1169), .B(u_alu_pre_sum_3a[6]), .C(n1141), .Q(n1142) );
  NAND22 U1042 ( .A(n1150), .B(u_alu_pre_sum_3b[6]), .Q(n1137) );
  NOR21 U1043 ( .A(u_alu_ashr_4_SH_3_), .B(n293), .Q(n360) );
  NAND22 U1044 ( .A(n1252), .B(u_alu_pre_suba[6]), .Q(n1143) );
  NAND22 U1045 ( .A(n1258), .B(u_alu_pre_subb[6]), .Q(n1144) );
  OAI2111 U1046 ( .A(n1261), .B(n1187), .C(n1186), .D(n1185), .Q(
        alu_o_data_AluRes[25]) );
  AOI211 U1047 ( .A(n1241), .B(u_alu_pre_sum_4b[1]), .C(n1184), .Q(n1185) );
  NAND41 U1048 ( .A(n1183), .B(n1182), .C(n1181), .D(n1180), .Q(n1184) );
  NOR21 U1049 ( .A(u_alu_ashr_4_SH_3_), .B(n454), .Q(n506) );
  MUX21 U1050 ( .A(n313), .B(n363), .S(i_data_immext[10]), .Q(u_alu_N218) );
  OAI2111 U1051 ( .A(n1261), .B(n97), .C(n1260), .D(n1259), .Q(
        alu_o_data_AluRes[31]) );
  AOI211 U1052 ( .A(n1258), .B(u_alu_pre_subb[15]), .C(n1257), .Q(n1259) );
  NAND31 U1053 ( .A(n450), .B(n520), .C(n379), .Q(n469) );
  IMUX20 U1054 ( .A(alu_i_data_B[31]), .B(alu_i_data_B[30]), .S(
        i_data_immext[6]), .Q(n350) );
  OAI2111 U1055 ( .A(n1261), .B(n1240), .C(n1239), .D(n1238), .Q(
        alu_o_data_AluRes[30]) );
  AOI211 U1056 ( .A(n1258), .B(u_alu_pre_subb[14]), .C(n1237), .Q(n1238) );
  NAND41 U1057 ( .A(n1236), .B(n1235), .C(n1234), .D(n1233), .Q(n1237) );
  IMUX20 U1058 ( .A(alu_i_data_B[28]), .B(alu_i_data_B[27]), .S(
        i_data_immext[6]), .Q(n341) );
  IMUX20 U1059 ( .A(alu_i_data_B[30]), .B(alu_i_data_B[29]), .S(
        i_data_immext[6]), .Q(n342) );
  INV3 U1060 ( .A(u_alu_pre_sum_4a[6]), .Q(n1240) );
  NAND31 U1061 ( .A(n447), .B(n520), .C(n379), .Q(n468) );
  NAND41 U1062 ( .A(n1028), .B(n1027), .C(n1026), .D(n1025), .Q(
        alu_o_data_AluRes[10]) );
  NOR21 U1063 ( .A(n378), .B(n374), .Q(u_alu_N203) );
  INV3 U1064 ( .A(n318), .Q(n374) );
  MUX21 U1065 ( .A(n398), .B(n455), .S(i_data_immext[10]), .Q(u_alu_N235) );
  NOR21 U1066 ( .A(u_alu_ashr_4_SH_3_), .B(n431), .Q(n455) );
  MUX21 U1067 ( .A(n399), .B(n456), .S(i_data_immext[10]), .Q(u_alu_N236) );
  NOR21 U1068 ( .A(u_alu_ashr_4_SH_3_), .B(n433), .Q(n456) );
  IMUX20 U1069 ( .A(alu_i_data_B[15]), .B(alu_i_data_B[16]), .S(
        i_data_immext[6]), .Q(n405) );
  IMUX20 U1070 ( .A(alu_i_data_B[13]), .B(alu_i_data_B[14]), .S(
        i_data_immext[6]), .Q(n406) );
  IMUX20 U1071 ( .A(alu_i_data_B[11]), .B(alu_i_data_B[12]), .S(
        i_data_immext[6]), .Q(n437) );
  OAI2111 U1072 ( .A(n1033), .B(n96), .C(n1032), .D(n1031), .Q(n1034) );
  NAND22 U1073 ( .A(n379), .B(n255), .Q(n277) );
  OAI2111 U1074 ( .A(n88), .B(n1168), .C(n1167), .D(n1166), .Q(n1172) );
  IMUX20 U1075 ( .A(n83), .B(alu_i_data_B[19]), .S(i_data_immext[6]), .Q(n290)
         );
  IMUX20 U1076 ( .A(alu_i_data_B[22]), .B(alu_i_data_B[21]), .S(
        i_data_immext[6]), .Q(n300) );
  IMUX20 U1077 ( .A(alu_i_data_B[24]), .B(alu_i_data_B[23]), .S(
        i_data_immext[6]), .Q(n314) );
  NOR21 U1078 ( .A(n378), .B(n512), .Q(u_alu_N249) );
  INV3 U1079 ( .A(u_alu_pre_sum_4a[0]), .Q(n223) );
  NOR21 U1080 ( .A(n95), .B(n1001), .Q(n1006) );
  NOR21 U1081 ( .A(u_alu_ashr_4_SH_3_), .B(n453), .Q(n502) );
  IMUX20 U1082 ( .A(alu_i_data_B[14]), .B(alu_i_data_B[15]), .S(
        i_data_immext[6]), .Q(n390) );
  IMUX20 U1083 ( .A(alu_i_data_B[12]), .B(alu_i_data_B[13]), .S(
        i_data_immext[6]), .Q(n387) );
  IMUX20 U1084 ( .A(alu_i_data_B[10]), .B(alu_i_data_B[11]), .S(
        i_data_immext[6]), .Q(n388) );
  IMUX20 U1085 ( .A(alu_i_data_B[8]), .B(alu_i_data_B[9]), .S(i_data_immext[6]), .Q(n461) );
  INV3 U1086 ( .A(n362), .Q(n372) );
  NAND22 U1087 ( .A(n1258), .B(u_alu_pre_subb[13]), .Q(n1224) );
  OAI2111 U1088 ( .A(n1261), .B(n1222), .C(n1221), .D(n1220), .Q(n1223) );
  MUX21 U1089 ( .A(n339), .B(n338), .S(i_data_immext[10]), .Q(u_alu_N222) );
  IMUX20 U1090 ( .A(alu_i_data_B[27]), .B(alu_i_data_B[26]), .S(
        i_data_immext[6]), .Q(n333) );
  IMUX20 U1091 ( .A(alu_i_data_B[29]), .B(alu_i_data_B[28]), .S(
        i_data_immext[6]), .Q(n349) );
  NOR21 U1092 ( .A(u_alu_ashr_4_SH_3_), .B(n445), .Q(n458) );
  NAND22 U1093 ( .A(n379), .B(n429), .Q(n445) );
  NAND22 U1094 ( .A(u_alu_pre_sum_4b[5]), .B(n1241), .Q(n1226) );
  INV3 U1095 ( .A(n1170), .Q(n225) );
  NAND31 U1096 ( .A(n1105), .B(n1104), .C(n1103), .Q(alu_o_data_AluRes[18]) );
  AOI211 U1097 ( .A(n1169), .B(u_alu_pre_sum_3a[2]), .C(n1102), .Q(n1103) );
  NAND41 U1098 ( .A(n1101), .B(n1100), .C(n1099), .D(n1098), .Q(n1102) );
  NAND22 U1099 ( .A(n1150), .B(u_alu_pre_sum_3b[2]), .Q(n1098) );
  NOR21 U1100 ( .A(u_alu_ashr_4_SH_3_), .B(n272), .Q(n340) );
  NAND22 U1101 ( .A(n379), .B(n251), .Q(n272) );
  IMUX20 U1102 ( .A(alu_i_data_B[18]), .B(alu_i_data_B[17]), .S(
        i_data_immext[6]), .Q(n280) );
  NOR21 U1103 ( .A(n381), .B(n397), .Q(n447) );
  NAND22 U1104 ( .A(n1252), .B(u_alu_pre_suba[2]), .Q(n1104) );
  NAND22 U1105 ( .A(n1258), .B(u_alu_pre_subb[2]), .Q(n1105) );
  NAND31 U1106 ( .A(n1158), .B(n1157), .C(n1156), .Q(alu_o_data_AluRes[23]) );
  AOI211 U1107 ( .A(n1169), .B(u_alu_pre_sum_3a[7]), .C(n1155), .Q(n1156) );
  NAND41 U1108 ( .A(n1154), .B(n1153), .C(n1152), .D(n1151), .Q(n1155) );
  NAND22 U1109 ( .A(n1150), .B(u_alu_pre_sum_3b[7]), .Q(n1151) );
  NOR21 U1110 ( .A(n381), .B(n413), .Q(n450) );
  NOR21 U1111 ( .A(u_alu_ashr_4_SH_3_), .B(n298), .Q(n361) );
  IMUX20 U1112 ( .A(alu_i_data_B[19]), .B(alu_i_data_B[18]), .S(
        i_data_immext[6]), .Q(n285) );
  IMUX20 U1113 ( .A(alu_i_data_B[21]), .B(n83), .S(i_data_immext[6]), .Q(n295)
         );
  IMUX20 U1114 ( .A(alu_i_data_B[23]), .B(alu_i_data_B[22]), .S(
        i_data_immext[6]), .Q(n307) );
  NAND22 U1115 ( .A(n1252), .B(u_alu_pre_suba[7]), .Q(n1157) );
  NAND22 U1116 ( .A(n1258), .B(u_alu_pre_subb[7]), .Q(n1158) );
  OAI2111 U1117 ( .A(n87), .B(n1075), .C(n1074), .D(n1073), .Q(n1076) );
  NAND22 U1118 ( .A(n81), .B(n382), .Q(n241) );
  IMUX20 U1119 ( .A(n112), .B(alu_i_data_B[5]), .S(i_data_immext[6]), .Q(n237)
         );
  IMUX20 U1120 ( .A(alu_i_data_B[10]), .B(alu_i_data_B[9]), .S(
        i_data_immext[6]), .Q(n236) );
  IMUX20 U1121 ( .A(alu_i_data_B[12]), .B(alu_i_data_B[11]), .S(
        i_data_immext[6]), .Q(n249) );
  IMUX20 U1122 ( .A(alu_i_data_B[14]), .B(alu_i_data_B[13]), .S(
        i_data_immext[6]), .Q(n257) );
  IMUX20 U1123 ( .A(alu_i_data_B[16]), .B(alu_i_data_B[15]), .S(
        i_data_immext[6]), .Q(n269) );
  INV3 U1124 ( .A(n1267), .Q(n1162) );
  IMUX20 U1125 ( .A(alu_i_data_B[28]), .B(alu_i_data_B[29]), .S(
        i_data_immext[6]), .Q(n395) );
  IMUX20 U1126 ( .A(alu_i_data_B[26]), .B(alu_i_data_B[27]), .S(
        i_data_immext[6]), .Q(n396) );
  IMUX20 U1127 ( .A(alu_i_data_B[22]), .B(alu_i_data_B[23]), .S(
        i_data_immext[6]), .Q(n394) );
  IMUX20 U1128 ( .A(n83), .B(alu_i_data_B[21]), .S(i_data_immext[6]), .Q(n391)
         );
  IMUX20 U1129 ( .A(alu_i_data_B[18]), .B(alu_i_data_B[19]), .S(
        i_data_immext[6]), .Q(n392) );
  IMUX20 U1130 ( .A(alu_i_data_B[16]), .B(alu_i_data_B[17]), .S(
        i_data_immext[6]), .Q(n389) );
  NOR31 U1131 ( .A(i_con_bop[2]), .B(n953), .C(n954), .Q(n958) );
  NAND22 U1132 ( .A(n811), .B(n810), .Q(compare_i_data_rs[27]) );
  NOR21 U1133 ( .A(n805), .B(n120), .Q(n809) );
  NAND22 U1134 ( .A(n118), .B(i_data_rs[27]), .Q(n811) );
  NAND22 U1135 ( .A(n825), .B(n824), .Q(compare_i_data_rs[25]) );
  NOR21 U1136 ( .A(n819), .B(n120), .Q(n823) );
  NAND22 U1137 ( .A(n118), .B(i_data_rs[25]), .Q(n825) );
  NAND41 U1138 ( .A(n940), .B(n939), .C(n938), .D(n937), .Q(n946) );
  NOR21 U1139 ( .A(n812), .B(n120), .Q(n816) );
  NAND22 U1140 ( .A(n118), .B(i_data_rs[30]), .Q(n791) );
  NAND22 U1141 ( .A(n896), .B(n895), .Q(compare_i_data_rs[24]) );
  NOR21 U1142 ( .A(n890), .B(n120), .Q(n894) );
  NAND22 U1143 ( .A(n118), .B(i_data_rs[24]), .Q(n896) );
  NAND41 U1144 ( .A(n936), .B(n935), .C(n934), .D(n933), .Q(n947) );
  NAND22 U1145 ( .A(n804), .B(n803), .Q(compare_i_data_rs[28]) );
  NOR21 U1146 ( .A(n798), .B(n120), .Q(n802) );
  NOR21 U1147 ( .A(n860), .B(n120), .Q(n864) );
  NAND22 U1148 ( .A(n118), .B(i_data_rs[18]), .Q(n866) );
  NAND41 U1149 ( .A(n932), .B(n931), .C(n930), .D(n929), .Q(n948) );
  NOR21 U1150 ( .A(n853), .B(n120), .Q(n857) );
  NAND22 U1151 ( .A(n118), .B(i_data_rs[19]), .Q(n859) );
  NAND22 U1152 ( .A(n832), .B(n831), .Q(compare_i_data_rs[23]) );
  NOR21 U1153 ( .A(n826), .B(n120), .Q(n830) );
  NAND22 U1154 ( .A(n118), .B(i_data_rs[23]), .Q(n832) );
  NAND41 U1155 ( .A(n924), .B(n923), .C(n922), .D(n921), .Q(n925) );
  NAND22 U1156 ( .A(n839), .B(n838), .Q(compare_i_data_rs[22]) );
  NOR21 U1157 ( .A(n833), .B(n120), .Q(n837) );
  NAND22 U1158 ( .A(n118), .B(i_data_rs[22]), .Q(n839) );
  NAND22 U1159 ( .A(n849), .B(n848), .Q(compare_i_data_rs[20]) );
  NOR21 U1160 ( .A(n843), .B(n120), .Q(n847) );
  NAND22 U1161 ( .A(n118), .B(i_data_rs[20]), .Q(n849) );
  NAND41 U1162 ( .A(n920), .B(n919), .C(n918), .D(n917), .Q(n926) );
  NAND41 U1163 ( .A(n916), .B(n915), .C(n914), .D(n913), .Q(n927) );
  NAND41 U1164 ( .A(n912), .B(n911), .C(n910), .D(n909), .Q(n928) );
  NOR21 U1165 ( .A(n778), .B(n119), .Q(n782) );
  NAND31 U1166 ( .A(n1091), .B(n1090), .C(n1089), .Q(alu_o_data_AluRes[17]) );
  NAND22 U1167 ( .A(n1150), .B(u_alu_pre_sum_3b[1]), .Q(n1084) );
  NOR21 U1168 ( .A(u_alu_ashr_4_SH_3_), .B(n311), .Q(n279) );
  NAND22 U1169 ( .A(n267), .B(n379), .Q(n311) );
  INV3 U1170 ( .A(i_data_immext[8]), .Q(n379) );
  NOR21 U1171 ( .A(n381), .B(n248), .Q(n267) );
  IMUX20 U1172 ( .A(alu_i_data_B[1]), .B(n81), .S(i_data_immext[6]), .Q(n248)
         );
  IMUX20 U1173 ( .A(u_alu_lt_x_11_B_7_), .B(n112), .S(i_data_immext[6]), .Q(
        n244) );
  IMUX20 U1174 ( .A(alu_i_data_B[11]), .B(alu_i_data_B[10]), .S(
        i_data_immext[6]), .Q(n243) );
  IMUX20 U1175 ( .A(alu_i_data_B[13]), .B(alu_i_data_B[12]), .S(
        i_data_immext[6]), .Q(n253) );
  IMUX20 U1176 ( .A(alu_i_data_B[15]), .B(alu_i_data_B[14]), .S(
        i_data_immext[6]), .Q(n263) );
  IMUX20 U1177 ( .A(alu_i_data_B[17]), .B(alu_i_data_B[16]), .S(
        i_data_immext[6]), .Q(n274) );
  NAND22 U1178 ( .A(alu_i_data_B[31]), .B(n382), .Q(n413) );
  NAND22 U1179 ( .A(n563), .B(n624), .Q(alu_i_data_B[31]) );
  IMUX20 U1180 ( .A(alu_i_data_B[29]), .B(alu_i_data_B[30]), .S(
        i_data_immext[6]), .Q(n414) );
  NAND22 U1181 ( .A(n567), .B(n624), .Q(alu_i_data_B[30]) );
  NAND31 U1182 ( .A(n566), .B(n565), .C(n564), .Q(compare_i_data_rt[30]) );
  NAND22 U1183 ( .A(n571), .B(n624), .Q(alu_i_data_B[29]) );
  NAND31 U1184 ( .A(n570), .B(n569), .C(n568), .Q(compare_i_data_rt[29]) );
  IMUX20 U1185 ( .A(alu_i_data_B[27]), .B(alu_i_data_B[28]), .S(
        i_data_immext[6]), .Q(n411) );
  NAND22 U1186 ( .A(n575), .B(n624), .Q(alu_i_data_B[28]) );
  NAND31 U1187 ( .A(n574), .B(n573), .C(n572), .Q(compare_i_data_rt[28]) );
  NAND22 U1188 ( .A(n579), .B(n624), .Q(alu_i_data_B[27]) );
  NAND31 U1189 ( .A(n578), .B(n577), .C(n576), .Q(compare_i_data_rt[27]) );
  NAND22 U1190 ( .A(n583), .B(n624), .Q(alu_i_data_B[26]) );
  NAND31 U1191 ( .A(n582), .B(n581), .C(n580), .Q(compare_i_data_rt[26]) );
  NAND31 U1192 ( .A(n586), .B(n585), .C(n584), .Q(compare_i_data_rt[25]) );
  INV3 U1193 ( .A(u_alu_ashr_4_SH_1_), .Q(n380) );
  IMUX20 U1194 ( .A(alu_i_data_B[23]), .B(alu_i_data_B[24]), .S(
        i_data_immext[6]), .Q(n409) );
  NAND22 U1195 ( .A(n591), .B(n624), .Q(alu_i_data_B[24]) );
  NAND31 U1196 ( .A(n590), .B(n589), .C(n588), .Q(compare_i_data_rt[24]) );
  NAND22 U1197 ( .A(n595), .B(n624), .Q(alu_i_data_B[23]) );
  NAND31 U1198 ( .A(n594), .B(n593), .C(n592), .Q(compare_i_data_rt[23]) );
  IMUX20 U1199 ( .A(alu_i_data_B[21]), .B(alu_i_data_B[22]), .S(
        i_data_immext[6]), .Q(n410) );
  NAND31 U1200 ( .A(n598), .B(n597), .C(n596), .Q(compare_i_data_rt[22]) );
  IMUX20 U1201 ( .A(alu_i_data_B[19]), .B(n83), .S(i_data_immext[6]), .Q(n407)
         );
  NAND22 U1202 ( .A(n607), .B(n624), .Q(alu_i_data_B[20]) );
  NAND31 U1203 ( .A(n610), .B(n609), .C(n608), .Q(compare_i_data_rt[19]) );
  NAND22 U1204 ( .A(n230), .B(i_data_rt[19]), .Q(n610) );
  IMUX20 U1205 ( .A(alu_i_data_B[17]), .B(alu_i_data_B[18]), .S(
        i_data_immext[6]), .Q(n408) );
  NAND31 U1206 ( .A(n614), .B(n613), .C(n612), .Q(compare_i_data_rt[18]) );
  NAND22 U1207 ( .A(n230), .B(i_data_rt[18]), .Q(n614) );
  NAND22 U1208 ( .A(alu_i_con_AluCtrl[3]), .B(n766), .Q(n1069) );
  NAND22 U1209 ( .A(u_alu_add_x_1_n20), .B(u_alu_add_x_1_n12), .Q(
        u_alu_add_x_1_n10) );
  NAND22 U1210 ( .A(n1252), .B(u_alu_pre_suba[1]), .Q(n1090) );
  NAND22 U1211 ( .A(n1258), .B(u_alu_pre_subb[1]), .Q(n1091) );
  NAND22 U1212 ( .A(n229), .B(i_data_rt[17]), .Q(n618) );
  NOR21 U1213 ( .A(n867), .B(n120), .Q(n871) );
  NAND22 U1214 ( .A(n118), .B(i_data_rs[17]), .Q(n873) );
  NOR21 U1215 ( .A(n899), .B(n120), .Q(n905) );
  NAND22 U1216 ( .A(n118), .B(i_data_rs[16]), .Q(n908) );
  NAND22 U1217 ( .A(n963), .B(n765), .Q(n1063) );
  OAI2112 U1218 ( .A(n1315), .B(n1322), .C(n1327), .D(n1314), .Q(
        alu_i_con_AluCtrl[0]) );
  OAI212 U1219 ( .A(i_data_immext[0]), .B(n880), .C(n1262), .Q(n888) );
  NOR21 U1220 ( .A(n879), .B(n889), .Q(n880) );
  NOR31 U1221 ( .A(n877), .B(n875), .C(n876), .Q(n889) );
  OAI212 U1222 ( .A(n1322), .B(n541), .C(n1321), .Q(n544) );
  NAND22 U1223 ( .A(n874), .B(i_data_immext[1]), .Q(n876) );
  NAND22 U1224 ( .A(i_data_immext[5]), .B(n1307), .Q(n1308) );
  AOI211 U1225 ( .A(i_con_Ealuop[1]), .B(n1310), .C(n1328), .Q(n1320) );
  NAND22 U1226 ( .A(n875), .B(i_data_immext[5]), .Q(n538) );
  NAND22 U1227 ( .A(n230), .B(i_data_rt[13]), .Q(n636) );
  NAND22 U1228 ( .A(n694), .B(n693), .Q(compare_i_data_rs[13]) );
  NOR21 U1229 ( .A(n688), .B(n120), .Q(n692) );
  NAND22 U1230 ( .A(n118), .B(i_data_rs[13]), .Q(n694) );
  NAND22 U1231 ( .A(n230), .B(i_data_rt[10]), .Q(n645) );
  NOR21 U1232 ( .A(n709), .B(n120), .Q(n713) );
  NAND22 U1233 ( .A(n118), .B(i_data_rs[10]), .Q(n715) );
  NOR21 U1234 ( .A(n716), .B(n120), .Q(n720) );
  NAND22 U1235 ( .A(n118), .B(i_data_rs[9]), .Q(n722) );
  NOR21 U1236 ( .A(n723), .B(n120), .Q(n727) );
  NAND22 U1237 ( .A(n118), .B(i_data_rs[8]), .Q(n729) );
  NAND22 U1238 ( .A(n708), .B(n707), .Q(compare_i_data_rs[11]) );
  NOR21 U1239 ( .A(n702), .B(n120), .Q(n706) );
  NAND22 U1240 ( .A(n118), .B(i_data_rs[11]), .Q(n708) );
  INV3 U1241 ( .A(alu_i_data_B[3]), .Q(n234) );
  NAND22 U1242 ( .A(n230), .B(i_data_rt[3]), .Q(n663) );
  NAND22 U1243 ( .A(n118), .B(i_data_rs[3]), .Q(n749) );
  NAND22 U1244 ( .A(n230), .B(i_data_rt[1]), .Q(n669) );
  NAND22 U1245 ( .A(n118), .B(i_data_rs[1]), .Q(n755) );
  MUX22 U1246 ( .A(compare_i_data_rt[0]), .B(i_data_immext[0]), .S(n235), .Q(
        alu_i_data_B[0]) );
  NAND22 U1247 ( .A(n762), .B(n761), .Q(compare_i_data_rs[0]) );
  INV3 U1248 ( .A(n233), .Q(u_alu_lt_x_11_B_7_) );
  INV3 U1249 ( .A(alu_i_data_B[7]), .Q(n233) );
  NAND31 U1250 ( .A(n654), .B(n653), .C(n652), .Q(compare_i_data_rt[7]) );
  NAND22 U1251 ( .A(n118), .B(i_data_rs[7]), .Q(n736) );
  NOR21 U1252 ( .A(n737), .B(n120), .Q(n741) );
  NAND22 U1253 ( .A(n118), .B(i_data_rs[6]), .Q(n743) );
  INV3 U1254 ( .A(alu_i_data_B[5]), .Q(n232) );
  NAND22 U1255 ( .A(n118), .B(i_data_rs[4]), .Q(n746) );
  MUX22 U1256 ( .A(compare_i_data_rt[12]), .B(i_data_immext[12]), .S(n235), 
        .Q(alu_i_data_B[12]) );
  NAND31 U1257 ( .A(n639), .B(n638), .C(n637), .Q(compare_i_data_rt[12]) );
  NAND22 U1258 ( .A(n701), .B(n700), .Q(compare_i_data_rs[12]) );
  NOR21 U1259 ( .A(n695), .B(n120), .Q(n699) );
  NAND22 U1260 ( .A(n118), .B(i_data_rs[12]), .Q(n701) );
  NAND31 U1261 ( .A(n633), .B(n632), .C(n631), .Q(compare_i_data_rt[14]) );
  NAND22 U1262 ( .A(n687), .B(n686), .Q(compare_i_data_rs[14]) );
  AOI2111 U1263 ( .A(n121), .B(i_data_FEalures[14]), .C(n685), .D(n684), .Q(
        n686) );
  NOR21 U1264 ( .A(n681), .B(n120), .Q(n685) );
  NAND22 U1265 ( .A(n118), .B(i_data_rs[14]), .Q(n687) );
  AOI211 U1266 ( .A(n118), .B(i_data_rs[15]), .C(n679), .Q(n680) );
  NAND22 U1267 ( .A(n678), .B(n677), .Q(n679) );
  NAND22 U1268 ( .A(n530), .B(n534), .Q(n898) );
  NOR21 U1269 ( .A(n227), .B(i_con_Efamux[2]), .Q(n530) );
  NAND22 U1270 ( .A(n534), .B(n533), .Q(n902) );
  INV3 U1271 ( .A(n532), .Q(n533) );
  NAND22 U1272 ( .A(i_con_Efamux[2]), .B(i_con_Efamux[0]), .Q(n532) );
  AOI211 U1273 ( .A(n229), .B(i_data_rt[15]), .C(n628), .Q(n629) );
  NAND22 U1274 ( .A(n627), .B(n626), .Q(n628) );
  IMUX20 U1275 ( .A(n383), .B(n460), .S(u_alu_ashr_4_SH_1_), .Q(n384) );
  IMUX20 U1276 ( .A(n483), .B(n482), .S(n378), .Q(u_alu_N229) );
  MUX21 U1277 ( .A(n467), .B(n466), .S(n378), .Q(u_alu_N227) );
  IMUX20 U1278 ( .A(n460), .B(n459), .S(u_alu_ashr_4_SH_1_), .Q(n463) );
  MUX21 U1279 ( .A(n489), .B(n488), .S(n378), .Q(u_alu_N230) );
  MUX21 U1280 ( .A(n478), .B(n477), .S(n378), .Q(u_alu_N228) );
  IMUX20 U1281 ( .A(n471), .B(n470), .S(n381), .Q(n474) );
  MUX21 U1282 ( .A(n441), .B(n440), .S(n378), .Q(u_alu_N226) );
  IMUX20 U1283 ( .A(n435), .B(n471), .S(n381), .Q(n436) );
  IMUX20 U1284 ( .A(n341), .B(n326), .S(n381), .Q(n328) );
  MUX21 U1285 ( .A(n278), .B(n357), .S(n378), .Q(u_alu_N212) );
  MUX21 U1286 ( .A(n284), .B(n358), .S(n378), .Q(u_alu_N213) );
  MUX21 U1287 ( .A(n294), .B(n360), .S(n378), .Q(u_alu_N215) );
  MUX21 U1288 ( .A(n356), .B(n355), .S(n378), .Q(u_alu_N224) );
  IMUX20 U1289 ( .A(n350), .B(n349), .S(n381), .Q(n352) );
  MUX21 U1290 ( .A(n348), .B(n347), .S(n378), .Q(u_alu_N223) );
  IMUX20 U1291 ( .A(n342), .B(n341), .S(u_alu_ashr_4_SH_1_), .Q(n344) );
  IMUX20 U1292 ( .A(n405), .B(n408), .S(u_alu_ashr_4_SH_1_), .Q(n422) );
  MUX21 U1293 ( .A(n306), .B(n362), .S(n378), .Q(u_alu_N217) );
  IMUX20 U1294 ( .A(n349), .B(n333), .S(n381), .Q(n335) );
  MUX21 U1295 ( .A(n273), .B(n340), .S(n378), .Q(u_alu_N211) );
  MUX21 U1296 ( .A(n299), .B(n361), .S(n378), .Q(u_alu_N216) );
  MUX21 U1297 ( .A(n262), .B(n261), .S(n378), .Q(u_alu_N209) );
  MUX21 U1298 ( .A(n268), .B(n279), .S(n378), .Q(u_alu_N210) );
  IMUX20 U1299 ( .A(n274), .B(n263), .S(u_alu_ashr_4_SH_1_), .Q(n286) );
  IMUX20 U1300 ( .A(n408), .B(n407), .S(u_alu_ashr_4_SH_1_), .Q(n428) );
  NAND22 U1301 ( .A(n963), .B(n1068), .Q(n1066) );
  NOR21 U1302 ( .A(alu_i_con_AluCtrl[2]), .B(alu_i_con_AluCtrl[0]), .Q(n1068)
         );
  NAND22 U1303 ( .A(u_alu_half_sub_16_), .B(n1064), .Q(n1065) );
  NAND22 U1304 ( .A(n978), .B(alu_i_con_AluCtrl[2]), .Q(n771) );
  INV3 U1305 ( .A(i_data_immext[5]), .Q(n877) );
  INV3 U1306 ( .A(i_data_immext[3]), .Q(n874) );
  INV3 U1307 ( .A(i_data_immext[2]), .Q(n875) );
  INV3 U1308 ( .A(n1325), .Q(n1322) );
  NOR21 U1309 ( .A(n549), .B(i_con_Efbmux[2]), .Q(n550) );
  BUF6 U1310 ( .A(n228), .Q(n229) );
  NAND22 U1311 ( .A(i_con_Efbmux[2]), .B(i_con_Efbmux[0]), .Q(n552) );
  OAI310 U1312 ( .A(n81), .B(n1247), .C(compare_i_data_rs[0]), .D(n969), .Q(
        n970) );
  AOI220 U1313 ( .A(n1064), .B(u_alu_half_sub_0_), .C(n1159), .D(
        u_alu_sum_1_0_), .Q(n969) );
  OAI210 U1314 ( .A(n81), .B(n1266), .C(n526), .Q(n971) );
  NAND20 U1315 ( .A(u_alu_N193), .B(n1250), .Q(n973) );
  AOI2110 U1316 ( .A(n1162), .B(compare_i_data_rs[0]), .C(n968), .D(n98), .Q(
        n974) );
  NOR20 U1317 ( .A(compare_i_data_rs[0]), .B(n1266), .Q(n968) );
  NAND20 U1318 ( .A(n1264), .B(n1190), .Q(n1191) );
  XNR21 U1319 ( .A(n1189), .B(alu_i_data_B[26]), .Q(n1190) );
  INV0 U1320 ( .A(compare_i_data_rs[26]), .Q(n1189) );
  OAI310 U1321 ( .A(n85), .B(n1293), .C(n1267), .D(n1188), .Q(n1192) );
  NAND20 U1322 ( .A(n1242), .B(alu_i_data_B[10]), .Q(n1188) );
  AOI220 U1323 ( .A(n1159), .B(u_alu_sum_1_4_), .C(u_alu_half_sub_4_), .D(
        n1064), .Q(n773) );
  AOI220 U1324 ( .A(n1159), .B(u_alu_sum_1_2_), .C(u_alu_half_sub_2_), .D(
        n1064), .Q(n793) );
  AOI220 U1325 ( .A(n1159), .B(u_alu_sum_1_3_), .C(u_alu_half_sub_3_), .D(
        n1064), .Q(n776) );
  AOI220 U1326 ( .A(n1064), .B(u_alu_half_sub_1_), .C(n1159), .D(
        u_alu_sum_1_1_), .Q(n851) );
  NAND20 U1327 ( .A(u_alu_N238), .B(n1251), .Q(n1048) );
  AOI2110 U1328 ( .A(n1162), .B(compare_i_data_rs[13]), .C(n1046), .D(n98), 
        .Q(n1049) );
  NOR20 U1329 ( .A(compare_i_data_rs[13]), .B(n1266), .Q(n1046) );
  NAND20 U1330 ( .A(u_alu_half_sub_12_), .B(n1064), .Q(n1040) );
  AOI2110 U1331 ( .A(n1162), .B(compare_i_data_rs[12]), .C(n1038), .D(n98), 
        .Q(n1041) );
  NOR20 U1332 ( .A(compare_i_data_rs[12]), .B(n1266), .Q(n1038) );
  OAI210 U1333 ( .A(u_alu_lt_x_11_B_7_), .B(n1266), .C(n526), .Q(n992) );
  AOI2110 U1334 ( .A(n1162), .B(compare_i_data_rs[7]), .C(n990), .D(n98), .Q(
        n995) );
  NOR20 U1335 ( .A(compare_i_data_rs[7]), .B(n1266), .Q(n990) );
  NOR30 U1336 ( .A(alu_i_data_B[9]), .B(compare_i_data_rs[9]), .C(n1247), .Q(
        n1011) );
  OAI210 U1337 ( .A(alu_i_data_B[9]), .B(n1266), .C(n526), .Q(n1012) );
  NAND20 U1338 ( .A(u_alu_N166), .B(n1159), .Q(n1014) );
  AOI2110 U1339 ( .A(n1162), .B(compare_i_data_rs[9]), .C(n1010), .D(n98), .Q(
        n1015) );
  NOR20 U1340 ( .A(compare_i_data_rs[9]), .B(n1266), .Q(n1010) );
  NOR30 U1341 ( .A(n112), .B(compare_i_data_rs[6]), .C(n1247), .Q(n981) );
  OAI210 U1342 ( .A(n112), .B(n1266), .C(n526), .Q(n982) );
  AOI2110 U1343 ( .A(n1162), .B(compare_i_data_rs[6]), .C(n980), .D(n98), .Q(
        n985) );
  NOR20 U1344 ( .A(compare_i_data_rs[6]), .B(n1266), .Q(n980) );
  NAND20 U1345 ( .A(u_alu_N240), .B(n1251), .Q(n1061) );
  AOI2110 U1346 ( .A(n1162), .B(n80), .C(n1059), .D(n98), .Q(n1062) );
  NOR20 U1347 ( .A(n80), .B(n1266), .Q(n1059) );
  NAND20 U1348 ( .A(n1242), .B(alu_i_data_B[11]), .Q(n1197) );
  NAND20 U1349 ( .A(u_alu_N253), .B(n1251), .Q(n1208) );
  AOI2110 U1350 ( .A(n98), .B(compare_i_data_rs[28]), .C(n1207), .D(n1206), 
        .Q(n1209) );
  OAI310 U1351 ( .A(compare_i_data_rs[28]), .B(alu_i_data_B[28]), .C(n1247), 
        .D(n1205), .Q(n1206) );
  NAND20 U1352 ( .A(n1264), .B(n1204), .Q(n1205) );
  XNR21 U1353 ( .A(n106), .B(alu_i_data_B[28]), .Q(n1204) );
  OAI310 U1354 ( .A(n113), .B(n1291), .C(n1267), .D(n1203), .Q(n1207) );
  NAND20 U1355 ( .A(n1242), .B(alu_i_data_B[12]), .Q(n1203) );
  AOI2110 U1356 ( .A(n98), .B(compare_i_data_rs[19]), .C(n1110), .D(n1109), 
        .Q(n1114) );
  OAI310 U1357 ( .A(compare_i_data_rs[19]), .B(alu_i_data_B[19]), .C(n1247), 
        .D(n1108), .Q(n1109) );
  NAND20 U1358 ( .A(n1264), .B(n1107), .Q(n1108) );
  XNR21 U1359 ( .A(n101), .B(alu_i_data_B[19]), .Q(n1107) );
  OAI310 U1360 ( .A(n105), .B(n1304), .C(n1267), .D(n1106), .Q(n1110) );
  OAI310 U1361 ( .A(compare_i_data_rs[20]), .B(n83), .C(n1247), .D(n1121), .Q(
        n1122) );
  NAND20 U1362 ( .A(n1264), .B(n1120), .Q(n1121) );
  XNR21 U1363 ( .A(n103), .B(n83), .Q(n1120) );
  OAI310 U1364 ( .A(n82), .B(n1298), .C(n1267), .D(n1119), .Q(n1123) );
  NAND20 U1365 ( .A(n1242), .B(alu_i_data_B[4]), .Q(n1119) );
  OAI310 U1366 ( .A(compare_i_data_rs[21]), .B(alu_i_data_B[21]), .C(n1247), 
        .D(n1128), .Q(n1129) );
  NAND20 U1367 ( .A(n1264), .B(n1127), .Q(n1128) );
  INV0 U1368 ( .A(compare_i_data_rs[21]), .Q(n1126) );
  OAI310 U1369 ( .A(n92), .B(n1297), .C(n1267), .D(n1125), .Q(n1130) );
  NAND20 U1370 ( .A(n1242), .B(alu_i_data_B[5]), .Q(n1125) );
  AOI2110 U1371 ( .A(n98), .B(compare_i_data_rs[22]), .C(n1136), .D(n1135), 
        .Q(n1140) );
  OAI310 U1372 ( .A(compare_i_data_rs[22]), .B(alu_i_data_B[22]), .C(n1247), 
        .D(n1134), .Q(n1135) );
  NAND20 U1373 ( .A(n1264), .B(n1133), .Q(n1134) );
  XNR21 U1374 ( .A(n100), .B(alu_i_data_B[22]), .Q(n1133) );
  OAI310 U1375 ( .A(n99), .B(n1296), .C(n1267), .D(n1132), .Q(n1136) );
  NAND20 U1376 ( .A(u_alu_N250), .B(n1251), .Q(n1180) );
  NOR20 U1377 ( .A(n1294), .B(n1267), .Q(n1178) );
  NOR20 U1378 ( .A(compare_i_data_rs[25]), .B(n1247), .Q(n1179) );
  AOI210 U1379 ( .A(n98), .B(compare_i_data_rs[25]), .C(n1177), .Q(n1183) );
  OAI220 U1380 ( .A(n1176), .B(n116), .C(n1266), .D(n1175), .Q(n1177) );
  XNR21 U1381 ( .A(compare_i_data_rs[25]), .B(alu_i_data_B[25]), .Q(n1175) );
  NAND20 U1382 ( .A(u_alu_N256), .B(n1251), .Q(n1254) );
  AOI2110 U1383 ( .A(n98), .B(compare_i_data_rs[31]), .C(n1249), .D(n1248), 
        .Q(n1256) );
  OAI310 U1384 ( .A(compare_i_data_rs[31]), .B(alu_i_data_B[31]), .C(n1247), 
        .D(n1246), .Q(n1248) );
  NAND20 U1385 ( .A(n1264), .B(n1245), .Q(n1246) );
  XNR21 U1386 ( .A(n91), .B(alu_i_data_B[31]), .Q(n1245) );
  OAI310 U1387 ( .A(n1244), .B(n1283), .C(n1267), .D(n1243), .Q(n1249) );
  NAND20 U1388 ( .A(n1242), .B(alu_i_data_B[15]), .Q(n1243) );
  NAND20 U1389 ( .A(u_alu_N255), .B(n1251), .Q(n1234) );
  AOI2110 U1390 ( .A(n98), .B(compare_i_data_rs[30]), .C(n1232), .D(n1231), 
        .Q(n1236) );
  OAI310 U1391 ( .A(compare_i_data_rs[30]), .B(alu_i_data_B[30]), .C(n1247), 
        .D(n1230), .Q(n1231) );
  NAND20 U1392 ( .A(n1264), .B(n1229), .Q(n1230) );
  INV0 U1393 ( .A(compare_i_data_rs[30]), .Q(n1228) );
  OAI310 U1394 ( .A(n89), .B(n1284), .C(n1267), .D(n1227), .Q(n1232) );
  NAND20 U1395 ( .A(n1242), .B(alu_i_data_B[14]), .Q(n1227) );
  OAI310 U1396 ( .A(alu_i_data_B[14]), .B(n1247), .C(compare_i_data_rs[14]), 
        .D(n1056), .Q(n1057) );
  NAND20 U1397 ( .A(n1055), .B(compare_i_data_rs[14]), .Q(n1056) );
  OAI210 U1398 ( .A(alu_i_data_B[14]), .B(n1266), .C(n526), .Q(n1055) );
  OAI210 U1399 ( .A(n1266), .B(compare_i_data_rs[14]), .C(n1054), .Q(n1058) );
  AOI210 U1400 ( .A(n1162), .B(compare_i_data_rs[14]), .C(n98), .Q(n1054) );
  OAI210 U1401 ( .A(alu_i_data_B[10]), .B(n1266), .C(n526), .Q(n1021) );
  AOI210 U1402 ( .A(n1162), .B(compare_i_data_rs[10]), .C(n98), .Q(n1020) );
  NAND30 U1403 ( .A(n1263), .B(n102), .C(n96), .Q(n1031) );
  OAI210 U1404 ( .A(n1030), .B(n98), .C(compare_i_data_rs[11]), .Q(n1032) );
  NOR20 U1405 ( .A(alu_i_data_B[11]), .B(n1266), .Q(n1030) );
  AOI2110 U1406 ( .A(n1264), .B(n102), .C(n1029), .D(n98), .Q(n1033) );
  NOR20 U1407 ( .A(n102), .B(n1267), .Q(n1029) );
  NAND20 U1408 ( .A(n1242), .B(alu_i_data_B[8]), .Q(n1163) );
  OAI210 U1409 ( .A(n1266), .B(alu_i_data_B[24]), .C(n526), .Q(n1165) );
  NOR20 U1410 ( .A(compare_i_data_rs[24]), .B(n1266), .Q(n1161) );
  AOI210 U1411 ( .A(n1264), .B(n95), .C(n98), .Q(n1004) );
  AOI2110 U1412 ( .A(n1264), .B(n1003), .C(n1000), .D(n98), .Q(n1001) );
  NOR20 U1413 ( .A(n1003), .B(n1267), .Q(n1000) );
  INV0 U1414 ( .A(compare_i_data_rs[29]), .Q(n1217) );
  AOI210 U1415 ( .A(n98), .B(compare_i_data_rs[29]), .C(n1216), .Q(n1219) );
  OAI310 U1416 ( .A(n90), .B(n1290), .C(n1267), .D(n1215), .Q(n1216) );
  NAND20 U1417 ( .A(n1242), .B(alu_i_data_B[13]), .Q(n1215) );
  OAI310 U1418 ( .A(compare_i_data_rs[18]), .B(alu_i_data_B[18]), .C(n1247), 
        .D(n1095), .Q(n1096) );
  NAND20 U1419 ( .A(n1264), .B(n1094), .Q(n1095) );
  INV0 U1420 ( .A(compare_i_data_rs[18]), .Q(n1093) );
  NAND20 U1421 ( .A(n1242), .B(u_alu_lt_x_11_B_2_), .Q(n1092) );
  OAI310 U1422 ( .A(compare_i_data_rs[23]), .B(alu_i_data_B[23]), .C(n1247), 
        .D(n1147), .Q(n1148) );
  NAND20 U1423 ( .A(n1264), .B(n1146), .Q(n1147) );
  XNR21 U1424 ( .A(n104), .B(alu_i_data_B[23]), .Q(n1146) );
  NAND20 U1425 ( .A(n1242), .B(n81), .Q(n1070) );
  OAI210 U1426 ( .A(n1266), .B(alu_i_data_B[16]), .C(n526), .Q(n1072) );
  NAND20 U1427 ( .A(u_alu_N209), .B(n1250), .Q(n1074) );
  NOR20 U1428 ( .A(compare_i_data_rs[16]), .B(n1266), .Q(n1067) );
  XNR21 U1429 ( .A(compare_i_data_rt[15]), .B(n80), .Q(n941) );
  XNR21 U1430 ( .A(compare_i_data_rs[27]), .B(compare_i_data_rt[27]), .Q(n942)
         );
  NAND20 U1431 ( .A(n122), .B(i_data_FMmemout[27]), .Q(n806) );
  INV0 U1432 ( .A(i_data_FMalures[27]), .Q(n805) );
  XNR21 U1433 ( .A(compare_i_data_rt[31]), .B(compare_i_data_rs[31]), .Q(n943)
         );
  XNR21 U1434 ( .A(compare_i_data_rs[25]), .B(compare_i_data_rt[25]), .Q(n944)
         );
  NAND20 U1435 ( .A(n122), .B(i_data_FMmemout[25]), .Q(n820) );
  INV0 U1436 ( .A(i_data_FMalures[25]), .Q(n819) );
  XNR21 U1437 ( .A(compare_i_data_rs[26]), .B(compare_i_data_rt[26]), .Q(n937)
         );
  NAND20 U1438 ( .A(n122), .B(i_data_FMmemout[26]), .Q(n813) );
  INV0 U1439 ( .A(i_data_FMalures[26]), .Q(n812) );
  XNR21 U1440 ( .A(compare_i_data_rs[30]), .B(compare_i_data_rt[30]), .Q(n938)
         );
  NAND20 U1441 ( .A(n122), .B(i_data_FMmemout[30]), .Q(n786) );
  INV0 U1442 ( .A(i_data_FMalures[30]), .Q(n785) );
  NAND20 U1443 ( .A(n122), .B(i_data_FMmemout[24]), .Q(n891) );
  INV0 U1444 ( .A(i_data_FMalures[24]), .Q(n890) );
  XNR21 U1445 ( .A(compare_i_data_rs[29]), .B(compare_i_data_rt[29]), .Q(n940)
         );
  NAND20 U1446 ( .A(n122), .B(i_data_FMmemout[29]), .Q(n796) );
  INV0 U1447 ( .A(i_data_FMalures[29]), .Q(n795) );
  XNR21 U1448 ( .A(compare_i_data_rt[2]), .B(compare_i_data_rs[2]), .Q(n933)
         );
  XNR21 U1449 ( .A(compare_i_data_rs[28]), .B(compare_i_data_rt[28]), .Q(n935)
         );
  NAND20 U1450 ( .A(n122), .B(i_data_FMmemout[28]), .Q(n799) );
  INV0 U1451 ( .A(i_data_FMalures[28]), .Q(n798) );
  XNR21 U1452 ( .A(compare_i_data_rs[18]), .B(compare_i_data_rt[18]), .Q(n936)
         );
  INV0 U1453 ( .A(i_data_FMalures[18]), .Q(n860) );
  XNR21 U1454 ( .A(compare_i_data_rs[19]), .B(compare_i_data_rt[19]), .Q(n929)
         );
  INV0 U1455 ( .A(i_data_FMalures[19]), .Q(n853) );
  XNR21 U1456 ( .A(compare_i_data_rs[23]), .B(compare_i_data_rt[23]), .Q(n930)
         );
  NAND20 U1457 ( .A(n122), .B(i_data_FMmemout[23]), .Q(n827) );
  INV0 U1458 ( .A(i_data_FMalures[23]), .Q(n826) );
  XNR21 U1459 ( .A(compare_i_data_rs[21]), .B(compare_i_data_rt[21]), .Q(n932)
         );
  INV0 U1460 ( .A(i_data_FMalures[21]), .Q(n840) );
  XNR21 U1461 ( .A(compare_i_data_rs[22]), .B(compare_i_data_rt[22]), .Q(n921)
         );
  NAND20 U1462 ( .A(n122), .B(i_data_FMmemout[22]), .Q(n834) );
  INV0 U1463 ( .A(i_data_FMalures[22]), .Q(n833) );
  XNR21 U1464 ( .A(compare_i_data_rs[20]), .B(compare_i_data_rt[20]), .Q(n923)
         );
  INV0 U1465 ( .A(i_data_FMalures[20]), .Q(n843) );
  XNR21 U1466 ( .A(compare_i_data_rs[8]), .B(compare_i_data_rt[8]), .Q(n924)
         );
  XNR21 U1467 ( .A(compare_i_data_rs[9]), .B(compare_i_data_rt[9]), .Q(n917)
         );
  XNR21 U1468 ( .A(compare_i_data_rs[6]), .B(compare_i_data_rt[6]), .Q(n918)
         );
  XNR21 U1469 ( .A(compare_i_data_rt[4]), .B(compare_i_data_rs[4]), .Q(n919)
         );
  XNR21 U1470 ( .A(compare_i_data_rs[7]), .B(compare_i_data_rt[7]), .Q(n920)
         );
  XNR21 U1471 ( .A(compare_i_data_rt[5]), .B(compare_i_data_rs[5]), .Q(n913)
         );
  XNR21 U1472 ( .A(compare_i_data_rs[11]), .B(compare_i_data_rt[11]), .Q(n914)
         );
  XNR21 U1473 ( .A(compare_i_data_rs[12]), .B(compare_i_data_rt[12]), .Q(n915)
         );
  XNR21 U1474 ( .A(compare_i_data_rs[10]), .B(compare_i_data_rt[10]), .Q(n909)
         );
  XNR21 U1475 ( .A(compare_i_data_rs[13]), .B(compare_i_data_rt[13]), .Q(n911)
         );
  XNR21 U1476 ( .A(compare_i_data_rs[14]), .B(compare_i_data_rt[14]), .Q(n912)
         );
  NAND22 U1477 ( .A(n562), .B(n561), .Q(compare_i_data_rt[31]) );
  OAI220 U1478 ( .A(n522), .B(n780), .C(n558), .D(n779), .Q(n559) );
  NOR20 U1479 ( .A(n778), .B(n630), .Q(n560) );
  AOI220 U1480 ( .A(n231), .B(i_data_FMmemout[30]), .C(n672), .D(
        i_data_FWmemout[30]), .Q(n564) );
  AOI220 U1481 ( .A(n671), .B(i_data_FMalures[30]), .C(n521), .D(
        i_data_FEalures[30]), .Q(n565) );
  AOI220 U1482 ( .A(n231), .B(i_data_FMmemout[29]), .C(n672), .D(
        i_data_FWmemout[29]), .Q(n568) );
  AOI220 U1483 ( .A(n671), .B(i_data_FMalures[29]), .C(n521), .D(
        i_data_FEalures[29]), .Q(n569) );
  AOI220 U1484 ( .A(n231), .B(i_data_FMmemout[28]), .C(n672), .D(
        i_data_FWmemout[28]), .Q(n572) );
  AOI220 U1485 ( .A(n671), .B(i_data_FMalures[28]), .C(n521), .D(
        i_data_FEalures[28]), .Q(n573) );
  NAND20 U1486 ( .A(n228), .B(i_data_rt[28]), .Q(n574) );
  AOI220 U1487 ( .A(n231), .B(i_data_FMmemout[27]), .C(n672), .D(
        i_data_FWmemout[27]), .Q(n576) );
  AOI220 U1488 ( .A(n671), .B(i_data_FMalures[27]), .C(n521), .D(
        i_data_FEalures[27]), .Q(n577) );
  AOI220 U1489 ( .A(n231), .B(i_data_FMmemout[26]), .C(n672), .D(
        i_data_FWmemout[26]), .Q(n580) );
  AOI220 U1490 ( .A(n671), .B(i_data_FMalures[26]), .C(n521), .D(
        i_data_FEalures[26]), .Q(n581) );
  AOI220 U1491 ( .A(n231), .B(i_data_FMmemout[25]), .C(n672), .D(
        i_data_FWmemout[25]), .Q(n584) );
  AOI220 U1492 ( .A(n671), .B(i_data_FMalures[25]), .C(n521), .D(
        i_data_FEalures[25]), .Q(n585) );
  AOI220 U1493 ( .A(n231), .B(i_data_FMmemout[24]), .C(n672), .D(
        i_data_FWmemout[24]), .Q(n588) );
  AOI220 U1494 ( .A(n231), .B(i_data_FMmemout[23]), .C(n672), .D(
        i_data_FWmemout[23]), .Q(n592) );
  AOI220 U1495 ( .A(n671), .B(i_data_FMalures[23]), .C(n521), .D(
        i_data_FEalures[23]), .Q(n593) );
  NAND20 U1496 ( .A(n228), .B(i_data_rt[23]), .Q(n594) );
  AOI220 U1497 ( .A(n231), .B(i_data_FMmemout[22]), .C(n672), .D(
        i_data_FWmemout[22]), .Q(n596) );
  AOI220 U1498 ( .A(n671), .B(i_data_FMalures[22]), .C(n521), .D(
        i_data_FEalures[22]), .Q(n597) );
  AOI220 U1499 ( .A(n671), .B(i_data_FMalures[21]), .C(n521), .D(
        i_data_FEalures[21]), .Q(n601) );
  AOI220 U1500 ( .A(n671), .B(i_data_FMalures[20]), .C(n521), .D(
        i_data_FEalures[20]), .Q(n605) );
  AOI220 U1501 ( .A(n671), .B(i_data_FMalures[19]), .C(n521), .D(
        i_data_FEalures[19]), .Q(n609) );
  AOI220 U1502 ( .A(n671), .B(i_data_FMalures[18]), .C(n521), .D(
        i_data_FEalures[18]), .Q(n613) );
  NAND20 U1503 ( .A(n1264), .B(n1080), .Q(n1081) );
  XNR21 U1504 ( .A(n107), .B(alu_i_data_B[17]), .Q(n1080) );
  NAND20 U1505 ( .A(n1242), .B(alu_i_data_B[1]), .Q(n1079) );
  INV0 U1506 ( .A(i_data_FMalures[17]), .Q(n867) );
  NAND20 U1507 ( .A(n122), .B(i_data_FMmemout[16]), .Q(n901) );
  INV0 U1508 ( .A(i_data_FMalures[16]), .Q(n899) );
  INV3 U1509 ( .A(n771), .Q(n765) );
  INV3 U1510 ( .A(alu_i_con_AluCtrl[0]), .Q(n978) );
  INV3 U1511 ( .A(n544), .Q(n766) );
  NAND20 U1512 ( .A(n122), .B(i_data_FMmemout[13]), .Q(n689) );
  INV0 U1513 ( .A(i_data_FMalures[13]), .Q(n688) );
  INV0 U1514 ( .A(i_data_FMalures[10]), .Q(n709) );
  INV0 U1515 ( .A(i_data_FMalures[9]), .Q(n716) );
  INV0 U1516 ( .A(i_data_FMalures[8]), .Q(n723) );
  INV0 U1517 ( .A(i_data_FMalures[11]), .Q(n702) );
  AOI220 U1518 ( .A(n523), .B(i_data_FMalures[3]), .C(n121), .D(
        i_data_FEalures[3]), .Q(n748) );
  AOI220 U1519 ( .A(n523), .B(i_data_FMalures[2]), .C(n121), .D(
        i_data_FEalures[2]), .Q(n751) );
  AOI220 U1520 ( .A(n671), .B(i_data_FMalures[0]), .C(n521), .D(
        i_data_FEalures[0]), .Q(n675) );
  NAND20 U1521 ( .A(n122), .B(i_data_FMmemout[0]), .Q(n757) );
  INV0 U1522 ( .A(i_data_FMalures[0]), .Q(n756) );
  NAND20 U1523 ( .A(n122), .B(i_data_FMmemout[7]), .Q(n731) );
  INV0 U1524 ( .A(i_data_FMalures[7]), .Q(n730) );
  INV0 U1525 ( .A(i_data_FMalures[6]), .Q(n737) );
  AOI220 U1526 ( .A(n523), .B(i_data_FMalures[5]), .C(n121), .D(
        i_data_FEalures[5]), .Q(n536) );
  AOI220 U1527 ( .A(n523), .B(i_data_FMalures[4]), .C(n121), .D(
        i_data_FEalures[4]), .Q(n745) );
  NAND20 U1528 ( .A(n122), .B(i_data_FMmemout[12]), .Q(n696) );
  INV0 U1529 ( .A(i_data_FMalures[12]), .Q(n695) );
  NAND20 U1530 ( .A(n122), .B(i_data_FMmemout[14]), .Q(n682) );
  AOI220 U1531 ( .A(n122), .B(i_data_FMmemout[15]), .C(n523), .D(
        i_data_FMalures[15]), .Q(n678) );
  AOI220 U1532 ( .A(n673), .B(i_data_FMmemout[15]), .C(n671), .D(
        i_data_FMalures[15]), .Q(n627) );
  INV3 U1533 ( .A(n552), .Q(n553) );
  AOI220 U1534 ( .A(n671), .B(i_data_FMalures[24]), .C(n521), .D(
        i_data_FEalures[24]), .Q(n589) );
  OAI310 U1535 ( .A(compare_i_data_rs[17]), .B(alu_i_data_B[17]), .C(n1247), 
        .D(n1081), .Q(n1082) );
  XNR21 U1536 ( .A(compare_i_data_rs[17]), .B(compare_i_data_rt[17]), .Q(n931)
         );
  AOI2110 U1537 ( .A(n1162), .B(compare_i_data_rs[24]), .C(n1161), .D(n98), 
        .Q(n1168) );
  AOI210 U1538 ( .A(n1165), .B(compare_i_data_rs[24]), .C(n1164), .Q(n1166) );
  OAI310 U1539 ( .A(alu_i_data_B[24]), .B(compare_i_data_rs[24]), .C(n1247), 
        .D(n1163), .Q(n1164) );
  XNR21 U1540 ( .A(compare_i_data_rs[24]), .B(compare_i_data_rt[24]), .Q(n939)
         );
  INV3 U1541 ( .A(n547), .Q(n546) );
  AOI2110 U1542 ( .A(n1162), .B(compare_i_data_rs[16]), .C(n1067), .D(n98), 
        .Q(n1075) );
  AOI210 U1543 ( .A(n1072), .B(compare_i_data_rs[16]), .C(n1071), .Q(n1073) );
  OAI310 U1544 ( .A(alu_i_data_B[16]), .B(compare_i_data_rs[16]), .C(n1247), 
        .D(n1070), .Q(n1071) );
  XNR21 U1545 ( .A(compare_i_data_rt[1]), .B(compare_i_data_rs[1]), .Q(n934)
         );
  AOI220 U1546 ( .A(n671), .B(i_data_FMalures[17]), .C(n521), .D(
        i_data_FEalures[17]), .Q(n617) );
  XNR21 U1547 ( .A(compare_i_data_rs[0]), .B(compare_i_data_rt[0]), .Q(n916)
         );
  XNR21 U1548 ( .A(compare_i_data_rs[16]), .B(compare_i_data_rt[16]), .Q(n910)
         );
  XNR21 U1549 ( .A(compare_i_data_rt[3]), .B(compare_i_data_rs[3]), .Q(n922)
         );
  NOR40 U1550 ( .A(u_alu_ashr_4_SH_3_), .B(i_data_immext[8]), .C(n381), .D(
        n241), .Q(n261) );
  IMUX20 U1551 ( .A(n236), .B(n238), .S(n381), .Q(n250) );
  IMUX20 U1552 ( .A(n253), .B(n243), .S(n381), .Q(n264) );
  IMUX20 U1553 ( .A(n302), .B(n305), .S(u_alu_ashr_4_SH_3_), .Q(n262) );
  IMUX20 U1554 ( .A(n286), .B(n264), .S(i_data_immext[8]), .Q(n309) );
  IMUX20 U1555 ( .A(n309), .B(n312), .S(u_alu_ashr_4_SH_3_), .Q(n268) );
  IMUX20 U1556 ( .A(n280), .B(n269), .S(n381), .Q(n291) );
  IMUX20 U1557 ( .A(n316), .B(n271), .S(u_alu_ashr_4_SH_3_), .Q(n273) );
  IMUX20 U1558 ( .A(n296), .B(n275), .S(i_data_immext[8]), .Q(n322) );
  IMUX20 U1559 ( .A(n322), .B(n276), .S(u_alu_ashr_4_SH_3_), .Q(n278) );
  IMUX20 U1560 ( .A(n329), .B(n282), .S(u_alu_ashr_4_SH_3_), .Q(n284) );
  IMUX20 U1561 ( .A(n336), .B(n287), .S(u_alu_ashr_4_SH_3_), .Q(n289) );
  IMUX20 U1562 ( .A(n345), .B(n292), .S(u_alu_ashr_4_SH_3_), .Q(n294) );
  IMUX20 U1563 ( .A(n353), .B(n297), .S(u_alu_ashr_4_SH_3_), .Q(n299) );
  IMUX20 U1564 ( .A(n314), .B(n300), .S(n381), .Q(n327) );
  IMUX20 U1565 ( .A(n327), .B(n301), .S(i_data_immext[8]), .Q(n303) );
  IMUX20 U1566 ( .A(n303), .B(n302), .S(u_alu_ashr_4_SH_3_), .Q(n306) );
  IMUX20 U1567 ( .A(alu_i_data_B[25]), .B(alu_i_data_B[24]), .S(
        i_data_immext[6]), .Q(n320) );
  IMUX20 U1568 ( .A(n320), .B(n307), .S(n381), .Q(n334) );
  IMUX20 U1569 ( .A(n334), .B(n308), .S(i_data_immext[8]), .Q(n310) );
  IMUX20 U1570 ( .A(n310), .B(n309), .S(u_alu_ashr_4_SH_3_), .Q(n313) );
  IMUX20 U1571 ( .A(alu_i_data_B[26]), .B(alu_i_data_B[25]), .S(
        i_data_immext[6]), .Q(n326) );
  IMUX20 U1572 ( .A(n343), .B(n315), .S(i_data_immext[8]), .Q(n317) );
  IMUX20 U1573 ( .A(n317), .B(n316), .S(u_alu_ashr_4_SH_3_), .Q(n319) );
  IMUX20 U1574 ( .A(n351), .B(n321), .S(i_data_immext[8]), .Q(n323) );
  IMUX20 U1575 ( .A(n323), .B(n322), .S(u_alu_ashr_4_SH_3_), .Q(n325) );
  IMUX20 U1576 ( .A(n328), .B(n327), .S(i_data_immext[8]), .Q(n330) );
  IMUX20 U1577 ( .A(n330), .B(n329), .S(u_alu_ashr_4_SH_3_), .Q(n332) );
  IMUX20 U1578 ( .A(n335), .B(n334), .S(i_data_immext[8]), .Q(n337) );
  IMUX20 U1579 ( .A(n337), .B(n336), .S(u_alu_ashr_4_SH_3_), .Q(n339) );
  IMUX20 U1580 ( .A(n344), .B(n343), .S(i_data_immext[8]), .Q(n346) );
  IMUX20 U1581 ( .A(n346), .B(n345), .S(u_alu_ashr_4_SH_3_), .Q(n348) );
  IMUX20 U1582 ( .A(n352), .B(n351), .S(i_data_immext[8]), .Q(n354) );
  IMUX20 U1583 ( .A(n354), .B(n353), .S(u_alu_ashr_4_SH_3_), .Q(n356) );
  NOR20 U1584 ( .A(i_data_immext[10]), .B(n367), .Q(u_alu_N196) );
  NOR20 U1585 ( .A(i_data_immext[10]), .B(n369), .Q(u_alu_N198) );
  IMUX20 U1586 ( .A(n384), .B(n481), .S(i_data_immext[8]), .Q(n385) );
  IMUX20 U1587 ( .A(n385), .B(n501), .S(u_alu_ashr_4_SH_3_), .Q(n386) );
  IMUX20 U1588 ( .A(alu_i_data_B[24]), .B(alu_i_data_B[25]), .S(
        i_data_immext[6]), .Q(n393) );
  IMUX20 U1589 ( .A(n390), .B(n389), .S(n381), .Q(n417) );
  IMUX20 U1590 ( .A(n392), .B(n391), .S(n381), .Q(n416) );
  IMUX20 U1591 ( .A(n394), .B(n393), .S(n381), .Q(n419) );
  IMUX20 U1592 ( .A(n416), .B(n419), .S(i_data_immext[8]), .Q(n432) );
  IMUX20 U1593 ( .A(n464), .B(n432), .S(u_alu_ashr_4_SH_3_), .Q(n398) );
  IMUX20 U1594 ( .A(n407), .B(n410), .S(n381), .Q(n421) );
  IMUX20 U1595 ( .A(alu_i_data_B[25]), .B(alu_i_data_B[26]), .S(
        i_data_immext[6]), .Q(n412) );
  IMUX20 U1596 ( .A(n409), .B(n412), .S(n381), .Q(n424) );
  IMUX20 U1597 ( .A(n475), .B(n434), .S(u_alu_ashr_4_SH_3_), .Q(n399) );
  IMUX20 U1598 ( .A(n411), .B(n414), .S(n381), .Q(n423) );
  MUX21 U1599 ( .A(n401), .B(n400), .S(i_data_immext[8]), .Q(n479) );
  IMUX20 U1600 ( .A(n406), .B(n405), .S(n381), .Q(n438) );
  IMUX20 U1601 ( .A(n438), .B(n428), .S(i_data_immext[8]), .Q(n486) );
  IMUX20 U1602 ( .A(n410), .B(n409), .S(n381), .Q(n427) );
  IMUX20 U1603 ( .A(n427), .B(n430), .S(i_data_immext[8]), .Q(n446) );
  IMUX20 U1604 ( .A(n486), .B(n446), .S(u_alu_ashr_4_SH_3_), .Q(n415) );
  MUX21 U1605 ( .A(n417), .B(n416), .S(i_data_immext[8]), .Q(n490) );
  MUX21 U1606 ( .A(n422), .B(n421), .S(i_data_immext[8]), .Q(n495) );
  MUX21 U1607 ( .A(n424), .B(n423), .S(i_data_immext[8]), .Q(n452) );
  IMUX20 U1608 ( .A(n495), .B(n452), .S(u_alu_ashr_4_SH_3_), .Q(n425) );
  IMUX20 U1609 ( .A(n436), .B(n485), .S(i_data_immext[8]), .Q(n439) );
  IMUX20 U1610 ( .A(n439), .B(n505), .S(u_alu_ashr_4_SH_3_), .Q(n441) );
  NOR20 U1611 ( .A(i_data_immext[10]), .B(n482), .Q(u_alu_N245) );
  NOR20 U1612 ( .A(i_data_immext[10]), .B(n493), .Q(u_alu_N247) );
  NOR20 U1613 ( .A(i_data_immext[10]), .B(n457), .Q(u_alu_N253) );
  IMUX20 U1614 ( .A(n463), .B(n492), .S(i_data_immext[8]), .Q(n465) );
  IMUX20 U1615 ( .A(n465), .B(n464), .S(u_alu_ashr_4_SH_3_), .Q(n467) );
  NOR20 U1616 ( .A(i_data_immext[10]), .B(n468), .Q(u_alu_N255) );
  IMUX20 U1617 ( .A(n474), .B(n497), .S(i_data_immext[8]), .Q(n476) );
  IMUX20 U1618 ( .A(n476), .B(n475), .S(u_alu_ashr_4_SH_3_), .Q(n478) );
  IMUX30 U1619 ( .A(n481), .B(n480), .C(n479), .S0(i_data_immext[8]), .S1(
        u_alu_ashr_4_SH_3_), .Q(n483) );
  IMUX20 U1620 ( .A(n485), .B(n484), .S(i_data_immext[8]), .Q(n487) );
  IMUX20 U1621 ( .A(n487), .B(n486), .S(u_alu_ashr_4_SH_3_), .Q(n489) );
  IMUX30 U1622 ( .A(n492), .B(n491), .C(n490), .S0(i_data_immext[8]), .S1(
        u_alu_ashr_4_SH_3_), .Q(n494) );
  IMUX30 U1623 ( .A(n497), .B(n496), .C(n495), .S0(i_data_immext[8]), .S1(
        u_alu_ashr_4_SH_3_), .Q(n499) );
  IMUX20 U1624 ( .A(n501), .B(n500), .S(u_alu_ashr_4_SH_3_), .Q(n503) );
  OAI212 U1625 ( .A(n630), .B(n1330), .C(n629), .Q(compare_i_data_rt[15]) );
  IMUX20 U1626 ( .A(n1266), .B(n1267), .S(alu_i_data_B[5]), .Q(n1271) );
  IMUX20 U1627 ( .A(n1266), .B(n1267), .S(alu_i_data_B[3]), .Q(n1281) );
  NOR20 U1628 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[31]), .Q(n1283)
         );
  NOR20 U1629 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[30]), .Q(n1284)
         );
  NOR20 U1630 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[29]), .Q(n1290)
         );
  NOR20 U1631 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[28]), .Q(n1291)
         );
  NOR20 U1632 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[27]), .Q(n1292)
         );
  NOR20 U1633 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[26]), .Q(n1293)
         );
  NOR20 U1634 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[25]), .Q(n1294)
         );
  NOR20 U1635 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[23]), .Q(n1295)
         );
  NOR20 U1636 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[22]), .Q(n1296)
         );
  NOR20 U1637 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[21]), .Q(n1297)
         );
  NOR20 U1638 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[20]), .Q(n1298)
         );
  NOR20 U1639 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[19]), .Q(n1304)
         );
  NOR20 U1640 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[18]), .Q(n1305)
         );
  NOR20 U1641 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[17]), .Q(n1306)
         );
  NOR30 U1642 ( .A(i_con_Ealuop[2]), .B(i_con_Ealuop[3]), .C(n1328), .Q(n1319)
         );
  IMUX20 U1643 ( .A(i_addr_rt[0]), .B(i_data_immext[11]), .S(i_con_Eregdst), 
        .Q(n1331) );
  IMUX20 U1644 ( .A(i_addr_rt[1]), .B(i_data_immext[12]), .S(i_con_Eregdst), 
        .Q(n1332) );
  IMUX20 U1645 ( .A(i_addr_rt[2]), .B(i_data_immext[13]), .S(i_con_Eregdst), 
        .Q(n1333) );
  IMUX20 U1646 ( .A(i_addr_rt[3]), .B(i_data_immext[14]), .S(i_con_Eregdst), 
        .Q(n1334) );
  IMUX20 U1647 ( .A(i_addr_rt[4]), .B(i_data_immext[15]), .S(i_con_Eregdst), 
        .Q(n1335) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_con_RegWr, i_addr_Rd, 
        i_data_Rd, o_data_Rs, o_data_Rt, i_addr_Rt_4_, i_addr_Rt_3_, 
        i_addr_Rt_2_, i_addr_Rt_1_, i_addr_Rt_0_ );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr, i_addr_Rt_4_, i_addr_Rt_3_, i_addr_Rt_2_,
         i_addr_Rt_1_, i_addr_Rt_0_;
  wire   n5, n6, n9, n11, n13, n15, n16, n17, n18, n20, n21, n22, n23, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n1, n2, n3, n4, n7, n8, n10, n12, n14, n19, n24,
         n33, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591;
  wire   [1023:0] regs;

  DFEC1 regs_reg_31__30_ ( .D(i_data_Rd[30]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(i_data_Rd[29]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(i_data_Rd[28]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(i_data_Rd[27]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(i_data_Rd[26]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(i_data_Rd[25]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(i_data_Rd[24]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(i_data_Rd[23]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(i_data_Rd[22]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(i_data_Rd[21]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(i_data_Rd[20]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(i_data_Rd[18]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(i_data_Rd[17]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(i_data_Rd[16]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(i_data_Rd[15]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(i_data_Rd[14]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(i_data_Rd[13]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(i_data_Rd[12]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(i_data_Rd[11]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(i_data_Rd[10]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(i_data_Rd[9]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(i_data_Rd[8]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(i_data_Rd[7]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(i_data_Rd[5]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(i_data_Rd[4]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(i_data_Rd[3]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(i_data_Rd[2]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(i_data_Rd[0]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[992]) );
  DFEC1 regs_reg_30__31_ ( .D(i_data_Rd[31]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(i_data_Rd[30]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(i_data_Rd[29]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(i_data_Rd[28]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(i_data_Rd[27]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(i_data_Rd[26]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(i_data_Rd[25]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(i_data_Rd[24]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(i_data_Rd[23]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(i_data_Rd[22]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(i_data_Rd[21]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(i_data_Rd[20]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(i_data_Rd[18]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(i_data_Rd[17]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(i_data_Rd[16]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(i_data_Rd[15]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(i_data_Rd[14]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(i_data_Rd[13]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(i_data_Rd[12]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(i_data_Rd[11]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(i_data_Rd[10]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(i_data_Rd[9]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(i_data_Rd[8]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(i_data_Rd[7]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(i_data_Rd[5]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(i_data_Rd[4]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(i_data_Rd[3]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(i_data_Rd[2]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(i_data_Rd[0]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[960]) );
  DFEC1 regs_reg_29__31_ ( .D(i_data_Rd[31]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(i_data_Rd[30]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(i_data_Rd[29]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(i_data_Rd[28]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[956]) );
  DFEC1 regs_reg_29__27_ ( .D(i_data_Rd[27]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(i_data_Rd[26]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(i_data_Rd[25]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(i_data_Rd[24]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(i_data_Rd[23]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(i_data_Rd[22]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(i_data_Rd[21]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(i_data_Rd[20]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(i_data_Rd[18]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(i_data_Rd[17]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(i_data_Rd[16]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(i_data_Rd[15]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(i_data_Rd[14]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(i_data_Rd[13]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(i_data_Rd[12]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(i_data_Rd[11]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(i_data_Rd[10]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(i_data_Rd[9]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(i_data_Rd[8]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(i_data_Rd[7]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(i_data_Rd[5]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(i_data_Rd[4]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(i_data_Rd[3]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(i_data_Rd[2]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(i_data_Rd[0]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[928]) );
  DFEC1 regs_reg_28__31_ ( .D(i_data_Rd[31]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(i_data_Rd[30]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(i_data_Rd[29]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(i_data_Rd[28]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(i_data_Rd[27]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(i_data_Rd[26]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(i_data_Rd[25]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(i_data_Rd[24]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(i_data_Rd[23]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(i_data_Rd[22]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(i_data_Rd[21]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(i_data_Rd[20]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(i_data_Rd[18]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(i_data_Rd[17]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(i_data_Rd[16]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(i_data_Rd[15]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(i_data_Rd[14]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(i_data_Rd[13]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(i_data_Rd[12]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(i_data_Rd[11]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(i_data_Rd[10]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(i_data_Rd[9]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(i_data_Rd[8]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(i_data_Rd[7]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(i_data_Rd[5]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(i_data_Rd[4]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(i_data_Rd[3]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(i_data_Rd[2]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(i_data_Rd[0]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(i_data_Rd[31]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(i_data_Rd[30]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(i_data_Rd[29]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(i_data_Rd[28]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(i_data_Rd[27]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(i_data_Rd[26]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(i_data_Rd[25]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(i_data_Rd[24]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(i_data_Rd[23]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(i_data_Rd[22]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(i_data_Rd[21]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(i_data_Rd[20]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(i_data_Rd[18]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(i_data_Rd[17]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(i_data_Rd[16]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(i_data_Rd[15]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(i_data_Rd[14]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(i_data_Rd[13]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(i_data_Rd[12]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(i_data_Rd[11]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(i_data_Rd[10]), .E(n123), .C(i_clk), .RN(i_rst_n), .Q(regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(i_data_Rd[9]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(i_data_Rd[8]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(i_data_Rd[7]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(i_data_Rd[5]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(i_data_Rd[4]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(i_data_Rd[3]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(i_data_Rd[2]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(i_data_Rd[1]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(i_data_Rd[0]), .E(n123), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[864]) );
  DFEC1 regs_reg_26__31_ ( .D(i_data_Rd[31]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(i_data_Rd[30]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(i_data_Rd[29]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(i_data_Rd[28]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(i_data_Rd[27]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(i_data_Rd[26]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(i_data_Rd[25]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(i_data_Rd[24]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(i_data_Rd[23]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(i_data_Rd[22]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(i_data_Rd[21]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(i_data_Rd[20]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(i_data_Rd[18]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(i_data_Rd[17]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(i_data_Rd[16]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(i_data_Rd[15]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(i_data_Rd[14]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(i_data_Rd[13]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(i_data_Rd[12]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(i_data_Rd[11]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(i_data_Rd[10]), .E(n124), .C(i_clk), .RN(i_rst_n), .Q(regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(i_data_Rd[9]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(i_data_Rd[8]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(i_data_Rd[7]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(i_data_Rd[5]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(i_data_Rd[4]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(i_data_Rd[3]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(i_data_Rd[2]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(i_data_Rd[0]), .E(n124), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[832]) );
  DFEC1 regs_reg_25__31_ ( .D(i_data_Rd[31]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(i_data_Rd[30]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(i_data_Rd[29]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(i_data_Rd[28]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(i_data_Rd[27]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(i_data_Rd[26]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(i_data_Rd[25]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(i_data_Rd[24]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(i_data_Rd[23]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(i_data_Rd[22]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(i_data_Rd[21]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(i_data_Rd[20]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(i_data_Rd[19]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(i_data_Rd[18]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(i_data_Rd[17]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(i_data_Rd[16]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(i_data_Rd[15]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(i_data_Rd[14]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(i_data_Rd[13]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(i_data_Rd[12]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(i_data_Rd[11]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(i_data_Rd[10]), .E(n125), .C(i_clk), .RN(i_rst_n), .Q(regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(i_data_Rd[9]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(i_data_Rd[8]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(i_data_Rd[7]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(i_data_Rd[6]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(i_data_Rd[5]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(i_data_Rd[4]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(i_data_Rd[3]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(i_data_Rd[2]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(i_data_Rd[1]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(i_data_Rd[0]), .E(n125), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[800]) );
  DFEC1 regs_reg_24__31_ ( .D(i_data_Rd[31]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(i_data_Rd[30]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(i_data_Rd[29]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(i_data_Rd[28]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(i_data_Rd[27]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(i_data_Rd[26]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(i_data_Rd[25]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(i_data_Rd[24]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(i_data_Rd[23]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(i_data_Rd[22]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(i_data_Rd[21]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(i_data_Rd[20]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(i_data_Rd[19]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(i_data_Rd[18]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(i_data_Rd[17]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(i_data_Rd[16]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(i_data_Rd[15]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(i_data_Rd[14]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(i_data_Rd[13]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(i_data_Rd[12]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(i_data_Rd[11]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(i_data_Rd[10]), .E(n126), .C(i_clk), .RN(i_rst_n), .Q(regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(i_data_Rd[9]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(i_data_Rd[8]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(i_data_Rd[7]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(i_data_Rd[6]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(i_data_Rd[5]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(i_data_Rd[4]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(i_data_Rd[3]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(i_data_Rd[2]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(i_data_Rd[1]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(i_data_Rd[0]), .E(n126), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(i_data_Rd[31]), .E(n22), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(i_data_Rd[30]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(i_data_Rd[29]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(i_data_Rd[28]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(i_data_Rd[27]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(i_data_Rd[26]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(i_data_Rd[25]), .E(n22), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(i_data_Rd[24]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(i_data_Rd[23]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(i_data_Rd[22]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(i_data_Rd[21]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(i_data_Rd[20]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(i_data_Rd[19]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(i_data_Rd[18]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(i_data_Rd[17]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(i_data_Rd[16]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(i_data_Rd[15]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(i_data_Rd[14]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(i_data_Rd[13]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(i_data_Rd[12]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(i_data_Rd[11]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(i_data_Rd[10]), .E(n127), .C(i_clk), .RN(i_rst_n), .Q(regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(i_data_Rd[9]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(i_data_Rd[8]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(i_data_Rd[7]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(i_data_Rd[6]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(i_data_Rd[5]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(i_data_Rd[4]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(i_data_Rd[3]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(i_data_Rd[2]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(i_data_Rd[1]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(i_data_Rd[0]), .E(n127), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[736]) );
  DFEC1 regs_reg_22__31_ ( .D(i_data_Rd[31]), .E(n21), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(i_data_Rd[30]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(i_data_Rd[29]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(i_data_Rd[28]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(i_data_Rd[27]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(i_data_Rd[26]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(i_data_Rd[25]), .E(n21), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(i_data_Rd[24]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(i_data_Rd[23]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(i_data_Rd[22]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(i_data_Rd[21]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(i_data_Rd[20]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(i_data_Rd[19]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(i_data_Rd[18]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(i_data_Rd[17]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(i_data_Rd[16]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(i_data_Rd[15]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(i_data_Rd[14]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(i_data_Rd[13]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(i_data_Rd[12]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(i_data_Rd[11]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(i_data_Rd[10]), .E(n128), .C(i_clk), .RN(i_rst_n), .Q(regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(i_data_Rd[9]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(i_data_Rd[8]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(i_data_Rd[7]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(i_data_Rd[6]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(i_data_Rd[5]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(i_data_Rd[4]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(i_data_Rd[3]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(i_data_Rd[2]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(i_data_Rd[1]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(i_data_Rd[0]), .E(n128), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[704]) );
  DFEC1 regs_reg_21__31_ ( .D(i_data_Rd[31]), .E(n20), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(i_data_Rd[30]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(i_data_Rd[29]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(i_data_Rd[28]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(i_data_Rd[27]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(i_data_Rd[26]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(i_data_Rd[25]), .E(n20), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(i_data_Rd[24]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(i_data_Rd[23]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(i_data_Rd[22]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(i_data_Rd[21]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(i_data_Rd[20]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(i_data_Rd[19]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(i_data_Rd[18]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(i_data_Rd[17]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(i_data_Rd[16]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(i_data_Rd[15]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(i_data_Rd[14]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(i_data_Rd[13]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(i_data_Rd[12]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(i_data_Rd[11]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(i_data_Rd[10]), .E(n129), .C(i_clk), .RN(i_rst_n), .Q(regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(i_data_Rd[9]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(i_data_Rd[8]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(i_data_Rd[7]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(i_data_Rd[6]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(i_data_Rd[5]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(i_data_Rd[4]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(i_data_Rd[3]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(i_data_Rd[2]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(i_data_Rd[1]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(i_data_Rd[0]), .E(n129), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[672]) );
  DFEC1 regs_reg_20__31_ ( .D(i_data_Rd[31]), .E(n18), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(i_data_Rd[30]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(i_data_Rd[29]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(i_data_Rd[28]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(i_data_Rd[27]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(i_data_Rd[26]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(i_data_Rd[25]), .E(n18), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(i_data_Rd[24]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(i_data_Rd[23]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(i_data_Rd[22]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(i_data_Rd[21]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(i_data_Rd[20]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(i_data_Rd[19]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(i_data_Rd[18]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(i_data_Rd[17]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(i_data_Rd[16]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(i_data_Rd[15]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(i_data_Rd[14]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(i_data_Rd[13]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(i_data_Rd[12]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(i_data_Rd[11]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(i_data_Rd[10]), .E(n130), .C(i_clk), .RN(i_rst_n), .Q(regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(i_data_Rd[9]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(i_data_Rd[8]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(i_data_Rd[7]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(i_data_Rd[6]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(i_data_Rd[5]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(i_data_Rd[4]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(i_data_Rd[3]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(i_data_Rd[2]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(i_data_Rd[1]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(i_data_Rd[0]), .E(n130), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(i_data_Rd[31]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(i_data_Rd[30]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(i_data_Rd[29]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(i_data_Rd[28]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(i_data_Rd[27]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(i_data_Rd[26]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(i_data_Rd[25]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(i_data_Rd[24]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(i_data_Rd[23]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(i_data_Rd[22]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(i_data_Rd[21]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(i_data_Rd[20]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(i_data_Rd[19]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(i_data_Rd[18]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(i_data_Rd[17]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(i_data_Rd[16]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(i_data_Rd[15]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(i_data_Rd[14]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(i_data_Rd[13]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(i_data_Rd[12]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(i_data_Rd[11]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(i_data_Rd[10]), .E(n131), .C(i_clk), .RN(i_rst_n), .Q(regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(i_data_Rd[9]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(i_data_Rd[8]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(i_data_Rd[7]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(i_data_Rd[6]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(i_data_Rd[5]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(i_data_Rd[4]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(i_data_Rd[3]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(i_data_Rd[2]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(i_data_Rd[1]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(i_data_Rd[0]), .E(n131), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[608]) );
  DFEC1 regs_reg_18__31_ ( .D(i_data_Rd[31]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(i_data_Rd[30]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(i_data_Rd[29]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(i_data_Rd[28]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(i_data_Rd[27]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(i_data_Rd[26]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(i_data_Rd[25]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(i_data_Rd[24]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(i_data_Rd[23]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(i_data_Rd[22]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(i_data_Rd[21]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(i_data_Rd[20]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(i_data_Rd[19]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(i_data_Rd[18]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(i_data_Rd[17]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(i_data_Rd[16]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(i_data_Rd[15]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(i_data_Rd[14]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(i_data_Rd[13]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(i_data_Rd[12]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(i_data_Rd[11]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(i_data_Rd[10]), .E(n132), .C(i_clk), .RN(i_rst_n), .Q(regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(i_data_Rd[9]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(i_data_Rd[8]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(i_data_Rd[7]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(i_data_Rd[6]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(i_data_Rd[5]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(i_data_Rd[4]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(i_data_Rd[3]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(i_data_Rd[2]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(i_data_Rd[1]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(i_data_Rd[0]), .E(n132), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[576]) );
  DFEC1 regs_reg_17__31_ ( .D(i_data_Rd[31]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(i_data_Rd[30]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(i_data_Rd[29]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(i_data_Rd[28]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(i_data_Rd[27]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(i_data_Rd[26]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(i_data_Rd[25]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(i_data_Rd[24]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(i_data_Rd[23]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(i_data_Rd[22]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(i_data_Rd[21]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(i_data_Rd[20]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(i_data_Rd[19]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(i_data_Rd[18]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(i_data_Rd[17]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(i_data_Rd[16]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(i_data_Rd[15]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(i_data_Rd[14]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(i_data_Rd[13]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(i_data_Rd[12]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(i_data_Rd[11]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(i_data_Rd[10]), .E(n133), .C(i_clk), .RN(i_rst_n), .Q(regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(i_data_Rd[9]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(i_data_Rd[8]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(i_data_Rd[7]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(i_data_Rd[6]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(i_data_Rd[5]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(i_data_Rd[4]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(i_data_Rd[3]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(i_data_Rd[2]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(i_data_Rd[1]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(i_data_Rd[0]), .E(n133), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(i_data_Rd[31]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(i_data_Rd[30]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(i_data_Rd[29]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(i_data_Rd[28]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(i_data_Rd[27]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(i_data_Rd[26]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(i_data_Rd[25]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(i_data_Rd[24]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(i_data_Rd[23]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(i_data_Rd[22]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(i_data_Rd[21]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(i_data_Rd[20]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(i_data_Rd[19]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(i_data_Rd[18]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(i_data_Rd[17]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(i_data_Rd[16]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(i_data_Rd[15]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(i_data_Rd[14]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(i_data_Rd[13]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(i_data_Rd[12]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(i_data_Rd[11]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(i_data_Rd[10]), .E(n134), .C(i_clk), .RN(i_rst_n), .Q(regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(i_data_Rd[9]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(i_data_Rd[8]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(i_data_Rd[7]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(i_data_Rd[6]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(i_data_Rd[5]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(i_data_Rd[4]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(i_data_Rd[3]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(i_data_Rd[2]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(i_data_Rd[1]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(i_data_Rd[0]), .E(n134), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[512]) );
  DFEC1 regs_reg_15__31_ ( .D(i_data_Rd[31]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(i_data_Rd[30]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(i_data_Rd[29]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(i_data_Rd[28]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(i_data_Rd[27]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(i_data_Rd[26]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(i_data_Rd[25]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(i_data_Rd[24]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(i_data_Rd[23]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(i_data_Rd[22]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(i_data_Rd[21]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(i_data_Rd[20]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(i_data_Rd[19]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(i_data_Rd[18]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(i_data_Rd[17]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(i_data_Rd[16]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(i_data_Rd[15]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(i_data_Rd[13]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(i_data_Rd[12]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(i_data_Rd[11]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(i_data_Rd[9]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(i_data_Rd[8]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(i_data_Rd[7]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(i_data_Rd[6]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(i_data_Rd[5]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(i_data_Rd[4]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(i_data_Rd[3]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(i_data_Rd[2]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(i_data_Rd[1]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(i_data_Rd[0]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[480]) );
  DFEC1 regs_reg_14__31_ ( .D(i_data_Rd[31]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(i_data_Rd[30]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(i_data_Rd[29]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(i_data_Rd[28]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(i_data_Rd[27]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(i_data_Rd[26]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(i_data_Rd[25]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(i_data_Rd[24]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(i_data_Rd[23]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(i_data_Rd[22]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(i_data_Rd[21]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(i_data_Rd[20]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(i_data_Rd[19]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(i_data_Rd[18]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(i_data_Rd[17]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(i_data_Rd[16]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(i_data_Rd[15]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(i_data_Rd[13]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(i_data_Rd[12]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(i_data_Rd[11]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(i_data_Rd[9]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(i_data_Rd[8]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(i_data_Rd[7]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(i_data_Rd[6]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(i_data_Rd[5]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(i_data_Rd[4]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(i_data_Rd[3]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(i_data_Rd[2]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(i_data_Rd[1]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(i_data_Rd[0]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[448]) );
  DFEC1 regs_reg_13__31_ ( .D(i_data_Rd[31]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(i_data_Rd[30]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(i_data_Rd[29]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(i_data_Rd[28]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[444]) );
  DFEC1 regs_reg_13__27_ ( .D(i_data_Rd[27]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(i_data_Rd[26]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(i_data_Rd[25]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(i_data_Rd[24]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(i_data_Rd[23]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(i_data_Rd[22]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(i_data_Rd[21]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(i_data_Rd[20]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(i_data_Rd[19]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(i_data_Rd[18]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(i_data_Rd[17]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(i_data_Rd[16]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(i_data_Rd[15]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(i_data_Rd[13]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(i_data_Rd[12]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(i_data_Rd[11]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(i_data_Rd[9]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(i_data_Rd[8]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(i_data_Rd[7]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(i_data_Rd[6]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(i_data_Rd[5]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(i_data_Rd[4]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(i_data_Rd[3]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(i_data_Rd[2]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(i_data_Rd[1]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(i_data_Rd[0]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[416]) );
  DFEC1 regs_reg_12__31_ ( .D(i_data_Rd[31]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(i_data_Rd[30]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(i_data_Rd[29]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(i_data_Rd[28]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(i_data_Rd[27]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(i_data_Rd[26]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(i_data_Rd[25]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(i_data_Rd[24]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(i_data_Rd[23]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(i_data_Rd[22]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(i_data_Rd[21]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(i_data_Rd[20]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(i_data_Rd[19]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(i_data_Rd[18]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(i_data_Rd[17]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(i_data_Rd[16]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(i_data_Rd[15]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(i_data_Rd[13]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(i_data_Rd[12]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(i_data_Rd[11]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(i_data_Rd[9]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(i_data_Rd[8]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(i_data_Rd[7]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(i_data_Rd[6]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(i_data_Rd[5]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(i_data_Rd[4]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(i_data_Rd[3]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(i_data_Rd[2]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(i_data_Rd[1]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(i_data_Rd[0]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[384]) );
  DFEC1 regs_reg_11__31_ ( .D(i_data_Rd[31]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(i_data_Rd[30]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(i_data_Rd[29]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(i_data_Rd[28]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(i_data_Rd[27]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(i_data_Rd[26]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(i_data_Rd[25]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(i_data_Rd[24]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(i_data_Rd[23]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(i_data_Rd[22]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(i_data_Rd[21]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(i_data_Rd[20]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(i_data_Rd[19]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(i_data_Rd[18]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(i_data_Rd[17]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(i_data_Rd[16]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(i_data_Rd[15]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(i_data_Rd[13]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(i_data_Rd[12]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(i_data_Rd[11]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(i_data_Rd[10]), .E(n115), .C(i_clk), .RN(i_rst_n), .Q(regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(i_data_Rd[9]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(i_data_Rd[8]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(i_data_Rd[7]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(i_data_Rd[6]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(i_data_Rd[5]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(i_data_Rd[4]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(i_data_Rd[3]), .E(n115), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(i_data_Rd[2]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(i_data_Rd[1]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(i_data_Rd[0]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[352]) );
  DFEC1 regs_reg_10__31_ ( .D(i_data_Rd[31]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(i_data_Rd[30]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(i_data_Rd[29]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(i_data_Rd[28]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(i_data_Rd[27]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(i_data_Rd[26]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(i_data_Rd[25]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(i_data_Rd[24]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(i_data_Rd[23]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(i_data_Rd[22]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(i_data_Rd[21]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(i_data_Rd[20]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(i_data_Rd[19]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(i_data_Rd[18]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(i_data_Rd[17]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(i_data_Rd[16]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(i_data_Rd[15]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(i_data_Rd[13]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(i_data_Rd[12]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(i_data_Rd[11]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n116), .C(i_clk), .RN(i_rst_n), .Q(regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(i_data_Rd[9]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(i_data_Rd[8]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(i_data_Rd[7]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(i_data_Rd[6]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(i_data_Rd[5]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(i_data_Rd[4]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(i_data_Rd[3]), .E(n116), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(i_data_Rd[2]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(i_data_Rd[1]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(i_data_Rd[0]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[320]) );
  DFEC1 regs_reg_9__31_ ( .D(i_data_Rd[31]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(i_data_Rd[30]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(i_data_Rd[29]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(i_data_Rd[28]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(i_data_Rd[27]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(i_data_Rd[26]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(i_data_Rd[25]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(i_data_Rd[24]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(i_data_Rd[23]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(i_data_Rd[22]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(i_data_Rd[21]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(i_data_Rd[20]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(i_data_Rd[19]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(i_data_Rd[18]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(i_data_Rd[17]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(i_data_Rd[16]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(i_data_Rd[15]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(i_data_Rd[14]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(i_data_Rd[13]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(i_data_Rd[12]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(i_data_Rd[11]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(i_data_Rd[10]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(i_data_Rd[9]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(i_data_Rd[8]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(i_data_Rd[7]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(i_data_Rd[6]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(i_data_Rd[5]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(i_data_Rd[4]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(i_data_Rd[3]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(i_data_Rd[2]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(i_data_Rd[1]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(i_data_Rd[0]), .E(n117), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[288]) );
  DFEC1 regs_reg_8__31_ ( .D(i_data_Rd[31]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(i_data_Rd[30]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(i_data_Rd[29]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(i_data_Rd[28]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(i_data_Rd[27]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(i_data_Rd[26]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(i_data_Rd[25]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(i_data_Rd[24]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(i_data_Rd[23]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(i_data_Rd[22]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(i_data_Rd[21]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(i_data_Rd[20]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(i_data_Rd[19]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(i_data_Rd[18]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(i_data_Rd[17]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(i_data_Rd[16]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(i_data_Rd[15]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(i_data_Rd[14]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(i_data_Rd[13]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(i_data_Rd[12]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(i_data_Rd[11]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(i_data_Rd[10]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(i_data_Rd[9]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(i_data_Rd[8]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(i_data_Rd[7]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(i_data_Rd[6]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(i_data_Rd[5]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(i_data_Rd[4]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(i_data_Rd[3]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(i_data_Rd[2]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(i_data_Rd[1]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(i_data_Rd[0]), .E(n118), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[256]) );
  DFEC1 regs_reg_7__31_ ( .D(i_data_Rd[31]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(i_data_Rd[30]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(i_data_Rd[29]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(i_data_Rd[28]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(i_data_Rd[27]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(i_data_Rd[26]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(i_data_Rd[25]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(i_data_Rd[24]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(i_data_Rd[23]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(i_data_Rd[22]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(i_data_Rd[21]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(i_data_Rd[20]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(i_data_Rd[19]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(i_data_Rd[18]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(i_data_Rd[17]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(i_data_Rd[16]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(i_data_Rd[15]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(i_data_Rd[14]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(i_data_Rd[13]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(i_data_Rd[12]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(i_data_Rd[11]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(i_data_Rd[10]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(i_data_Rd[9]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(i_data_Rd[8]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(i_data_Rd[7]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(i_data_Rd[6]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(i_data_Rd[5]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(i_data_Rd[4]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(i_data_Rd[3]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(i_data_Rd[2]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(i_data_Rd[1]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(i_data_Rd[0]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[224]) );
  DFEC1 regs_reg_6__31_ ( .D(i_data_Rd[31]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(i_data_Rd[30]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(i_data_Rd[29]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(i_data_Rd[28]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(i_data_Rd[27]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(i_data_Rd[26]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(i_data_Rd[25]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(i_data_Rd[24]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(i_data_Rd[23]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(i_data_Rd[22]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(i_data_Rd[21]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(i_data_Rd[20]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(i_data_Rd[19]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(i_data_Rd[18]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(i_data_Rd[17]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(i_data_Rd[16]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(i_data_Rd[15]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(i_data_Rd[14]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(i_data_Rd[13]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(i_data_Rd[12]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(i_data_Rd[11]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(i_data_Rd[10]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(i_data_Rd[9]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(i_data_Rd[8]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(i_data_Rd[7]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(i_data_Rd[6]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(i_data_Rd[5]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(i_data_Rd[4]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(i_data_Rd[3]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(i_data_Rd[2]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(i_data_Rd[1]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(i_data_Rd[0]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[192]) );
  DFEC1 regs_reg_5__31_ ( .D(i_data_Rd[31]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(i_data_Rd[30]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(i_data_Rd[29]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(i_data_Rd[28]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[188]) );
  DFEC1 regs_reg_5__27_ ( .D(i_data_Rd[27]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(i_data_Rd[26]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(i_data_Rd[25]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(i_data_Rd[24]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(i_data_Rd[23]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(i_data_Rd[22]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(i_data_Rd[21]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(i_data_Rd[20]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(i_data_Rd[19]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(i_data_Rd[18]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(i_data_Rd[17]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(i_data_Rd[16]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(i_data_Rd[15]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(i_data_Rd[14]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(i_data_Rd[13]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(i_data_Rd[12]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(i_data_Rd[11]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(i_data_Rd[10]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(i_data_Rd[9]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(i_data_Rd[8]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(i_data_Rd[7]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(i_data_Rd[6]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(i_data_Rd[5]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(i_data_Rd[4]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(i_data_Rd[3]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(i_data_Rd[2]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(i_data_Rd[1]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(i_data_Rd[0]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[160]) );
  DFEC1 regs_reg_4__31_ ( .D(i_data_Rd[31]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(i_data_Rd[30]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(i_data_Rd[29]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(i_data_Rd[28]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(i_data_Rd[27]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(i_data_Rd[26]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(i_data_Rd[25]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(i_data_Rd[24]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(i_data_Rd[23]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(i_data_Rd[22]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(i_data_Rd[21]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(i_data_Rd[20]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(i_data_Rd[19]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(i_data_Rd[18]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(i_data_Rd[17]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(i_data_Rd[16]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(i_data_Rd[15]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(i_data_Rd[14]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(i_data_Rd[13]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(i_data_Rd[12]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(i_data_Rd[11]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(i_data_Rd[10]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(i_data_Rd[9]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(i_data_Rd[8]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(i_data_Rd[7]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(i_data_Rd[6]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(i_data_Rd[5]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(i_data_Rd[4]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(i_data_Rd[3]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(i_data_Rd[2]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(i_data_Rd[1]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(i_data_Rd[0]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[128]) );
  DFEC1 regs_reg_3__31_ ( .D(i_data_Rd[31]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(i_data_Rd[30]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(i_data_Rd[29]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(i_data_Rd[28]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(i_data_Rd[27]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(i_data_Rd[26]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(i_data_Rd[25]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(i_data_Rd[24]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(i_data_Rd[23]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(i_data_Rd[22]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(i_data_Rd[21]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(i_data_Rd[20]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(i_data_Rd[19]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(i_data_Rd[18]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(i_data_Rd[17]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(i_data_Rd[16]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(i_data_Rd[15]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(i_data_Rd[14]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(i_data_Rd[13]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(i_data_Rd[12]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(i_data_Rd[11]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(i_data_Rd[10]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(i_data_Rd[9]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(i_data_Rd[8]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(i_data_Rd[7]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(i_data_Rd[6]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(i_data_Rd[5]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(i_data_Rd[4]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(i_data_Rd[3]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(i_data_Rd[2]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(i_data_Rd[1]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(i_data_Rd[0]), .E(n119), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[96]) );
  DFEC1 regs_reg_2__31_ ( .D(i_data_Rd[31]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(i_data_Rd[30]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(i_data_Rd[29]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(i_data_Rd[28]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(i_data_Rd[27]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(i_data_Rd[26]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(i_data_Rd[25]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(i_data_Rd[24]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(i_data_Rd[23]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(i_data_Rd[22]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(i_data_Rd[21]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(i_data_Rd[20]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(i_data_Rd[19]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(i_data_Rd[18]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(i_data_Rd[17]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(i_data_Rd[16]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(i_data_Rd[15]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(i_data_Rd[14]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(i_data_Rd[13]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(i_data_Rd[12]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(i_data_Rd[11]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(i_data_Rd[10]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(i_data_Rd[9]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(i_data_Rd[8]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(i_data_Rd[7]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(i_data_Rd[6]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(i_data_Rd[5]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(i_data_Rd[4]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(i_data_Rd[3]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(i_data_Rd[2]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(i_data_Rd[1]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(i_data_Rd[0]), .E(n120), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[64]) );
  DFEC1 regs_reg_1__31_ ( .D(n1), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(n64), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(n63), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(n62), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(n61), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(n60), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(n59), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(n58), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(n57), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(n56), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(n55), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(n54), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(n53), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(n52), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(n51), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(n50), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(n49), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(n48), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(n47), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(n46), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(n45), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(n33), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(n24), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(n19), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(n14), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(n12), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(n10), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(n8), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(n7), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(n4), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(n3), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(n2), .E(n121), .C(i_clk), .RN(i_rst_n), .Q(
        regs[32]) );
  DFEC1 regs_reg_0__31_ ( .D(n1), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(n64), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(n63), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(n62), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(n61), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(n60), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(n59), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(n58), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(n57), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(n56), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(n55), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(n54), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(n53), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(n52), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(n51), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(n50), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(n49), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(n48), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(n47), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(n46), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(n45), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(n33), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(n24), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(n19), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(n14), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(n12), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(n10), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(
        regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(n8), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(n7), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(n4), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(n3), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(n2), .E(n122), .C(i_clk), .RN(i_rst_n), .Q(regs[0]) );
  MUX21 regs_reg_31__31__U4 ( .A(regs[1023]), .B(i_data_Rd[31]), .S(n31), .Q(
        n65) );
  DFC1 regs_reg_31__31_ ( .D(n65), .C(i_clk), .RN(i_rst_n), .Q(regs[1023]) );
  BUF6 U2 ( .A(n846), .Q(n68) );
  BUF6 U3 ( .A(n1568), .Q(n75) );
  NOR33 U4 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[2]), .C(n860), .Q(n1568) );
  BUF6 U5 ( .A(n1563), .Q(n72) );
  BUF6 U6 ( .A(n843), .Q(n70) );
  NOR32 U7 ( .A(i_addr_Rs[1]), .B(i_addr_Rs[2]), .C(n859), .Q(n1565) );
  BUF6 U8 ( .A(n1565), .Q(n74) );
  BUF6 U9 ( .A(n1562), .Q(n112) );
  BUF6 U10 ( .A(n1564), .Q(n113) );
  NOR31 U11 ( .A(i_addr_Rs[1]), .B(n859), .C(n857), .Q(n1561) );
  BUF6 U12 ( .A(n839), .Q(n66) );
  BUF6 U13 ( .A(n842), .Q(n111) );
  BUF2 U14 ( .A(i_data_Rd[31]), .Q(n1) );
  BUF2 U15 ( .A(i_data_Rd[0]), .Q(n2) );
  BUF2 U16 ( .A(i_data_Rd[1]), .Q(n3) );
  BUF2 U17 ( .A(i_data_Rd[2]), .Q(n4) );
  BUF2 U18 ( .A(i_data_Rd[3]), .Q(n7) );
  BUF2 U19 ( .A(i_data_Rd[4]), .Q(n8) );
  BUF2 U20 ( .A(i_data_Rd[5]), .Q(n10) );
  BUF2 U21 ( .A(i_data_Rd[6]), .Q(n12) );
  BUF2 U22 ( .A(i_data_Rd[7]), .Q(n14) );
  BUF2 U23 ( .A(i_data_Rd[8]), .Q(n19) );
  BUF2 U24 ( .A(i_data_Rd[9]), .Q(n24) );
  BUF2 U25 ( .A(i_data_Rd[10]), .Q(n33) );
  BUF2 U26 ( .A(i_data_Rd[11]), .Q(n45) );
  BUF2 U27 ( .A(i_data_Rd[12]), .Q(n46) );
  BUF2 U28 ( .A(i_data_Rd[13]), .Q(n47) );
  BUF2 U29 ( .A(i_data_Rd[14]), .Q(n48) );
  BUF2 U30 ( .A(i_data_Rd[15]), .Q(n49) );
  BUF2 U31 ( .A(i_data_Rd[16]), .Q(n50) );
  BUF2 U32 ( .A(i_data_Rd[17]), .Q(n51) );
  BUF2 U33 ( .A(i_data_Rd[18]), .Q(n52) );
  BUF2 U34 ( .A(i_data_Rd[19]), .Q(n53) );
  BUF2 U35 ( .A(i_data_Rd[20]), .Q(n54) );
  BUF2 U36 ( .A(i_data_Rd[21]), .Q(n55) );
  BUF2 U37 ( .A(i_data_Rd[22]), .Q(n56) );
  BUF2 U38 ( .A(i_data_Rd[23]), .Q(n57) );
  BUF2 U39 ( .A(i_data_Rd[24]), .Q(n58) );
  BUF2 U40 ( .A(i_data_Rd[25]), .Q(n59) );
  BUF2 U41 ( .A(i_data_Rd[26]), .Q(n60) );
  BUF2 U42 ( .A(i_data_Rd[27]), .Q(n61) );
  BUF2 U43 ( .A(i_data_Rd[28]), .Q(n62) );
  BUF2 U44 ( .A(i_data_Rd[29]), .Q(n63) );
  BUF2 U45 ( .A(i_data_Rd[30]), .Q(n64) );
  AOI221 U46 ( .A(n834), .B(n216), .C(n832), .D(n215), .Q(n228) );
  AOI221 U47 ( .A(n834), .B(n282), .C(n832), .D(n281), .Q(n294) );
  AOI220 U48 ( .A(n834), .B(n260), .C(n832), .D(n259), .Q(n272) );
  AOI221 U49 ( .A(n834), .B(n502), .C(n832), .D(n501), .Q(n514) );
  AOI221 U50 ( .A(n834), .B(n788), .C(n832), .D(n787), .Q(n800) );
  AOI221 U51 ( .A(n834), .B(n238), .C(n832), .D(n237), .Q(n250) );
  AOI221 U52 ( .A(n1556), .B(n1158), .C(n1554), .D(n1157), .Q(n1170) );
  AOI221 U53 ( .A(n1556), .B(n938), .C(n1554), .D(n937), .Q(n950) );
  AOI221 U54 ( .A(n834), .B(n370), .C(n832), .D(n369), .Q(n382) );
  AOI221 U55 ( .A(n1556), .B(n1378), .C(n1554), .D(n1377), .Q(n1390) );
  AOI220 U56 ( .A(n834), .B(n590), .C(n832), .D(n589), .Q(n602) );
  AOI221 U57 ( .A(n1556), .B(n916), .C(n1554), .D(n915), .Q(n928) );
  AOI221 U58 ( .A(n1556), .B(n1532), .C(n1554), .D(n1531), .Q(n1544) );
  AOI220 U59 ( .A(n834), .B(n568), .C(n832), .D(n567), .Q(n580) );
  AOI220 U60 ( .A(n834), .B(n700), .C(n832), .D(n699), .Q(n712) );
  AOI221 U61 ( .A(n834), .B(n304), .C(n832), .D(n303), .Q(n316) );
  AOI221 U62 ( .A(n1556), .B(n1555), .C(n1554), .D(n1553), .Q(n1578) );
  AOI221 U63 ( .A(n1556), .B(n1114), .C(n1554), .D(n1113), .Q(n1126) );
  AOI221 U64 ( .A(n1556), .B(n1356), .C(n1554), .D(n1355), .Q(n1368) );
  AOI221 U65 ( .A(n834), .B(n634), .C(n832), .D(n633), .Q(n646) );
  AOI221 U66 ( .A(n1556), .B(n1224), .C(n1554), .D(n1223), .Q(n1236) );
  AOI220 U67 ( .A(n834), .B(n172), .C(n832), .D(n171), .Q(n184) );
  AOI220 U68 ( .A(n834), .B(n149), .C(n832), .D(n148), .Q(n162) );
  AOI220 U69 ( .A(n834), .B(n194), .C(n832), .D(n193), .Q(n206) );
  AOI220 U70 ( .A(n1556), .B(n1004), .C(n1554), .D(n1003), .Q(n1016) );
  AOI221 U71 ( .A(n834), .B(n833), .C(n832), .D(n831), .Q(n856) );
  AOI221 U72 ( .A(n1556), .B(n1048), .C(n1554), .D(n1047), .Q(n1060) );
  AOI221 U73 ( .A(n1556), .B(n1444), .C(n1554), .D(n1443), .Q(n1456) );
  AOI221 U74 ( .A(n1556), .B(n1422), .C(n1554), .D(n1421), .Q(n1434) );
  AOI221 U75 ( .A(n1556), .B(n1466), .C(n1554), .D(n1465), .Q(n1478) );
  AOI221 U76 ( .A(n1556), .B(n1026), .C(n1554), .D(n1025), .Q(n1038) );
  AOI221 U77 ( .A(n1556), .B(n1180), .C(n1554), .D(n1179), .Q(n1192) );
  AOI220 U78 ( .A(n111), .B(regs[478]), .C(n67), .D(regs[414]), .Q(n807) );
  AOI221 U79 ( .A(n842), .B(regs[963]), .C(n67), .D(regs[899]), .Q(n209) );
  AOI220 U80 ( .A(regs[86]), .B(n1568), .C(regs[22]), .D(n114), .Q(n1361) );
  AOI220 U81 ( .A(n111), .B(regs[732]), .C(n67), .D(regs[668]), .Q(n769) );
  AOI220 U82 ( .A(regs[590]), .B(n1568), .C(regs[526]), .D(n114), .Q(n1181) );
  AOI221 U83 ( .A(n842), .B(regs[452]), .C(n67), .D(regs[388]), .Q(n235) );
  AOI221 U84 ( .A(n111), .B(regs[964]), .C(n67), .D(regs[900]), .Q(n231) );
  AOI220 U85 ( .A(n111), .B(regs[723]), .C(n841), .D(regs[659]), .Q(n571) );
  AOI220 U86 ( .A(n111), .B(regs[211]), .C(n67), .D(regs[147]), .Q(n575) );
  AOI220 U87 ( .A(regs[855]), .B(n1568), .C(regs[791]), .D(n114), .Q(n1369) );
  AOI220 U88 ( .A(n111), .B(regs[220]), .C(n67), .D(regs[156]), .Q(n773) );
  AOI220 U89 ( .A(n111), .B(regs[960]), .C(n841), .D(regs[896]), .Q(n141) );
  AOI221 U90 ( .A(n111), .B(regs[707]), .C(n67), .D(regs[643]), .Q(n219) );
  AOI220 U91 ( .A(regs[704]), .B(n111), .C(regs[640]), .D(n67), .Q(n153) );
  AOI220 U92 ( .A(n111), .B(regs[985]), .C(n841), .D(regs[921]), .Q(n693) );
  AOI220 U93 ( .A(n111), .B(regs[980]), .C(n67), .D(regs[916]), .Q(n583) );
  AOI221 U94 ( .A(regs[250]), .B(n112), .C(regs[186]), .D(n76), .Q(n1452) );
  AOI220 U95 ( .A(regs[735]), .B(n113), .C(regs[671]), .D(n72), .Q(n1559) );
  AOI220 U96 ( .A(regs[205]), .B(n113), .C(regs[141]), .D(n72), .Q(n1165) );
  AOI220 U97 ( .A(n111), .B(regs[467]), .C(n67), .D(regs[403]), .Q(n565) );
  AOI220 U98 ( .A(n111), .B(regs[728]), .C(n67), .D(regs[664]), .Q(n681) );
  AOI220 U99 ( .A(n111), .B(regs[729]), .C(n67), .D(regs[665]), .Q(n703) );
  AOI221 U100 ( .A(regs[996]), .B(n112), .C(regs[932]), .D(n76), .Q(n954) );
  AOI220 U101 ( .A(n111), .B(regs[979]), .C(n67), .D(regs[915]), .Q(n561) );
  AOI221 U102 ( .A(regs[1019]), .B(n112), .C(regs[955]), .D(n76), .Q(n1460) );
  AOI220 U103 ( .A(n111), .B(regs[734]), .C(n841), .D(regs[670]), .Q(n813) );
  AOI220 U104 ( .A(regs[249]), .B(n112), .C(regs[185]), .D(n1561), .Q(n1430)
         );
  AOI220 U105 ( .A(regs[760]), .B(n112), .C(regs[696]), .D(n76), .Q(n1404) );
  AOI220 U106 ( .A(n111), .B(regs[222]), .C(n67), .D(regs[158]), .Q(n817) );
  AOI221 U107 ( .A(regs[507]), .B(n112), .C(regs[443]), .D(n76), .Q(n1464) );
  AOI220 U108 ( .A(n111), .B(regs[991]), .C(n67), .D(regs[927]), .Q(n825) );
  AOI220 U109 ( .A(n111), .B(regs[479]), .C(n67), .D(regs[415]), .Q(n829) );
  NOR22 U110 ( .A(n1588), .B(n1581), .Q(n40) );
  NOR22 U111 ( .A(n1584), .B(n1581), .Q(n37) );
  AOI220 U112 ( .A(n111), .B(regs[735]), .C(n841), .D(regs[671]), .Q(n837) );
  AOI220 U113 ( .A(n111), .B(regs[210]), .C(n67), .D(regs[146]), .Q(n553) );
  AOI220 U114 ( .A(n111), .B(regs[722]), .C(n841), .D(regs[658]), .Q(n549) );
  AOI220 U115 ( .A(n111), .B(regs[466]), .C(n67), .D(regs[402]), .Q(n543) );
  AOI220 U116 ( .A(n111), .B(regs[986]), .C(n841), .D(regs[922]), .Q(n715) );
  BUF6 U117 ( .A(n844), .Q(n69) );
  AOI221 U118 ( .A(regs[224]), .B(n112), .C(regs[160]), .D(n76), .Q(n880) );
  NOR22 U119 ( .A(n1584), .B(n1582), .Q(n28) );
  BUF8 U120 ( .A(n845), .Q(n71) );
  NOR22 U121 ( .A(n1588), .B(n1582), .Q(n31) );
  NOR22 U122 ( .A(n1590), .B(n1582), .Q(n29) );
  NOR22 U123 ( .A(n1589), .B(n1582), .Q(n30) );
  BUF6 U124 ( .A(n841), .Q(n67) );
  AOI220 U125 ( .A(n834), .B(n458), .C(n832), .D(n457), .Q(n470) );
  AOI220 U126 ( .A(n834), .B(n480), .C(n832), .D(n479), .Q(n492) );
  AOI220 U127 ( .A(n834), .B(n436), .C(n832), .D(n435), .Q(n448) );
  AOI220 U128 ( .A(n834), .B(n766), .C(n832), .D(n765), .Q(n778) );
  AOI220 U129 ( .A(n1556), .B(n1246), .C(n1554), .D(n1245), .Q(n1258) );
  AOI220 U130 ( .A(n1556), .B(n1510), .C(n1554), .D(n1509), .Q(n1522) );
  AOI220 U131 ( .A(n1556), .B(n1290), .C(n1554), .D(n1289), .Q(n1302) );
  AOI220 U132 ( .A(n834), .B(n612), .C(n832), .D(n611), .Q(n624) );
  AOI220 U133 ( .A(n834), .B(n722), .C(n832), .D(n721), .Q(n734) );
  AOI220 U134 ( .A(n1556), .B(n1334), .C(n1554), .D(n1333), .Q(n1346) );
  AOI220 U135 ( .A(n834), .B(n656), .C(n832), .D(n655), .Q(n668) );
  AOI220 U136 ( .A(n1556), .B(n1268), .C(n1554), .D(n1267), .Q(n1280) );
  AOI220 U137 ( .A(n834), .B(n744), .C(n832), .D(n743), .Q(n756) );
  AOI220 U138 ( .A(n1556), .B(n1312), .C(n1554), .D(n1311), .Q(n1324) );
  AOI220 U139 ( .A(regs[490]), .B(n112), .C(regs[426]), .D(n76), .Q(n1090) );
  AOI220 U140 ( .A(regs[1002]), .B(n112), .C(regs[938]), .D(n76), .Q(n1086) );
  AOI220 U141 ( .A(regs[232]), .B(n112), .C(regs[168]), .D(n76), .Q(n1056) );
  AOI220 U142 ( .A(regs[764]), .B(n112), .C(regs[700]), .D(n76), .Q(n1492) );
  NOR22 U143 ( .A(n1591), .B(n1589), .Q(n9) );
  NOR22 U144 ( .A(n1591), .B(n1590), .Q(n6) );
  NOR22 U145 ( .A(n1581), .B(n1590), .Q(n38) );
  NOR22 U146 ( .A(n1581), .B(n1589), .Q(n39) );
  NOR22 U147 ( .A(n1591), .B(n1588), .Q(n11) );
  NOR22 U148 ( .A(n1591), .B(n1584), .Q(n5) );
  NOR22 U149 ( .A(i_addr_Rs[4]), .B(n865), .Q(n1554) );
  NOR22 U150 ( .A(i_addr_Rt_3_), .B(n150), .Q(n854) );
  NOR22 U151 ( .A(i_addr_Rt_4_), .B(n143), .Q(n832) );
  BUF6 U152 ( .A(n1566), .Q(n73) );
  BUF8 U153 ( .A(n1567), .Q(n114) );
  NOR22 U154 ( .A(n143), .B(n150), .Q(n834) );
  NAND22 U155 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[1]), .Q(n858) );
  INV3 U156 ( .A(i_addr_Rs[4]), .Q(n872) );
  NOR22 U157 ( .A(i_addr_Rs[3]), .B(i_addr_Rs[4]), .Q(n1574) );
  AOI220 U158 ( .A(n1556), .B(n1400), .C(n1554), .D(n1399), .Q(n1412) );
  AOI220 U159 ( .A(n1556), .B(n1488), .C(n1554), .D(n1487), .Q(n1500) );
  AOI220 U160 ( .A(n834), .B(n678), .C(n832), .D(n677), .Q(n690) );
  AOI220 U161 ( .A(n1556), .B(n1202), .C(n1554), .D(n1201), .Q(n1214) );
  AOI220 U162 ( .A(regs[1003]), .B(n112), .C(regs[939]), .D(n76), .Q(n1108) );
  AOI220 U163 ( .A(regs[234]), .B(n112), .C(regs[170]), .D(n76), .Q(n1100) );
  AOI220 U164 ( .A(regs[202]), .B(n113), .C(regs[138]), .D(n72), .Q(n1099) );
  AOI220 U165 ( .A(regs[1004]), .B(n112), .C(regs[940]), .D(n76), .Q(n1130) );
  AOI220 U166 ( .A(regs[972]), .B(n113), .C(regs[908]), .D(n1563), .Q(n1129)
         );
  AOI220 U167 ( .A(regs[997]), .B(n112), .C(regs[933]), .D(n76), .Q(n976) );
  AOI220 U168 ( .A(n110), .B(regs[1000]), .C(n66), .D(regs[936]), .Q(n320) );
  AOI220 U169 ( .A(regs[971]), .B(n113), .C(regs[907]), .D(n1563), .Q(n1107)
         );
  AOI220 U170 ( .A(regs[714]), .B(n113), .C(regs[650]), .D(n72), .Q(n1095) );
  AOI220 U171 ( .A(n110), .B(regs[999]), .C(n66), .D(regs[935]), .Q(n298) );
  AOI220 U172 ( .A(regs[459]), .B(n113), .C(regs[395]), .D(n1563), .Q(n1111)
         );
  AOI220 U173 ( .A(regs[746]), .B(n112), .C(regs[682]), .D(n76), .Q(n1096) );
  AOI220 U174 ( .A(regs[715]), .B(n113), .C(regs[651]), .D(n72), .Q(n1117) );
  AOI220 U175 ( .A(regs[203]), .B(n113), .C(regs[139]), .D(n1563), .Q(n1121)
         );
  AOI220 U176 ( .A(n110), .B(regs[743]), .C(n66), .D(regs[679]), .Q(n308) );
  AOI220 U177 ( .A(regs[1018]), .B(n112), .C(regs[954]), .D(n76), .Q(n1438) );
  AOI220 U178 ( .A(regs[706]), .B(n1564), .C(regs[642]), .D(n72), .Q(n919) );
  AOI220 U179 ( .A(regs[731]), .B(n113), .C(regs[667]), .D(n72), .Q(n1469) );
  AOI220 U180 ( .A(n110), .B(regs[511]), .C(n66), .D(regs[447]), .Q(n830) );
  AOI220 U181 ( .A(n110), .B(regs[1023]), .C(n66), .D(regs[959]), .Q(n826) );
  AOI220 U182 ( .A(n110), .B(regs[742]), .C(n66), .D(regs[678]), .Q(n286) );
  AOI220 U183 ( .A(regs[736]), .B(n110), .C(regs[672]), .D(n66), .Q(n154) );
  AOI220 U184 ( .A(n840), .B(regs[254]), .C(n66), .D(regs[190]), .Q(n818) );
  AOI220 U185 ( .A(n110), .B(regs[766]), .C(n66), .D(regs[702]), .Q(n814) );
  AOI220 U186 ( .A(regs[248]), .B(n112), .C(regs[184]), .D(n76), .Q(n1408) );
  AOI220 U187 ( .A(regs[217]), .B(n113), .C(regs[153]), .D(n72), .Q(n1429) );
  AOI220 U188 ( .A(n110), .B(regs[510]), .C(n66), .D(regs[446]), .Q(n808) );
  AOI220 U189 ( .A(regs[761]), .B(n112), .C(regs[697]), .D(n76), .Q(n1426) );
  AOI220 U190 ( .A(regs[730]), .B(n113), .C(regs[666]), .D(n72), .Q(n1447) );
  AOI220 U191 ( .A(regs[762]), .B(n112), .C(regs[698]), .D(n76), .Q(n1448) );
  AOI220 U192 ( .A(regs[505]), .B(n112), .C(regs[441]), .D(n76), .Q(n1420) );
  AOI220 U193 ( .A(n111), .B(regs[464]), .C(n67), .D(regs[400]), .Q(n499) );
  AOI221 U194 ( .A(regs[601]), .B(n75), .C(regs[537]), .D(n114), .Q(n1423) );
  AOI220 U195 ( .A(n111), .B(regs[977]), .C(n67), .D(regs[913]), .Q(n517) );
  AOI220 U196 ( .A(n111), .B(regs[961]), .C(n841), .D(regs[897]), .Q(n165) );
  AOI220 U197 ( .A(regs[504]), .B(n1562), .C(regs[440]), .D(n76), .Q(n1398) );
  AOI220 U198 ( .A(regs[1016]), .B(n112), .C(regs[952]), .D(n76), .Q(n1394) );
  AOI220 U199 ( .A(n111), .B(regs[203]), .C(n67), .D(regs[139]), .Q(n399) );
  AOI220 U200 ( .A(regs[611]), .B(n73), .C(regs[547]), .D(n74), .Q(n940) );
  AOI220 U201 ( .A(n840), .B(regs[1012]), .C(n66), .D(regs[948]), .Q(n584) );
  AOI220 U202 ( .A(regs[247]), .B(n112), .C(regs[183]), .D(n1561), .Q(n1386)
         );
  AOI220 U203 ( .A(n840), .B(regs[246]), .C(n66), .D(regs[182]), .Q(n642) );
  AOI220 U204 ( .A(n111), .B(regs[721]), .C(n67), .D(regs[657]), .Q(n527) );
  AOI220 U205 ( .A(n111), .B(regs[214]), .C(n67), .D(regs[150]), .Q(n641) );
  AOI220 U206 ( .A(n111), .B(regs[450]), .C(n67), .D(regs[386]), .Q(n191) );
  AOI220 U207 ( .A(n111), .B(regs[970]), .C(n67), .D(regs[906]), .Q(n363) );
  AOI220 U208 ( .A(n111), .B(regs[981]), .C(n67), .D(regs[917]), .Q(n605) );
  AOI220 U209 ( .A(regs[759]), .B(n112), .C(regs[695]), .D(n76), .Q(n1382) );
  AOI220 U210 ( .A(n111), .B(regs[465]), .C(n67), .D(regs[401]), .Q(n521) );
  AOI220 U211 ( .A(n111), .B(regs[209]), .C(n67), .D(regs[145]), .Q(n531) );
  AOI220 U212 ( .A(regs[612]), .B(n1566), .C(regs[548]), .D(n74), .Q(n962) );
  AOI220 U213 ( .A(n111), .B(regs[194]), .C(n67), .D(regs[130]), .Q(n201) );
  AOI220 U214 ( .A(n111), .B(regs[725]), .C(n67), .D(regs[661]), .Q(n615) );
  AOI220 U215 ( .A(n110), .B(regs[498]), .C(n66), .D(regs[434]), .Q(n544) );
  AOI220 U216 ( .A(n840), .B(regs[1011]), .C(n66), .D(regs[947]), .Q(n562) );
  AOI220 U217 ( .A(n111), .B(regs[199]), .C(n67), .D(regs[135]), .Q(n311) );
  AOI220 U218 ( .A(n842), .B(regs[459]), .C(n67), .D(regs[395]), .Q(n389) );
  AOI220 U219 ( .A(n111), .B(regs[978]), .C(n67), .D(regs[914]), .Q(n539) );
  AOI220 U220 ( .A(n842), .B(regs[971]), .C(n67), .D(regs[907]), .Q(n385) );
  AOI220 U221 ( .A(n110), .B(regs[499]), .C(n66), .D(regs[435]), .Q(n566) );
  AOI220 U222 ( .A(n111), .B(regs[448]), .C(n67), .D(regs[384]), .Q(n146) );
  AOI220 U223 ( .A(n842), .B(regs[460]), .C(n67), .D(regs[396]), .Q(n411) );
  AOI220 U224 ( .A(n110), .B(regs[755]), .C(n66), .D(regs[691]), .Q(n572) );
  AOI220 U225 ( .A(n842), .B(regs[972]), .C(n67), .D(regs[908]), .Q(n407) );
  AOI220 U226 ( .A(n111), .B(regs[192]), .C(n67), .D(regs[128]), .Q(n157) );
  AOI220 U227 ( .A(n840), .B(regs[243]), .C(n66), .D(regs[179]), .Q(n576) );
  AOI220 U228 ( .A(regs[605]), .B(n75), .C(regs[541]), .D(n114), .Q(n1511) );
  AOI220 U229 ( .A(n111), .B(regs[720]), .C(n67), .D(regs[656]), .Q(n505) );
  AOI220 U230 ( .A(n111), .B(regs[449]), .C(n67), .D(regs[385]), .Q(n169) );
  AOI220 U231 ( .A(regs[865]), .B(n73), .C(regs[801]), .D(n74), .Q(n886) );
  AOI220 U232 ( .A(n840), .B(regs[242]), .C(n66), .D(regs[178]), .Q(n554) );
  AOI220 U233 ( .A(n111), .B(regs[208]), .C(n67), .D(regs[144]), .Q(n509) );
  AOI220 U234 ( .A(n111), .B(regs[710]), .C(n67), .D(regs[646]), .Q(n285) );
  AOI220 U235 ( .A(n111), .B(regs[724]), .C(n67), .D(regs[660]), .Q(n593) );
  AOI220 U236 ( .A(regs[97]), .B(n73), .C(regs[33]), .D(n1565), .Q(n900) );
  AOI220 U237 ( .A(n110), .B(regs[754]), .C(n66), .D(regs[690]), .Q(n550) );
  AOI220 U238 ( .A(n111), .B(regs[193]), .C(n67), .D(regs[129]), .Q(n179) );
  AOI220 U239 ( .A(n111), .B(regs[715]), .C(n67), .D(regs[651]), .Q(n395) );
  AOI220 U240 ( .A(n111), .B(regs[711]), .C(n67), .D(regs[647]), .Q(n307) );
  AOI220 U241 ( .A(n111), .B(regs[212]), .C(n67), .D(regs[148]), .Q(n597) );
  AOI220 U242 ( .A(regs[106]), .B(n1566), .C(regs[42]), .D(n74), .Q(n1098) );
  AOI220 U243 ( .A(n111), .B(regs[456]), .C(n67), .D(regs[392]), .Q(n323) );
  AOI220 U244 ( .A(n111), .B(regs[968]), .C(n67), .D(regs[904]), .Q(n319) );
  AOI220 U245 ( .A(n840), .B(regs[1015]), .C(n66), .D(regs[951]), .Q(n650) );
  AOI220 U246 ( .A(n111), .B(regs[198]), .C(n67), .D(regs[134]), .Q(n289) );
  AOI220 U247 ( .A(n111), .B(regs[983]), .C(n67), .D(regs[919]), .Q(n649) );
  AOI220 U248 ( .A(n111), .B(regs[201]), .C(n67), .D(regs[137]), .Q(n355) );
  AOI220 U249 ( .A(regs[617]), .B(n73), .C(regs[553]), .D(n74), .Q(n1072) );
  AOI220 U250 ( .A(n111), .B(regs[713]), .C(n67), .D(regs[649]), .Q(n351) );
  AOI220 U251 ( .A(n110), .B(regs[503]), .C(n66), .D(regs[439]), .Q(n654) );
  AOI220 U252 ( .A(n842), .B(regs[451]), .C(n67), .D(regs[387]), .Q(n213) );
  AOI220 U253 ( .A(n111), .B(regs[471]), .C(n67), .D(regs[407]), .Q(n653) );
  AOI220 U254 ( .A(n111), .B(regs[457]), .C(n67), .D(regs[393]), .Q(n345) );
  AOI220 U255 ( .A(n111), .B(regs[969]), .C(n67), .D(regs[905]), .Q(n341) );
  AOI220 U256 ( .A(n840), .B(regs[759]), .C(n66), .D(regs[695]), .Q(n660) );
  AOI220 U257 ( .A(n842), .B(regs[202]), .C(n67), .D(regs[138]), .Q(n377) );
  AOI220 U258 ( .A(n111), .B(regs[727]), .C(n67), .D(regs[663]), .Q(n659) );
  AOI220 U259 ( .A(n111), .B(regs[714]), .C(n67), .D(regs[650]), .Q(n373) );
  AOI220 U260 ( .A(n840), .B(regs[1016]), .C(n66), .D(regs[952]), .Q(n672) );
  AOI220 U261 ( .A(n111), .B(regs[967]), .C(n67), .D(regs[903]), .Q(n297) );
  AOI220 U262 ( .A(n111), .B(regs[984]), .C(n67), .D(regs[920]), .Q(n671) );
  AOI220 U263 ( .A(regs[589]), .B(n75), .C(regs[525]), .D(n114), .Q(n1159) );
  AOI220 U264 ( .A(n111), .B(regs[200]), .C(n67), .D(regs[136]), .Q(n333) );
  AOI220 U265 ( .A(n111), .B(regs[455]), .C(n67), .D(regs[391]), .Q(n301) );
  AOI220 U266 ( .A(regs[874]), .B(n73), .C(regs[810]), .D(n1565), .Q(n1084) );
  AOI220 U267 ( .A(n111), .B(regs[712]), .C(n67), .D(regs[648]), .Q(n329) );
  AOI220 U268 ( .A(regs[362]), .B(n73), .C(regs[298]), .D(n1565), .Q(n1088) );
  AOI220 U269 ( .A(regs[618]), .B(n1566), .C(regs[554]), .D(n74), .Q(n1094) );
  AOI220 U270 ( .A(n111), .B(regs[982]), .C(n67), .D(regs[918]), .Q(n627) );
  AOI220 U271 ( .A(regs[81]), .B(n75), .C(regs[17]), .D(n114), .Q(n1251) );
  AOI220 U272 ( .A(n110), .B(regs[502]), .C(n66), .D(regs[438]), .Q(n632) );
  AOI220 U273 ( .A(regs[593]), .B(n1568), .C(regs[529]), .D(n114), .Q(n1247)
         );
  AOI220 U274 ( .A(n111), .B(regs[470]), .C(n67), .D(regs[406]), .Q(n631) );
  AOI220 U275 ( .A(n111), .B(regs[458]), .C(n67), .D(regs[394]), .Q(n367) );
  AOI220 U276 ( .A(regs[864]), .B(n73), .C(regs[800]), .D(n1565), .Q(n862) );
  AOI220 U277 ( .A(n111), .B(regs[962]), .C(n841), .D(regs[898]), .Q(n187) );
  AOI220 U278 ( .A(n840), .B(regs[758]), .C(n66), .D(regs[694]), .Q(n638) );
  AOI220 U279 ( .A(n111), .B(regs[726]), .C(n67), .D(regs[662]), .Q(n637) );
  AOI220 U280 ( .A(regs[876]), .B(n1566), .C(regs[812]), .D(n74), .Q(n1128) );
  AOI220 U281 ( .A(n840), .B(regs[247]), .C(n66), .D(regs[183]), .Q(n664) );
  AOI220 U282 ( .A(n111), .B(regs[215]), .C(n67), .D(regs[151]), .Q(n663) );
  AOI220 U283 ( .A(regs[104]), .B(n73), .C(regs[40]), .D(n1565), .Q(n1054) );
  AOI220 U284 ( .A(n111), .B(regs[195]), .C(n67), .D(regs[131]), .Q(n223) );
  NOR21 U285 ( .A(n1589), .B(n1587), .Q(n21) );
  NOR21 U286 ( .A(n1588), .B(n1587), .Q(n22) );
  NOR21 U287 ( .A(n1590), .B(n1587), .Q(n20) );
  NAND31 U288 ( .A(i_addr_Rd[0]), .B(n109), .C(n1585), .Q(n1590) );
  NOR21 U289 ( .A(i_addr_Rd[4]), .B(n1579), .Q(n1580) );
  NOR22 U290 ( .A(i_addr_Rs[3]), .B(n872), .Q(n1576) );
  NAND31 U291 ( .A(i_con_RegWr), .B(i_addr_Rd[4]), .C(n1583), .Q(n1587) );
  NAND31 U292 ( .A(i_addr_Rd[1]), .B(n109), .C(n1586), .Q(n1589) );
  NOR32 U293 ( .A(i_addr_Rs[0]), .B(n860), .C(n857), .Q(n1564) );
  NOR22 U294 ( .A(n858), .B(n857), .Q(n1562) );
  NOR22 U295 ( .A(n865), .B(n872), .Q(n1556) );
  NAND31 U296 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n109), .Q(n1588) );
  NOR23 U297 ( .A(i_addr_Rs[2]), .B(n858), .Q(n1566) );
  BUF6 U298 ( .A(n1561), .Q(n76) );
  INV3 U299 ( .A(i_addr_Rd[3]), .Q(n1583) );
  INV2 U300 ( .A(i_con_RegWr), .Q(n1579) );
  INV2 U301 ( .A(i_addr_Rs[1]), .Q(n860) );
  INV2 U302 ( .A(i_addr_Rs[0]), .Q(n859) );
  NOR22 U303 ( .A(i_addr_Rt_3_), .B(i_addr_Rt_4_), .Q(n852) );
  INV3 U304 ( .A(i_addr_Rt_4_), .Q(n150) );
  INV3 U305 ( .A(i_addr_Rt_3_), .Q(n143) );
  INV3 U306 ( .A(i_addr_Rs[3]), .Q(n865) );
  NAND31 U307 ( .A(i_addr_Rd[4]), .B(i_con_RegWr), .C(i_addr_Rd[3]), .Q(n1582)
         );
  BUF6 U308 ( .A(n840), .Q(n110) );
  NAND22 U309 ( .A(n1580), .B(i_addr_Rd[3]), .Q(n1591) );
  INV3 U310 ( .A(i_addr_Rd[1]), .Q(n1585) );
  INV3 U311 ( .A(i_addr_Rd[0]), .Q(n1586) );
  AOI220 U312 ( .A(n68), .B(regs[89]), .C(n71), .D(regs[25]), .Q(n705) );
  AOI220 U313 ( .A(n68), .B(regs[601]), .C(n71), .D(regs[537]), .Q(n701) );
  AOI220 U314 ( .A(n68), .B(regs[345]), .C(n71), .D(regs[281]), .Q(n695) );
  AOI220 U315 ( .A(n68), .B(regs[857]), .C(n71), .D(regs[793]), .Q(n691) );
  AOI220 U316 ( .A(n69), .B(regs[371]), .C(n70), .D(regs[307]), .Q(n564) );
  AOI220 U317 ( .A(n69), .B(regs[883]), .C(n70), .D(regs[819]), .Q(n560) );
  AOI220 U318 ( .A(n69), .B(regs[117]), .C(n70), .D(regs[53]), .Q(n618) );
  AOI220 U319 ( .A(n69), .B(regs[629]), .C(n70), .D(regs[565]), .Q(n614) );
  AOI220 U320 ( .A(n68), .B(regs[88]), .C(n71), .D(regs[24]), .Q(n683) );
  AOI220 U321 ( .A(n68), .B(regs[600]), .C(n71), .D(regs[536]), .Q(n679) );
  AOI220 U322 ( .A(n68), .B(regs[344]), .C(n71), .D(regs[280]), .Q(n673) );
  AOI220 U323 ( .A(n69), .B(regs[122]), .C(n70), .D(regs[58]), .Q(n728) );
  AOI220 U324 ( .A(n69), .B(regs[378]), .C(n70), .D(regs[314]), .Q(n718) );
  AOI220 U325 ( .A(n68), .B(regs[858]), .C(n71), .D(regs[794]), .Q(n713) );
  AOI220 U326 ( .A(n68), .B(regs[75]), .C(n71), .D(regs[11]), .Q(n397) );
  AOI220 U327 ( .A(n69), .B(regs[107]), .C(n70), .D(regs[43]), .Q(n398) );
  AOI220 U328 ( .A(n68), .B(regs[587]), .C(n71), .D(regs[523]), .Q(n393) );
  AOI220 U329 ( .A(n69), .B(regs[619]), .C(n70), .D(regs[555]), .Q(n394) );
  AOI220 U330 ( .A(n68), .B(regs[331]), .C(n71), .D(regs[267]), .Q(n387) );
  AOI220 U331 ( .A(n69), .B(regs[363]), .C(n843), .D(regs[299]), .Q(n388) );
  AOI220 U332 ( .A(n68), .B(regs[843]), .C(n71), .D(regs[779]), .Q(n383) );
  AOI220 U333 ( .A(n69), .B(regs[875]), .C(n70), .D(regs[811]), .Q(n384) );
  AOI220 U334 ( .A(n69), .B(regs[108]), .C(n70), .D(regs[44]), .Q(n420) );
  AOI220 U335 ( .A(n69), .B(regs[620]), .C(n70), .D(regs[556]), .Q(n416) );
  AOI220 U336 ( .A(n68), .B(regs[332]), .C(n71), .D(regs[268]), .Q(n409) );
  AOI220 U337 ( .A(n69), .B(regs[364]), .C(n843), .D(regs[300]), .Q(n410) );
  AOI220 U338 ( .A(n68), .B(regs[844]), .C(n71), .D(regs[780]), .Q(n405) );
  AOI220 U339 ( .A(n69), .B(regs[876]), .C(n70), .D(regs[812]), .Q(n406) );
  AOI220 U340 ( .A(n69), .B(regs[109]), .C(n70), .D(regs[45]), .Q(n442) );
  AOI220 U341 ( .A(n69), .B(regs[621]), .C(n70), .D(regs[557]), .Q(n438) );
  AOI220 U342 ( .A(n69), .B(regs[365]), .C(n70), .D(regs[301]), .Q(n432) );
  AOI220 U343 ( .A(n69), .B(regs[877]), .C(n70), .D(regs[813]), .Q(n428) );
  AOI220 U344 ( .A(n69), .B(regs[628]), .C(n70), .D(regs[564]), .Q(n592) );
  AOI220 U345 ( .A(n69), .B(regs[372]), .C(n70), .D(regs[308]), .Q(n586) );
  AOI220 U346 ( .A(n69), .B(regs[884]), .C(n70), .D(regs[820]), .Q(n582) );
  AOI220 U347 ( .A(n69), .B(regs[111]), .C(n70), .D(regs[47]), .Q(n486) );
  AOI221 U348 ( .A(n68), .B(regs[591]), .C(n71), .D(regs[527]), .Q(n481) );
  AOI220 U349 ( .A(n69), .B(regs[623]), .C(n70), .D(regs[559]), .Q(n482) );
  AOI221 U350 ( .A(n68), .B(regs[335]), .C(n71), .D(regs[271]), .Q(n475) );
  AOI220 U351 ( .A(n69), .B(regs[367]), .C(n70), .D(regs[303]), .Q(n476) );
  AOI221 U352 ( .A(n68), .B(regs[847]), .C(n71), .D(regs[783]), .Q(n471) );
  AOI220 U353 ( .A(n69), .B(regs[879]), .C(n70), .D(regs[815]), .Q(n472) );
  AOI220 U354 ( .A(n69), .B(regs[886]), .C(n70), .D(regs[822]), .Q(n626) );
  AOI220 U355 ( .A(n69), .B(regs[114]), .C(n70), .D(regs[50]), .Q(n552) );
  AOI220 U356 ( .A(n69), .B(regs[626]), .C(n70), .D(regs[562]), .Q(n548) );
  AOI220 U357 ( .A(n69), .B(regs[370]), .C(n70), .D(regs[306]), .Q(n542) );
  AOI220 U358 ( .A(n69), .B(regs[882]), .C(n70), .D(regs[818]), .Q(n538) );
  AOI220 U359 ( .A(n68), .B(regs[73]), .C(n71), .D(regs[9]), .Q(n353) );
  AOI220 U360 ( .A(n68), .B(regs[585]), .C(n71), .D(regs[521]), .Q(n349) );
  AOI220 U361 ( .A(n69), .B(regs[617]), .C(n70), .D(regs[553]), .Q(n350) );
  AOI220 U362 ( .A(n68), .B(regs[329]), .C(n71), .D(regs[265]), .Q(n343) );
  AOI220 U363 ( .A(n68), .B(regs[841]), .C(n71), .D(regs[777]), .Q(n339) );
  AOI220 U364 ( .A(n69), .B(regs[112]), .C(n70), .D(regs[48]), .Q(n508) );
  AOI220 U365 ( .A(n69), .B(regs[624]), .C(n70), .D(regs[560]), .Q(n504) );
  AOI220 U366 ( .A(n69), .B(regs[368]), .C(n70), .D(regs[304]), .Q(n498) );
  AOI220 U367 ( .A(n69), .B(regs[880]), .C(n70), .D(regs[816]), .Q(n494) );
  AOI220 U368 ( .A(n68), .B(regs[72]), .C(n71), .D(regs[8]), .Q(n331) );
  AOI220 U369 ( .A(n68), .B(regs[584]), .C(n71), .D(regs[520]), .Q(n327) );
  AOI220 U370 ( .A(n69), .B(regs[616]), .C(n70), .D(regs[552]), .Q(n328) );
  AOI221 U371 ( .A(n68), .B(regs[328]), .C(n71), .D(regs[264]), .Q(n321) );
  AOI220 U372 ( .A(n69), .B(regs[360]), .C(n70), .D(regs[296]), .Q(n322) );
  AOI221 U373 ( .A(n68), .B(regs[840]), .C(n71), .D(regs[776]), .Q(n317) );
  AOI220 U374 ( .A(n69), .B(regs[872]), .C(n843), .D(regs[808]), .Q(n318) );
  AOI220 U375 ( .A(n68), .B(regs[330]), .C(n71), .D(regs[266]), .Q(n365) );
  AOI220 U376 ( .A(n68), .B(regs[842]), .C(n71), .D(regs[778]), .Q(n361) );
  AOI220 U377 ( .A(n68), .B(regs[92]), .C(n71), .D(regs[28]), .Q(n771) );
  AOI220 U378 ( .A(n69), .B(regs[124]), .C(n70), .D(regs[60]), .Q(n772) );
  AOI220 U379 ( .A(n68), .B(regs[604]), .C(n71), .D(regs[540]), .Q(n767) );
  AOI220 U380 ( .A(n69), .B(regs[636]), .C(n70), .D(regs[572]), .Q(n768) );
  AOI220 U381 ( .A(n68), .B(regs[348]), .C(n71), .D(regs[284]), .Q(n761) );
  AOI220 U382 ( .A(n69), .B(regs[380]), .C(n70), .D(regs[316]), .Q(n762) );
  AOI220 U383 ( .A(n69), .B(regs[892]), .C(n70), .D(regs[828]), .Q(n758) );
  AOI221 U384 ( .A(n68), .B(regs[71]), .C(n71), .D(regs[7]), .Q(n309) );
  AOI221 U385 ( .A(n68), .B(regs[583]), .C(n71), .D(regs[519]), .Q(n305) );
  AOI221 U386 ( .A(n68), .B(regs[327]), .C(n71), .D(regs[263]), .Q(n299) );
  AOI221 U387 ( .A(n68), .B(regs[839]), .C(n71), .D(regs[775]), .Q(n295) );
  AOI220 U388 ( .A(n69), .B(regs[871]), .C(n70), .D(regs[807]), .Q(n296) );
  AOI220 U389 ( .A(n69), .B(regs[356]), .C(n70), .D(regs[292]), .Q(n234) );
  AOI220 U390 ( .A(n68), .B(regs[93]), .C(n71), .D(regs[29]), .Q(n793) );
  AOI220 U391 ( .A(n69), .B(regs[125]), .C(n70), .D(regs[61]), .Q(n794) );
  AOI220 U392 ( .A(n68), .B(regs[605]), .C(n71), .D(regs[541]), .Q(n789) );
  AOI220 U393 ( .A(n69), .B(regs[637]), .C(n70), .D(regs[573]), .Q(n790) );
  AOI220 U394 ( .A(n68), .B(regs[349]), .C(n71), .D(regs[285]), .Q(n783) );
  AOI220 U395 ( .A(n69), .B(regs[381]), .C(n70), .D(regs[317]), .Q(n784) );
  AOI220 U396 ( .A(n68), .B(regs[861]), .C(n71), .D(regs[797]), .Q(n779) );
  AOI220 U397 ( .A(n69), .B(regs[893]), .C(n70), .D(regs[829]), .Q(n780) );
  AOI220 U398 ( .A(n68), .B(regs[65]), .C(n71), .D(regs[1]), .Q(n177) );
  AOI220 U399 ( .A(n69), .B(regs[97]), .C(n70), .D(regs[33]), .Q(n178) );
  AOI220 U400 ( .A(n68), .B(regs[577]), .C(n71), .D(regs[513]), .Q(n173) );
  AOI220 U401 ( .A(n69), .B(regs[609]), .C(n70), .D(regs[545]), .Q(n174) );
  AOI220 U402 ( .A(n68), .B(regs[321]), .C(n71), .D(regs[257]), .Q(n167) );
  AOI220 U403 ( .A(n69), .B(regs[353]), .C(n70), .D(regs[289]), .Q(n168) );
  AOI220 U404 ( .A(n68), .B(regs[833]), .C(n71), .D(regs[769]), .Q(n163) );
  AOI220 U405 ( .A(n69), .B(regs[865]), .C(n70), .D(regs[801]), .Q(n164) );
  AOI220 U406 ( .A(regs[193]), .B(n113), .C(regs[129]), .D(n72), .Q(n901) );
  AOI220 U407 ( .A(regs[225]), .B(n112), .C(regs[161]), .D(n1561), .Q(n902) );
  AOI220 U408 ( .A(regs[993]), .B(n112), .C(regs[929]), .D(n76), .Q(n888) );
  AOI220 U409 ( .A(regs[207]), .B(n113), .C(regs[143]), .D(n72), .Q(n1209) );
  AOI221 U410 ( .A(n68), .B(regs[70]), .C(n71), .D(regs[6]), .Q(n287) );
  AOI220 U411 ( .A(n69), .B(regs[102]), .C(n70), .D(regs[38]), .Q(n288) );
  AOI221 U412 ( .A(n68), .B(regs[582]), .C(n71), .D(regs[518]), .Q(n283) );
  AOI220 U413 ( .A(n69), .B(regs[614]), .C(n70), .D(regs[550]), .Q(n284) );
  AOI220 U414 ( .A(n69), .B(regs[99]), .C(n70), .D(regs[35]), .Q(n222) );
  AOI220 U415 ( .A(n69), .B(regs[611]), .C(n70), .D(regs[547]), .Q(n218) );
  AOI220 U416 ( .A(n69), .B(regs[867]), .C(n70), .D(regs[803]), .Q(n208) );
  AOI220 U417 ( .A(regs[107]), .B(n1566), .C(regs[43]), .D(n74), .Q(n1120) );
  AOI220 U418 ( .A(regs[235]), .B(n112), .C(regs[171]), .D(n76), .Q(n1122) );
  AOI220 U419 ( .A(regs[619]), .B(n1566), .C(regs[555]), .D(n74), .Q(n1116) );
  AOI220 U420 ( .A(regs[747]), .B(n112), .C(regs[683]), .D(n76), .Q(n1118) );
  AOI220 U421 ( .A(regs[363]), .B(n1566), .C(regs[299]), .D(n74), .Q(n1110) );
  AOI220 U422 ( .A(regs[491]), .B(n112), .C(regs[427]), .D(n76), .Q(n1112) );
  AOI220 U423 ( .A(regs[875]), .B(n1566), .C(regs[811]), .D(n74), .Q(n1106) );
  AOI220 U424 ( .A(regs[102]), .B(n1566), .C(regs[38]), .D(n1565), .Q(n1010)
         );
  AOI220 U425 ( .A(regs[230]), .B(n1562), .C(regs[166]), .D(n76), .Q(n1012) );
  AOI220 U426 ( .A(regs[614]), .B(n73), .C(regs[550]), .D(n74), .Q(n1006) );
  AOI220 U427 ( .A(regs[742]), .B(n1562), .C(regs[678]), .D(n1561), .Q(n1008)
         );
  AOI220 U428 ( .A(regs[358]), .B(n1566), .C(regs[294]), .D(n1565), .Q(n1000)
         );
  AOI220 U429 ( .A(regs[486]), .B(n1562), .C(regs[422]), .D(n76), .Q(n1002) );
  AOI220 U430 ( .A(regs[998]), .B(n1562), .C(regs[934]), .D(n1561), .Q(n998)
         );
  AOI220 U431 ( .A(regs[237]), .B(n112), .C(regs[173]), .D(n76), .Q(n1166) );
  AOI220 U432 ( .A(regs[717]), .B(n113), .C(regs[653]), .D(n72), .Q(n1161) );
  AOI220 U433 ( .A(regs[973]), .B(n113), .C(regs[909]), .D(n72), .Q(n1151) );
  AOI220 U434 ( .A(regs[1005]), .B(n112), .C(regs[941]), .D(n76), .Q(n1152) );
  AOI220 U435 ( .A(n68), .B(regs[66]), .C(n71), .D(regs[2]), .Q(n199) );
  AOI220 U436 ( .A(n68), .B(regs[578]), .C(n71), .D(regs[514]), .Q(n195) );
  AOI220 U437 ( .A(n69), .B(regs[610]), .C(n70), .D(regs[546]), .Q(n196) );
  AOI220 U438 ( .A(n68), .B(regs[322]), .C(n71), .D(regs[258]), .Q(n189) );
  AOI220 U439 ( .A(n69), .B(regs[354]), .C(n70), .D(regs[290]), .Q(n190) );
  AOI220 U440 ( .A(n68), .B(regs[834]), .C(n71), .D(regs[770]), .Q(n185) );
  AOI220 U441 ( .A(n69), .B(regs[866]), .C(n70), .D(regs[802]), .Q(n186) );
  AOI220 U442 ( .A(n69), .B(regs[101]), .C(n70), .D(regs[37]), .Q(n266) );
  AOI220 U443 ( .A(n69), .B(regs[869]), .C(n70), .D(regs[805]), .Q(n252) );
  AOI220 U444 ( .A(regs[721]), .B(n1564), .C(regs[657]), .D(n72), .Q(n1249) );
  AOI220 U445 ( .A(regs[465]), .B(n113), .C(regs[401]), .D(n72), .Q(n1243) );
  AOI220 U446 ( .A(regs[497]), .B(n112), .C(regs[433]), .D(n76), .Q(n1244) );
  AOI220 U447 ( .A(regs[103]), .B(n1566), .C(regs[39]), .D(n74), .Q(n1032) );
  AOI220 U448 ( .A(regs[199]), .B(n113), .C(regs[135]), .D(n1563), .Q(n1033)
         );
  AOI220 U449 ( .A(regs[231]), .B(n112), .C(regs[167]), .D(n76), .Q(n1034) );
  AOI220 U450 ( .A(regs[615]), .B(n1566), .C(regs[551]), .D(n74), .Q(n1028) );
  AOI220 U451 ( .A(regs[711]), .B(n113), .C(regs[647]), .D(n1563), .Q(n1029)
         );
  AOI220 U452 ( .A(regs[743]), .B(n1562), .C(regs[679]), .D(n76), .Q(n1030) );
  AOI220 U453 ( .A(regs[455]), .B(n113), .C(regs[391]), .D(n72), .Q(n1023) );
  AOI220 U454 ( .A(regs[487]), .B(n112), .C(regs[423]), .D(n76), .Q(n1024) );
  AOI220 U455 ( .A(regs[871]), .B(n1566), .C(regs[807]), .D(n74), .Q(n1018) );
  AOI220 U456 ( .A(regs[999]), .B(n112), .C(regs[935]), .D(n76), .Q(n1020) );
  AOI220 U457 ( .A(regs[616]), .B(n1566), .C(regs[552]), .D(n74), .Q(n1050) );
  AOI220 U458 ( .A(regs[712]), .B(n113), .C(regs[648]), .D(n1563), .Q(n1051)
         );
  AOI220 U459 ( .A(regs[744]), .B(n1562), .C(regs[680]), .D(n76), .Q(n1052) );
  AOI220 U460 ( .A(regs[360]), .B(n73), .C(regs[296]), .D(n74), .Q(n1044) );
  AOI220 U461 ( .A(regs[456]), .B(n113), .C(regs[392]), .D(n72), .Q(n1045) );
  AOI220 U462 ( .A(regs[488]), .B(n112), .C(regs[424]), .D(n76), .Q(n1046) );
  AOI220 U463 ( .A(regs[872]), .B(n1566), .C(regs[808]), .D(n74), .Q(n1040) );
  AOI220 U464 ( .A(regs[968]), .B(n113), .C(regs[904]), .D(n1563), .Q(n1041)
         );
  AOI220 U465 ( .A(regs[1000]), .B(n112), .C(regs[936]), .D(n76), .Q(n1042) );
  AOI220 U466 ( .A(n69), .B(regs[127]), .C(n70), .D(regs[63]), .Q(n848) );
  AOI220 U467 ( .A(n69), .B(regs[895]), .C(n70), .D(regs[831]), .Q(n824) );
  AOI220 U468 ( .A(n69), .B(regs[625]), .C(n70), .D(regs[561]), .Q(n526) );
  AOI221 U469 ( .A(n68), .B(regs[337]), .C(n71), .D(regs[273]), .Q(n519) );
  AOI220 U470 ( .A(n69), .B(regs[369]), .C(n70), .D(regs[305]), .Q(n520) );
  AOI220 U471 ( .A(n69), .B(regs[881]), .C(n70), .D(regs[817]), .Q(n516) );
  AOI220 U472 ( .A(n69), .B(regs[638]), .C(n70), .D(regs[574]), .Q(n812) );
  AOI220 U473 ( .A(n68), .B(regs[862]), .C(n71), .D(regs[798]), .Q(n801) );
  AOI220 U474 ( .A(n69), .B(regs[894]), .C(n70), .D(regs[830]), .Q(n802) );
  AOI220 U475 ( .A(n69), .B(regs[366]), .C(n70), .D(regs[302]), .Q(n454) );
  AOI220 U476 ( .A(regs[101]), .B(n1566), .C(regs[37]), .D(n74), .Q(n988) );
  AOI220 U477 ( .A(regs[229]), .B(n1562), .C(regs[165]), .D(n76), .Q(n990) );
  AOI220 U478 ( .A(regs[613]), .B(n73), .C(regs[549]), .D(n74), .Q(n984) );
  AOI220 U479 ( .A(regs[741]), .B(n1562), .C(regs[677]), .D(n1561), .Q(n986)
         );
  AOI220 U480 ( .A(regs[357]), .B(n73), .C(regs[293]), .D(n1565), .Q(n978) );
  AOI220 U481 ( .A(regs[485]), .B(n112), .C(regs[421]), .D(n76), .Q(n980) );
  AOI220 U482 ( .A(regs[469]), .B(n113), .C(regs[405]), .D(n72), .Q(n1331) );
  AOI220 U483 ( .A(regs[501]), .B(n112), .C(regs[437]), .D(n76), .Q(n1332) );
  AOI220 U484 ( .A(regs[981]), .B(n113), .C(regs[917]), .D(n72), .Q(n1327) );
  AOI220 U485 ( .A(regs[1013]), .B(n112), .C(regs[949]), .D(n76), .Q(n1328) );
  AOI220 U486 ( .A(regs[210]), .B(n113), .C(regs[146]), .D(n72), .Q(n1275) );
  AOI220 U487 ( .A(regs[242]), .B(n112), .C(regs[178]), .D(n76), .Q(n1276) );
  AOI220 U488 ( .A(regs[978]), .B(n113), .C(regs[914]), .D(n72), .Q(n1261) );
  AOI220 U489 ( .A(regs[1010]), .B(n112), .C(regs[946]), .D(n76), .Q(n1262) );
  AOI220 U490 ( .A(regs[223]), .B(n113), .C(regs[159]), .D(n72), .Q(n1571) );
  AOI220 U491 ( .A(regs[255]), .B(n112), .C(regs[191]), .D(n76), .Q(n1572) );
  AOI220 U492 ( .A(regs[767]), .B(n112), .C(regs[703]), .D(n76), .Q(n1560) );
  AOI220 U493 ( .A(regs[991]), .B(n113), .C(regs[927]), .D(n72), .Q(n1547) );
  AOI220 U494 ( .A(regs[222]), .B(n113), .C(regs[158]), .D(n72), .Q(n1539) );
  AOI220 U495 ( .A(regs[734]), .B(n113), .C(regs[670]), .D(n72), .Q(n1535) );
  AOI220 U496 ( .A(regs[478]), .B(n113), .C(regs[414]), .D(n72), .Q(n1529) );
  AOI220 U497 ( .A(regs[510]), .B(n112), .C(regs[446]), .D(n76), .Q(n1530) );
  AOI220 U498 ( .A(regs[105]), .B(n73), .C(regs[41]), .D(n1565), .Q(n1076) );
  AOI220 U499 ( .A(regs[233]), .B(n112), .C(regs[169]), .D(n76), .Q(n1078) );
  AOI220 U500 ( .A(regs[745]), .B(n1562), .C(regs[681]), .D(n76), .Q(n1074) );
  AOI220 U501 ( .A(regs[361]), .B(n73), .C(regs[297]), .D(n1565), .Q(n1066) );
  AOI220 U502 ( .A(regs[489]), .B(n112), .C(regs[425]), .D(n76), .Q(n1068) );
  AOI220 U503 ( .A(regs[873]), .B(n73), .C(regs[809]), .D(n1565), .Q(n1062) );
  AOI220 U504 ( .A(regs[1001]), .B(n112), .C(regs[937]), .D(n76), .Q(n1064) );
  AOI220 U505 ( .A(regs[732]), .B(n113), .C(regs[668]), .D(n72), .Q(n1491) );
  AOI220 U506 ( .A(n68), .B(regs[64]), .C(n71), .D(regs[0]), .Q(n155) );
  AOI220 U507 ( .A(n69), .B(regs[96]), .C(n70), .D(regs[32]), .Q(n156) );
  AOI220 U508 ( .A(regs[608]), .B(n69), .C(regs[544]), .D(n70), .Q(n152) );
  AOI220 U509 ( .A(n68), .B(regs[320]), .C(n71), .D(regs[256]), .Q(n144) );
  AOI220 U510 ( .A(n69), .B(regs[352]), .C(n70), .D(regs[288]), .Q(n145) );
  NOR31 U511 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .C(i_addr_Rt_2_), .Q(n845)
         );
  AOI220 U512 ( .A(n69), .B(regs[864]), .C(n70), .D(regs[800]), .Q(n140) );
  INV3 U513 ( .A(i_addr_Rt_1_), .Q(n138) );
  NAND22 U514 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .Q(n136) );
  AOI220 U515 ( .A(regs[221]), .B(n1564), .C(regs[157]), .D(n72), .Q(n1517) );
  AOI220 U516 ( .A(regs[733]), .B(n113), .C(regs[669]), .D(n72), .Q(n1513) );
  AOI220 U517 ( .A(regs[765]), .B(n112), .C(regs[701]), .D(n76), .Q(n1514) );
  AOI220 U518 ( .A(regs[477]), .B(n113), .C(regs[413]), .D(n72), .Q(n1507) );
  AOI220 U519 ( .A(regs[509]), .B(n112), .C(regs[445]), .D(n76), .Q(n1508) );
  AOI220 U520 ( .A(regs[989]), .B(n1564), .C(regs[925]), .D(n72), .Q(n1503) );
  AOI220 U521 ( .A(regs[99]), .B(n73), .C(regs[35]), .D(n74), .Q(n944) );
  AOI220 U522 ( .A(regs[483]), .B(n112), .C(regs[419]), .D(n1561), .Q(n936) );
  AOI220 U523 ( .A(regs[867]), .B(n73), .C(regs[803]), .D(n1565), .Q(n930) );
  AOI220 U524 ( .A(regs[995]), .B(n112), .C(regs[931]), .D(n76), .Q(n932) );
  AOI220 U525 ( .A(regs[100]), .B(n1566), .C(regs[36]), .D(n74), .Q(n966) );
  AOI220 U526 ( .A(regs[228]), .B(n112), .C(regs[164]), .D(n76), .Q(n968) );
  AOI220 U527 ( .A(regs[868]), .B(n73), .C(regs[804]), .D(n74), .Q(n952) );
  AOI220 U528 ( .A(regs[226]), .B(n1562), .C(regs[162]), .D(n76), .Q(n924) );
  AOI220 U529 ( .A(regs[738]), .B(n1562), .C(regs[674]), .D(n1561), .Q(n920)
         );
  AOI220 U530 ( .A(regs[482]), .B(n112), .C(regs[418]), .D(n76), .Q(n914) );
  AOI220 U531 ( .A(regs[994]), .B(n112), .C(regs[930]), .D(n76), .Q(n910) );
  AOI220 U532 ( .A(regs[736]), .B(n112), .C(regs[672]), .D(n76), .Q(n876) );
  AOI220 U533 ( .A(regs[480]), .B(n112), .C(regs[416]), .D(n76), .Q(n869) );
  AOI220 U534 ( .A(regs[992]), .B(n112), .C(regs[928]), .D(n76), .Q(n864) );
  AOI220 U535 ( .A(regs[467]), .B(n113), .C(regs[403]), .D(n72), .Q(n1287) );
  AOI220 U536 ( .A(regs[499]), .B(n112), .C(regs[435]), .D(n76), .Q(n1288) );
  AOI220 U537 ( .A(regs[979]), .B(n113), .C(regs[915]), .D(n72), .Q(n1283) );
  AOI220 U538 ( .A(regs[1011]), .B(n112), .C(regs[947]), .D(n76), .Q(n1284) );
  AOI220 U539 ( .A(regs[468]), .B(n1564), .C(regs[404]), .D(n72), .Q(n1309) );
  AOI220 U540 ( .A(regs[500]), .B(n1562), .C(regs[436]), .D(n76), .Q(n1310) );
  AOI220 U541 ( .A(regs[980]), .B(n1564), .C(regs[916]), .D(n72), .Q(n1305) );
  AOI220 U542 ( .A(regs[208]), .B(n113), .C(regs[144]), .D(n72), .Q(n1231) );
  AOI220 U543 ( .A(regs[240]), .B(n112), .C(regs[176]), .D(n76), .Q(n1232) );
  AOI220 U544 ( .A(regs[632]), .B(n73), .C(regs[568]), .D(n74), .Q(n1402) );
  AOI220 U545 ( .A(regs[728]), .B(n113), .C(regs[664]), .D(n72), .Q(n1403) );
  AOI220 U546 ( .A(regs[506]), .B(n112), .C(regs[442]), .D(n76), .Q(n1442) );
  AOI220 U547 ( .A(regs[251]), .B(n112), .C(regs[187]), .D(n76), .Q(n1474) );
  AOI220 U548 ( .A(regs[763]), .B(n112), .C(regs[699]), .D(n76), .Q(n1470) );
  AOI220 U549 ( .A(regs[475]), .B(n113), .C(regs[411]), .D(n72), .Q(n1463) );
  AOI220 U550 ( .A(n111), .B(regs[219]), .C(n67), .D(regs[155]), .Q(n751) );
  AOI220 U551 ( .A(n111), .B(regs[731]), .C(n841), .D(regs[667]), .Q(n747) );
  AOI220 U552 ( .A(n111), .B(regs[475]), .C(n67), .D(regs[411]), .Q(n741) );
  AOI220 U553 ( .A(n111), .B(regs[987]), .C(n841), .D(regs[923]), .Q(n737) );
  AOI220 U554 ( .A(n111), .B(regs[218]), .C(n67), .D(regs[154]), .Q(n729) );
  AOI220 U555 ( .A(n111), .B(regs[730]), .C(n841), .D(regs[666]), .Q(n725) );
  AOI220 U556 ( .A(n111), .B(regs[474]), .C(n67), .D(regs[410]), .Q(n719) );
  AOI220 U557 ( .A(n111), .B(regs[988]), .C(n841), .D(regs[924]), .Q(n759) );
  AOI220 U558 ( .A(n111), .B(regs[196]), .C(n67), .D(regs[132]), .Q(n245) );
  AOI220 U559 ( .A(n111), .B(regs[708]), .C(n67), .D(regs[644]), .Q(n241) );
  AOI220 U560 ( .A(n111), .B(regs[454]), .C(n67), .D(regs[390]), .Q(n279) );
  AOI220 U561 ( .A(n111), .B(regs[966]), .C(n67), .D(regs[902]), .Q(n275) );
  AOI220 U562 ( .A(n111), .B(regs[197]), .C(n67), .D(regs[133]), .Q(n267) );
  AOI220 U563 ( .A(n111), .B(regs[709]), .C(n841), .D(regs[645]), .Q(n263) );
  AOI220 U564 ( .A(n111), .B(regs[453]), .C(n67), .D(regs[389]), .Q(n257) );
  AOI220 U565 ( .A(n111), .B(regs[965]), .C(n841), .D(regs[901]), .Q(n253) );
  AOI220 U566 ( .A(n111), .B(regs[718]), .C(n67), .D(regs[654]), .Q(n461) );
  AOI221 U567 ( .A(n854), .B(n578), .C(n852), .D(n577), .Q(n579) );
  AOI221 U568 ( .A(n69), .B(regs[115]), .C(n70), .D(regs[51]), .Q(n574) );
  AOI221 U569 ( .A(n69), .B(regs[627]), .C(n70), .D(regs[563]), .Q(n570) );
  AOI221 U570 ( .A(n69), .B(regs[373]), .C(n70), .D(regs[309]), .Q(n608) );
  AOI221 U571 ( .A(n69), .B(regs[885]), .C(n70), .D(regs[821]), .Q(n604) );
  AOI221 U572 ( .A(n69), .B(regs[888]), .C(n70), .D(regs[824]), .Q(n670) );
  AOI221 U573 ( .A(n854), .B(n402), .C(n852), .D(n401), .Q(n403) );
  AOI221 U574 ( .A(n854), .B(n424), .C(n852), .D(n423), .Q(n425) );
  AOI221 U575 ( .A(n854), .B(n446), .C(n852), .D(n445), .Q(n447) );
  AOI221 U576 ( .A(n69), .B(regs[116]), .C(n70), .D(regs[52]), .Q(n596) );
  AOI221 U577 ( .A(n69), .B(regs[118]), .C(n70), .D(regs[54]), .Q(n640) );
  AOI221 U578 ( .A(n69), .B(regs[630]), .C(n70), .D(regs[566]), .Q(n636) );
  AOI221 U579 ( .A(n69), .B(regs[374]), .C(n70), .D(regs[310]), .Q(n630) );
  AOI221 U580 ( .A(n69), .B(regs[119]), .C(n70), .D(regs[55]), .Q(n662) );
  AOI221 U581 ( .A(n69), .B(regs[631]), .C(n70), .D(regs[567]), .Q(n658) );
  AOI221 U582 ( .A(n69), .B(regs[375]), .C(n70), .D(regs[311]), .Q(n652) );
  AOI221 U583 ( .A(n69), .B(regs[887]), .C(n70), .D(regs[823]), .Q(n648) );
  AOI221 U584 ( .A(n854), .B(n380), .C(n852), .D(n379), .Q(n381) );
  AOI221 U585 ( .A(n68), .B(regs[74]), .C(n71), .D(regs[10]), .Q(n375) );
  AOI221 U586 ( .A(n69), .B(regs[106]), .C(n843), .D(regs[42]), .Q(n376) );
  AOI221 U587 ( .A(n69), .B(regs[618]), .C(n70), .D(regs[554]), .Q(n372) );
  AOI220 U588 ( .A(regs[961]), .B(n113), .C(regs[897]), .D(n72), .Q(n887) );
  AOI221 U589 ( .A(n68), .B(regs[326]), .C(n71), .D(regs[262]), .Q(n277) );
  AOI221 U590 ( .A(n68), .B(regs[835]), .C(n71), .D(regs[771]), .Q(n207) );
  AOI221 U591 ( .A(n68), .B(regs[581]), .C(n71), .D(regs[517]), .Q(n261) );
  AOI221 U592 ( .A(n69), .B(regs[613]), .C(n70), .D(regs[549]), .Q(n262) );
  AOI221 U593 ( .A(n69), .B(regs[110]), .C(n70), .D(regs[46]), .Q(n464) );
  AOI221 U594 ( .A(n69), .B(regs[878]), .C(n70), .D(regs[814]), .Q(n450) );
  AOI220 U595 ( .A(regs[965]), .B(n113), .C(regs[901]), .D(n72), .Q(n975) );
  AOI221 U596 ( .A(regs[213]), .B(n113), .C(regs[149]), .D(n72), .Q(n1341) );
  AOI221 U597 ( .A(regs[245]), .B(n112), .C(regs[181]), .D(n76), .Q(n1342) );
  AOI221 U598 ( .A(regs[725]), .B(n113), .C(regs[661]), .D(n72), .Q(n1337) );
  AOI221 U599 ( .A(regs[757]), .B(n112), .C(regs[693]), .D(n76), .Q(n1338) );
  AOI220 U600 ( .A(regs[970]), .B(n1564), .C(regs[906]), .D(n72), .Q(n1085) );
  AOI220 U601 ( .A(regs[196]), .B(n113), .C(regs[132]), .D(n72), .Q(n967) );
  AOI220 U602 ( .A(regs[704]), .B(n113), .C(regs[640]), .D(n72), .Q(n875) );
  AOI220 U603 ( .A(regs[960]), .B(n113), .C(regs[896]), .D(n72), .Q(n863) );
  BUF2 U604 ( .A(n16), .Q(n132) );
  AOI221 U605 ( .A(n110), .B(regs[757]), .C(n66), .D(regs[693]), .Q(n616) );
  AOI220 U606 ( .A(regs[200]), .B(n113), .C(regs[136]), .D(n72), .Q(n1055) );
  AOI221 U607 ( .A(n68), .B(regs[351]), .C(n71), .D(regs[287]), .Q(n827) );
  AOI221 U608 ( .A(n68), .B(regs[863]), .C(n71), .D(regs[799]), .Q(n823) );
  AOI221 U609 ( .A(n69), .B(regs[622]), .C(n70), .D(regs[558]), .Q(n460) );
  AOI220 U610 ( .A(regs[201]), .B(n113), .C(regs[137]), .D(n72), .Q(n1077) );
  AOI220 U611 ( .A(regs[713]), .B(n1564), .C(regs[649]), .D(n72), .Q(n1073) );
  AOI220 U612 ( .A(regs[457]), .B(n113), .C(regs[393]), .D(n72), .Q(n1067) );
  AOI220 U613 ( .A(regs[969]), .B(n113), .C(regs[905]), .D(n72), .Q(n1063) );
  AOI221 U614 ( .A(n854), .B(n160), .C(n852), .D(n159), .Q(n161) );
  AOI220 U615 ( .A(regs[195]), .B(n113), .C(regs[131]), .D(n72), .Q(n945) );
  AOI220 U616 ( .A(regs[707]), .B(n113), .C(regs[643]), .D(n72), .Q(n941) );
  AOI220 U617 ( .A(regs[963]), .B(n113), .C(regs[899]), .D(n1563), .Q(n931) );
  AOI220 U618 ( .A(regs[458]), .B(n113), .C(regs[394]), .D(n72), .Q(n1089) );
  AOI220 U619 ( .A(regs[708]), .B(n113), .C(regs[644]), .D(n72), .Q(n963) );
  AOI220 U620 ( .A(regs[64]), .B(n1568), .C(regs[0]), .D(n114), .Q(n877) );
  AOI220 U621 ( .A(regs[448]), .B(n113), .C(regs[384]), .D(n72), .Q(n868) );
  AOI220 U622 ( .A(regs[592]), .B(n75), .C(regs[528]), .D(n114), .Q(n1225) );
  AOI220 U623 ( .A(regs[336]), .B(n1568), .C(regs[272]), .D(n114), .Q(n1219)
         );
  AOI221 U624 ( .A(regs[1017]), .B(n112), .C(regs[953]), .D(n76), .Q(n1416) );
  BUF2 U625 ( .A(n21), .Q(n128) );
  BUF2 U626 ( .A(n20), .Q(n129) );
  BUF2 U627 ( .A(n18), .Q(n130) );
  BUF2 U628 ( .A(n25), .Q(n125) );
  BUF2 U629 ( .A(n23), .Q(n126) );
  BUF2 U630 ( .A(n26), .Q(n124) );
  BUF2 U631 ( .A(n15), .Q(n133) );
  BUF2 U632 ( .A(n13), .Q(n134) );
  BUF2 U633 ( .A(n42), .Q(n117) );
  BUF2 U634 ( .A(n41), .Q(n118) );
  BUF2 U635 ( .A(n43), .Q(n116) );
  BUF2 U636 ( .A(n32), .Q(n122) );
  BUF2 U637 ( .A(n35), .Q(n120) );
  BUF2 U638 ( .A(n34), .Q(n121) );
  AOI221 U639 ( .A(n68), .B(regs[83]), .C(n71), .D(regs[19]), .Q(n573) );
  AOI221 U640 ( .A(n110), .B(regs[245]), .C(n66), .D(regs[181]), .Q(n620) );
  AOI221 U641 ( .A(n68), .B(regs[597]), .C(n71), .D(regs[533]), .Q(n613) );
  AOI221 U642 ( .A(n68), .B(regs[341]), .C(n71), .D(regs[277]), .Q(n607) );
  AOI221 U643 ( .A(n110), .B(regs[501]), .C(n66), .D(regs[437]), .Q(n610) );
  AOI221 U644 ( .A(n110), .B(regs[1013]), .C(n66), .D(regs[949]), .Q(n606) );
  AOI221 U645 ( .A(n68), .B(regs[856]), .C(n71), .D(regs[792]), .Q(n669) );
  AOI221 U646 ( .A(n110), .B(regs[244]), .C(n66), .D(regs[180]), .Q(n598) );
  AOI221 U647 ( .A(n68), .B(regs[596]), .C(n71), .D(regs[532]), .Q(n591) );
  AOI221 U648 ( .A(n110), .B(regs[756]), .C(n66), .D(regs[692]), .Q(n594) );
  AOI221 U649 ( .A(n110), .B(regs[500]), .C(n66), .D(regs[436]), .Q(n588) );
  AOI221 U650 ( .A(n68), .B(regs[852]), .C(n71), .D(regs[788]), .Q(n581) );
  AOI221 U651 ( .A(n110), .B(regs[239]), .C(n66), .D(regs[175]), .Q(n488) );
  AOI221 U652 ( .A(n110), .B(regs[751]), .C(n66), .D(regs[687]), .Q(n484) );
  AOI221 U653 ( .A(n68), .B(regs[86]), .C(n71), .D(regs[22]), .Q(n639) );
  AOI221 U654 ( .A(n68), .B(regs[598]), .C(n71), .D(regs[534]), .Q(n635) );
  AOI221 U655 ( .A(n68), .B(regs[342]), .C(n71), .D(regs[278]), .Q(n629) );
  AOI221 U656 ( .A(n110), .B(regs[1014]), .C(n66), .D(regs[950]), .Q(n628) );
  AOI221 U657 ( .A(n68), .B(regs[599]), .C(n71), .D(regs[535]), .Q(n657) );
  AOI221 U658 ( .A(n68), .B(regs[343]), .C(n71), .D(regs[279]), .Q(n651) );
  AOI221 U659 ( .A(n68), .B(regs[855]), .C(n71), .D(regs[791]), .Q(n647) );
  AOI221 U660 ( .A(n68), .B(regs[82]), .C(n71), .D(regs[18]), .Q(n551) );
  AOI221 U661 ( .A(n68), .B(regs[594]), .C(n71), .D(regs[530]), .Q(n547) );
  AOI221 U662 ( .A(n68), .B(regs[338]), .C(n71), .D(regs[274]), .Q(n541) );
  AOI221 U663 ( .A(n842), .B(regs[476]), .C(n67), .D(regs[412]), .Q(n763) );
  AOI221 U664 ( .A(n842), .B(regs[989]), .C(n67), .D(regs[925]), .Q(n781) );
  AOI220 U665 ( .A(regs[76]), .B(n1568), .C(regs[12]), .D(n114), .Q(n1141) );
  AOI220 U666 ( .A(regs[588]), .B(n1568), .C(regs[524]), .D(n114), .Q(n1137)
         );
  AOI220 U667 ( .A(regs[716]), .B(n1564), .C(regs[652]), .D(n72), .Q(n1139) );
  AOI220 U668 ( .A(regs[333]), .B(n1568), .C(regs[269]), .D(n114), .Q(n1153)
         );
  AOI220 U669 ( .A(regs[209]), .B(n1564), .C(regs[145]), .D(n72), .Q(n1253) );
  AOI220 U670 ( .A(regs[625]), .B(n1566), .C(regs[561]), .D(n74), .Q(n1248) );
  AOI220 U671 ( .A(regs[753]), .B(n1562), .C(regs[689]), .D(n76), .Q(n1250) );
  AOI220 U672 ( .A(regs[967]), .B(n113), .C(regs[903]), .D(n1563), .Q(n1019)
         );
  AOI221 U673 ( .A(n68), .B(regs[94]), .C(n71), .D(regs[30]), .Q(n815) );
  AOI221 U674 ( .A(n68), .B(regs[606]), .C(n71), .D(regs[542]), .Q(n811) );
  AOI221 U675 ( .A(n68), .B(regs[350]), .C(n71), .D(regs[286]), .Q(n805) );
  AOI221 U676 ( .A(n842), .B(regs[990]), .C(n67), .D(regs[926]), .Q(n803) );
  AOI220 U677 ( .A(n68), .B(regs[78]), .C(n71), .D(regs[14]), .Q(n463) );
  AOI220 U678 ( .A(regs[869]), .B(n1566), .C(regs[805]), .D(n74), .Q(n974) );
  AOI220 U679 ( .A(regs[117]), .B(n1566), .C(regs[53]), .D(n74), .Q(n1340) );
  AOI220 U680 ( .A(regs[629]), .B(n1566), .C(regs[565]), .D(n74), .Q(n1336) );
  AOI220 U681 ( .A(regs[373]), .B(n1566), .C(regs[309]), .D(n74), .Q(n1330) );
  AOI220 U682 ( .A(regs[885]), .B(n1566), .C(regs[821]), .D(n74), .Q(n1326) );
  AOI220 U683 ( .A(regs[114]), .B(n1566), .C(regs[50]), .D(n74), .Q(n1274) );
  AOI220 U684 ( .A(regs[626]), .B(n73), .C(regs[562]), .D(n74), .Q(n1270) );
  AOI220 U685 ( .A(regs[722]), .B(n1564), .C(regs[658]), .D(n72), .Q(n1271) );
  AOI220 U686 ( .A(regs[754]), .B(n1562), .C(regs[690]), .D(n76), .Q(n1272) );
  AOI220 U687 ( .A(regs[370]), .B(n73), .C(regs[306]), .D(n74), .Q(n1264) );
  AOI220 U688 ( .A(regs[466]), .B(n1564), .C(regs[402]), .D(n72), .Q(n1265) );
  AOI220 U689 ( .A(regs[498]), .B(n1562), .C(regs[434]), .D(n76), .Q(n1266) );
  AOI220 U690 ( .A(regs[882]), .B(n73), .C(regs[818]), .D(n74), .Q(n1260) );
  AOI220 U691 ( .A(regs[351]), .B(n1568), .C(regs[287]), .D(n114), .Q(n1549)
         );
  AOI220 U692 ( .A(regs[94]), .B(n1568), .C(regs[30]), .D(n114), .Q(n1537) );
  AOI220 U693 ( .A(regs[124]), .B(n73), .C(regs[60]), .D(n74), .Q(n1494) );
  AOI220 U694 ( .A(regs[220]), .B(n1564), .C(regs[156]), .D(n72), .Q(n1495) );
  AOI220 U695 ( .A(regs[252]), .B(n1562), .C(regs[188]), .D(n76), .Q(n1496) );
  AOI220 U696 ( .A(regs[636]), .B(n73), .C(regs[572]), .D(n74), .Q(n1490) );
  AOI220 U697 ( .A(regs[380]), .B(n1566), .C(regs[316]), .D(n74), .Q(n1484) );
  AOI220 U698 ( .A(regs[476]), .B(n1564), .C(regs[412]), .D(n72), .Q(n1485) );
  AOI220 U699 ( .A(regs[508]), .B(n1562), .C(regs[444]), .D(n76), .Q(n1486) );
  AOI220 U700 ( .A(regs[892]), .B(n73), .C(regs[828]), .D(n74), .Q(n1480) );
  AOI220 U701 ( .A(regs[988]), .B(n1564), .C(regs[924]), .D(n72), .Q(n1481) );
  AOI220 U702 ( .A(regs[1020]), .B(n1562), .C(regs[956]), .D(n76), .Q(n1482)
         );
  AOI221 U703 ( .A(regs[576]), .B(n68), .C(regs[512]), .D(n71), .Q(n151) );
  NOR31 U704 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_2_), .C(n138), .Q(n846) );
  NOR31 U705 ( .A(i_addr_Rt_1_), .B(i_addr_Rt_2_), .C(n137), .Q(n843) );
  NOR21 U706 ( .A(i_addr_Rt_2_), .B(n136), .Q(n844) );
  NOR31 U707 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .C(n135), .Q(n841) );
  NOR31 U708 ( .A(i_addr_Rt_0_), .B(n138), .C(n135), .Q(n842) );
  NOR21 U709 ( .A(n136), .B(n135), .Q(n840) );
  AOI220 U710 ( .A(regs[637]), .B(n1566), .C(regs[573]), .D(n74), .Q(n1512) );
  AOI220 U711 ( .A(regs[893]), .B(n1566), .C(regs[829]), .D(n74), .Q(n1502) );
  AOI220 U712 ( .A(regs[1021]), .B(n1562), .C(regs[957]), .D(n76), .Q(n1504)
         );
  AOI220 U713 ( .A(regs[451]), .B(n113), .C(regs[387]), .D(n72), .Q(n935) );
  AOI220 U714 ( .A(regs[74]), .B(n1568), .C(regs[10]), .D(n114), .Q(n1097) );
  AOI220 U715 ( .A(regs[586]), .B(n75), .C(regs[522]), .D(n114), .Q(n1093) );
  AOI220 U716 ( .A(regs[194]), .B(n1564), .C(regs[130]), .D(n72), .Q(n923) );
  AOI220 U717 ( .A(regs[450]), .B(n113), .C(regs[386]), .D(n1563), .Q(n913) );
  AOI220 U718 ( .A(regs[962]), .B(n113), .C(regs[898]), .D(n1563), .Q(n909) );
  AOI220 U719 ( .A(regs[352]), .B(n73), .C(regs[288]), .D(n74), .Q(n867) );
  AOI220 U720 ( .A(regs[115]), .B(n73), .C(regs[51]), .D(n74), .Q(n1296) );
  AOI220 U721 ( .A(regs[211]), .B(n1564), .C(regs[147]), .D(n72), .Q(n1297) );
  AOI220 U722 ( .A(regs[243]), .B(n1562), .C(regs[179]), .D(n76), .Q(n1298) );
  AOI220 U723 ( .A(regs[627]), .B(n73), .C(regs[563]), .D(n74), .Q(n1292) );
  AOI220 U724 ( .A(regs[723]), .B(n1564), .C(regs[659]), .D(n72), .Q(n1293) );
  AOI220 U725 ( .A(regs[755]), .B(n1562), .C(regs[691]), .D(n76), .Q(n1294) );
  AOI220 U726 ( .A(regs[371]), .B(n73), .C(regs[307]), .D(n74), .Q(n1286) );
  AOI220 U727 ( .A(regs[883]), .B(n1566), .C(regs[819]), .D(n74), .Q(n1282) );
  AOI220 U728 ( .A(regs[630]), .B(n1566), .C(regs[566]), .D(n74), .Q(n1358) );
  AOI220 U729 ( .A(regs[726]), .B(n1564), .C(regs[662]), .D(n72), .Q(n1359) );
  AOI220 U730 ( .A(regs[758]), .B(n1562), .C(regs[694]), .D(n76), .Q(n1360) );
  AOI220 U731 ( .A(regs[374]), .B(n1566), .C(regs[310]), .D(n74), .Q(n1352) );
  AOI220 U732 ( .A(regs[470]), .B(n113), .C(regs[406]), .D(n72), .Q(n1353) );
  AOI220 U733 ( .A(regs[502]), .B(n112), .C(regs[438]), .D(n76), .Q(n1354) );
  AOI220 U734 ( .A(regs[886]), .B(n1566), .C(regs[822]), .D(n74), .Q(n1348) );
  AOI220 U735 ( .A(regs[982]), .B(n113), .C(regs[918]), .D(n72), .Q(n1349) );
  AOI220 U736 ( .A(regs[1014]), .B(n1562), .C(regs[950]), .D(n76), .Q(n1350)
         );
  AOI220 U737 ( .A(regs[116]), .B(n1566), .C(regs[52]), .D(n74), .Q(n1318) );
  AOI220 U738 ( .A(regs[212]), .B(n1564), .C(regs[148]), .D(n72), .Q(n1319) );
  AOI220 U739 ( .A(regs[244]), .B(n1562), .C(regs[180]), .D(n76), .Q(n1320) );
  AOI220 U740 ( .A(regs[628]), .B(n1566), .C(regs[564]), .D(n74), .Q(n1314) );
  AOI220 U741 ( .A(regs[724]), .B(n1564), .C(regs[660]), .D(n72), .Q(n1315) );
  AOI220 U742 ( .A(regs[756]), .B(n1562), .C(regs[692]), .D(n76), .Q(n1316) );
  AOI220 U743 ( .A(regs[884]), .B(n1566), .C(regs[820]), .D(n74), .Q(n1304) );
  AOI220 U744 ( .A(regs[1012]), .B(n1562), .C(regs[948]), .D(n76), .Q(n1306)
         );
  AOI220 U745 ( .A(regs[720]), .B(n1564), .C(regs[656]), .D(n72), .Q(n1227) );
  AOI220 U746 ( .A(regs[464]), .B(n113), .C(regs[400]), .D(n72), .Q(n1221) );
  AOI220 U747 ( .A(regs[976]), .B(n113), .C(regs[912]), .D(n72), .Q(n1217) );
  AOI220 U748 ( .A(regs[344]), .B(n1568), .C(regs[280]), .D(n114), .Q(n1395)
         );
  AOI220 U749 ( .A(regs[599]), .B(n75), .C(regs[535]), .D(n114), .Q(n1379) );
  AOI220 U750 ( .A(regs[121]), .B(n73), .C(regs[57]), .D(n74), .Q(n1428) );
  AOI220 U751 ( .A(regs[729]), .B(n113), .C(regs[665]), .D(n72), .Q(n1425) );
  AOI220 U752 ( .A(regs[345]), .B(n1568), .C(regs[281]), .D(n114), .Q(n1417)
         );
  AOI220 U753 ( .A(regs[889]), .B(n73), .C(regs[825]), .D(n74), .Q(n1414) );
  AOI220 U754 ( .A(regs[602]), .B(n75), .C(regs[538]), .D(n114), .Q(n1445) );
  AOI220 U755 ( .A(regs[219]), .B(n113), .C(regs[155]), .D(n72), .Q(n1473) );
  AOI220 U756 ( .A(regs[635]), .B(n73), .C(regs[571]), .D(n74), .Q(n1468) );
  NOR31 U757 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[1]), .C(n857), .Q(n1563) );
  BUF2 U758 ( .A(n22), .Q(n127) );
  BUF2 U759 ( .A(n27), .Q(n123) );
  BUF2 U760 ( .A(n17), .Q(n131) );
  BUF2 U761 ( .A(i_addr_Rd[2]), .Q(n109) );
  AOI221 U762 ( .A(n68), .B(regs[595]), .C(n71), .D(regs[531]), .Q(n569) );
  AOI221 U763 ( .A(n68), .B(regs[339]), .C(n71), .D(regs[275]), .Q(n563) );
  AOI221 U764 ( .A(n68), .B(regs[851]), .C(n71), .D(regs[787]), .Q(n559) );
  AOI221 U765 ( .A(n834), .B(n392), .C(n832), .D(n391), .Q(n404) );
  AOI221 U766 ( .A(n834), .B(n414), .C(n832), .D(n413), .Q(n426) );
  AOI221 U767 ( .A(n110), .B(regs[495]), .C(n839), .D(regs[431]), .Q(n478) );
  AOI221 U768 ( .A(n110), .B(regs[1007]), .C(n66), .D(regs[943]), .Q(n474) );
  AOI221 U769 ( .A(n68), .B(regs[87]), .C(n71), .D(regs[23]), .Q(n661) );
  AOI221 U770 ( .A(n834), .B(n348), .C(n832), .D(n347), .Q(n360) );
  AOI221 U771 ( .A(n110), .B(regs[240]), .C(n66), .D(regs[176]), .Q(n510) );
  AOI221 U772 ( .A(n110), .B(regs[752]), .C(n66), .D(regs[688]), .Q(n506) );
  AOI221 U773 ( .A(n110), .B(regs[496]), .C(n839), .D(regs[432]), .Q(n500) );
  AOI221 U774 ( .A(n110), .B(regs[1008]), .C(n839), .D(regs[944]), .Q(n496) );
  AOI221 U775 ( .A(n68), .B(regs[586]), .C(n71), .D(regs[522]), .Q(n371) );
  AOI221 U776 ( .A(n111), .B(regs[221]), .C(n67), .D(regs[157]), .Q(n795) );
  AOI221 U777 ( .A(n111), .B(regs[733]), .C(n67), .D(regs[669]), .Q(n791) );
  AOI220 U778 ( .A(regs[622]), .B(n73), .C(regs[558]), .D(n74), .Q(n1182) );
  AOI220 U779 ( .A(regs[878]), .B(n73), .C(regs[814]), .D(n74), .Q(n1172) );
  AOI220 U780 ( .A(regs[577]), .B(n1568), .C(regs[513]), .D(n114), .Q(n895) );
  AOI220 U781 ( .A(regs[833]), .B(n1568), .C(regs[769]), .D(n114), .Q(n885) );
  AOI220 U782 ( .A(regs[111]), .B(n73), .C(regs[47]), .D(n74), .Q(n1208) );
  AOI220 U783 ( .A(regs[239]), .B(n112), .C(regs[175]), .D(n76), .Q(n1210) );
  AOI220 U784 ( .A(regs[623]), .B(n73), .C(regs[559]), .D(n74), .Q(n1204) );
  AOI220 U785 ( .A(regs[879]), .B(n73), .C(regs[815]), .D(n74), .Q(n1194) );
  AOI220 U786 ( .A(regs[108]), .B(n1566), .C(regs[44]), .D(n74), .Q(n1142) );
  AOI220 U787 ( .A(regs[620]), .B(n1566), .C(regs[556]), .D(n74), .Q(n1138) );
  AOI220 U788 ( .A(regs[748]), .B(n1562), .C(regs[684]), .D(n76), .Q(n1140) );
  AOI220 U789 ( .A(regs[332]), .B(n75), .C(regs[268]), .D(n114), .Q(n1131) );
  AOI220 U790 ( .A(regs[364]), .B(n73), .C(regs[300]), .D(n74), .Q(n1132) );
  AOI220 U791 ( .A(regs[844]), .B(n1568), .C(regs[780]), .D(n114), .Q(n1127)
         );
  AOI220 U792 ( .A(regs[109]), .B(n1566), .C(regs[45]), .D(n74), .Q(n1164) );
  AOI220 U793 ( .A(regs[621]), .B(n1566), .C(regs[557]), .D(n74), .Q(n1160) );
  AOI220 U794 ( .A(regs[749]), .B(n1562), .C(regs[685]), .D(n76), .Q(n1162) );
  AOI220 U795 ( .A(regs[365]), .B(n73), .C(regs[301]), .D(n74), .Q(n1154) );
  AOI220 U796 ( .A(regs[877]), .B(n1566), .C(regs[813]), .D(n74), .Q(n1150) );
  AOI220 U797 ( .A(regs[369]), .B(n1566), .C(regs[305]), .D(n74), .Q(n1242) );
  AOI220 U798 ( .A(regs[584]), .B(n1568), .C(regs[520]), .D(n114), .Q(n1049)
         );
  AOI221 U799 ( .A(n110), .B(regs[255]), .C(n66), .D(regs[191]), .Q(n850) );
  AOI220 U800 ( .A(regs[895]), .B(n73), .C(regs[831]), .D(n74), .Q(n1546) );
  AOI220 U801 ( .A(regs[1023]), .B(n112), .C(regs[959]), .D(n76), .Q(n1548) );
  AOI220 U802 ( .A(regs[126]), .B(n73), .C(regs[62]), .D(n74), .Q(n1538) );
  AOI220 U803 ( .A(regs[254]), .B(n112), .C(regs[190]), .D(n76), .Q(n1540) );
  AOI220 U804 ( .A(regs[638]), .B(n73), .C(regs[574]), .D(n74), .Q(n1534) );
  AOI220 U805 ( .A(regs[766]), .B(n112), .C(regs[702]), .D(n76), .Q(n1536) );
  AOI220 U806 ( .A(regs[382]), .B(n73), .C(regs[318]), .D(n74), .Q(n1528) );
  NOR31 U807 ( .A(i_addr_Rt_1_), .B(n137), .C(n135), .Q(n839) );
  AOI220 U808 ( .A(regs[125]), .B(n1566), .C(regs[61]), .D(n74), .Q(n1516) );
  AOI220 U809 ( .A(regs[253]), .B(n1562), .C(regs[189]), .D(n76), .Q(n1518) );
  AOI220 U810 ( .A(regs[579]), .B(n1568), .C(regs[515]), .D(n114), .Q(n939) );
  AOI220 U811 ( .A(regs[323]), .B(n75), .C(regs[259]), .D(n114), .Q(n933) );
  AOI220 U812 ( .A(regs[835]), .B(n75), .C(regs[771]), .D(n114), .Q(n929) );
  AOI220 U813 ( .A(regs[580]), .B(n75), .C(regs[516]), .D(n114), .Q(n961) );
  AOI220 U814 ( .A(regs[66]), .B(n75), .C(regs[2]), .D(n114), .Q(n921) );
  AOI220 U815 ( .A(regs[578]), .B(n75), .C(regs[514]), .D(n114), .Q(n917) );
  AOI220 U816 ( .A(regs[576]), .B(n75), .C(regs[512]), .D(n114), .Q(n873) );
  AOI220 U817 ( .A(regs[832]), .B(n75), .C(regs[768]), .D(n114), .Q(n861) );
  AOI220 U818 ( .A(regs[112]), .B(n1566), .C(regs[48]), .D(n74), .Q(n1230) );
  AOI220 U819 ( .A(regs[624]), .B(n73), .C(regs[560]), .D(n74), .Q(n1226) );
  AOI220 U820 ( .A(regs[752]), .B(n1562), .C(regs[688]), .D(n76), .Q(n1228) );
  AOI220 U821 ( .A(regs[368]), .B(n73), .C(regs[304]), .D(n74), .Q(n1220) );
  AOI220 U822 ( .A(regs[496]), .B(n112), .C(regs[432]), .D(n76), .Q(n1222) );
  AOI220 U823 ( .A(regs[880]), .B(n73), .C(regs[816]), .D(n74), .Q(n1216) );
  AOI220 U824 ( .A(regs[1008]), .B(n112), .C(regs[944]), .D(n76), .Q(n1218) );
  AOI220 U825 ( .A(regs[600]), .B(n75), .C(regs[536]), .D(n114), .Q(n1401) );
  AOI221 U826 ( .A(regs[503]), .B(n112), .C(regs[439]), .D(n76), .Q(n1376) );
  AOI221 U827 ( .A(regs[1015]), .B(n112), .C(regs[951]), .D(n76), .Q(n1372) );
  AOI220 U828 ( .A(regs[858]), .B(n1568), .C(regs[794]), .D(n114), .Q(n1435)
         );
  NOR40 U829 ( .A(i_addr_Rd[0]), .B(n109), .C(n1591), .D(n1585), .Q(n43) );
  BUF2 U830 ( .A(n44), .Q(n115) );
  NOR40 U831 ( .A(n109), .B(n1586), .C(n1591), .D(n1585), .Q(n44) );
  NOR40 U832 ( .A(i_addr_Rd[0]), .B(n109), .C(n1585), .D(n1581), .Q(n35) );
  BUF2 U833 ( .A(n36), .Q(n119) );
  NOR40 U834 ( .A(n109), .B(i_addr_Rd[1]), .C(n1586), .D(n1581), .Q(n34) );
  AOI220 U835 ( .A(n68), .B(regs[838]), .C(n71), .D(regs[774]), .Q(n273) );
  AOI220 U836 ( .A(regs[75]), .B(n1568), .C(regs[11]), .D(n114), .Q(n1119) );
  AOI220 U837 ( .A(regs[587]), .B(n1568), .C(regs[523]), .D(n114), .Q(n1115)
         );
  AOI220 U838 ( .A(regs[331]), .B(n1568), .C(regs[267]), .D(n114), .Q(n1109)
         );
  AOI220 U839 ( .A(regs[843]), .B(n1568), .C(regs[779]), .D(n114), .Q(n1105)
         );
  AOI220 U840 ( .A(regs[70]), .B(n75), .C(regs[6]), .D(n114), .Q(n1009) );
  AOI220 U841 ( .A(regs[582]), .B(n75), .C(regs[518]), .D(n114), .Q(n1005) );
  AOI220 U842 ( .A(regs[326]), .B(n75), .C(regs[262]), .D(n114), .Q(n999) );
  AOI220 U843 ( .A(regs[838]), .B(n75), .C(regs[774]), .D(n114), .Q(n995) );
  AOI220 U844 ( .A(regs[77]), .B(n75), .C(regs[13]), .D(n114), .Q(n1163) );
  AOI220 U845 ( .A(regs[71]), .B(n1568), .C(regs[7]), .D(n114), .Q(n1031) );
  AOI220 U846 ( .A(regs[583]), .B(n1568), .C(regs[519]), .D(n114), .Q(n1027)
         );
  AOI220 U847 ( .A(regs[327]), .B(n1568), .C(regs[263]), .D(n114), .Q(n1021)
         );
  AOI220 U848 ( .A(regs[359]), .B(n73), .C(regs[295]), .D(n74), .Q(n1022) );
  AOI220 U849 ( .A(regs[839]), .B(n1568), .C(regs[775]), .D(n114), .Q(n1017)
         );
  AOI220 U850 ( .A(regs[328]), .B(n1568), .C(regs[264]), .D(n114), .Q(n1043)
         );
  AOI220 U851 ( .A(regs[840]), .B(n1568), .C(regs[776]), .D(n114), .Q(n1039)
         );
  AOI221 U852 ( .A(n854), .B(n468), .C(n852), .D(n467), .Q(n469) );
  AOI220 U853 ( .A(n68), .B(regs[334]), .C(n71), .D(regs[270]), .Q(n453) );
  AOI220 U854 ( .A(n111), .B(regs[462]), .C(n67), .D(regs[398]), .Q(n455) );
  AOI220 U855 ( .A(n68), .B(regs[846]), .C(n71), .D(regs[782]), .Q(n449) );
  AOI220 U856 ( .A(n111), .B(regs[974]), .C(n67), .D(regs[910]), .Q(n451) );
  AOI220 U857 ( .A(regs[69]), .B(n1568), .C(regs[5]), .D(n114), .Q(n987) );
  AOI220 U858 ( .A(regs[581]), .B(n75), .C(regs[517]), .D(n114), .Q(n983) );
  AOI220 U859 ( .A(regs[325]), .B(n75), .C(regs[261]), .D(n114), .Q(n977) );
  AOI220 U860 ( .A(regs[95]), .B(n1568), .C(regs[31]), .D(n114), .Q(n1569) );
  AOI221 U861 ( .A(n1576), .B(n1542), .C(n1574), .D(n1541), .Q(n1543) );
  AOI220 U862 ( .A(regs[350]), .B(n75), .C(regs[286]), .D(n114), .Q(n1527) );
  AOI221 U863 ( .A(n1576), .B(n1498), .C(n1574), .D(n1497), .Q(n1499) );
  INV3 U864 ( .A(i_addr_Rt_2_), .Q(n135) );
  AOI221 U865 ( .A(n1576), .B(n1520), .C(n1574), .D(n1519), .Q(n1521) );
  AOI221 U866 ( .A(n1576), .B(n948), .C(n1574), .D(n947), .Q(n949) );
  AOI220 U867 ( .A(regs[355]), .B(n73), .C(regs[291]), .D(n1565), .Q(n934) );
  AOI221 U868 ( .A(n1576), .B(n1102), .C(n1574), .D(n1101), .Q(n1103) );
  AOI221 U869 ( .A(n1576), .B(n970), .C(n1574), .D(n969), .Q(n971) );
  AOI220 U870 ( .A(regs[356]), .B(n73), .C(regs[292]), .D(n74), .Q(n956) );
  AOI220 U871 ( .A(regs[836]), .B(n1568), .C(regs[772]), .D(n114), .Q(n951) );
  AOI221 U872 ( .A(n1576), .B(n926), .C(n1574), .D(n925), .Q(n927) );
  AOI220 U873 ( .A(regs[98]), .B(n73), .C(regs[34]), .D(n1565), .Q(n922) );
  AOI220 U874 ( .A(regs[610]), .B(n73), .C(regs[546]), .D(n1565), .Q(n918) );
  AOI220 U875 ( .A(regs[322]), .B(n75), .C(regs[258]), .D(n114), .Q(n911) );
  AOI220 U876 ( .A(regs[354]), .B(n73), .C(regs[290]), .D(n1565), .Q(n912) );
  AOI220 U877 ( .A(regs[834]), .B(n1568), .C(regs[770]), .D(n114), .Q(n907) );
  AOI220 U878 ( .A(regs[866]), .B(n73), .C(regs[802]), .D(n1565), .Q(n908) );
  AOI220 U879 ( .A(regs[320]), .B(n1568), .C(regs[256]), .D(n114), .Q(n866) );
  AOI220 U880 ( .A(regs[856]), .B(n75), .C(regs[792]), .D(n114), .Q(n1391) );
  AOI220 U881 ( .A(regs[87]), .B(n75), .C(regs[23]), .D(n114), .Q(n1383) );
  AOI220 U882 ( .A(regs[343]), .B(n75), .C(regs[279]), .D(n114), .Q(n1373) );
  AOI221 U883 ( .A(n1576), .B(n1432), .C(n1574), .D(n1431), .Q(n1433) );
  AOI220 U884 ( .A(regs[89]), .B(n75), .C(regs[25]), .D(n114), .Q(n1427) );
  AOI220 U885 ( .A(regs[633]), .B(n73), .C(regs[569]), .D(n74), .Q(n1424) );
  AOI221 U886 ( .A(n1576), .B(n1454), .C(n1574), .D(n1453), .Q(n1455) );
  AOI220 U887 ( .A(regs[122]), .B(n73), .C(regs[58]), .D(n74), .Q(n1450) );
  AOI220 U888 ( .A(regs[634]), .B(n73), .C(regs[570]), .D(n74), .Q(n1446) );
  AOI220 U889 ( .A(regs[378]), .B(n73), .C(regs[314]), .D(n74), .Q(n1440) );
  AOI220 U890 ( .A(regs[890]), .B(n1566), .C(regs[826]), .D(n74), .Q(n1436) );
  AOI221 U891 ( .A(n1576), .B(n1476), .C(n1574), .D(n1475), .Q(n1477) );
  AOI220 U892 ( .A(regs[91]), .B(n1568), .C(regs[27]), .D(n114), .Q(n1471) );
  AOI220 U893 ( .A(regs[123]), .B(n73), .C(regs[59]), .D(n1565), .Q(n1472) );
  AOI220 U894 ( .A(regs[347]), .B(n1568), .C(regs[283]), .D(n114), .Q(n1461)
         );
  AOI220 U895 ( .A(regs[891]), .B(n73), .C(regs[827]), .D(n74), .Q(n1458) );
  AOI220 U896 ( .A(regs[987]), .B(n113), .C(regs[923]), .D(n72), .Q(n1459) );
  NOR40 U897 ( .A(n109), .B(n1585), .C(n1586), .D(n1582), .Q(n27) );
  NOR40 U898 ( .A(n109), .B(i_addr_Rd[1]), .C(n1586), .D(n1582), .Q(n25) );
  NOR40 U899 ( .A(n109), .B(n1585), .C(n1586), .D(n1587), .Q(n17) );
  NOR40 U900 ( .A(n109), .B(i_addr_Rd[1]), .C(n1586), .D(n1587), .Q(n15) );
  NOR40 U901 ( .A(i_addr_Rd[1]), .B(n109), .C(n1586), .D(n1591), .Q(n42) );
  NOR40 U902 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n109), .D(n1581), .Q(n32) );
  NOR40 U903 ( .A(n109), .B(n1585), .C(n1586), .D(n1581), .Q(n36) );
  NAND22 U904 ( .A(n1580), .B(n1583), .Q(n1581) );
  AOI220 U905 ( .A(n69), .B(regs[633]), .C(n70), .D(regs[569]), .Q(n702) );
  AOI220 U906 ( .A(n69), .B(regs[377]), .C(n70), .D(regs[313]), .Q(n696) );
  AOI220 U907 ( .A(n69), .B(regs[889]), .C(n70), .D(regs[825]), .Q(n692) );
  AOI220 U908 ( .A(n68), .B(regs[91]), .C(n71), .D(regs[27]), .Q(n749) );
  AOI220 U909 ( .A(n68), .B(regs[603]), .C(n71), .D(regs[539]), .Q(n745) );
  AOI220 U910 ( .A(n69), .B(regs[635]), .C(n70), .D(regs[571]), .Q(n746) );
  AOI220 U911 ( .A(n68), .B(regs[347]), .C(n71), .D(regs[283]), .Q(n739) );
  AOI220 U912 ( .A(n69), .B(regs[379]), .C(n70), .D(regs[315]), .Q(n740) );
  AOI220 U913 ( .A(n68), .B(regs[859]), .C(n71), .D(regs[795]), .Q(n735) );
  AOI220 U914 ( .A(n69), .B(regs[120]), .C(n70), .D(regs[56]), .Q(n684) );
  AOI220 U915 ( .A(n69), .B(regs[632]), .C(n70), .D(regs[568]), .Q(n680) );
  AOI220 U916 ( .A(n69), .B(regs[376]), .C(n70), .D(regs[312]), .Q(n674) );
  AOI220 U917 ( .A(n68), .B(regs[90]), .C(n71), .D(regs[26]), .Q(n727) );
  AOI220 U918 ( .A(n68), .B(regs[602]), .C(n71), .D(regs[538]), .Q(n723) );
  AOI220 U919 ( .A(n69), .B(regs[634]), .C(n70), .D(regs[570]), .Q(n724) );
  AOI220 U920 ( .A(n68), .B(regs[346]), .C(n71), .D(regs[282]), .Q(n717) );
  AOI220 U921 ( .A(n69), .B(regs[890]), .C(n70), .D(regs[826]), .Q(n714) );
  AOI220 U922 ( .A(n68), .B(regs[76]), .C(n71), .D(regs[12]), .Q(n419) );
  AOI220 U923 ( .A(n68), .B(regs[588]), .C(n71), .D(regs[524]), .Q(n415) );
  AOI220 U924 ( .A(n68), .B(regs[77]), .C(n71), .D(regs[13]), .Q(n441) );
  AOI220 U925 ( .A(n68), .B(regs[589]), .C(n71), .D(regs[525]), .Q(n437) );
  AOI220 U926 ( .A(n68), .B(regs[333]), .C(n71), .D(regs[269]), .Q(n431) );
  AOI220 U927 ( .A(n68), .B(regs[845]), .C(n71), .D(regs[781]), .Q(n427) );
  AOI220 U928 ( .A(n68), .B(regs[79]), .C(n71), .D(regs[15]), .Q(n485) );
  AOI220 U929 ( .A(n69), .B(regs[361]), .C(n70), .D(regs[297]), .Q(n344) );
  AOI220 U930 ( .A(n69), .B(regs[873]), .C(n70), .D(regs[809]), .Q(n340) );
  AOI220 U931 ( .A(n68), .B(regs[592]), .C(n71), .D(regs[528]), .Q(n503) );
  AOI220 U932 ( .A(n68), .B(regs[848]), .C(n71), .D(regs[784]), .Q(n493) );
  AOI220 U933 ( .A(n69), .B(regs[362]), .C(n70), .D(regs[298]), .Q(n366) );
  AOI220 U934 ( .A(n69), .B(regs[874]), .C(n70), .D(regs[810]), .Q(n362) );
  AOI220 U935 ( .A(n68), .B(regs[860]), .C(n71), .D(regs[796]), .Q(n757) );
  AOI220 U936 ( .A(n69), .B(regs[103]), .C(n70), .D(regs[39]), .Q(n310) );
  AOI220 U937 ( .A(n69), .B(regs[359]), .C(n70), .D(regs[295]), .Q(n300) );
  AOI220 U938 ( .A(n69), .B(regs[100]), .C(n70), .D(regs[36]), .Q(n244) );
  AOI220 U939 ( .A(n68), .B(regs[580]), .C(n71), .D(regs[516]), .Q(n239) );
  AOI220 U940 ( .A(n68), .B(regs[324]), .C(n71), .D(regs[260]), .Q(n233) );
  AOI220 U941 ( .A(regs[65]), .B(n75), .C(regs[1]), .D(n114), .Q(n899) );
  AOI221 U942 ( .A(n1556), .B(n894), .C(n1554), .D(n893), .Q(n906) );
  AOI220 U943 ( .A(regs[321]), .B(n75), .C(regs[257]), .D(n114), .Q(n889) );
  AOI220 U944 ( .A(regs[79]), .B(n75), .C(regs[15]), .D(n114), .Q(n1207) );
  AOI220 U945 ( .A(regs[591]), .B(n75), .C(regs[527]), .D(n114), .Q(n1203) );
  AOI220 U946 ( .A(n68), .B(regs[67]), .C(n71), .D(regs[3]), .Q(n221) );
  AOI220 U947 ( .A(n68), .B(regs[579]), .C(n71), .D(regs[515]), .Q(n217) );
  AOI220 U948 ( .A(n68), .B(regs[323]), .C(n71), .D(regs[259]), .Q(n211) );
  AOI220 U949 ( .A(regs[845]), .B(n75), .C(regs[781]), .D(n114), .Q(n1149) );
  AOI220 U950 ( .A(n69), .B(regs[98]), .C(n70), .D(regs[34]), .Q(n200) );
  AOI220 U951 ( .A(n68), .B(regs[325]), .C(n71), .D(regs[261]), .Q(n255) );
  AOI220 U952 ( .A(n69), .B(regs[357]), .C(n70), .D(regs[293]), .Q(n256) );
  AOI220 U953 ( .A(regs[337]), .B(n75), .C(regs[273]), .D(n114), .Q(n1241) );
  AOI220 U954 ( .A(regs[849]), .B(n75), .C(regs[785]), .D(n114), .Q(n1237) );
  AOI220 U955 ( .A(regs[72]), .B(n75), .C(regs[8]), .D(n114), .Q(n1053) );
  AOI220 U956 ( .A(n68), .B(regs[95]), .C(n71), .D(regs[31]), .Q(n847) );
  AOI220 U957 ( .A(n68), .B(regs[81]), .C(n71), .D(regs[17]), .Q(n529) );
  AOI220 U958 ( .A(regs[837]), .B(n75), .C(regs[773]), .D(n114), .Q(n973) );
  AOI220 U959 ( .A(regs[85]), .B(n75), .C(regs[21]), .D(n114), .Q(n1339) );
  AOI220 U960 ( .A(regs[597]), .B(n1568), .C(regs[533]), .D(n114), .Q(n1335)
         );
  AOI220 U961 ( .A(regs[341]), .B(n75), .C(regs[277]), .D(n114), .Q(n1329) );
  AOI220 U962 ( .A(regs[853]), .B(n75), .C(regs[789]), .D(n114), .Q(n1325) );
  AOI220 U963 ( .A(regs[82]), .B(n1568), .C(regs[18]), .D(n114), .Q(n1273) );
  AOI220 U964 ( .A(regs[594]), .B(n75), .C(regs[530]), .D(n114), .Q(n1269) );
  AOI220 U965 ( .A(regs[338]), .B(n1568), .C(regs[274]), .D(n114), .Q(n1263)
         );
  AOI220 U966 ( .A(regs[607]), .B(n75), .C(regs[543]), .D(n114), .Q(n1557) );
  AOI220 U967 ( .A(regs[863]), .B(n75), .C(regs[799]), .D(n114), .Q(n1545) );
  AOI220 U968 ( .A(regs[73]), .B(n75), .C(regs[9]), .D(n114), .Q(n1075) );
  AOI220 U969 ( .A(regs[585]), .B(n75), .C(regs[521]), .D(n114), .Q(n1071) );
  AOI220 U970 ( .A(regs[329]), .B(n75), .C(regs[265]), .D(n114), .Q(n1065) );
  AOI220 U971 ( .A(regs[841]), .B(n75), .C(regs[777]), .D(n114), .Q(n1061) );
  AOI220 U972 ( .A(regs[604]), .B(n1568), .C(regs[540]), .D(n114), .Q(n1489)
         );
  AOI220 U973 ( .A(regs[860]), .B(n75), .C(regs[796]), .D(n114), .Q(n1479) );
  AOI220 U974 ( .A(regs[349]), .B(n75), .C(regs[285]), .D(n114), .Q(n1505) );
  AOI220 U975 ( .A(regs[861]), .B(n75), .C(regs[797]), .D(n114), .Q(n1501) );
  AOI221 U976 ( .A(n1556), .B(n1092), .C(n1554), .D(n1091), .Q(n1104) );
  AOI220 U977 ( .A(regs[330]), .B(n75), .C(regs[266]), .D(n114), .Q(n1087) );
  AOI220 U978 ( .A(regs[842]), .B(n75), .C(regs[778]), .D(n114), .Q(n1083) );
  AOI221 U979 ( .A(n1556), .B(n871), .C(n1554), .D(n870), .Q(n884) );
  AOI220 U980 ( .A(regs[83]), .B(n75), .C(regs[19]), .D(n114), .Q(n1295) );
  AOI220 U981 ( .A(regs[595]), .B(n1568), .C(regs[531]), .D(n114), .Q(n1291)
         );
  AOI220 U982 ( .A(regs[851]), .B(n75), .C(regs[787]), .D(n114), .Q(n1281) );
  AOI220 U983 ( .A(regs[214]), .B(n1564), .C(regs[150]), .D(n72), .Q(n1363) );
  AOI220 U984 ( .A(regs[598]), .B(n1568), .C(regs[534]), .D(n114), .Q(n1357)
         );
  AOI220 U985 ( .A(regs[342]), .B(n75), .C(regs[278]), .D(n114), .Q(n1351) );
  AOI220 U986 ( .A(regs[854]), .B(n75), .C(regs[790]), .D(n114), .Q(n1347) );
  AOI220 U987 ( .A(regs[84]), .B(n75), .C(regs[20]), .D(n114), .Q(n1317) );
  AOI220 U988 ( .A(regs[596]), .B(n1568), .C(regs[532]), .D(n114), .Q(n1313)
         );
  AOI220 U989 ( .A(regs[340]), .B(n75), .C(regs[276]), .D(n114), .Q(n1307) );
  AOI220 U990 ( .A(regs[848]), .B(n75), .C(regs[784]), .D(n114), .Q(n1215) );
  AOI220 U991 ( .A(regs[472]), .B(n1564), .C(regs[408]), .D(n72), .Q(n1397) );
  AOI220 U992 ( .A(regs[984]), .B(n113), .C(regs[920]), .D(n72), .Q(n1393) );
  AOI220 U993 ( .A(regs[215]), .B(n113), .C(regs[151]), .D(n72), .Q(n1385) );
  AOI220 U994 ( .A(regs[727]), .B(n113), .C(regs[663]), .D(n72), .Q(n1381) );
  AOI220 U995 ( .A(regs[471]), .B(n1564), .C(regs[407]), .D(n72), .Q(n1375) );
  AOI220 U996 ( .A(regs[983]), .B(n1564), .C(regs[919]), .D(n72), .Q(n1371) );
  AOI220 U997 ( .A(regs[90]), .B(n75), .C(regs[26]), .D(n114), .Q(n1449) );
  AOI220 U998 ( .A(regs[346]), .B(n75), .C(regs[282]), .D(n114), .Q(n1439) );
  AOI220 U999 ( .A(regs[986]), .B(n113), .C(regs[922]), .D(n72), .Q(n1437) );
  NOR40 U1000 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n109), .D(n1582), .Q(
        n23) );
  NOR40 U1001 ( .A(i_addr_Rd[0]), .B(n109), .C(n1585), .D(n1582), .Q(n26) );
  NOR40 U1002 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n109), .D(n1587), .Q(
        n13) );
  NOR40 U1003 ( .A(i_addr_Rd[0]), .B(n109), .C(n1585), .D(n1587), .Q(n16) );
  NOR40 U1004 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[0]), .C(n109), .D(n1591), .Q(
        n41) );
  NAND31 U1005 ( .A(n109), .B(n1586), .C(n1585), .Q(n1584) );
  NAND22 U1006 ( .A(n712), .B(n711), .Q(o_data_Rt[25]) );
  AOI221 U1007 ( .A(n854), .B(n710), .C(n852), .D(n709), .Q(n711) );
  NAND41 U1008 ( .A(n708), .B(n707), .C(n706), .D(n705), .Q(n709) );
  AOI221 U1009 ( .A(n110), .B(regs[249]), .C(n66), .D(regs[185]), .Q(n708) );
  NAND41 U1010 ( .A(n704), .B(n703), .C(n702), .D(n701), .Q(n710) );
  AOI221 U1011 ( .A(n110), .B(regs[761]), .C(n66), .D(regs[697]), .Q(n704) );
  NAND41 U1012 ( .A(n698), .B(n697), .C(n696), .D(n695), .Q(n699) );
  AOI221 U1013 ( .A(n110), .B(regs[505]), .C(n66), .D(regs[441]), .Q(n698) );
  NAND41 U1014 ( .A(n694), .B(n693), .C(n692), .D(n691), .Q(n700) );
  AOI221 U1015 ( .A(n110), .B(regs[1017]), .C(n66), .D(regs[953]), .Q(n694) );
  NAND22 U1016 ( .A(n756), .B(n755), .Q(o_data_Rt[27]) );
  AOI221 U1017 ( .A(n854), .B(n754), .C(n852), .D(n753), .Q(n755) );
  NAND41 U1018 ( .A(n752), .B(n751), .C(n750), .D(n749), .Q(n753) );
  NAND41 U1019 ( .A(n748), .B(n747), .C(n746), .D(n745), .Q(n754) );
  NAND41 U1020 ( .A(n742), .B(n741), .C(n740), .D(n739), .Q(n743) );
  NAND41 U1021 ( .A(n738), .B(n737), .C(n736), .D(n735), .Q(n744) );
  NAND22 U1022 ( .A(n580), .B(n579), .Q(o_data_Rt[19]) );
  NAND41 U1023 ( .A(n576), .B(n575), .C(n574), .D(n573), .Q(n577) );
  NAND41 U1024 ( .A(n572), .B(n571), .C(n570), .D(n569), .Q(n578) );
  NAND41 U1025 ( .A(n566), .B(n565), .C(n564), .D(n563), .Q(n567) );
  NAND41 U1026 ( .A(n562), .B(n561), .C(n560), .D(n559), .Q(n568) );
  NAND22 U1027 ( .A(n624), .B(n623), .Q(o_data_Rt[21]) );
  AOI221 U1028 ( .A(n854), .B(n622), .C(n852), .D(n621), .Q(n623) );
  NAND41 U1029 ( .A(n620), .B(n619), .C(n618), .D(n617), .Q(n621) );
  NAND41 U1030 ( .A(n616), .B(n615), .C(n614), .D(n613), .Q(n622) );
  NAND41 U1031 ( .A(n610), .B(n609), .C(n608), .D(n607), .Q(n611) );
  NAND41 U1032 ( .A(n606), .B(n605), .C(n604), .D(n603), .Q(n612) );
  NAND22 U1033 ( .A(n690), .B(n689), .Q(o_data_Rt[24]) );
  AOI221 U1034 ( .A(n854), .B(n688), .C(n852), .D(n687), .Q(n689) );
  NAND41 U1035 ( .A(n686), .B(n685), .C(n684), .D(n683), .Q(n687) );
  AOI221 U1036 ( .A(n110), .B(regs[248]), .C(n66), .D(regs[184]), .Q(n686) );
  NAND41 U1037 ( .A(n682), .B(n681), .C(n680), .D(n679), .Q(n688) );
  AOI221 U1038 ( .A(n110), .B(regs[760]), .C(n66), .D(regs[696]), .Q(n682) );
  NAND41 U1039 ( .A(n676), .B(n675), .C(n674), .D(n673), .Q(n677) );
  AOI221 U1040 ( .A(n110), .B(regs[504]), .C(n66), .D(regs[440]), .Q(n676) );
  NAND41 U1041 ( .A(n672), .B(n671), .C(n670), .D(n669), .Q(n678) );
  NAND22 U1042 ( .A(n734), .B(n733), .Q(o_data_Rt[26]) );
  AOI221 U1043 ( .A(n854), .B(n732), .C(n852), .D(n731), .Q(n733) );
  NAND41 U1044 ( .A(n730), .B(n729), .C(n728), .D(n727), .Q(n731) );
  NAND41 U1045 ( .A(n726), .B(n725), .C(n724), .D(n723), .Q(n732) );
  NAND41 U1046 ( .A(n720), .B(n719), .C(n718), .D(n717), .Q(n721) );
  NAND41 U1047 ( .A(n716), .B(n715), .C(n714), .D(n713), .Q(n722) );
  AOI221 U1048 ( .A(n110), .B(regs[1018]), .C(n66), .D(regs[954]), .Q(n716) );
  NAND22 U1049 ( .A(n404), .B(n403), .Q(o_data_Rt[11]) );
  NAND41 U1050 ( .A(n400), .B(n399), .C(n398), .D(n397), .Q(n401) );
  NAND41 U1051 ( .A(n396), .B(n395), .C(n394), .D(n393), .Q(n402) );
  NAND41 U1052 ( .A(n390), .B(n389), .C(n388), .D(n387), .Q(n391) );
  NAND41 U1053 ( .A(n386), .B(n385), .C(n384), .D(n383), .Q(n392) );
  NAND22 U1054 ( .A(n426), .B(n425), .Q(o_data_Rt[12]) );
  NAND41 U1055 ( .A(n422), .B(n421), .C(n420), .D(n419), .Q(n423) );
  AOI221 U1056 ( .A(n110), .B(regs[236]), .C(n66), .D(regs[172]), .Q(n422) );
  NAND41 U1057 ( .A(n418), .B(n417), .C(n416), .D(n415), .Q(n424) );
  AOI221 U1058 ( .A(n110), .B(regs[748]), .C(n66), .D(regs[684]), .Q(n418) );
  NAND41 U1059 ( .A(n412), .B(n411), .C(n410), .D(n409), .Q(n413) );
  NAND41 U1060 ( .A(n408), .B(n407), .C(n406), .D(n405), .Q(n414) );
  NAND22 U1061 ( .A(n448), .B(n447), .Q(o_data_Rt[13]) );
  NAND41 U1062 ( .A(n444), .B(n443), .C(n442), .D(n441), .Q(n445) );
  AOI221 U1063 ( .A(n110), .B(regs[237]), .C(n839), .D(regs[173]), .Q(n444) );
  NAND41 U1064 ( .A(n440), .B(n439), .C(n438), .D(n437), .Q(n446) );
  AOI221 U1065 ( .A(n110), .B(regs[749]), .C(n66), .D(regs[685]), .Q(n440) );
  NAND41 U1066 ( .A(n434), .B(n433), .C(n432), .D(n431), .Q(n435) );
  AOI221 U1067 ( .A(n110), .B(regs[493]), .C(n839), .D(regs[429]), .Q(n434) );
  NAND41 U1068 ( .A(n430), .B(n429), .C(n428), .D(n427), .Q(n436) );
  AOI221 U1069 ( .A(n110), .B(regs[1005]), .C(n66), .D(regs[941]), .Q(n430) );
  NAND22 U1070 ( .A(n602), .B(n601), .Q(o_data_Rt[20]) );
  AOI221 U1071 ( .A(n854), .B(n600), .C(n852), .D(n599), .Q(n601) );
  NAND41 U1072 ( .A(n598), .B(n597), .C(n596), .D(n595), .Q(n599) );
  NAND41 U1073 ( .A(n594), .B(n593), .C(n592), .D(n591), .Q(n600) );
  NAND41 U1074 ( .A(n588), .B(n587), .C(n586), .D(n585), .Q(n589) );
  NAND41 U1075 ( .A(n584), .B(n583), .C(n582), .D(n581), .Q(n590) );
  NAND22 U1076 ( .A(n492), .B(n491), .Q(o_data_Rt[15]) );
  AOI221 U1077 ( .A(n854), .B(n490), .C(n852), .D(n489), .Q(n491) );
  NAND41 U1078 ( .A(n488), .B(n487), .C(n486), .D(n485), .Q(n489) );
  NAND41 U1079 ( .A(n484), .B(n483), .C(n482), .D(n481), .Q(n490) );
  NAND41 U1080 ( .A(n478), .B(n477), .C(n476), .D(n475), .Q(n479) );
  NAND41 U1081 ( .A(n474), .B(n473), .C(n472), .D(n471), .Q(n480) );
  NAND22 U1082 ( .A(n646), .B(n645), .Q(o_data_Rt[22]) );
  AOI221 U1083 ( .A(n854), .B(n644), .C(n852), .D(n643), .Q(n645) );
  NAND41 U1084 ( .A(n642), .B(n641), .C(n640), .D(n639), .Q(n643) );
  NAND41 U1085 ( .A(n638), .B(n637), .C(n636), .D(n635), .Q(n644) );
  NAND41 U1086 ( .A(n632), .B(n631), .C(n630), .D(n629), .Q(n633) );
  NAND41 U1087 ( .A(n628), .B(n627), .C(n626), .D(n625), .Q(n634) );
  NAND22 U1088 ( .A(n668), .B(n667), .Q(o_data_Rt[23]) );
  AOI221 U1089 ( .A(n854), .B(n666), .C(n852), .D(n665), .Q(n667) );
  NAND41 U1090 ( .A(n664), .B(n663), .C(n662), .D(n661), .Q(n665) );
  NAND41 U1091 ( .A(n660), .B(n659), .C(n658), .D(n657), .Q(n666) );
  NAND41 U1092 ( .A(n654), .B(n653), .C(n652), .D(n651), .Q(n655) );
  NAND41 U1093 ( .A(n650), .B(n649), .C(n648), .D(n647), .Q(n656) );
  NAND22 U1094 ( .A(n558), .B(n557), .Q(o_data_Rt[18]) );
  AOI221 U1095 ( .A(n854), .B(n556), .C(n852), .D(n555), .Q(n557) );
  NAND41 U1096 ( .A(n554), .B(n553), .C(n552), .D(n551), .Q(n555) );
  NAND41 U1097 ( .A(n550), .B(n549), .C(n548), .D(n547), .Q(n556) );
  AOI221 U1098 ( .A(n834), .B(n546), .C(n832), .D(n545), .Q(n558) );
  NAND41 U1099 ( .A(n544), .B(n543), .C(n542), .D(n541), .Q(n545) );
  NAND41 U1100 ( .A(n540), .B(n539), .C(n538), .D(n537), .Q(n546) );
  AOI221 U1101 ( .A(n110), .B(regs[1010]), .C(n66), .D(regs[946]), .Q(n540) );
  NAND22 U1102 ( .A(n360), .B(n359), .Q(o_data_Rt[9]) );
  AOI221 U1103 ( .A(n854), .B(n358), .C(n852), .D(n357), .Q(n359) );
  NAND41 U1104 ( .A(n356), .B(n355), .C(n354), .D(n353), .Q(n357) );
  NAND41 U1105 ( .A(n352), .B(n351), .C(n350), .D(n349), .Q(n358) );
  NAND41 U1106 ( .A(n346), .B(n345), .C(n344), .D(n343), .Q(n347) );
  NAND41 U1107 ( .A(n342), .B(n341), .C(n340), .D(n339), .Q(n348) );
  NAND22 U1108 ( .A(n514), .B(n513), .Q(o_data_Rt[16]) );
  AOI221 U1109 ( .A(n854), .B(n512), .C(n852), .D(n511), .Q(n513) );
  NAND41 U1110 ( .A(n510), .B(n509), .C(n508), .D(n507), .Q(n511) );
  NAND41 U1111 ( .A(n506), .B(n505), .C(n504), .D(n503), .Q(n512) );
  NAND41 U1112 ( .A(n500), .B(n499), .C(n498), .D(n497), .Q(n501) );
  NAND41 U1113 ( .A(n496), .B(n495), .C(n494), .D(n493), .Q(n502) );
  NAND22 U1114 ( .A(n338), .B(n337), .Q(o_data_Rt[8]) );
  AOI221 U1115 ( .A(n854), .B(n336), .C(n852), .D(n335), .Q(n337) );
  NAND41 U1116 ( .A(n334), .B(n333), .C(n332), .D(n331), .Q(n335) );
  NAND41 U1117 ( .A(n330), .B(n329), .C(n328), .D(n327), .Q(n336) );
  AOI221 U1118 ( .A(n834), .B(n326), .C(n832), .D(n325), .Q(n338) );
  NAND41 U1119 ( .A(n324), .B(n323), .C(n322), .D(n321), .Q(n325) );
  NAND41 U1120 ( .A(n320), .B(n319), .C(n318), .D(n317), .Q(n326) );
  NAND22 U1121 ( .A(n382), .B(n381), .Q(o_data_Rt[10]) );
  NAND41 U1122 ( .A(n378), .B(n377), .C(n376), .D(n375), .Q(n379) );
  NAND41 U1123 ( .A(n374), .B(n373), .C(n372), .D(n371), .Q(n380) );
  NAND41 U1124 ( .A(n368), .B(n367), .C(n366), .D(n365), .Q(n369) );
  NAND41 U1125 ( .A(n364), .B(n363), .C(n362), .D(n361), .Q(n370) );
  NAND22 U1126 ( .A(n778), .B(n777), .Q(o_data_Rt[28]) );
  AOI221 U1127 ( .A(n854), .B(n776), .C(n852), .D(n775), .Q(n777) );
  NAND41 U1128 ( .A(n774), .B(n773), .C(n772), .D(n771), .Q(n775) );
  AOI221 U1129 ( .A(n110), .B(regs[252]), .C(n66), .D(regs[188]), .Q(n774) );
  NAND41 U1130 ( .A(n770), .B(n769), .C(n768), .D(n767), .Q(n776) );
  AOI221 U1131 ( .A(n110), .B(regs[764]), .C(n66), .D(regs[700]), .Q(n770) );
  NAND41 U1132 ( .A(n764), .B(n763), .C(n762), .D(n761), .Q(n765) );
  AOI221 U1133 ( .A(n110), .B(regs[508]), .C(n66), .D(regs[444]), .Q(n764) );
  NAND41 U1134 ( .A(n760), .B(n759), .C(n758), .D(n757), .Q(n766) );
  NAND22 U1135 ( .A(n316), .B(n315), .Q(o_data_Rt[7]) );
  AOI221 U1136 ( .A(n854), .B(n314), .C(n852), .D(n313), .Q(n315) );
  NAND41 U1137 ( .A(n312), .B(n311), .C(n310), .D(n309), .Q(n313) );
  NAND41 U1138 ( .A(n308), .B(n307), .C(n306), .D(n305), .Q(n314) );
  NAND41 U1139 ( .A(n302), .B(n301), .C(n300), .D(n299), .Q(n303) );
  NAND41 U1140 ( .A(n298), .B(n297), .C(n296), .D(n295), .Q(n304) );
  NAND22 U1141 ( .A(n250), .B(n249), .Q(o_data_Rt[4]) );
  AOI221 U1142 ( .A(n854), .B(n248), .C(n852), .D(n247), .Q(n249) );
  NAND41 U1143 ( .A(n246), .B(n245), .C(n244), .D(n243), .Q(n247) );
  AOI221 U1144 ( .A(n110), .B(regs[228]), .C(n66), .D(regs[164]), .Q(n246) );
  NAND41 U1145 ( .A(n242), .B(n241), .C(n240), .D(n239), .Q(n248) );
  AOI221 U1146 ( .A(n110), .B(regs[740]), .C(n66), .D(regs[676]), .Q(n242) );
  NAND41 U1147 ( .A(n236), .B(n235), .C(n234), .D(n233), .Q(n237) );
  AOI221 U1148 ( .A(n110), .B(regs[484]), .C(n66), .D(regs[420]), .Q(n236) );
  NAND41 U1149 ( .A(n232), .B(n231), .C(n230), .D(n229), .Q(n238) );
  AOI221 U1150 ( .A(n110), .B(regs[996]), .C(n66), .D(regs[932]), .Q(n232) );
  NAND22 U1151 ( .A(n800), .B(n799), .Q(o_data_Rt[29]) );
  AOI221 U1152 ( .A(n854), .B(n798), .C(n852), .D(n797), .Q(n799) );
  NAND41 U1153 ( .A(n796), .B(n795), .C(n794), .D(n793), .Q(n797) );
  AOI221 U1154 ( .A(n110), .B(regs[253]), .C(n66), .D(regs[189]), .Q(n796) );
  NAND41 U1155 ( .A(n792), .B(n791), .C(n790), .D(n789), .Q(n798) );
  AOI221 U1156 ( .A(n110), .B(regs[765]), .C(n66), .D(regs[701]), .Q(n792) );
  NAND41 U1157 ( .A(n786), .B(n785), .C(n784), .D(n783), .Q(n787) );
  AOI221 U1158 ( .A(n110), .B(regs[509]), .C(n66), .D(regs[445]), .Q(n786) );
  NAND41 U1159 ( .A(n782), .B(n781), .C(n780), .D(n779), .Q(n788) );
  AOI221 U1160 ( .A(n110), .B(regs[1021]), .C(n66), .D(regs[957]), .Q(n782) );
  NAND22 U1161 ( .A(n184), .B(n183), .Q(o_data_Rt[1]) );
  AOI221 U1162 ( .A(n854), .B(n182), .C(n852), .D(n181), .Q(n183) );
  NAND41 U1163 ( .A(n180), .B(n179), .C(n178), .D(n177), .Q(n181) );
  NAND41 U1164 ( .A(n176), .B(n175), .C(n174), .D(n173), .Q(n182) );
  NAND41 U1165 ( .A(n170), .B(n169), .C(n168), .D(n167), .Q(n171) );
  NAND41 U1166 ( .A(n166), .B(n165), .C(n164), .D(n163), .Q(n172) );
  NAND22 U1167 ( .A(n1192), .B(n1191), .Q(o_data_Rs[14]) );
  AOI221 U1168 ( .A(n1576), .B(n1190), .C(n1574), .D(n1189), .Q(n1191) );
  NAND41 U1169 ( .A(n1188), .B(n1187), .C(n1186), .D(n1185), .Q(n1189) );
  NAND41 U1170 ( .A(n1184), .B(n1183), .C(n1182), .D(n1181), .Q(n1190) );
  NAND41 U1171 ( .A(n1178), .B(n1177), .C(n1176), .D(n1175), .Q(n1179) );
  NAND41 U1172 ( .A(n1174), .B(n1173), .C(n1172), .D(n1171), .Q(n1180) );
  NAND22 U1173 ( .A(n906), .B(n905), .Q(o_data_Rs[1]) );
  AOI221 U1174 ( .A(n1576), .B(n904), .C(n1574), .D(n903), .Q(n905) );
  NAND41 U1175 ( .A(n902), .B(n901), .C(n900), .D(n899), .Q(n903) );
  NAND41 U1176 ( .A(n898), .B(n897), .C(n896), .D(n895), .Q(n904) );
  NAND41 U1177 ( .A(n892), .B(n891), .C(n890), .D(n889), .Q(n893) );
  NAND41 U1178 ( .A(n888), .B(n887), .C(n886), .D(n885), .Q(n894) );
  NAND22 U1179 ( .A(n1214), .B(n1213), .Q(o_data_Rs[15]) );
  AOI221 U1180 ( .A(n1576), .B(n1212), .C(n1574), .D(n1211), .Q(n1213) );
  NAND41 U1181 ( .A(n1210), .B(n1209), .C(n1208), .D(n1207), .Q(n1211) );
  NAND41 U1182 ( .A(n1206), .B(n1205), .C(n1204), .D(n1203), .Q(n1212) );
  NAND41 U1183 ( .A(n1200), .B(n1199), .C(n1198), .D(n1197), .Q(n1201) );
  NAND41 U1184 ( .A(n1196), .B(n1195), .C(n1194), .D(n1193), .Q(n1202) );
  NAND22 U1185 ( .A(n294), .B(n293), .Q(o_data_Rt[6]) );
  AOI221 U1186 ( .A(n854), .B(n292), .C(n852), .D(n291), .Q(n293) );
  NAND41 U1187 ( .A(n290), .B(n289), .C(n288), .D(n287), .Q(n291) );
  NAND41 U1188 ( .A(n286), .B(n285), .C(n284), .D(n283), .Q(n292) );
  NAND41 U1189 ( .A(n280), .B(n279), .C(n278), .D(n277), .Q(n281) );
  AOI221 U1190 ( .A(n110), .B(regs[486]), .C(n839), .D(regs[422]), .Q(n280) );
  NAND41 U1191 ( .A(n276), .B(n275), .C(n274), .D(n273), .Q(n282) );
  AOI221 U1192 ( .A(n110), .B(regs[998]), .C(n839), .D(regs[934]), .Q(n276) );
  NAND22 U1193 ( .A(n228), .B(n227), .Q(o_data_Rt[3]) );
  AOI221 U1194 ( .A(n854), .B(n226), .C(n852), .D(n225), .Q(n227) );
  NAND41 U1195 ( .A(n224), .B(n223), .C(n222), .D(n221), .Q(n225) );
  NAND41 U1196 ( .A(n220), .B(n219), .C(n218), .D(n217), .Q(n226) );
  AOI221 U1197 ( .A(n110), .B(regs[739]), .C(n66), .D(regs[675]), .Q(n220) );
  NAND41 U1198 ( .A(n214), .B(n213), .C(n212), .D(n211), .Q(n215) );
  AOI221 U1199 ( .A(n110), .B(regs[483]), .C(n66), .D(regs[419]), .Q(n214) );
  NAND41 U1200 ( .A(n210), .B(n209), .C(n208), .D(n207), .Q(n216) );
  AOI221 U1201 ( .A(n110), .B(regs[995]), .C(n66), .D(regs[931]), .Q(n210) );
  NAND22 U1202 ( .A(n1126), .B(n1125), .Q(o_data_Rs[11]) );
  AOI221 U1203 ( .A(n1576), .B(n1124), .C(n1574), .D(n1123), .Q(n1125) );
  NAND41 U1204 ( .A(n1122), .B(n1121), .C(n1120), .D(n1119), .Q(n1123) );
  NAND41 U1205 ( .A(n1118), .B(n1117), .C(n1116), .D(n1115), .Q(n1124) );
  NAND41 U1206 ( .A(n1112), .B(n1111), .C(n1110), .D(n1109), .Q(n1113) );
  NAND41 U1207 ( .A(n1108), .B(n1107), .C(n1106), .D(n1105), .Q(n1114) );
  NAND22 U1208 ( .A(n1148), .B(n1147), .Q(o_data_Rs[12]) );
  AOI221 U1209 ( .A(n1576), .B(n1146), .C(n1574), .D(n1145), .Q(n1147) );
  NAND41 U1210 ( .A(n1144), .B(n1143), .C(n1142), .D(n1141), .Q(n1145) );
  NAND41 U1211 ( .A(n1140), .B(n1139), .C(n1138), .D(n1137), .Q(n1146) );
  AOI221 U1212 ( .A(n1556), .B(n1136), .C(n1554), .D(n1135), .Q(n1148) );
  NAND41 U1213 ( .A(n1134), .B(n1133), .C(n1132), .D(n1131), .Q(n1135) );
  NAND41 U1214 ( .A(n1130), .B(n1129), .C(n1128), .D(n1127), .Q(n1136) );
  NAND22 U1215 ( .A(n1016), .B(n1015), .Q(o_data_Rs[6]) );
  AOI221 U1216 ( .A(n1576), .B(n1014), .C(n1574), .D(n1013), .Q(n1015) );
  NAND41 U1217 ( .A(n1012), .B(n1011), .C(n1010), .D(n1009), .Q(n1013) );
  NAND41 U1218 ( .A(n1008), .B(n1007), .C(n1006), .D(n1005), .Q(n1014) );
  NAND41 U1219 ( .A(n1002), .B(n1001), .C(n1000), .D(n999), .Q(n1003) );
  NAND41 U1220 ( .A(n998), .B(n997), .C(n996), .D(n995), .Q(n1004) );
  NAND22 U1221 ( .A(n1170), .B(n1169), .Q(o_data_Rs[13]) );
  AOI221 U1222 ( .A(n1576), .B(n1168), .C(n1574), .D(n1167), .Q(n1169) );
  NAND41 U1223 ( .A(n1166), .B(n1165), .C(n1164), .D(n1163), .Q(n1167) );
  NAND41 U1224 ( .A(n1162), .B(n1161), .C(n1160), .D(n1159), .Q(n1168) );
  NAND41 U1225 ( .A(n1156), .B(n1155), .C(n1154), .D(n1153), .Q(n1157) );
  NAND41 U1226 ( .A(n1152), .B(n1151), .C(n1150), .D(n1149), .Q(n1158) );
  NAND22 U1227 ( .A(n206), .B(n205), .Q(o_data_Rt[2]) );
  AOI221 U1228 ( .A(n854), .B(n204), .C(n852), .D(n203), .Q(n205) );
  NAND41 U1229 ( .A(n202), .B(n201), .C(n200), .D(n199), .Q(n203) );
  AOI221 U1230 ( .A(n110), .B(regs[226]), .C(n66), .D(regs[162]), .Q(n202) );
  NAND41 U1231 ( .A(n198), .B(n197), .C(n196), .D(n195), .Q(n204) );
  AOI221 U1232 ( .A(n110), .B(regs[738]), .C(n66), .D(regs[674]), .Q(n198) );
  NAND41 U1233 ( .A(n192), .B(n191), .C(n190), .D(n189), .Q(n193) );
  NAND41 U1234 ( .A(n188), .B(n187), .C(n186), .D(n185), .Q(n194) );
  NAND22 U1235 ( .A(n272), .B(n271), .Q(o_data_Rt[5]) );
  AOI221 U1236 ( .A(n854), .B(n270), .C(n852), .D(n269), .Q(n271) );
  NAND41 U1237 ( .A(n268), .B(n267), .C(n266), .D(n265), .Q(n269) );
  AOI221 U1238 ( .A(n110), .B(regs[229]), .C(n66), .D(regs[165]), .Q(n268) );
  NAND41 U1239 ( .A(n264), .B(n263), .C(n262), .D(n261), .Q(n270) );
  AOI221 U1240 ( .A(n110), .B(regs[741]), .C(n66), .D(regs[677]), .Q(n264) );
  NAND41 U1241 ( .A(n258), .B(n257), .C(n256), .D(n255), .Q(n259) );
  AOI221 U1242 ( .A(n110), .B(regs[485]), .C(n839), .D(regs[421]), .Q(n258) );
  NAND41 U1243 ( .A(n254), .B(n253), .C(n252), .D(n251), .Q(n260) );
  AOI221 U1244 ( .A(n110), .B(regs[997]), .C(n66), .D(regs[933]), .Q(n254) );
  NAND22 U1245 ( .A(n1258), .B(n1257), .Q(o_data_Rs[17]) );
  AOI221 U1246 ( .A(n1576), .B(n1256), .C(n1574), .D(n1255), .Q(n1257) );
  NAND41 U1247 ( .A(n1254), .B(n1253), .C(n1252), .D(n1251), .Q(n1255) );
  NAND41 U1248 ( .A(n1250), .B(n1249), .C(n1248), .D(n1247), .Q(n1256) );
  NAND41 U1249 ( .A(n1244), .B(n1243), .C(n1242), .D(n1241), .Q(n1245) );
  NAND41 U1250 ( .A(n1240), .B(n1239), .C(n1238), .D(n1237), .Q(n1246) );
  NAND22 U1251 ( .A(n1038), .B(n1037), .Q(o_data_Rs[7]) );
  AOI221 U1252 ( .A(n1576), .B(n1036), .C(n1574), .D(n1035), .Q(n1037) );
  NAND41 U1253 ( .A(n1034), .B(n1033), .C(n1032), .D(n1031), .Q(n1035) );
  NAND41 U1254 ( .A(n1030), .B(n1029), .C(n1028), .D(n1027), .Q(n1036) );
  NAND41 U1255 ( .A(n1024), .B(n1023), .C(n1022), .D(n1021), .Q(n1025) );
  NAND41 U1256 ( .A(n1020), .B(n1019), .C(n1018), .D(n1017), .Q(n1026) );
  NAND22 U1257 ( .A(n1060), .B(n1059), .Q(o_data_Rs[8]) );
  AOI221 U1258 ( .A(n1576), .B(n1058), .C(n1574), .D(n1057), .Q(n1059) );
  NAND41 U1259 ( .A(n1056), .B(n1055), .C(n1054), .D(n1053), .Q(n1057) );
  NAND41 U1260 ( .A(n1052), .B(n1051), .C(n1050), .D(n1049), .Q(n1058) );
  NAND41 U1261 ( .A(n1046), .B(n1045), .C(n1044), .D(n1043), .Q(n1047) );
  NAND41 U1262 ( .A(n1042), .B(n1041), .C(n1040), .D(n1039), .Q(n1048) );
  NAND22 U1263 ( .A(n856), .B(n855), .Q(o_data_Rt[31]) );
  AOI221 U1264 ( .A(n854), .B(n853), .C(n852), .D(n851), .Q(n855) );
  NAND41 U1265 ( .A(n850), .B(n849), .C(n848), .D(n847), .Q(n851) );
  NAND41 U1266 ( .A(n838), .B(n837), .C(n836), .D(n835), .Q(n853) );
  AOI221 U1267 ( .A(n68), .B(regs[607]), .C(n71), .D(regs[543]), .Q(n835) );
  AOI221 U1268 ( .A(n110), .B(regs[767]), .C(n66), .D(regs[703]), .Q(n838) );
  NAND41 U1269 ( .A(n830), .B(n829), .C(n828), .D(n827), .Q(n831) );
  NAND41 U1270 ( .A(n826), .B(n825), .C(n824), .D(n823), .Q(n833) );
  NAND22 U1271 ( .A(n536), .B(n535), .Q(o_data_Rt[17]) );
  AOI221 U1272 ( .A(n854), .B(n534), .C(n852), .D(n533), .Q(n535) );
  NAND41 U1273 ( .A(n532), .B(n531), .C(n530), .D(n529), .Q(n533) );
  AOI221 U1274 ( .A(n110), .B(regs[241]), .C(n66), .D(regs[177]), .Q(n532) );
  NAND41 U1275 ( .A(n528), .B(n527), .C(n526), .D(n525), .Q(n534) );
  AOI221 U1276 ( .A(n68), .B(regs[593]), .C(n71), .D(regs[529]), .Q(n525) );
  AOI221 U1277 ( .A(n110), .B(regs[753]), .C(n66), .D(regs[689]), .Q(n528) );
  AOI221 U1278 ( .A(n834), .B(n524), .C(n832), .D(n523), .Q(n536) );
  NAND41 U1279 ( .A(n522), .B(n521), .C(n520), .D(n519), .Q(n523) );
  AOI221 U1280 ( .A(n110), .B(regs[497]), .C(n839), .D(regs[433]), .Q(n522) );
  NAND41 U1281 ( .A(n518), .B(n517), .C(n516), .D(n515), .Q(n524) );
  AOI221 U1282 ( .A(n110), .B(regs[1009]), .C(n839), .D(regs[945]), .Q(n518)
         );
  NAND22 U1283 ( .A(n822), .B(n821), .Q(o_data_Rt[30]) );
  AOI221 U1284 ( .A(n854), .B(n820), .C(n852), .D(n819), .Q(n821) );
  NAND41 U1285 ( .A(n818), .B(n817), .C(n816), .D(n815), .Q(n819) );
  NAND41 U1286 ( .A(n814), .B(n813), .C(n812), .D(n811), .Q(n820) );
  AOI221 U1287 ( .A(n834), .B(n810), .C(n832), .D(n809), .Q(n822) );
  NAND41 U1288 ( .A(n808), .B(n807), .C(n806), .D(n805), .Q(n809) );
  NAND41 U1289 ( .A(n804), .B(n803), .C(n802), .D(n801), .Q(n810) );
  AOI221 U1290 ( .A(n110), .B(regs[1022]), .C(n66), .D(regs[958]), .Q(n804) );
  NAND22 U1291 ( .A(n470), .B(n469), .Q(o_data_Rt[14]) );
  NAND41 U1292 ( .A(n466), .B(n465), .C(n464), .D(n463), .Q(n467) );
  AOI221 U1293 ( .A(n110), .B(regs[238]), .C(n839), .D(regs[174]), .Q(n466) );
  NAND41 U1294 ( .A(n462), .B(n461), .C(n460), .D(n459), .Q(n468) );
  AOI221 U1295 ( .A(n68), .B(regs[590]), .C(n71), .D(regs[526]), .Q(n459) );
  AOI221 U1296 ( .A(n110), .B(regs[750]), .C(n66), .D(regs[686]), .Q(n462) );
  NAND41 U1297 ( .A(n456), .B(n455), .C(n454), .D(n453), .Q(n457) );
  AOI221 U1298 ( .A(n110), .B(regs[494]), .C(n839), .D(regs[430]), .Q(n456) );
  NAND41 U1299 ( .A(n452), .B(n451), .C(n450), .D(n449), .Q(n458) );
  AOI221 U1300 ( .A(n110), .B(regs[1006]), .C(n66), .D(regs[942]), .Q(n452) );
  NAND22 U1301 ( .A(n994), .B(n993), .Q(o_data_Rs[5]) );
  AOI221 U1302 ( .A(n1576), .B(n992), .C(n1574), .D(n991), .Q(n993) );
  NAND41 U1303 ( .A(n990), .B(n989), .C(n988), .D(n987), .Q(n991) );
  NAND41 U1304 ( .A(n986), .B(n985), .C(n984), .D(n983), .Q(n992) );
  AOI221 U1305 ( .A(n1556), .B(n982), .C(n1554), .D(n981), .Q(n994) );
  NAND41 U1306 ( .A(n980), .B(n979), .C(n978), .D(n977), .Q(n981) );
  NAND41 U1307 ( .A(n976), .B(n975), .C(n974), .D(n973), .Q(n982) );
  NAND22 U1308 ( .A(n1346), .B(n1345), .Q(o_data_Rs[21]) );
  AOI221 U1309 ( .A(n1576), .B(n1344), .C(n1574), .D(n1343), .Q(n1345) );
  NAND41 U1310 ( .A(n1342), .B(n1341), .C(n1340), .D(n1339), .Q(n1343) );
  NAND41 U1311 ( .A(n1338), .B(n1337), .C(n1336), .D(n1335), .Q(n1344) );
  NAND41 U1312 ( .A(n1332), .B(n1331), .C(n1330), .D(n1329), .Q(n1333) );
  NAND41 U1313 ( .A(n1328), .B(n1327), .C(n1326), .D(n1325), .Q(n1334) );
  NAND22 U1314 ( .A(n1280), .B(n1279), .Q(o_data_Rs[18]) );
  AOI221 U1315 ( .A(n1576), .B(n1278), .C(n1574), .D(n1277), .Q(n1279) );
  NAND41 U1316 ( .A(n1276), .B(n1275), .C(n1274), .D(n1273), .Q(n1277) );
  NAND41 U1317 ( .A(n1272), .B(n1271), .C(n1270), .D(n1269), .Q(n1278) );
  NAND41 U1318 ( .A(n1266), .B(n1265), .C(n1264), .D(n1263), .Q(n1267) );
  NAND41 U1319 ( .A(n1262), .B(n1261), .C(n1260), .D(n1259), .Q(n1268) );
  NAND22 U1320 ( .A(n1578), .B(n1577), .Q(o_data_Rs[31]) );
  AOI221 U1321 ( .A(n1576), .B(n1575), .C(n1574), .D(n1573), .Q(n1577) );
  NAND41 U1322 ( .A(n1572), .B(n1571), .C(n1570), .D(n1569), .Q(n1573) );
  NAND41 U1323 ( .A(n1560), .B(n1559), .C(n1558), .D(n1557), .Q(n1575) );
  NAND41 U1324 ( .A(n1552), .B(n1551), .C(n1550), .D(n1549), .Q(n1553) );
  NAND41 U1325 ( .A(n1548), .B(n1547), .C(n1546), .D(n1545), .Q(n1555) );
  NAND22 U1326 ( .A(n1544), .B(n1543), .Q(o_data_Rs[30]) );
  NAND41 U1327 ( .A(n1540), .B(n1539), .C(n1538), .D(n1537), .Q(n1541) );
  NAND41 U1328 ( .A(n1536), .B(n1535), .C(n1534), .D(n1533), .Q(n1542) );
  NAND41 U1329 ( .A(n1530), .B(n1529), .C(n1528), .D(n1527), .Q(n1531) );
  NAND41 U1330 ( .A(n1526), .B(n1525), .C(n1524), .D(n1523), .Q(n1532) );
  NAND22 U1331 ( .A(n1082), .B(n1081), .Q(o_data_Rs[9]) );
  AOI221 U1332 ( .A(n1576), .B(n1080), .C(n1574), .D(n1079), .Q(n1081) );
  NAND41 U1333 ( .A(n1078), .B(n1077), .C(n1076), .D(n1075), .Q(n1079) );
  NAND41 U1334 ( .A(n1074), .B(n1073), .C(n1072), .D(n1071), .Q(n1080) );
  AOI221 U1335 ( .A(n1556), .B(n1070), .C(n1554), .D(n1069), .Q(n1082) );
  NAND41 U1336 ( .A(n1068), .B(n1067), .C(n1066), .D(n1065), .Q(n1069) );
  NAND41 U1337 ( .A(n1064), .B(n1063), .C(n1062), .D(n1061), .Q(n1070) );
  NAND22 U1338 ( .A(n1500), .B(n1499), .Q(o_data_Rs[28]) );
  NAND41 U1339 ( .A(n1496), .B(n1495), .C(n1494), .D(n1493), .Q(n1497) );
  NAND41 U1340 ( .A(n1492), .B(n1491), .C(n1490), .D(n1489), .Q(n1498) );
  NAND41 U1341 ( .A(n1486), .B(n1485), .C(n1484), .D(n1483), .Q(n1487) );
  NAND41 U1342 ( .A(n1482), .B(n1481), .C(n1480), .D(n1479), .Q(n1488) );
  NAND22 U1343 ( .A(n162), .B(n161), .Q(o_data_Rt[0]) );
  NAND41 U1344 ( .A(n158), .B(n157), .C(n156), .D(n155), .Q(n159) );
  NAND41 U1345 ( .A(n154), .B(n153), .C(n152), .D(n151), .Q(n160) );
  NAND41 U1346 ( .A(n147), .B(n146), .C(n145), .D(n144), .Q(n148) );
  NAND41 U1347 ( .A(n142), .B(n141), .C(n140), .D(n139), .Q(n149) );
  AOI221 U1348 ( .A(n68), .B(regs[832]), .C(n71), .D(regs[768]), .Q(n139) );
  AOI221 U1349 ( .A(n110), .B(regs[992]), .C(n66), .D(regs[928]), .Q(n142) );
  NAND22 U1350 ( .A(n1522), .B(n1521), .Q(o_data_Rs[29]) );
  NAND41 U1351 ( .A(n1518), .B(n1517), .C(n1516), .D(n1515), .Q(n1519) );
  NAND41 U1352 ( .A(n1514), .B(n1513), .C(n1512), .D(n1511), .Q(n1520) );
  NAND41 U1353 ( .A(n1508), .B(n1507), .C(n1506), .D(n1505), .Q(n1509) );
  NAND41 U1354 ( .A(n1504), .B(n1503), .C(n1502), .D(n1501), .Q(n1510) );
  NAND22 U1355 ( .A(n950), .B(n949), .Q(o_data_Rs[3]) );
  NAND41 U1356 ( .A(n946), .B(n945), .C(n944), .D(n943), .Q(n947) );
  NAND41 U1357 ( .A(n942), .B(n941), .C(n940), .D(n939), .Q(n948) );
  NAND41 U1358 ( .A(n936), .B(n935), .C(n934), .D(n933), .Q(n937) );
  NAND41 U1359 ( .A(n932), .B(n931), .C(n930), .D(n929), .Q(n938) );
  NAND22 U1360 ( .A(n1104), .B(n1103), .Q(o_data_Rs[10]) );
  NAND41 U1361 ( .A(n1100), .B(n1099), .C(n1098), .D(n1097), .Q(n1101) );
  NAND41 U1362 ( .A(n1096), .B(n1095), .C(n1094), .D(n1093), .Q(n1102) );
  NAND41 U1363 ( .A(n1090), .B(n1089), .C(n1088), .D(n1087), .Q(n1091) );
  NAND41 U1364 ( .A(n1086), .B(n1085), .C(n1084), .D(n1083), .Q(n1092) );
  NAND22 U1365 ( .A(n972), .B(n971), .Q(o_data_Rs[4]) );
  NAND41 U1366 ( .A(n968), .B(n967), .C(n966), .D(n965), .Q(n969) );
  NAND41 U1367 ( .A(n964), .B(n963), .C(n962), .D(n961), .Q(n970) );
  AOI221 U1368 ( .A(n1556), .B(n960), .C(n1554), .D(n959), .Q(n972) );
  NAND41 U1369 ( .A(n958), .B(n957), .C(n956), .D(n955), .Q(n959) );
  NAND41 U1370 ( .A(n954), .B(n953), .C(n952), .D(n951), .Q(n960) );
  NAND22 U1371 ( .A(n928), .B(n927), .Q(o_data_Rs[2]) );
  NAND41 U1372 ( .A(n924), .B(n923), .C(n922), .D(n921), .Q(n925) );
  NAND41 U1373 ( .A(n920), .B(n919), .C(n918), .D(n917), .Q(n926) );
  NAND41 U1374 ( .A(n914), .B(n913), .C(n912), .D(n911), .Q(n915) );
  NAND41 U1375 ( .A(n910), .B(n909), .C(n908), .D(n907), .Q(n916) );
  NAND22 U1376 ( .A(n884), .B(n883), .Q(o_data_Rs[0]) );
  AOI221 U1377 ( .A(n1576), .B(n882), .C(n1574), .D(n881), .Q(n883) );
  NAND41 U1378 ( .A(n880), .B(n879), .C(n878), .D(n877), .Q(n881) );
  NAND41 U1379 ( .A(n876), .B(n875), .C(n874), .D(n873), .Q(n882) );
  NAND41 U1380 ( .A(n869), .B(n868), .C(n867), .D(n866), .Q(n870) );
  NAND41 U1381 ( .A(n864), .B(n863), .C(n862), .D(n861), .Q(n871) );
  NAND22 U1382 ( .A(n1302), .B(n1301), .Q(o_data_Rs[19]) );
  AOI221 U1383 ( .A(n1576), .B(n1300), .C(n1574), .D(n1299), .Q(n1301) );
  NAND41 U1384 ( .A(n1298), .B(n1297), .C(n1296), .D(n1295), .Q(n1299) );
  NAND41 U1385 ( .A(n1294), .B(n1293), .C(n1292), .D(n1291), .Q(n1300) );
  NAND41 U1386 ( .A(n1288), .B(n1287), .C(n1286), .D(n1285), .Q(n1289) );
  NAND41 U1387 ( .A(n1284), .B(n1283), .C(n1282), .D(n1281), .Q(n1290) );
  NAND22 U1388 ( .A(n1368), .B(n1367), .Q(o_data_Rs[22]) );
  AOI221 U1389 ( .A(n1576), .B(n1366), .C(n1574), .D(n1365), .Q(n1367) );
  NAND41 U1390 ( .A(n1364), .B(n1363), .C(n1362), .D(n1361), .Q(n1365) );
  AOI221 U1391 ( .A(regs[246]), .B(n112), .C(regs[182]), .D(n76), .Q(n1364) );
  NAND41 U1392 ( .A(n1360), .B(n1359), .C(n1358), .D(n1357), .Q(n1366) );
  NAND41 U1393 ( .A(n1354), .B(n1353), .C(n1352), .D(n1351), .Q(n1355) );
  NAND41 U1394 ( .A(n1350), .B(n1349), .C(n1348), .D(n1347), .Q(n1356) );
  NAND22 U1395 ( .A(n1324), .B(n1323), .Q(o_data_Rs[20]) );
  AOI221 U1396 ( .A(n1576), .B(n1322), .C(n1574), .D(n1321), .Q(n1323) );
  NAND41 U1397 ( .A(n1320), .B(n1319), .C(n1318), .D(n1317), .Q(n1321) );
  NAND41 U1398 ( .A(n1316), .B(n1315), .C(n1314), .D(n1313), .Q(n1322) );
  NAND41 U1399 ( .A(n1310), .B(n1309), .C(n1308), .D(n1307), .Q(n1311) );
  NAND41 U1400 ( .A(n1306), .B(n1305), .C(n1304), .D(n1303), .Q(n1312) );
  NAND22 U1401 ( .A(n1236), .B(n1235), .Q(o_data_Rs[16]) );
  AOI221 U1402 ( .A(n1576), .B(n1234), .C(n1574), .D(n1233), .Q(n1235) );
  NAND41 U1403 ( .A(n1232), .B(n1231), .C(n1230), .D(n1229), .Q(n1233) );
  NAND41 U1404 ( .A(n1228), .B(n1227), .C(n1226), .D(n1225), .Q(n1234) );
  NAND41 U1405 ( .A(n1222), .B(n1221), .C(n1220), .D(n1219), .Q(n1223) );
  NAND41 U1406 ( .A(n1218), .B(n1217), .C(n1216), .D(n1215), .Q(n1224) );
  NAND22 U1407 ( .A(n1412), .B(n1411), .Q(o_data_Rs[24]) );
  AOI221 U1408 ( .A(n1576), .B(n1410), .C(n1574), .D(n1409), .Q(n1411) );
  NAND41 U1409 ( .A(n1408), .B(n1407), .C(n1406), .D(n1405), .Q(n1409) );
  NAND41 U1410 ( .A(n1404), .B(n1403), .C(n1402), .D(n1401), .Q(n1410) );
  NAND41 U1411 ( .A(n1398), .B(n1397), .C(n1396), .D(n1395), .Q(n1399) );
  NAND41 U1412 ( .A(n1394), .B(n1393), .C(n1392), .D(n1391), .Q(n1400) );
  NAND22 U1413 ( .A(n1390), .B(n1389), .Q(o_data_Rs[23]) );
  AOI221 U1414 ( .A(n1576), .B(n1388), .C(n1574), .D(n1387), .Q(n1389) );
  NAND41 U1415 ( .A(n1386), .B(n1385), .C(n1384), .D(n1383), .Q(n1387) );
  NAND41 U1416 ( .A(n1382), .B(n1381), .C(n1380), .D(n1379), .Q(n1388) );
  NAND41 U1417 ( .A(n1376), .B(n1375), .C(n1374), .D(n1373), .Q(n1377) );
  NAND41 U1418 ( .A(n1372), .B(n1371), .C(n1370), .D(n1369), .Q(n1378) );
  NAND22 U1419 ( .A(n1434), .B(n1433), .Q(o_data_Rs[25]) );
  NAND41 U1420 ( .A(n1430), .B(n1429), .C(n1428), .D(n1427), .Q(n1431) );
  NAND41 U1421 ( .A(n1426), .B(n1425), .C(n1424), .D(n1423), .Q(n1432) );
  NAND41 U1422 ( .A(n1420), .B(n1419), .C(n1418), .D(n1417), .Q(n1421) );
  NAND41 U1423 ( .A(n1416), .B(n1415), .C(n1414), .D(n1413), .Q(n1422) );
  NAND22 U1424 ( .A(n1456), .B(n1455), .Q(o_data_Rs[26]) );
  NAND41 U1425 ( .A(n1452), .B(n1451), .C(n1450), .D(n1449), .Q(n1453) );
  NAND41 U1426 ( .A(n1448), .B(n1447), .C(n1446), .D(n1445), .Q(n1454) );
  NAND41 U1427 ( .A(n1442), .B(n1441), .C(n1440), .D(n1439), .Q(n1443) );
  NAND41 U1428 ( .A(n1438), .B(n1437), .C(n1436), .D(n1435), .Q(n1444) );
  NAND22 U1429 ( .A(n1478), .B(n1477), .Q(o_data_Rs[27]) );
  NAND41 U1430 ( .A(n1474), .B(n1473), .C(n1472), .D(n1471), .Q(n1475) );
  NAND41 U1431 ( .A(n1470), .B(n1469), .C(n1468), .D(n1467), .Q(n1476) );
  NAND41 U1432 ( .A(n1464), .B(n1463), .C(n1462), .D(n1461), .Q(n1465) );
  NAND41 U1433 ( .A(n1460), .B(n1459), .C(n1458), .D(n1457), .Q(n1466) );
  INV3 U1434 ( .A(i_addr_Rs[2]), .Q(n857) );
  NOR21 U1435 ( .A(n1584), .B(n1587), .Q(n18) );
  INV3 U1436 ( .A(i_addr_Rt_0_), .Q(n137) );
  NOR31 U1437 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[1]), .C(i_addr_Rs[2]), .Q(n1567) );
  AOI220 U1438 ( .A(n110), .B(regs[480]), .C(n66), .D(regs[416]), .Q(n147) );
  AOI220 U1439 ( .A(n110), .B(regs[224]), .C(n66), .D(regs[160]), .Q(n158) );
  AOI220 U1440 ( .A(n110), .B(regs[993]), .C(n66), .D(regs[929]), .Q(n166) );
  AOI220 U1441 ( .A(n110), .B(regs[481]), .C(n66), .D(regs[417]), .Q(n170) );
  AOI220 U1442 ( .A(n110), .B(regs[737]), .C(n66), .D(regs[673]), .Q(n176) );
  AOI220 U1443 ( .A(n842), .B(regs[705]), .C(n67), .D(regs[641]), .Q(n175) );
  AOI220 U1444 ( .A(n110), .B(regs[225]), .C(n66), .D(regs[161]), .Q(n180) );
  AOI220 U1445 ( .A(n110), .B(regs[994]), .C(n66), .D(regs[930]), .Q(n188) );
  AOI220 U1446 ( .A(n110), .B(regs[482]), .C(n66), .D(regs[418]), .Q(n192) );
  AOI220 U1447 ( .A(n111), .B(regs[706]), .C(n841), .D(regs[642]), .Q(n197) );
  AOI220 U1448 ( .A(n69), .B(regs[355]), .C(n843), .D(regs[291]), .Q(n212) );
  AOI220 U1449 ( .A(n840), .B(regs[227]), .C(n66), .D(regs[163]), .Q(n224) );
  AOI220 U1450 ( .A(n69), .B(regs[868]), .C(n843), .D(regs[804]), .Q(n230) );
  AOI220 U1451 ( .A(n846), .B(regs[836]), .C(n71), .D(regs[772]), .Q(n229) );
  AOI220 U1452 ( .A(n69), .B(regs[612]), .C(n843), .D(regs[548]), .Q(n240) );
  AOI220 U1453 ( .A(n846), .B(regs[68]), .C(n71), .D(regs[4]), .Q(n243) );
  AOI220 U1454 ( .A(n846), .B(regs[837]), .C(n71), .D(regs[773]), .Q(n251) );
  AOI220 U1455 ( .A(n846), .B(regs[69]), .C(n71), .D(regs[5]), .Q(n265) );
  AOI220 U1456 ( .A(n844), .B(regs[870]), .C(n70), .D(regs[806]), .Q(n274) );
  AOI220 U1457 ( .A(n844), .B(regs[358]), .C(n70), .D(regs[294]), .Q(n278) );
  AOI220 U1458 ( .A(n840), .B(regs[230]), .C(n66), .D(regs[166]), .Q(n290) );
  AOI220 U1459 ( .A(n840), .B(regs[487]), .C(n66), .D(regs[423]), .Q(n302) );
  AOI220 U1460 ( .A(n69), .B(regs[615]), .C(n843), .D(regs[551]), .Q(n306) );
  AOI220 U1461 ( .A(n840), .B(regs[231]), .C(n66), .D(regs[167]), .Q(n312) );
  AOI220 U1462 ( .A(n840), .B(regs[488]), .C(n66), .D(regs[424]), .Q(n324) );
  AOI220 U1463 ( .A(n110), .B(regs[744]), .C(n66), .D(regs[680]), .Q(n330) );
  AOI220 U1464 ( .A(n110), .B(regs[232]), .C(n66), .D(regs[168]), .Q(n334) );
  AOI220 U1465 ( .A(n69), .B(regs[104]), .C(n843), .D(regs[40]), .Q(n332) );
  AOI220 U1466 ( .A(n110), .B(regs[1001]), .C(n839), .D(regs[937]), .Q(n342)
         );
  AOI220 U1467 ( .A(n110), .B(regs[489]), .C(n66), .D(regs[425]), .Q(n346) );
  AOI220 U1468 ( .A(n110), .B(regs[745]), .C(n66), .D(regs[681]), .Q(n352) );
  AOI220 U1469 ( .A(n110), .B(regs[233]), .C(n66), .D(regs[169]), .Q(n356) );
  AOI220 U1470 ( .A(n69), .B(regs[105]), .C(n843), .D(regs[41]), .Q(n354) );
  AOI220 U1471 ( .A(n110), .B(regs[1002]), .C(n66), .D(regs[938]), .Q(n364) );
  AOI220 U1472 ( .A(n110), .B(regs[490]), .C(n66), .D(regs[426]), .Q(n368) );
  AOI220 U1473 ( .A(n110), .B(regs[746]), .C(n66), .D(regs[682]), .Q(n374) );
  AOI220 U1474 ( .A(n110), .B(regs[234]), .C(n839), .D(regs[170]), .Q(n378) );
  AOI220 U1475 ( .A(n110), .B(regs[1003]), .C(n839), .D(regs[939]), .Q(n386)
         );
  AOI220 U1476 ( .A(n110), .B(regs[491]), .C(n66), .D(regs[427]), .Q(n390) );
  AOI220 U1477 ( .A(n110), .B(regs[747]), .C(n66), .D(regs[683]), .Q(n396) );
  AOI220 U1478 ( .A(n110), .B(regs[235]), .C(n839), .D(regs[171]), .Q(n400) );
  AOI220 U1479 ( .A(n110), .B(regs[1004]), .C(n839), .D(regs[940]), .Q(n408)
         );
  AOI220 U1480 ( .A(n110), .B(regs[492]), .C(n66), .D(regs[428]), .Q(n412) );
  AOI220 U1481 ( .A(n111), .B(regs[716]), .C(n67), .D(regs[652]), .Q(n417) );
  AOI220 U1482 ( .A(n111), .B(regs[204]), .C(n67), .D(regs[140]), .Q(n421) );
  AOI220 U1483 ( .A(n111), .B(regs[973]), .C(n67), .D(regs[909]), .Q(n429) );
  AOI220 U1484 ( .A(n111), .B(regs[461]), .C(n67), .D(regs[397]), .Q(n433) );
  AOI220 U1485 ( .A(n111), .B(regs[717]), .C(n67), .D(regs[653]), .Q(n439) );
  AOI220 U1486 ( .A(n111), .B(regs[205]), .C(n67), .D(regs[141]), .Q(n443) );
  AOI220 U1487 ( .A(n842), .B(regs[206]), .C(n67), .D(regs[142]), .Q(n465) );
  AOI220 U1488 ( .A(n111), .B(regs[975]), .C(n67), .D(regs[911]), .Q(n473) );
  AOI220 U1489 ( .A(n111), .B(regs[463]), .C(n67), .D(regs[399]), .Q(n477) );
  AOI220 U1490 ( .A(n111), .B(regs[719]), .C(n67), .D(regs[655]), .Q(n483) );
  AOI220 U1491 ( .A(n842), .B(regs[207]), .C(n67), .D(regs[143]), .Q(n487) );
  AOI220 U1492 ( .A(n111), .B(regs[976]), .C(n67), .D(regs[912]), .Q(n495) );
  AOI220 U1493 ( .A(n68), .B(regs[336]), .C(n845), .D(regs[272]), .Q(n497) );
  AOI220 U1494 ( .A(n846), .B(regs[80]), .C(n71), .D(regs[16]), .Q(n507) );
  AOI220 U1495 ( .A(n846), .B(regs[849]), .C(n71), .D(regs[785]), .Q(n515) );
  AOI220 U1496 ( .A(n844), .B(regs[113]), .C(n70), .D(regs[49]), .Q(n530) );
  AOI220 U1497 ( .A(n846), .B(regs[850]), .C(n71), .D(regs[786]), .Q(n537) );
  AOI220 U1498 ( .A(n842), .B(regs[468]), .C(n67), .D(regs[404]), .Q(n587) );
  AOI220 U1499 ( .A(n68), .B(regs[340]), .C(n845), .D(regs[276]), .Q(n585) );
  AOI220 U1500 ( .A(n68), .B(regs[84]), .C(n845), .D(regs[20]), .Q(n595) );
  AOI220 U1501 ( .A(n68), .B(regs[853]), .C(n845), .D(regs[789]), .Q(n603) );
  AOI220 U1502 ( .A(n842), .B(regs[469]), .C(n67), .D(regs[405]), .Q(n609) );
  AOI220 U1503 ( .A(n842), .B(regs[213]), .C(n67), .D(regs[149]), .Q(n619) );
  AOI220 U1504 ( .A(n68), .B(regs[85]), .C(n845), .D(regs[21]), .Q(n617) );
  AOI220 U1505 ( .A(n68), .B(regs[854]), .C(n845), .D(regs[790]), .Q(n625) );
  AOI220 U1506 ( .A(n111), .B(regs[472]), .C(n841), .D(regs[408]), .Q(n675) );
  AOI220 U1507 ( .A(n111), .B(regs[216]), .C(n841), .D(regs[152]), .Q(n685) );
  AOI220 U1508 ( .A(n111), .B(regs[473]), .C(n841), .D(regs[409]), .Q(n697) );
  AOI220 U1509 ( .A(n111), .B(regs[217]), .C(n841), .D(regs[153]), .Q(n707) );
  AOI220 U1510 ( .A(n844), .B(regs[121]), .C(n70), .D(regs[57]), .Q(n706) );
  AOI220 U1511 ( .A(n840), .B(regs[506]), .C(n66), .D(regs[442]), .Q(n720) );
  AOI220 U1512 ( .A(n110), .B(regs[762]), .C(n66), .D(regs[698]), .Q(n726) );
  AOI220 U1513 ( .A(n840), .B(regs[250]), .C(n66), .D(regs[186]), .Q(n730) );
  AOI220 U1514 ( .A(n840), .B(regs[1019]), .C(n66), .D(regs[955]), .Q(n738) );
  AOI220 U1515 ( .A(n69), .B(regs[891]), .C(n843), .D(regs[827]), .Q(n736) );
  AOI220 U1516 ( .A(n110), .B(regs[507]), .C(n66), .D(regs[443]), .Q(n742) );
  AOI220 U1517 ( .A(n110), .B(regs[763]), .C(n66), .D(regs[699]), .Q(n748) );
  AOI220 U1518 ( .A(n840), .B(regs[251]), .C(n66), .D(regs[187]), .Q(n752) );
  AOI220 U1519 ( .A(n69), .B(regs[123]), .C(n843), .D(regs[59]), .Q(n750) );
  AOI220 U1520 ( .A(n840), .B(regs[1020]), .C(n66), .D(regs[956]), .Q(n760) );
  AOI220 U1521 ( .A(n111), .B(regs[477]), .C(n841), .D(regs[413]), .Q(n785) );
  AOI220 U1522 ( .A(n844), .B(regs[382]), .C(n70), .D(regs[318]), .Q(n806) );
  AOI220 U1523 ( .A(n844), .B(regs[126]), .C(n70), .D(regs[62]), .Q(n816) );
  AOI220 U1524 ( .A(n844), .B(regs[383]), .C(n70), .D(regs[319]), .Q(n828) );
  AOI220 U1525 ( .A(n844), .B(regs[639]), .C(n70), .D(regs[575]), .Q(n836) );
  AOI220 U1526 ( .A(n111), .B(regs[223]), .C(n67), .D(regs[159]), .Q(n849) );
  AOI220 U1527 ( .A(regs[608]), .B(n73), .C(regs[544]), .D(n74), .Q(n874) );
  AOI220 U1528 ( .A(regs[192]), .B(n113), .C(regs[128]), .D(n72), .Q(n879) );
  AOI220 U1529 ( .A(regs[96]), .B(n73), .C(regs[32]), .D(n74), .Q(n878) );
  AOI220 U1530 ( .A(regs[481]), .B(n1562), .C(regs[417]), .D(n1561), .Q(n892)
         );
  AOI220 U1531 ( .A(regs[449]), .B(n1564), .C(regs[385]), .D(n72), .Q(n891) );
  AOI220 U1532 ( .A(regs[353]), .B(n73), .C(regs[289]), .D(n74), .Q(n890) );
  AOI220 U1533 ( .A(regs[737]), .B(n1562), .C(regs[673]), .D(n1561), .Q(n898)
         );
  AOI220 U1534 ( .A(regs[705]), .B(n1564), .C(regs[641]), .D(n72), .Q(n897) );
  AOI220 U1535 ( .A(regs[609]), .B(n1566), .C(regs[545]), .D(n1565), .Q(n896)
         );
  AOI220 U1536 ( .A(regs[739]), .B(n112), .C(regs[675]), .D(n76), .Q(n942) );
  AOI220 U1537 ( .A(regs[227]), .B(n112), .C(regs[163]), .D(n76), .Q(n946) );
  AOI220 U1538 ( .A(regs[67]), .B(n75), .C(regs[3]), .D(n1567), .Q(n943) );
  AOI220 U1539 ( .A(regs[964]), .B(n113), .C(regs[900]), .D(n72), .Q(n953) );
  AOI220 U1540 ( .A(regs[484]), .B(n1562), .C(regs[420]), .D(n1561), .Q(n958)
         );
  AOI220 U1541 ( .A(regs[452]), .B(n1564), .C(regs[388]), .D(n72), .Q(n957) );
  AOI220 U1542 ( .A(regs[324]), .B(n1568), .C(regs[260]), .D(n1567), .Q(n955)
         );
  AOI220 U1543 ( .A(regs[740]), .B(n112), .C(regs[676]), .D(n76), .Q(n964) );
  AOI220 U1544 ( .A(regs[68]), .B(n1568), .C(regs[4]), .D(n1567), .Q(n965) );
  AOI220 U1545 ( .A(regs[453]), .B(n113), .C(regs[389]), .D(n72), .Q(n979) );
  AOI220 U1546 ( .A(regs[709]), .B(n1564), .C(regs[645]), .D(n72), .Q(n985) );
  AOI220 U1547 ( .A(regs[197]), .B(n1564), .C(regs[133]), .D(n72), .Q(n989) );
  AOI220 U1548 ( .A(regs[966]), .B(n1564), .C(regs[902]), .D(n72), .Q(n997) );
  AOI220 U1549 ( .A(regs[870]), .B(n1566), .C(regs[806]), .D(n74), .Q(n996) );
  AOI220 U1550 ( .A(regs[454]), .B(n1564), .C(regs[390]), .D(n72), .Q(n1001)
         );
  AOI220 U1551 ( .A(regs[710]), .B(n1564), .C(regs[646]), .D(n72), .Q(n1007)
         );
  AOI220 U1552 ( .A(regs[198]), .B(n1564), .C(regs[134]), .D(n72), .Q(n1011)
         );
  AOI220 U1553 ( .A(regs[492]), .B(n1562), .C(regs[428]), .D(n76), .Q(n1134)
         );
  AOI220 U1554 ( .A(regs[460]), .B(n1564), .C(regs[396]), .D(n72), .Q(n1133)
         );
  AOI220 U1555 ( .A(regs[236]), .B(n1562), .C(regs[172]), .D(n76), .Q(n1144)
         );
  AOI220 U1556 ( .A(regs[204]), .B(n1564), .C(regs[140]), .D(n72), .Q(n1143)
         );
  AOI220 U1557 ( .A(regs[493]), .B(n1562), .C(regs[429]), .D(n76), .Q(n1156)
         );
  AOI220 U1558 ( .A(regs[461]), .B(n1564), .C(regs[397]), .D(n72), .Q(n1155)
         );
  AOI220 U1559 ( .A(regs[1006]), .B(n112), .C(regs[942]), .D(n76), .Q(n1174)
         );
  AOI220 U1560 ( .A(regs[974]), .B(n113), .C(regs[910]), .D(n72), .Q(n1173) );
  AOI220 U1561 ( .A(regs[846]), .B(n1568), .C(regs[782]), .D(n114), .Q(n1171)
         );
  AOI220 U1562 ( .A(regs[494]), .B(n112), .C(regs[430]), .D(n1561), .Q(n1178)
         );
  AOI220 U1563 ( .A(regs[462]), .B(n113), .C(regs[398]), .D(n1563), .Q(n1177)
         );
  AOI220 U1564 ( .A(regs[366]), .B(n73), .C(regs[302]), .D(n1565), .Q(n1176)
         );
  AOI220 U1565 ( .A(regs[334]), .B(n1568), .C(regs[270]), .D(n114), .Q(n1175)
         );
  AOI220 U1566 ( .A(regs[750]), .B(n112), .C(regs[686]), .D(n76), .Q(n1184) );
  AOI220 U1567 ( .A(regs[718]), .B(n113), .C(regs[654]), .D(n72), .Q(n1183) );
  AOI220 U1568 ( .A(regs[238]), .B(n112), .C(regs[174]), .D(n1561), .Q(n1188)
         );
  AOI220 U1569 ( .A(regs[206]), .B(n113), .C(regs[142]), .D(n1563), .Q(n1187)
         );
  AOI220 U1570 ( .A(regs[110]), .B(n73), .C(regs[46]), .D(n1565), .Q(n1186) );
  AOI220 U1571 ( .A(regs[78]), .B(n1568), .C(regs[14]), .D(n114), .Q(n1185) );
  AOI220 U1572 ( .A(regs[1007]), .B(n112), .C(regs[943]), .D(n76), .Q(n1196)
         );
  AOI220 U1573 ( .A(regs[975]), .B(n113), .C(regs[911]), .D(n72), .Q(n1195) );
  AOI220 U1574 ( .A(regs[847]), .B(n1568), .C(regs[783]), .D(n114), .Q(n1193)
         );
  AOI220 U1575 ( .A(regs[495]), .B(n112), .C(regs[431]), .D(n1561), .Q(n1200)
         );
  AOI220 U1576 ( .A(regs[463]), .B(n113), .C(regs[399]), .D(n1563), .Q(n1199)
         );
  AOI220 U1577 ( .A(regs[367]), .B(n73), .C(regs[303]), .D(n1565), .Q(n1198)
         );
  AOI220 U1578 ( .A(regs[335]), .B(n1568), .C(regs[271]), .D(n114), .Q(n1197)
         );
  AOI220 U1579 ( .A(regs[751]), .B(n112), .C(regs[687]), .D(n76), .Q(n1206) );
  AOI220 U1580 ( .A(regs[719]), .B(n113), .C(regs[655]), .D(n72), .Q(n1205) );
  AOI220 U1581 ( .A(regs[80]), .B(n1568), .C(regs[16]), .D(n1567), .Q(n1229)
         );
  AOI220 U1582 ( .A(regs[1009]), .B(n1562), .C(regs[945]), .D(n1561), .Q(n1240) );
  AOI220 U1583 ( .A(regs[977]), .B(n1564), .C(regs[913]), .D(n1563), .Q(n1239)
         );
  AOI220 U1584 ( .A(regs[881]), .B(n1566), .C(regs[817]), .D(n1565), .Q(n1238)
         );
  AOI220 U1585 ( .A(regs[241]), .B(n1562), .C(regs[177]), .D(n1561), .Q(n1254)
         );
  AOI220 U1586 ( .A(regs[113]), .B(n73), .C(regs[49]), .D(n1565), .Q(n1252) );
  AOI220 U1587 ( .A(regs[850]), .B(n1568), .C(regs[786]), .D(n1567), .Q(n1259)
         );
  AOI220 U1588 ( .A(regs[339]), .B(n75), .C(regs[275]), .D(n114), .Q(n1285) );
  AOI220 U1589 ( .A(regs[852]), .B(n75), .C(regs[788]), .D(n114), .Q(n1303) );
  AOI220 U1590 ( .A(regs[372]), .B(n1566), .C(regs[308]), .D(n74), .Q(n1308)
         );
  AOI220 U1591 ( .A(regs[118]), .B(n1566), .C(regs[54]), .D(n1565), .Q(n1362)
         );
  AOI220 U1592 ( .A(regs[887]), .B(n1566), .C(regs[823]), .D(n74), .Q(n1370)
         );
  AOI220 U1593 ( .A(regs[375]), .B(n1566), .C(regs[311]), .D(n74), .Q(n1374)
         );
  AOI220 U1594 ( .A(regs[631]), .B(n1566), .C(regs[567]), .D(n74), .Q(n1380)
         );
  AOI220 U1595 ( .A(regs[119]), .B(n1566), .C(regs[55]), .D(n74), .Q(n1384) );
  AOI220 U1596 ( .A(regs[888]), .B(n1566), .C(regs[824]), .D(n74), .Q(n1392)
         );
  AOI220 U1597 ( .A(regs[376]), .B(n1566), .C(regs[312]), .D(n74), .Q(n1396)
         );
  AOI220 U1598 ( .A(regs[216]), .B(n113), .C(regs[152]), .D(n72), .Q(n1407) );
  AOI220 U1599 ( .A(regs[120]), .B(n1566), .C(regs[56]), .D(n74), .Q(n1406) );
  AOI220 U1600 ( .A(regs[88]), .B(n75), .C(regs[24]), .D(n114), .Q(n1405) );
  AOI220 U1601 ( .A(regs[985]), .B(n113), .C(regs[921]), .D(n72), .Q(n1415) );
  AOI220 U1602 ( .A(regs[857]), .B(n75), .C(regs[793]), .D(n114), .Q(n1413) );
  AOI220 U1603 ( .A(regs[473]), .B(n113), .C(regs[409]), .D(n72), .Q(n1419) );
  AOI220 U1604 ( .A(regs[377]), .B(n1566), .C(regs[313]), .D(n74), .Q(n1418)
         );
  AOI220 U1605 ( .A(regs[474]), .B(n113), .C(regs[410]), .D(n72), .Q(n1441) );
  AOI220 U1606 ( .A(regs[218]), .B(n113), .C(regs[154]), .D(n72), .Q(n1451) );
  AOI220 U1607 ( .A(regs[859]), .B(n75), .C(regs[795]), .D(n114), .Q(n1457) );
  AOI220 U1608 ( .A(regs[379]), .B(n73), .C(regs[315]), .D(n74), .Q(n1462) );
  AOI220 U1609 ( .A(regs[603]), .B(n75), .C(regs[539]), .D(n114), .Q(n1467) );
  AOI220 U1610 ( .A(regs[348]), .B(n75), .C(regs[284]), .D(n1567), .Q(n1483)
         );
  AOI220 U1611 ( .A(regs[92]), .B(n75), .C(regs[28]), .D(n1567), .Q(n1493) );
  AOI220 U1612 ( .A(regs[381]), .B(n1566), .C(regs[317]), .D(n74), .Q(n1506)
         );
  AOI220 U1613 ( .A(regs[93]), .B(n75), .C(regs[29]), .D(n1567), .Q(n1515) );
  AOI220 U1614 ( .A(regs[1022]), .B(n112), .C(regs[958]), .D(n1561), .Q(n1526)
         );
  AOI220 U1615 ( .A(regs[990]), .B(n113), .C(regs[926]), .D(n1563), .Q(n1525)
         );
  AOI220 U1616 ( .A(regs[894]), .B(n73), .C(regs[830]), .D(n1565), .Q(n1524)
         );
  AOI220 U1617 ( .A(regs[862]), .B(n1568), .C(regs[798]), .D(n114), .Q(n1523)
         );
  AOI220 U1618 ( .A(regs[606]), .B(n1568), .C(regs[542]), .D(n114), .Q(n1533)
         );
  AOI220 U1619 ( .A(regs[511]), .B(n112), .C(regs[447]), .D(n1561), .Q(n1552)
         );
  AOI220 U1620 ( .A(regs[479]), .B(n113), .C(regs[415]), .D(n1563), .Q(n1551)
         );
  AOI220 U1621 ( .A(regs[383]), .B(n73), .C(regs[319]), .D(n1565), .Q(n1550)
         );
  AOI220 U1622 ( .A(regs[639]), .B(n1566), .C(regs[575]), .D(n74), .Q(n1558)
         );
  AOI220 U1623 ( .A(regs[127]), .B(n1566), .C(regs[63]), .D(n74), .Q(n1570) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Mmemread, ex_con_Mmemwrite, ex_con_Malupc8, ex_con_Wmemtoreg,
         mem_con_Malupc8, mem_con_Wmemtoreg, wb_con_Wmemtoreg,
         u_fetch_jmux_i_addr_pc4_3_, u_fetch_jmux_i_addr_pc4_4_,
         u_fetch_jmux_i_addr_pc4_5_, u_fetch_jmux_i_addr_pc4_6_,
         u_fetch_jmux_i_addr_pc4_7_, u_fetch_jmux_i_addr_pc4_8_,
         u_fetch_jmux_i_addr_pc4_9_, u_fetch_jmux_i_addr_pc4_10_,
         u_fetch_jmux_i_addr_pc4_11_, u_fetch_jmux_i_addr_pc4_12_,
         u_fetch_jmux_i_addr_pc4_13_, u_fetch_jmux_i_addr_pc4_14_,
         u_fetch_jmux_i_addr_pc4_15_, u_fetch_jmux_i_addr_pc4_16_,
         u_fetch_jmux_i_addr_pc4_17_, u_fetch_jmux_i_addr_pc4_18_,
         u_fetch_jmux_i_addr_pc4_19_, u_fetch_jmux_i_addr_pc4_20_,
         u_fetch_jmux_i_addr_pc4_21_, u_fetch_jmux_i_addr_pc4_22_,
         u_fetch_jmux_i_addr_pc4_23_, u_fetch_jmux_i_addr_pc4_24_,
         u_fetch_jmux_i_addr_pc4_25_, u_fetch_jmux_i_addr_pc4_26_,
         u_fetch_jmux_i_addr_pc4_27_, u_fetch_jmux_i_addr_pc4_28_,
         u_fetch_jmux_i_addr_pc4_29_, u_fetch_jmux_i_addr_pc4_30_,
         u_fetch_jmux_i_addr_pc4_31_, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, u_decode_n6, u_decode_n1, u_decode_for_o_con_fa_0_,
         u_decode_for_o_con_fa_1_, u_decode_for_o_con_fa_2_,
         u_decode_control_o_con_regwrite, u_decode_control_o_con_memtoreg,
         u_decode_control_o_con_memwrite, u_decode_control_o_con_memread,
         u_decode_jbcon_o_con_aluPC4, u_decode_control_o_con_regdst,
         u_decode_control_o_con_alusrc, u_decode_control_o_con_aluop_0_,
         u_decode_control_o_con_aluop_1_, u_decode_control_o_con_aluop_2_,
         u_decode_control_o_con_aluop_3_, u_decode_control_o_con_aluop_4_,
         u_decode_control_o_con_aluop_5_, u_decode_add_x_16_n182,
         u_decode_add_x_16_n181, u_decode_add_x_16_n178,
         u_decode_add_x_16_n176, u_decode_add_x_16_n175,
         u_decode_add_x_16_n158, u_decode_add_x_16_n156,
         u_decode_add_x_16_n155, u_decode_add_x_16_n154,
         u_decode_add_x_16_n153, u_decode_add_x_16_n152,
         u_decode_add_x_16_n151, u_decode_add_x_16_n150,
         u_decode_add_x_16_n149, u_decode_add_x_16_n148,
         u_decode_add_x_16_n147, u_decode_add_x_16_n146,
         u_decode_add_x_16_n145, u_decode_add_x_16_n144,
         u_decode_add_x_16_n143, u_decode_add_x_16_n142,
         u_decode_add_x_16_n138, u_decode_add_x_16_n137,
         u_decode_add_x_16_n136, u_decode_add_x_16_n135,
         u_decode_add_x_16_n134, u_decode_add_x_16_n133,
         u_decode_add_x_16_n132, u_decode_add_x_16_n131,
         u_decode_add_x_16_n130, u_decode_add_x_16_n129,
         u_decode_add_x_16_n128, u_decode_add_x_16_n127,
         u_decode_add_x_16_n126, u_decode_add_x_16_n125,
         u_decode_add_x_16_n124, u_decode_add_x_16_n123,
         u_decode_add_x_16_n122, u_decode_add_x_16_n121,
         u_decode_add_x_16_n120, u_decode_add_x_16_n119,
         u_decode_add_x_16_n118, u_decode_add_x_16_n117,
         u_decode_add_x_16_n116, u_decode_add_x_16_n115,
         u_decode_add_x_16_n114, u_decode_add_x_16_n113,
         u_decode_add_x_16_n112, u_decode_add_x_16_n111,
         u_decode_add_x_16_n107, u_decode_add_x_16_n106,
         u_decode_add_x_16_n105, u_decode_add_x_16_n104,
         u_decode_add_x_16_n103, u_decode_add_x_16_n102,
         u_decode_add_x_16_n101, u_decode_add_x_16_n100, u_decode_add_x_16_n99,
         u_decode_add_x_16_n98, u_decode_add_x_16_n96, u_decode_add_x_16_n94,
         u_decode_add_x_16_n93, u_decode_add_x_16_n92, u_decode_add_x_16_n91,
         u_decode_add_x_16_n90, u_decode_add_x_16_n89, u_decode_add_x_16_n88,
         u_decode_add_x_16_n87, u_decode_add_x_16_n86, u_decode_add_x_16_n84,
         u_decode_add_x_16_n82, u_decode_add_x_16_n81, u_decode_add_x_16_n80,
         u_decode_add_x_16_n79, u_decode_add_x_16_n78, u_decode_add_x_16_n77,
         u_decode_add_x_16_n76, u_decode_add_x_16_n75, u_decode_add_x_16_n74,
         u_decode_add_x_16_n73, u_decode_add_x_16_n72, u_decode_add_x_16_n71,
         u_decode_add_x_16_n70, u_decode_add_x_16_n69, u_decode_add_x_16_n68,
         u_decode_add_x_16_n67, u_decode_add_x_16_n66, u_decode_add_x_16_n65,
         u_decode_add_x_16_n64, u_decode_add_x_16_n63, u_decode_add_x_16_n62,
         u_decode_add_x_16_n61, u_decode_add_x_16_n60, u_decode_add_x_16_n59,
         u_decode_add_x_16_n58, u_decode_add_x_16_n57, u_decode_add_x_16_n56,
         u_decode_add_x_16_n55, u_decode_add_x_16_n54, u_decode_add_x_16_n53,
         u_decode_add_x_16_n52, u_decode_add_x_16_n51, u_decode_add_x_16_n50,
         u_decode_add_x_16_n49, u_decode_add_x_16_n48, u_decode_add_x_16_n47,
         u_decode_add_x_16_n46, u_decode_add_x_16_n45, u_decode_add_x_16_n44,
         u_decode_add_x_16_n43, u_decode_add_x_16_n42, u_decode_add_x_16_n41,
         u_decode_add_x_16_n40, u_decode_add_x_16_n39, u_decode_add_x_16_n38,
         u_decode_add_x_16_n37, u_decode_add_x_16_n36, u_decode_add_x_16_n35,
         u_decode_add_x_16_n34, u_decode_add_x_16_n33, u_decode_add_x_16_n32,
         u_decode_add_x_16_n31, u_decode_add_x_16_n30, u_decode_add_x_16_n29,
         u_decode_add_x_16_n25, u_decode_add_x_16_n24, u_decode_add_x_16_n21,
         u_decode_add_x_16_n19, u_decode_add_x_16_n18, u_decode_add_x_16_n16,
         u_decode_add_x_16_n14, u_decode_add_x_16_n11, u_decode_add_x_16_n9,
         u_decode_add_x_16_n7, u_decode_add_x_16_n5, u_decode_add_x_16_n3,
         add_x_4_n77, add_x_4_n76, add_x_4_n73, add_x_4_n70, add_x_4_n69,
         add_x_4_n68, add_x_4_n64, add_x_4_n61, add_x_4_n60, add_x_4_n57,
         add_x_4_n54, add_x_4_n53, add_x_4_n52, add_x_4_n51, add_x_4_n48,
         add_x_4_n45, add_x_4_n44, add_x_4_n43, add_x_4_n39, add_x_4_n36,
         add_x_4_n35, add_x_4_n34, add_x_4_n33, add_x_4_n29, add_x_4_n26,
         add_x_4_n25, add_x_4_n24, add_x_4_n20, add_x_4_n17, add_x_4_n16,
         add_x_4_n15, add_x_4_n14, add_x_4_n13, add_x_4_n12, add_x_4_n11,
         add_x_4_n10, add_x_4_n9, add_x_4_n8, add_x_4_n7, add_x_4_n6,
         add_x_4_n5, add_x_4_n4, add_x_4_n3, add_x_4_n2, add_x_4_n1,
         add_x_1_n72, add_x_1_n71, add_x_1_n65, add_x_1_n64, add_x_1_n63,
         add_x_1_n62, add_x_1_n56, add_x_1_n55, add_x_1_n49, add_x_1_n48,
         add_x_1_n47, add_x_1_n46, add_x_1_n40, add_x_1_n39, add_x_1_n38,
         add_x_1_n37, add_x_1_n31, add_x_1_n30, add_x_1_n29, add_x_1_n28,
         add_x_1_n27, add_x_1_n21, add_x_1_n17, add_x_1_n16, add_x_1_n15,
         add_x_1_n14, add_x_1_n13, add_x_1_n12, add_x_1_n11, add_x_1_n10,
         add_x_1_n9, add_x_1_n8, add_x_1_n7, add_x_1_n6, add_x_1_n5,
         add_x_1_n4, add_x_1_n3, add_x_1_n2, add_x_1_n1, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449;
  wire   [31:2] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [27:2] id_addr_pc4;
  wire   [31:26] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] wb_data_memout;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] mem_data_alures;
  wire   [31:2] mem_data_pc4;
  wire   [31:0] u_mem_resmux_o_data_alu;
  wire   [31:0] u_mem_pc8;
  wire   [1:0] u_decode_jbcon_o_con_bop;
  wire   [31:0] u_decode_pcadd_o_addr_pcbranchE;
  wire   [2:0] u_decode_for_o_con_fb;
  wire   [31:0] u_decode_regbank_o_data_Rt;

  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext({n242, 
        n242, n242, n242, n242, n242, n242, n242, n242, n242, n242, n242, n242, 
        n242, n242, ex_data_immext[31], ex_addr_rd, ex_data_immext[10:9], n246, 
        ex_data_immext[7], n245, ex_data_immext[5:0]}), .i_addr_rt(ex_addr_rt), 
        .i_addr_rd({n242, n242, n242, n242, n242}), .i_data_FEalures(
        data_address), .i_data_FMalures(mem_data_alures), .i_data_FMmemout(
        wb_data_memout), .i_data_FWmemout(for_memout), .i_con_Efamux(
        for_o_con_Efamux), .i_con_Efbmux(for_o_con_Efbmux), .i_con_Ealuop(
        ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), .i_con_Eregdst(
        ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), .i_con_Mmemwrite(
        ex_con_Mmemwrite), .i_con_Malupc8(ex_con_Malupc8), .i_con_Wmemtoreg(
        ex_con_Wmemtoreg), .i_con_Wregwrite(ex_con_Wregwrite), .i_con_bop(
        ex_con_bop), .o_data_alures(data_address), .o_data_rt(write_data), 
        .o_addr_regdst(mem_addr_regdst), .o_con_Mmemread(mem_read), 
        .o_con_Mmemwrite(mem_write), .o_con_Malupc8(mem_con_Malupc8), 
        .o_con_Wmemtoreg(mem_con_Wmemtoreg), .o_con_Wregwrite(
        mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), .o_addr_Mrt(
        for_addr_rtM), .o_con_ifbranch(if_con_b), .o_data_pc4_31_(
        mem_data_pc4[31]), .o_data_pc4_30_(mem_data_pc4[30]), .o_data_pc4_29_(
        mem_data_pc4[29]), .o_data_pc4_28_(mem_data_pc4[28]), .o_data_pc4_27_(
        mem_data_pc4[27]), .o_data_pc4_26_(mem_data_pc4[26]), .o_data_pc4_25_(
        mem_data_pc4[25]), .o_data_pc4_24_(mem_data_pc4[24]), .o_data_pc4_23_(
        mem_data_pc4[23]), .o_data_pc4_22_(mem_data_pc4[22]), .o_data_pc4_21_(
        mem_data_pc4[21]), .o_data_pc4_20_(mem_data_pc4[20]), .o_data_pc4_19_(
        mem_data_pc4[19]), .o_data_pc4_18_(mem_data_pc4[18]), .o_data_pc4_17_(
        mem_data_pc4[17]), .o_data_pc4_16__BAR(mem_data_pc4[16]), 
        .o_data_pc4_15_(mem_data_pc4[15]), .o_data_pc4_14_(mem_data_pc4[14]), 
        .o_data_pc4_13_(mem_data_pc4[13]), .o_data_pc4_12_(mem_data_pc4[12]), 
        .o_data_pc4_11_(mem_data_pc4[11]), .o_data_pc4_10_(mem_data_pc4[10]), 
        .o_data_pc4_9_(mem_data_pc4[9]), .o_data_pc4_8_(mem_data_pc4[8]), 
        .o_data_pc4_7_(mem_data_pc4[7]), .o_data_pc4_6_(mem_data_pc4[6]), 
        .o_data_pc4_5_(mem_data_pc4[5]), .o_data_pc4_4_(mem_data_pc4[4]), 
        .o_data_pc4_3_(mem_data_pc4[3]), .o_data_pc4_2_(mem_data_pc4[2]), 
        .o_data_pc4_1_(u_mem_pc8[1]), .o_data_pc4_0_(u_mem_pc8[0]) );
  DFC1 u_fetch_pipe_pc4_reg_0_ ( .D(instruction_address[0]), .C(clk), .RN(
        rst_n), .Q(u_decode_pcadd_o_addr_pcbranchE[0]) );
  DFC1 u_fetch_pipe_pc4_reg_1_ ( .D(instruction_address[1]), .C(clk), .RN(
        rst_n), .Q(u_decode_pcadd_o_addr_pcbranchE[1]) );
  DFC1 u_fetch_pipe_pc4_reg_2_ ( .D(n228), .C(clk), .RN(rst_n), .Q(
        id_addr_pc4[2]) );
  DFC1 u_fetch_pipe_pc4_reg_3_ ( .D(u_fetch_jmux_i_addr_pc4_3_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[3]) );
  DFC1 u_fetch_pipe_pc4_reg_4_ ( .D(u_fetch_jmux_i_addr_pc4_4_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[4]) );
  DFC1 u_fetch_pipe_pc4_reg_5_ ( .D(u_fetch_jmux_i_addr_pc4_5_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[5]) );
  DFC1 u_fetch_pipe_pc4_reg_6_ ( .D(u_fetch_jmux_i_addr_pc4_6_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[6]) );
  DFC1 u_fetch_pipe_pc4_reg_7_ ( .D(u_fetch_jmux_i_addr_pc4_7_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[7]) );
  DFC1 u_fetch_pipe_pc4_reg_8_ ( .D(u_fetch_jmux_i_addr_pc4_8_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[8]) );
  DFC1 u_fetch_pipe_pc4_reg_9_ ( .D(u_fetch_jmux_i_addr_pc4_9_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[9]) );
  DFC1 u_fetch_pipe_pc4_reg_10_ ( .D(u_fetch_jmux_i_addr_pc4_10_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[10]) );
  DFC1 u_fetch_pipe_pc4_reg_11_ ( .D(u_fetch_jmux_i_addr_pc4_11_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[11]) );
  DFC1 u_fetch_pipe_pc4_reg_12_ ( .D(u_fetch_jmux_i_addr_pc4_12_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[12]) );
  DFC1 u_fetch_pipe_pc4_reg_13_ ( .D(u_fetch_jmux_i_addr_pc4_13_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[13]) );
  DFC1 u_fetch_pipe_pc4_reg_14_ ( .D(u_fetch_jmux_i_addr_pc4_14_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[14]) );
  DFC1 u_fetch_pipe_pc4_reg_15_ ( .D(u_fetch_jmux_i_addr_pc4_15_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[15]) );
  DFC1 u_fetch_pipe_pc4_reg_16_ ( .D(u_fetch_jmux_i_addr_pc4_16_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[16]) );
  DFC1 u_fetch_pipe_pc4_reg_17_ ( .D(u_fetch_jmux_i_addr_pc4_17_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[17]) );
  DFC1 u_fetch_pipe_pc4_reg_18_ ( .D(u_fetch_jmux_i_addr_pc4_18_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[18]) );
  DFC1 u_fetch_pipe_pc4_reg_19_ ( .D(u_fetch_jmux_i_addr_pc4_19_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[19]) );
  DFC1 u_fetch_pipe_pc4_reg_20_ ( .D(u_fetch_jmux_i_addr_pc4_20_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[20]) );
  DFC1 u_fetch_pipe_pc4_reg_21_ ( .D(u_fetch_jmux_i_addr_pc4_21_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[21]) );
  DFC1 u_fetch_pipe_pc4_reg_22_ ( .D(u_fetch_jmux_i_addr_pc4_22_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[22]) );
  DFC1 u_fetch_pipe_pc4_reg_23_ ( .D(u_fetch_jmux_i_addr_pc4_23_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[23]) );
  DFC1 u_fetch_pipe_pc4_reg_24_ ( .D(u_fetch_jmux_i_addr_pc4_24_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[24]) );
  DFC1 u_fetch_pipe_pc4_reg_25_ ( .D(u_fetch_jmux_i_addr_pc4_25_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[25]) );
  DFC1 u_fetch_pipe_pc4_reg_26_ ( .D(u_fetch_jmux_i_addr_pc4_26_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[26]) );
  DFC1 u_fetch_pipe_pc4_reg_27_ ( .D(u_fetch_jmux_i_addr_pc4_27_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[27]) );
  DFC1 u_fetch_pipe_pc4_reg_28_ ( .D(u_fetch_jmux_i_addr_pc4_28_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[28]) );
  DFC1 u_fetch_pipe_pc4_reg_29_ ( .D(u_fetch_jmux_i_addr_pc4_29_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[29]), .QN(n238) );
  DFC1 u_fetch_pipe_pc4_reg_30_ ( .D(u_fetch_jmux_i_addr_pc4_30_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[30]), .QN(n237) );
  DFC1 u_fetch_pipe_pc4_reg_31_ ( .D(u_fetch_jmux_i_addr_pc4_31_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[31]), .QN(n239) );
  DFC1 u_fetch_pipe_instr_reg_0_ ( .D(read_instruction[0]), .C(clk), .RN(rst_n), .Q(if_addr_j[2]) );
  DFC1 u_fetch_pipe_instr_reg_1_ ( .D(read_instruction[1]), .C(clk), .RN(rst_n), .Q(if_addr_j[3]) );
  DFC1 u_fetch_pipe_instr_reg_2_ ( .D(read_instruction[2]), .C(clk), .RN(rst_n), .Q(if_addr_j[4]) );
  DFC1 u_fetch_pipe_instr_reg_3_ ( .D(read_instruction[3]), .C(clk), .RN(rst_n), .Q(if_addr_j[5]) );
  DFC1 u_fetch_pipe_instr_reg_4_ ( .D(read_instruction[4]), .C(clk), .RN(rst_n), .Q(if_addr_j[6]) );
  DFC1 u_fetch_pipe_instr_reg_5_ ( .D(read_instruction[5]), .C(clk), .RN(rst_n), .Q(if_addr_j[7]), .QN(n218) );
  DFC1 u_fetch_pipe_instr_reg_6_ ( .D(read_instruction[6]), .C(clk), .RN(rst_n), .Q(if_addr_j[8]) );
  DFC1 u_fetch_pipe_instr_reg_7_ ( .D(read_instruction[7]), .C(clk), .RN(rst_n), .Q(if_addr_j[9]) );
  DFC1 u_fetch_pipe_instr_reg_8_ ( .D(read_instruction[8]), .C(clk), .RN(rst_n), .Q(if_addr_j[10]) );
  DFC1 u_fetch_pipe_instr_reg_9_ ( .D(read_instruction[9]), .C(clk), .RN(rst_n), .Q(if_addr_j[11]) );
  DFC1 u_fetch_pipe_instr_reg_10_ ( .D(read_instruction[10]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[12]) );
  DFC1 u_fetch_pipe_instr_reg_11_ ( .D(read_instruction[11]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[13]) );
  DFC1 u_fetch_pipe_instr_reg_12_ ( .D(read_instruction[12]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[14]) );
  DFC1 u_fetch_pipe_instr_reg_13_ ( .D(read_instruction[13]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[15]) );
  DFC1 u_fetch_pipe_instr_reg_14_ ( .D(read_instruction[14]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[16]) );
  DFC1 u_fetch_pipe_instr_reg_21_ ( .D(read_instruction[21]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[23]), .QN(n211) );
  DFC1 u_fetch_pipe_instr_reg_22_ ( .D(read_instruction[22]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[24]), .QN(n210) );
  DFC1 u_fetch_pipe_instr_reg_23_ ( .D(read_instruction[23]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[25]), .QN(n209) );
  DFC1 u_fetch_pipe_instr_reg_24_ ( .D(read_instruction[24]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[26]), .QN(n217) );
  DFC1 u_fetch_pipe_instr_reg_25_ ( .D(read_instruction[25]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[27]), .QN(n213) );
  DFC1 u_fetch_pipe_instr_reg_26_ ( .D(read_instruction[26]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[26]), .QN(n204) );
  DFC1 u_fetch_pipe_instr_reg_27_ ( .D(read_instruction[27]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[27]), .QN(n212) );
  DFC1 u_fetch_pipe_instr_reg_28_ ( .D(read_instruction[28]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[28]), .QN(n208) );
  DFC1 u_fetch_pipe_instr_reg_29_ ( .D(read_instruction[29]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[29]), .QN(n205) );
  DFC1 u_fetch_pipe_instr_reg_30_ ( .D(read_instruction[30]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[30]) );
  DFC1 u_fetch_pipe_instr_reg_31_ ( .D(read_instruction[31]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[31]), .QN(n219) );
  DFC1 u_mem_pipe_data_memout_reg_0_ ( .D(read_data[0]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[0]) );
  DFC1 u_mem_pipe_data_memout_reg_1_ ( .D(read_data[1]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[1]) );
  DFC1 u_mem_pipe_data_memout_reg_2_ ( .D(read_data[2]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[2]) );
  DFC1 u_mem_pipe_data_memout_reg_3_ ( .D(read_data[3]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[3]) );
  DFC1 u_mem_pipe_data_memout_reg_4_ ( .D(read_data[4]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[4]) );
  DFC1 u_mem_pipe_data_memout_reg_5_ ( .D(read_data[5]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[5]) );
  DFC1 u_mem_pipe_data_memout_reg_6_ ( .D(read_data[6]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[6]) );
  DFC1 u_mem_pipe_data_memout_reg_7_ ( .D(read_data[7]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[7]) );
  DFC1 u_mem_pipe_data_memout_reg_8_ ( .D(read_data[8]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[8]) );
  DFC1 u_mem_pipe_data_memout_reg_9_ ( .D(read_data[9]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[9]) );
  DFC1 u_mem_pipe_data_memout_reg_10_ ( .D(read_data[10]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[10]) );
  DFC1 u_mem_pipe_data_memout_reg_11_ ( .D(read_data[11]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[11]) );
  DFC1 u_mem_pipe_data_memout_reg_12_ ( .D(read_data[12]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[12]) );
  DFC1 u_mem_pipe_data_memout_reg_13_ ( .D(read_data[13]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[13]) );
  DFC1 u_mem_pipe_data_memout_reg_14_ ( .D(read_data[14]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[14]) );
  DFC1 u_mem_pipe_data_memout_reg_15_ ( .D(read_data[15]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[15]) );
  DFC1 u_mem_pipe_data_memout_reg_16_ ( .D(read_data[16]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[16]) );
  DFC1 u_mem_pipe_data_memout_reg_17_ ( .D(read_data[17]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[17]) );
  DFC1 u_mem_pipe_data_memout_reg_18_ ( .D(read_data[18]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[18]) );
  DFC1 u_mem_pipe_data_memout_reg_19_ ( .D(read_data[19]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[19]) );
  DFC1 u_mem_pipe_data_memout_reg_20_ ( .D(read_data[20]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[20]) );
  DFC1 u_mem_pipe_data_memout_reg_21_ ( .D(read_data[21]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[21]) );
  DFC1 u_mem_pipe_data_memout_reg_22_ ( .D(read_data[22]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[22]) );
  DFC1 u_mem_pipe_data_memout_reg_23_ ( .D(read_data[23]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[23]) );
  DFC1 u_mem_pipe_data_memout_reg_24_ ( .D(read_data[24]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[24]) );
  DFC1 u_mem_pipe_data_memout_reg_25_ ( .D(read_data[25]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[25]) );
  DFC1 u_mem_pipe_data_memout_reg_26_ ( .D(read_data[26]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[26]) );
  DFC1 u_mem_pipe_data_memout_reg_27_ ( .D(read_data[27]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[27]) );
  DFC1 u_mem_pipe_data_memout_reg_28_ ( .D(read_data[28]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[28]) );
  DFC1 u_mem_pipe_data_memout_reg_29_ ( .D(read_data[29]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[29]) );
  DFC1 u_mem_pipe_data_memout_reg_30_ ( .D(read_data[30]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[30]) );
  DFC1 u_mem_pipe_data_memout_reg_31_ ( .D(read_data[31]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[31]) );
  DFC1 u_mem_pipe_rt_reg_4_ ( .D(for_addr_rtM[4]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[4]) );
  DFC1 u_mem_pipe_con_FWmemread_reg ( .D(ex_con_Mmemread), .C(clk), .RN(rst_n), 
        .Q(for_FWmemread) );
  DFC1 u_mem_pipe_rt_reg_0_ ( .D(for_addr_rtM[0]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[0]) );
  DFC1 u_mem_pipe_rt_reg_1_ ( .D(for_addr_rtM[1]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[1]) );
  DFC1 u_mem_pipe_rt_reg_2_ ( .D(for_addr_rtM[2]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[2]) );
  DFC1 u_mem_pipe_rt_reg_3_ ( .D(for_addr_rtM[3]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[3]) );
  DFC1 u_mem_pipe_con_Wregwrite_reg ( .D(mem_con_Wregwrite), .C(clk), .RN(
        rst_n), .Q(id_con_Wregwrite) );
  DFC1 u_mem_pipe_addr_regdst_reg_0_ ( .D(mem_addr_regdst[0]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[0]) );
  DFC1 u_mem_pipe_addr_regdst_reg_1_ ( .D(mem_addr_regdst[1]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[1]) );
  DFC1 u_mem_pipe_addr_regdst_reg_2_ ( .D(mem_addr_regdst[2]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[2]) );
  DFC1 u_mem_pipe_addr_regdst_reg_4_ ( .D(mem_addr_regdst[4]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[4]) );
  DFC1 u_mem_pipe_data_alures_reg_0_ ( .D(u_mem_resmux_o_data_alu[0]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[0]) );
  DFC1 u_mem_pipe_data_alures_reg_1_ ( .D(u_mem_resmux_o_data_alu[1]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[1]) );
  DFC1 u_mem_pipe_data_alures_reg_2_ ( .D(u_mem_resmux_o_data_alu[2]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[2]) );
  DFC1 u_mem_pipe_data_alures_reg_3_ ( .D(u_mem_resmux_o_data_alu[3]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[3]) );
  DFC1 u_mem_pipe_data_alures_reg_4_ ( .D(u_mem_resmux_o_data_alu[4]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[4]) );
  DFC1 u_mem_pipe_data_alures_reg_5_ ( .D(u_mem_resmux_o_data_alu[5]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[5]) );
  DFC1 u_mem_pipe_data_alures_reg_6_ ( .D(u_mem_resmux_o_data_alu[6]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[6]) );
  DFC1 u_mem_pipe_data_alures_reg_7_ ( .D(u_mem_resmux_o_data_alu[7]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[7]) );
  DFC1 u_mem_pipe_data_alures_reg_8_ ( .D(u_mem_resmux_o_data_alu[8]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[8]) );
  DFC1 u_mem_pipe_data_alures_reg_9_ ( .D(u_mem_resmux_o_data_alu[9]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[9]) );
  DFC1 u_mem_pipe_data_alures_reg_10_ ( .D(u_mem_resmux_o_data_alu[10]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[10]) );
  DFC1 u_mem_pipe_data_alures_reg_11_ ( .D(u_mem_resmux_o_data_alu[11]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[11]) );
  DFC1 u_mem_pipe_data_alures_reg_12_ ( .D(u_mem_resmux_o_data_alu[12]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[12]) );
  DFC1 u_mem_pipe_data_alures_reg_13_ ( .D(u_mem_resmux_o_data_alu[13]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[13]) );
  DFC1 u_mem_pipe_data_alures_reg_14_ ( .D(u_mem_resmux_o_data_alu[14]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[14]) );
  DFC1 u_mem_pipe_data_alures_reg_15_ ( .D(u_mem_resmux_o_data_alu[15]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[15]) );
  DFC1 u_mem_pipe_data_alures_reg_16_ ( .D(u_mem_resmux_o_data_alu[16]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[16]) );
  DFC1 u_mem_pipe_data_alures_reg_17_ ( .D(u_mem_resmux_o_data_alu[17]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[17]) );
  DFC1 u_mem_pipe_data_alures_reg_18_ ( .D(u_mem_resmux_o_data_alu[18]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[18]) );
  DFC1 u_mem_pipe_data_alures_reg_19_ ( .D(u_mem_resmux_o_data_alu[19]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[19]) );
  DFC1 u_mem_pipe_data_alures_reg_20_ ( .D(u_mem_resmux_o_data_alu[20]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[20]) );
  DFC1 u_mem_pipe_data_alures_reg_21_ ( .D(u_mem_resmux_o_data_alu[21]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[21]) );
  DFC1 u_mem_pipe_data_alures_reg_22_ ( .D(u_mem_resmux_o_data_alu[22]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[22]) );
  DFC1 u_mem_pipe_data_alures_reg_23_ ( .D(u_mem_resmux_o_data_alu[23]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[23]) );
  DFC1 u_mem_pipe_data_alures_reg_24_ ( .D(u_mem_resmux_o_data_alu[24]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[24]) );
  DFC1 u_mem_pipe_data_alures_reg_25_ ( .D(u_mem_resmux_o_data_alu[25]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[25]) );
  DFC1 u_mem_pipe_data_alures_reg_26_ ( .D(u_mem_resmux_o_data_alu[26]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[26]) );
  DFC1 u_mem_pipe_data_alures_reg_27_ ( .D(u_mem_resmux_o_data_alu[27]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[27]) );
  DFC1 u_mem_pipe_data_alures_reg_28_ ( .D(u_mem_resmux_o_data_alu[28]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[28]) );
  DFC1 u_mem_pipe_data_alures_reg_29_ ( .D(u_mem_resmux_o_data_alu[29]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[29]) );
  DFC1 u_mem_pipe_data_alures_reg_30_ ( .D(u_mem_resmux_o_data_alu[30]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[30]) );
  DFC1 u_mem_pipe_data_alures_reg_31_ ( .D(u_mem_resmux_o_data_alu[31]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[31]) );
  DFC1 u_fetch_u_pc_program_counter_reg_0_ ( .D(n137), .C(clk), .RN(rst_n), 
        .Q(instruction_address[0]), .QN(n241) );
  DFC1 u_fetch_u_pc_program_counter_reg_1_ ( .D(n136), .C(clk), .RN(rst_n), 
        .Q(instruction_address[1]), .QN(n240) );
  DFC1 u_fetch_u_pc_program_counter_reg_2_ ( .D(n135), .C(clk), .RN(rst_n), 
        .Q(instruction_address[2]), .QN(n228) );
  DFC1 u_fetch_u_pc_program_counter_reg_3_ ( .D(n134), .C(clk), .RN(rst_n), 
        .Q(instruction_address[3]), .QN(n236) );
  DFC1 u_fetch_u_pc_program_counter_reg_4_ ( .D(n133), .C(clk), .RN(rst_n), 
        .Q(instruction_address[4]), .QN(n223) );
  DFC1 u_fetch_u_pc_program_counter_reg_5_ ( .D(n132), .C(clk), .RN(rst_n), 
        .Q(instruction_address[5]), .QN(n235) );
  DFC1 u_fetch_u_pc_program_counter_reg_6_ ( .D(n131), .C(clk), .RN(rst_n), 
        .Q(instruction_address[6]), .QN(n227) );
  DFC1 u_fetch_u_pc_program_counter_reg_7_ ( .D(n130), .C(clk), .RN(rst_n), 
        .Q(instruction_address[7]), .QN(n232) );
  DFC1 u_fetch_u_pc_program_counter_reg_8_ ( .D(n129), .C(clk), .RN(rst_n), 
        .Q(instruction_address[8]), .QN(n222) );
  DFC1 u_fetch_u_pc_program_counter_reg_9_ ( .D(n128), .C(clk), .RN(rst_n), 
        .Q(instruction_address[9]), .QN(n234) );
  DFC1 u_fetch_u_pc_program_counter_reg_10_ ( .D(n127), .C(clk), .RN(rst_n), 
        .Q(instruction_address[10]), .QN(n221) );
  DFC1 u_fetch_u_pc_program_counter_reg_11_ ( .D(n126), .C(clk), .RN(rst_n), 
        .Q(instruction_address[11]), .QN(n233) );
  DFC1 u_fetch_u_pc_program_counter_reg_12_ ( .D(n125), .C(clk), .RN(rst_n), 
        .Q(instruction_address[12]), .QN(n226) );
  DFC1 u_fetch_u_pc_program_counter_reg_13_ ( .D(n124), .C(clk), .RN(rst_n), 
        .Q(instruction_address[13]), .QN(n231) );
  DFC1 u_fetch_u_pc_program_counter_reg_14_ ( .D(n123), .C(clk), .RN(rst_n), 
        .Q(instruction_address[14]), .QN(n224) );
  DFC1 u_fetch_u_pc_program_counter_reg_15_ ( .D(n122), .C(clk), .RN(rst_n), 
        .Q(instruction_address[15]), .QN(n230) );
  DFC1 u_fetch_u_pc_program_counter_reg_16_ ( .D(n121), .C(clk), .RN(rst_n), 
        .Q(instruction_address[16]), .QN(n225) );
  DFC1 u_fetch_u_pc_program_counter_reg_17_ ( .D(n120), .C(clk), .RN(rst_n), 
        .Q(instruction_address[17]), .QN(n229) );
  DFC1 u_fetch_u_pc_program_counter_reg_18_ ( .D(n119), .C(clk), .RN(rst_n), 
        .Q(instruction_address[18]) );
  DFC1 u_fetch_u_pc_program_counter_reg_19_ ( .D(n118), .C(clk), .RN(rst_n), 
        .Q(instruction_address[19]) );
  DFC1 u_fetch_u_pc_program_counter_reg_20_ ( .D(n117), .C(clk), .RN(rst_n), 
        .Q(instruction_address[20]) );
  DFC1 u_fetch_u_pc_program_counter_reg_21_ ( .D(n116), .C(clk), .RN(rst_n), 
        .Q(instruction_address[21]) );
  DFC1 u_fetch_u_pc_program_counter_reg_22_ ( .D(n115), .C(clk), .RN(rst_n), 
        .Q(instruction_address[22]) );
  DFC1 u_fetch_u_pc_program_counter_reg_23_ ( .D(n114), .C(clk), .RN(rst_n), 
        .Q(instruction_address[23]) );
  DFC1 u_fetch_u_pc_program_counter_reg_24_ ( .D(n113), .C(clk), .RN(rst_n), 
        .Q(instruction_address[24]) );
  DFC1 u_fetch_u_pc_program_counter_reg_25_ ( .D(n112), .C(clk), .RN(rst_n), 
        .Q(instruction_address[25]) );
  DFC1 u_fetch_u_pc_program_counter_reg_26_ ( .D(n111), .C(clk), .RN(rst_n), 
        .Q(instruction_address[26]) );
  DFC1 u_fetch_u_pc_program_counter_reg_27_ ( .D(n110), .C(clk), .RN(rst_n), 
        .Q(instruction_address[27]) );
  DFC1 u_fetch_u_pc_program_counter_reg_28_ ( .D(n109), .C(clk), .RN(rst_n), 
        .Q(instruction_address[28]) );
  DFC1 u_fetch_u_pc_program_counter_reg_29_ ( .D(n108), .C(clk), .RN(rst_n), 
        .Q(instruction_address[29]) );
  DFC1 u_fetch_u_pc_program_counter_reg_30_ ( .D(n107), .C(clk), .RN(rst_n), 
        .Q(instruction_address[30]) );
  DFC1 u_fetch_u_pc_program_counter_reg_31_ ( .D(n138), .C(clk), .RN(rst_n), 
        .Q(instruction_address[31]) );
  DFC1 u_decode_pipe_addr_branch_reg_0_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[0]), .C(clk), .RN(rst_n), .Q(
        ex_data_pc4[0]) );
  DFC1 u_decode_pipe_addr_branch_reg_1_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[1]), .C(clk), .RN(rst_n), .Q(
        ex_data_pc4[1]) );
  DFC1 u_decode_pipe_addr_branch_reg_2_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[2]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[2]) );
  DFC1 u_decode_pipe_addr_branch_reg_3_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[3]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[3]) );
  DFC1 u_decode_pipe_addr_branch_reg_4_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[4]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[4]) );
  DFC1 u_decode_pipe_addr_branch_reg_5_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[5]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[5]) );
  DFC1 u_decode_pipe_addr_branch_reg_6_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[6]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[6]) );
  DFC1 u_decode_pipe_addr_branch_reg_7_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[7]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[7]) );
  DFC1 u_decode_pipe_addr_branch_reg_8_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[8]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[8]) );
  DFC1 u_decode_pipe_addr_branch_reg_9_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[9]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[9]) );
  DFC1 u_decode_pipe_addr_branch_reg_10_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[10]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[10]) );
  DFC1 u_decode_pipe_addr_branch_reg_11_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[11]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[11]) );
  DFC1 u_decode_pipe_addr_branch_reg_12_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[12]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[12]) );
  DFC1 u_decode_pipe_addr_branch_reg_13_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[13]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[13]) );
  DFC1 u_decode_pipe_addr_branch_reg_14_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[14]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[14]) );
  DFC1 u_decode_pipe_addr_branch_reg_15_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[15]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[15]) );
  DFC1 u_decode_pipe_addr_branch_reg_16_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[16]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[16]) );
  DFC1 u_decode_pipe_addr_branch_reg_17_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[17]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[17]) );
  DFC1 u_decode_pipe_addr_branch_reg_18_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[18]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[18]) );
  DFC1 u_decode_pipe_addr_branch_reg_19_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[19]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[19]) );
  DFC1 u_decode_pipe_addr_branch_reg_20_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[20]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[20]) );
  DFC1 u_decode_pipe_addr_branch_reg_21_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[21]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[21]) );
  DFC1 u_decode_pipe_addr_branch_reg_22_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[22]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[22]) );
  DFC1 u_decode_pipe_addr_branch_reg_23_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[23]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[23]) );
  DFC1 u_decode_pipe_addr_branch_reg_24_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[24]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[24]) );
  DFC1 u_decode_pipe_addr_branch_reg_25_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[25]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[25]) );
  DFC1 u_decode_pipe_addr_branch_reg_26_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[26]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[26]) );
  DFC1 u_decode_pipe_addr_branch_reg_27_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[27]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[27]) );
  DFC1 u_decode_pipe_addr_branch_reg_28_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[28]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[28]) );
  DFC1 u_decode_pipe_addr_branch_reg_29_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[29]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[29]) );
  DFC1 u_decode_pipe_addr_branch_reg_30_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[30]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[30]) );
  DFC1 u_decode_pipe_addr_branch_reg_31_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[31]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[31]) );
  DFC1 u_decode_pipe_FWmemout_reg_0_ ( .D(wb_data_memout[0]), .C(clk), .RN(
        rst_n), .Q(for_memout[0]) );
  DFC1 u_decode_pipe_FWmemout_reg_1_ ( .D(wb_data_memout[1]), .C(clk), .RN(
        rst_n), .Q(for_memout[1]) );
  DFC1 u_decode_pipe_FWmemout_reg_2_ ( .D(wb_data_memout[2]), .C(clk), .RN(
        rst_n), .Q(for_memout[2]) );
  DFC1 u_decode_pipe_FWmemout_reg_3_ ( .D(wb_data_memout[3]), .C(clk), .RN(
        rst_n), .Q(for_memout[3]) );
  DFC1 u_decode_pipe_FWmemout_reg_4_ ( .D(wb_data_memout[4]), .C(clk), .RN(
        rst_n), .Q(for_memout[4]) );
  DFC1 u_decode_pipe_FWmemout_reg_5_ ( .D(wb_data_memout[5]), .C(clk), .RN(
        rst_n), .Q(for_memout[5]) );
  DFC1 u_decode_pipe_FWmemout_reg_6_ ( .D(wb_data_memout[6]), .C(clk), .RN(
        rst_n), .Q(for_memout[6]) );
  DFC1 u_decode_pipe_FWmemout_reg_7_ ( .D(wb_data_memout[7]), .C(clk), .RN(
        rst_n), .Q(for_memout[7]) );
  DFC1 u_decode_pipe_FWmemout_reg_8_ ( .D(wb_data_memout[8]), .C(clk), .RN(
        rst_n), .Q(for_memout[8]) );
  DFC1 u_decode_pipe_FWmemout_reg_9_ ( .D(wb_data_memout[9]), .C(clk), .RN(
        rst_n), .Q(for_memout[9]) );
  DFC1 u_decode_pipe_FWmemout_reg_10_ ( .D(wb_data_memout[10]), .C(clk), .RN(
        rst_n), .Q(for_memout[10]) );
  DFC1 u_decode_pipe_FWmemout_reg_11_ ( .D(wb_data_memout[11]), .C(clk), .RN(
        rst_n), .Q(for_memout[11]) );
  DFC1 u_decode_pipe_FWmemout_reg_12_ ( .D(wb_data_memout[12]), .C(clk), .RN(
        rst_n), .Q(for_memout[12]) );
  DFC1 u_decode_pipe_FWmemout_reg_13_ ( .D(wb_data_memout[13]), .C(clk), .RN(
        rst_n), .Q(for_memout[13]) );
  DFC1 u_decode_pipe_FWmemout_reg_14_ ( .D(wb_data_memout[14]), .C(clk), .RN(
        rst_n), .Q(for_memout[14]) );
  DFC1 u_decode_pipe_FWmemout_reg_15_ ( .D(wb_data_memout[15]), .C(clk), .RN(
        rst_n), .Q(for_memout[15]) );
  DFC1 u_decode_pipe_FWmemout_reg_16_ ( .D(wb_data_memout[16]), .C(clk), .RN(
        rst_n), .Q(for_memout[16]) );
  DFC1 u_decode_pipe_FWmemout_reg_17_ ( .D(wb_data_memout[17]), .C(clk), .RN(
        rst_n), .Q(for_memout[17]) );
  DFC1 u_decode_pipe_FWmemout_reg_18_ ( .D(wb_data_memout[18]), .C(clk), .RN(
        rst_n), .Q(for_memout[18]) );
  DFC1 u_decode_pipe_FWmemout_reg_19_ ( .D(wb_data_memout[19]), .C(clk), .RN(
        rst_n), .Q(for_memout[19]) );
  DFC1 u_decode_pipe_FWmemout_reg_20_ ( .D(wb_data_memout[20]), .C(clk), .RN(
        rst_n), .Q(for_memout[20]) );
  DFC1 u_decode_pipe_FWmemout_reg_21_ ( .D(wb_data_memout[21]), .C(clk), .RN(
        rst_n), .Q(for_memout[21]) );
  DFC1 u_decode_pipe_FWmemout_reg_22_ ( .D(wb_data_memout[22]), .C(clk), .RN(
        rst_n), .Q(for_memout[22]) );
  DFC1 u_decode_pipe_FWmemout_reg_23_ ( .D(wb_data_memout[23]), .C(clk), .RN(
        rst_n), .Q(for_memout[23]) );
  DFC1 u_decode_pipe_FWmemout_reg_24_ ( .D(wb_data_memout[24]), .C(clk), .RN(
        rst_n), .Q(for_memout[24]) );
  DFC1 u_decode_pipe_FWmemout_reg_25_ ( .D(wb_data_memout[25]), .C(clk), .RN(
        rst_n), .Q(for_memout[25]) );
  DFC1 u_decode_pipe_FWmemout_reg_26_ ( .D(wb_data_memout[26]), .C(clk), .RN(
        rst_n), .Q(for_memout[26]) );
  DFC1 u_decode_pipe_FWmemout_reg_27_ ( .D(wb_data_memout[27]), .C(clk), .RN(
        rst_n), .Q(for_memout[27]) );
  DFC1 u_decode_pipe_FWmemout_reg_28_ ( .D(wb_data_memout[28]), .C(clk), .RN(
        rst_n), .Q(for_memout[28]) );
  DFC1 u_decode_pipe_FWmemout_reg_29_ ( .D(wb_data_memout[29]), .C(clk), .RN(
        rst_n), .Q(for_memout[29]) );
  DFC1 u_decode_pipe_FWmemout_reg_30_ ( .D(wb_data_memout[30]), .C(clk), .RN(
        rst_n), .Q(for_memout[30]) );
  DFC1 u_decode_pipe_FWmemout_reg_31_ ( .D(wb_data_memout[31]), .C(clk), .RN(
        rst_n), .Q(for_memout[31]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_0_ ( .D(if_addr_j[2]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[0]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_3_ ( .D(if_addr_j[5]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[3]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_4_ ( .D(if_addr_j[6]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[4]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_5_ ( .D(if_addr_j[7]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[5]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_6_ ( .D(if_addr_j[8]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[6]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_7_ ( .D(if_addr_j[9]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[7]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_8_ ( .D(if_addr_j[10]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[8]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_9_ ( .D(if_addr_j[11]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[9]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_11_ ( .D(if_addr_j[13]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[0]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_12_ ( .D(if_addr_j[14]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[1]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_13_ ( .D(if_addr_j[15]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[2]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_14_ ( .D(if_addr_j[16]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[3]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_15_ ( .D(if_addr_j[17]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[4]) );
  DFC1 u_decode_pipe_con_Wregwrite_reg ( .D(u_decode_control_o_con_regwrite), 
        .C(clk), .RN(rst_n), .Q(ex_con_Wregwrite) );
  DFC1 u_decode_pipe_con_Wmemtoreg_reg ( .D(u_decode_control_o_con_memtoreg), 
        .C(clk), .RN(rst_n), .Q(ex_con_Wmemtoreg) );
  DFC1 u_decode_pipe_con_Mmemwrite_reg ( .D(u_decode_control_o_con_memwrite), 
        .C(clk), .RN(rst_n), .Q(ex_con_Mmemwrite) );
  DFC1 u_decode_pipe_con_Mmemread_reg ( .D(u_decode_control_o_con_memread), 
        .C(clk), .RN(rst_n), .Q(ex_con_Mmemread) );
  DFC1 u_decode_pipe_con_MaluPC4_reg ( .D(u_decode_jbcon_o_con_aluPC4), .C(clk), .RN(rst_n), .Q(ex_con_Malupc8) );
  DFC1 u_decode_pipe_con_Eregdst_reg ( .D(u_decode_control_o_con_regdst), .C(
        clk), .RN(rst_n), .Q(ex_con_Eregdst) );
  DFC1 u_decode_pipe_con_Ealusrc_reg ( .D(u_decode_control_o_con_alusrc), .C(
        clk), .RN(rst_n), .Q(ex_con_Ealusrc) );
  DFC1 u_decode_pipe_con_Ealuop_reg_0_ ( .D(u_decode_control_o_con_aluop_0_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[0]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_1_ ( .D(u_decode_control_o_con_aluop_1_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[1]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_2_ ( .D(u_decode_control_o_con_aluop_2_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[2]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_3_ ( .D(u_decode_control_o_con_aluop_3_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[3]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_4_ ( .D(u_decode_control_o_con_aluop_4_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[4]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_5_ ( .D(u_decode_control_o_con_aluop_5_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[5]) );
  DFC1 u_decode_pipe_addr_pc4_reg_2_ ( .D(id_addr_pc4[2]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[2]) );
  DFC1 u_decode_pipe_addr_pc4_reg_3_ ( .D(id_addr_pc4[3]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[3]) );
  DFC1 u_decode_pipe_addr_pc4_reg_4_ ( .D(id_addr_pc4[4]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[4]) );
  DFC1 u_decode_pipe_addr_pc4_reg_5_ ( .D(id_addr_pc4[5]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[5]) );
  DFC1 u_decode_pipe_addr_pc4_reg_6_ ( .D(id_addr_pc4[6]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[6]) );
  DFC1 u_decode_pipe_addr_pc4_reg_7_ ( .D(id_addr_pc4[7]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[7]) );
  DFC1 u_decode_pipe_addr_pc4_reg_8_ ( .D(id_addr_pc4[8]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[8]) );
  DFC1 u_decode_pipe_addr_pc4_reg_9_ ( .D(id_addr_pc4[9]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[9]) );
  DFC1 u_decode_pipe_addr_pc4_reg_10_ ( .D(id_addr_pc4[10]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[10]) );
  DFC1 u_decode_pipe_addr_pc4_reg_11_ ( .D(id_addr_pc4[11]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[11]) );
  DFC1 u_decode_pipe_addr_pc4_reg_12_ ( .D(id_addr_pc4[12]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[12]) );
  DFC1 u_decode_pipe_addr_pc4_reg_13_ ( .D(id_addr_pc4[13]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[13]) );
  DFC1 u_decode_pipe_addr_pc4_reg_14_ ( .D(id_addr_pc4[14]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[14]) );
  DFC1 u_decode_pipe_addr_pc4_reg_15_ ( .D(id_addr_pc4[15]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[15]) );
  DFC1 u_decode_pipe_addr_pc4_reg_16_ ( .D(id_addr_pc4[16]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[16]) );
  DFC1 u_decode_pipe_addr_pc4_reg_17_ ( .D(id_addr_pc4[17]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[17]) );
  DFC1 u_decode_pipe_addr_pc4_reg_18_ ( .D(id_addr_pc4[18]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[18]) );
  DFC1 u_decode_pipe_addr_pc4_reg_19_ ( .D(id_addr_pc4[19]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[19]) );
  DFC1 u_decode_pipe_addr_pc4_reg_20_ ( .D(id_addr_pc4[20]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[20]) );
  DFC1 u_decode_pipe_addr_pc4_reg_21_ ( .D(id_addr_pc4[21]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[21]) );
  DFC1 u_decode_pipe_addr_pc4_reg_22_ ( .D(id_addr_pc4[22]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[22]) );
  DFC1 u_decode_pipe_addr_pc4_reg_23_ ( .D(id_addr_pc4[23]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[23]) );
  DFC1 u_decode_pipe_addr_pc4_reg_24_ ( .D(id_addr_pc4[24]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[24]) );
  DFC1 u_decode_pipe_addr_pc4_reg_25_ ( .D(id_addr_pc4[25]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[25]) );
  DFC1 u_decode_pipe_addr_pc4_reg_26_ ( .D(id_addr_pc4[26]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[26]) );
  DFC1 u_decode_pipe_addr_pc4_reg_27_ ( .D(id_addr_pc4[27]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[27]) );
  DFC1 u_decode_pipe_addr_pc4_reg_28_ ( .D(if_addr_j[28]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[28]) );
  DFC1 u_decode_pipe_addr_pc4_reg_29_ ( .D(if_addr_j[29]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[29]) );
  DFC1 u_decode_pipe_addr_pc4_reg_30_ ( .D(if_addr_j[30]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[30]) );
  DFC1 u_decode_pipe_addr_pc4_reg_31_ ( .D(if_addr_j[31]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[31]) );
  DFC1 u_decode_pipe_addr_rt_reg_0_ ( .D(if_addr_j[18]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[0]) );
  DFC1 u_decode_pipe_addr_rt_reg_1_ ( .D(if_addr_j[19]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[1]) );
  DFC1 u_decode_pipe_addr_rt_reg_2_ ( .D(if_addr_j[20]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[2]) );
  DFC1 u_decode_pipe_addr_rt_reg_3_ ( .D(if_addr_j[21]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[3]) );
  DFC1 u_decode_pipe_addr_rt_reg_4_ ( .D(if_addr_j[22]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[4]) );
  DFC1 u_decode_pipe_data_rt_reg_0_ ( .D(u_decode_regbank_o_data_Rt[0]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[0]) );
  DFC1 u_decode_pipe_data_rt_reg_1_ ( .D(u_decode_regbank_o_data_Rt[1]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[1]) );
  DFC1 u_decode_pipe_data_rt_reg_2_ ( .D(u_decode_regbank_o_data_Rt[2]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[2]) );
  DFC1 u_decode_pipe_data_rt_reg_3_ ( .D(u_decode_regbank_o_data_Rt[3]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[3]) );
  DFC1 u_decode_pipe_data_rt_reg_4_ ( .D(u_decode_regbank_o_data_Rt[4]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[4]) );
  DFC1 u_decode_pipe_data_rt_reg_5_ ( .D(u_decode_regbank_o_data_Rt[5]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[5]) );
  DFC1 u_decode_pipe_data_rt_reg_6_ ( .D(u_decode_regbank_o_data_Rt[6]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[6]) );
  DFC1 u_decode_pipe_data_rt_reg_7_ ( .D(u_decode_regbank_o_data_Rt[7]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[7]) );
  DFC1 u_decode_pipe_data_rt_reg_8_ ( .D(u_decode_regbank_o_data_Rt[8]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[8]) );
  DFC1 u_decode_pipe_data_rt_reg_9_ ( .D(u_decode_regbank_o_data_Rt[9]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[9]) );
  DFC1 u_decode_pipe_data_rt_reg_10_ ( .D(u_decode_regbank_o_data_Rt[10]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[10]) );
  DFC1 u_decode_pipe_data_rt_reg_11_ ( .D(u_decode_regbank_o_data_Rt[11]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[11]) );
  DFC1 u_decode_pipe_data_rt_reg_12_ ( .D(u_decode_regbank_o_data_Rt[12]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[12]) );
  DFC1 u_decode_pipe_data_rt_reg_13_ ( .D(u_decode_regbank_o_data_Rt[13]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[13]) );
  DFC1 u_decode_pipe_data_rt_reg_14_ ( .D(u_decode_regbank_o_data_Rt[14]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[14]) );
  DFC1 u_decode_pipe_data_rt_reg_15_ ( .D(u_decode_regbank_o_data_Rt[15]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[15]) );
  DFC1 u_decode_pipe_data_rt_reg_16_ ( .D(u_decode_regbank_o_data_Rt[16]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[16]) );
  DFC1 u_decode_pipe_data_rt_reg_17_ ( .D(u_decode_regbank_o_data_Rt[17]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[17]) );
  DFC1 u_decode_pipe_data_rt_reg_18_ ( .D(u_decode_regbank_o_data_Rt[18]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[18]) );
  DFC1 u_decode_pipe_data_rt_reg_19_ ( .D(u_decode_regbank_o_data_Rt[19]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[19]) );
  DFC1 u_decode_pipe_data_rt_reg_20_ ( .D(u_decode_regbank_o_data_Rt[20]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[20]) );
  DFC1 u_decode_pipe_data_rt_reg_21_ ( .D(u_decode_regbank_o_data_Rt[21]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[21]) );
  DFC1 u_decode_pipe_data_rt_reg_22_ ( .D(u_decode_regbank_o_data_Rt[22]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[22]) );
  DFC1 u_decode_pipe_data_rt_reg_23_ ( .D(u_decode_regbank_o_data_Rt[23]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[23]) );
  DFC1 u_decode_pipe_data_rt_reg_24_ ( .D(u_decode_regbank_o_data_Rt[24]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[24]) );
  DFC1 u_decode_pipe_data_rt_reg_25_ ( .D(u_decode_regbank_o_data_Rt[25]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[25]) );
  DFC1 u_decode_pipe_data_rt_reg_26_ ( .D(u_decode_regbank_o_data_Rt[26]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[26]) );
  DFC1 u_decode_pipe_data_rt_reg_27_ ( .D(u_decode_regbank_o_data_Rt[27]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[27]) );
  DFC1 u_decode_pipe_data_rt_reg_28_ ( .D(u_decode_regbank_o_data_Rt[28]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[28]) );
  DFC1 u_decode_pipe_data_rt_reg_29_ ( .D(u_decode_regbank_o_data_Rt[29]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[29]) );
  DFC1 u_decode_pipe_data_rt_reg_30_ ( .D(u_decode_regbank_o_data_Rt[30]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[30]) );
  DFC1 u_decode_pipe_data_rt_reg_31_ ( .D(u_decode_regbank_o_data_Rt[31]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[31]) );
  DFC1 u_decode_pipe_data_rs_reg_0_ ( .D(id_data_jr[0]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[0]) );
  DFC1 u_decode_pipe_data_rs_reg_1_ ( .D(id_data_jr[1]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[1]) );
  DFC1 u_decode_pipe_data_rs_reg_2_ ( .D(id_data_jr[2]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[2]) );
  DFC1 u_decode_pipe_data_rs_reg_3_ ( .D(id_data_jr[3]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[3]) );
  DFC1 u_decode_pipe_data_rs_reg_4_ ( .D(id_data_jr[4]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[4]) );
  DFC1 u_decode_pipe_data_rs_reg_5_ ( .D(id_data_jr[5]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[5]) );
  DFC1 u_decode_pipe_data_rs_reg_6_ ( .D(id_data_jr[6]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[6]) );
  DFC1 u_decode_pipe_data_rs_reg_7_ ( .D(id_data_jr[7]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[7]) );
  DFC1 u_decode_pipe_data_rs_reg_8_ ( .D(id_data_jr[8]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[8]) );
  DFC1 u_decode_pipe_data_rs_reg_9_ ( .D(id_data_jr[9]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[9]) );
  DFC1 u_decode_pipe_data_rs_reg_10_ ( .D(id_data_jr[10]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[10]) );
  DFC1 u_decode_pipe_data_rs_reg_11_ ( .D(id_data_jr[11]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[11]) );
  DFC1 u_decode_pipe_data_rs_reg_12_ ( .D(id_data_jr[12]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[12]) );
  DFC1 u_decode_pipe_data_rs_reg_13_ ( .D(id_data_jr[13]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[13]) );
  DFC1 u_decode_pipe_data_rs_reg_14_ ( .D(id_data_jr[14]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[14]) );
  DFC1 u_decode_pipe_data_rs_reg_15_ ( .D(id_data_jr[15]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[15]) );
  DFC1 u_decode_pipe_data_rs_reg_16_ ( .D(id_data_jr[16]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[16]) );
  DFC1 u_decode_pipe_data_rs_reg_17_ ( .D(id_data_jr[17]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[17]) );
  DFC1 u_decode_pipe_data_rs_reg_18_ ( .D(id_data_jr[18]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[18]) );
  DFC1 u_decode_pipe_data_rs_reg_19_ ( .D(id_data_jr[19]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[19]) );
  DFC1 u_decode_pipe_data_rs_reg_20_ ( .D(id_data_jr[20]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[20]) );
  DFC1 u_decode_pipe_data_rs_reg_21_ ( .D(id_data_jr[21]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[21]) );
  DFC1 u_decode_pipe_data_rs_reg_22_ ( .D(id_data_jr[22]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[22]) );
  DFC1 u_decode_pipe_data_rs_reg_23_ ( .D(id_data_jr[23]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[23]) );
  DFC1 u_decode_pipe_data_rs_reg_24_ ( .D(id_data_jr[24]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[24]) );
  DFC1 u_decode_pipe_data_rs_reg_25_ ( .D(id_data_jr[25]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[25]) );
  DFC1 u_decode_pipe_data_rs_reg_26_ ( .D(id_data_jr[26]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[26]) );
  DFC1 u_decode_pipe_data_rs_reg_27_ ( .D(id_data_jr[27]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[27]) );
  DFC1 u_decode_pipe_data_rs_reg_28_ ( .D(id_data_jr[28]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[28]) );
  DFC1 u_decode_pipe_data_rs_reg_29_ ( .D(id_data_jr[29]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[29]) );
  DFC1 u_decode_pipe_data_rs_reg_30_ ( .D(id_data_jr[30]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[30]) );
  DFC1 u_decode_pipe_data_rs_reg_31_ ( .D(id_data_jr[31]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[31]) );
  DFC1 u_decode_pipe_bop_reg_0_ ( .D(u_decode_jbcon_o_con_bop[0]), .C(clk), 
        .RN(rst_n), .Q(ex_con_bop[0]) );
  DFC1 u_decode_pipe_bop_reg_1_ ( .D(u_decode_jbcon_o_con_bop[1]), .C(clk), 
        .RN(rst_n), .Q(ex_con_bop[1]) );
  DFC1 u_decode_pipe_bop_reg_2_ ( .D(u_decode_n6), .C(clk), .RN(rst_n), .Q(
        ex_con_bop[2]) );
  D_register_bank u_decode_u_regbank ( .i_clk(clk), .i_rst_n(rst_n), 
        .i_addr_Rs(if_addr_j[27:23]), .i_con_RegWr(id_con_Wregwrite), 
        .i_addr_Rd(id_addr_Wregwrite), .i_data_Rd(id_data_Wregwrite), 
        .o_data_Rs(id_data_jr), .o_data_Rt(u_decode_regbank_o_data_Rt), 
        .i_addr_Rt_4_(if_addr_j[22]), .i_addr_Rt_3_(if_addr_j[21]), 
        .i_addr_Rt_2_(if_addr_j[20]), .i_addr_Rt_1_(if_addr_j[19]), 
        .i_addr_Rt_0_(if_addr_j[18]) );
  DFC3 u_fetch_pipe_instr_reg_16_ ( .D(read_instruction[16]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[18]), .QN(n216) );
  DFC3 u_fetch_pipe_instr_reg_17_ ( .D(read_instruction[17]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[19]), .QN(n206) );
  DFC3 u_fetch_pipe_instr_reg_18_ ( .D(read_instruction[18]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[20]), .QN(n214) );
  DFC3 u_fetch_pipe_instr_reg_19_ ( .D(read_instruction[19]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[21]), .QN(n220) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_16_ ( .D(u_decode_n1), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[31]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_1_ ( .D(if_addr_j[3]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[1]) );
  DFC3 u_decode_pipe_con_Efbmux_reg_0_ ( .D(u_decode_for_o_con_fb[0]), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[0]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_2_ ( .D(if_addr_j[4]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[2]) );
  DFC3 u_decode_pipe_con_Efbmux_reg_2_ ( .D(u_decode_for_o_con_fb[2]), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[2]) );
  DFC3 u_decode_pipe_con_Efamux_reg_2_ ( .D(u_decode_for_o_con_fa_2_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[2]) );
  DFC3 u_decode_pipe_con_Efamux_reg_1_ ( .D(u_decode_for_o_con_fa_1_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[1]) );
  DFC3 u_decode_pipe_con_Efbmux_reg_1_ ( .D(u_decode_for_o_con_fb[1]), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[1]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_10_ ( .D(if_addr_j[12]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[10]) );
  DFC3 u_mem_pipe_con_Wmemtoreg_reg ( .D(mem_con_Wmemtoreg), .C(clk), .RN(
        rst_n), .Q(wb_con_Wmemtoreg) );
  XNR21 add_x_4_U71 ( .A(n232), .B(add_x_4_n64), .Q(u_fetch_jmux_i_addr_pc4_7_) );
  XNR21 add_x_4_U15 ( .A(n229), .B(add_x_4_n20), .Q(
        u_fetch_jmux_i_addr_pc4_17_) );
  XNR21 add_x_4_U38 ( .A(n231), .B(add_x_4_n39), .Q(
        u_fetch_jmux_i_addr_pc4_13_) );
  XNR21 add_x_4_U27 ( .A(n230), .B(add_x_4_n29), .Q(
        u_fetch_jmux_i_addr_pc4_15_) );
  OAI210 u_decode_add_x_16_U125 ( .A(u_decode_add_x_16_n112), .B(
        u_decode_add_x_16_n106), .C(u_decode_add_x_16_n107), .Q(
        u_decode_add_x_16_n105) );
  OAI210 u_decode_add_x_16_U88 ( .A(u_decode_add_x_16_n87), .B(
        u_decode_add_x_16_n81), .C(u_decode_add_x_16_n82), .Q(
        u_decode_add_x_16_n80) );
  XNR21 u_decode_add_x_16_U11 ( .A(u_decode_add_x_16_n3), .B(
        u_decode_add_x_16_n39), .Q(u_decode_pcadd_o_addr_pcbranchE[27]) );
  XNR21 u_decode_add_x_16_U25 ( .A(u_decode_add_x_16_n5), .B(
        u_decode_add_x_16_n47), .Q(u_decode_pcadd_o_addr_pcbranchE[25]) );
  XNR21 u_decode_add_x_16_U39 ( .A(u_decode_add_x_16_n7), .B(
        u_decode_add_x_16_n55), .Q(u_decode_pcadd_o_addr_pcbranchE[23]) );
  XNR21 u_decode_add_x_16_U53 ( .A(u_decode_add_x_16_n9), .B(
        u_decode_add_x_16_n63), .Q(u_decode_pcadd_o_addr_pcbranchE[21]) );
  XNR21 add_x_1_U27 ( .A(add_x_1_n27), .B(add_x_1_n28), .Q(u_mem_pc8[14]) );
  XNR21 u_decode_add_x_16_U67 ( .A(u_decode_add_x_16_n11), .B(
        u_decode_add_x_16_n71), .Q(u_decode_pcadd_o_addr_pcbranchE[19]) );
  XNR21 u_decode_add_x_16_U93 ( .A(u_decode_add_x_16_n14), .B(
        u_decode_add_x_16_n88), .Q(u_decode_pcadd_o_addr_pcbranchE[16]) );
  XNR21 u_decode_add_x_16_U130 ( .A(u_decode_add_x_16_n18), .B(
        u_decode_add_x_16_n113), .Q(u_decode_pcadd_o_addr_pcbranchE[12]) );
  XNR21 u_decode_add_x_16_U138 ( .A(u_decode_add_x_16_n19), .B(
        u_decode_add_x_16_n120), .Q(u_decode_pcadd_o_addr_pcbranchE[11]) );
  XNR21 u_decode_add_x_16_U154 ( .A(u_decode_add_x_16_n21), .B(
        u_decode_add_x_16_n131), .Q(u_decode_pcadd_o_addr_pcbranchE[9]) );
  XNR21 u_decode_add_x_16_U179 ( .A(u_decode_add_x_16_n24), .B(
        u_decode_add_x_16_n144), .Q(u_decode_pcadd_o_addr_pcbranchE[6]) );
  XNR21 u_decode_add_x_16_U187 ( .A(u_decode_add_x_16_n25), .B(
        u_decode_add_x_16_n150), .Q(u_decode_pcadd_o_addr_pcbranchE[5]) );
  NAND22 add_x_4_U84 ( .A(instruction_address[4]), .B(instruction_address[5]), 
        .Q(add_x_4_n70) );
  NAND22 add_x_4_U53 ( .A(instruction_address[10]), .B(instruction_address[11]), .Q(add_x_4_n45) );
  XNR21 add_x_4_U87 ( .A(n223), .B(add_x_4_n76), .Q(u_fetch_jmux_i_addr_pc4_4_) );
  XNR21 add_x_4_U56 ( .A(n221), .B(add_x_4_n51), .Q(
        u_fetch_jmux_i_addr_pc4_10_) );
  XNR21 add_x_4_U91 ( .A(instruction_address[2]), .B(n236), .Q(
        u_fetch_jmux_i_addr_pc4_3_) );
  XOR21 add_x_4_U1 ( .A(instruction_address[31]), .B(add_x_4_n1), .Q(
        u_fetch_jmux_i_addr_pc4_31_) );
  XNR21 add_x_4_U67 ( .A(n222), .B(add_x_4_n60), .Q(u_fetch_jmux_i_addr_pc4_8_) );
  NAND22 add_x_4_U51 ( .A(add_x_4_n51), .B(add_x_4_n44), .Q(add_x_4_n43) );
  XNR21 add_x_4_U33 ( .A(n224), .B(add_x_4_n33), .Q(
        u_fetch_jmux_i_addr_pc4_14_) );
  NOR21 add_x_4_U63 ( .A(add_x_4_n54), .B(add_x_4_n61), .Q(add_x_4_n53) );
  NAND22 add_x_4_U42 ( .A(instruction_address[12]), .B(instruction_address[13]), .Q(add_x_4_n36) );
  NAND22 add_x_4_U19 ( .A(instruction_address[16]), .B(instruction_address[17]), .Q(add_x_4_n17) );
  NAND22 add_x_4_U30 ( .A(instruction_address[14]), .B(instruction_address[15]), .Q(add_x_4_n26) );
  NOR21 add_x_4_U18 ( .A(add_x_4_n17), .B(add_x_4_n26), .Q(add_x_4_n16) );
  NAND22 add_x_4_U17 ( .A(add_x_4_n35), .B(add_x_4_n16), .Q(add_x_4_n15) );
  NAND22 add_x_4_U28 ( .A(add_x_4_n33), .B(add_x_4_n25), .Q(add_x_4_n24) );
  NOR21 u_decode_add_x_16_U173 ( .A(u_decode_add_x_16_n137), .B(
        u_decode_add_x_16_n142), .Q(u_decode_add_x_16_n135) );
  NOR21 u_decode_add_x_16_U159 ( .A(u_decode_add_x_16_n129), .B(
        u_decode_add_x_16_n132), .Q(u_decode_add_x_16_n127) );
  NAND22 u_decode_add_x_16_U157 ( .A(u_decode_add_x_16_n135), .B(
        u_decode_add_x_16_n127), .Q(u_decode_add_x_16_n125) );
  OAI212 u_decode_add_x_16_U204 ( .A(u_decode_add_x_16_n158), .B(
        u_decode_add_x_16_n155), .C(u_decode_add_x_16_n156), .Q(
        u_decode_add_x_16_n154) );
  NOR21 u_decode_add_x_16_U190 ( .A(u_decode_add_x_16_n148), .B(
        u_decode_add_x_16_n151), .Q(u_decode_add_x_16_n146) );
  AOI211 u_decode_add_x_16_U158 ( .A(u_decode_add_x_16_n136), .B(
        u_decode_add_x_16_n127), .C(u_decode_add_x_16_n128), .Q(
        u_decode_add_x_16_n126) );
  OAI212 u_decode_add_x_16_U156 ( .A(u_decode_add_x_16_n125), .B(
        u_decode_add_x_16_n145), .C(u_decode_add_x_16_n126), .Q(
        u_decode_add_x_16_n124) );
  NOR21 u_decode_add_x_16_U142 ( .A(u_decode_add_x_16_n118), .B(
        u_decode_add_x_16_n121), .Q(u_decode_add_x_16_n116) );
  NOR21 u_decode_add_x_16_U124 ( .A(u_decode_add_x_16_n106), .B(
        u_decode_add_x_16_n111), .Q(u_decode_add_x_16_n104) );
  NAND22 u_decode_add_x_16_U122 ( .A(u_decode_add_x_16_n116), .B(
        u_decode_add_x_16_n104), .Q(u_decode_add_x_16_n102) );
  NOR21 u_decode_add_x_16_U91 ( .A(id_addr_pc4[17]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n81) );
  NOR21 u_decode_add_x_16_U87 ( .A(u_decode_add_x_16_n86), .B(
        u_decode_add_x_16_n81), .Q(u_decode_add_x_16_n79) );
  NOR21 u_decode_add_x_16_U105 ( .A(u_decode_add_x_16_n93), .B(
        u_decode_add_x_16_n98), .Q(u_decode_add_x_16_n91) );
  NAND22 u_decode_add_x_16_U85 ( .A(u_decode_add_x_16_n79), .B(
        u_decode_add_x_16_n91), .Q(u_decode_add_x_16_n77) );
  NOR21 u_decode_add_x_16_U83 ( .A(u_decode_add_x_16_n102), .B(
        u_decode_add_x_16_n77), .Q(u_decode_add_x_16_n75) );
  AOI211 u_decode_add_x_16_U123 ( .A(u_decode_add_x_16_n117), .B(
        u_decode_add_x_16_n104), .C(u_decode_add_x_16_n105), .Q(
        u_decode_add_x_16_n103) );
  OAI212 u_decode_add_x_16_U76 ( .A(u_decode_add_x_16_n72), .B(
        u_decode_add_x_16_n74), .C(u_decode_add_x_16_n73), .Q(
        u_decode_add_x_16_n71) );
  OAI212 u_decode_add_x_16_U62 ( .A(u_decode_add_x_16_n64), .B(
        u_decode_add_x_16_n66), .C(u_decode_add_x_16_n65), .Q(
        u_decode_add_x_16_n63) );
  OAI212 u_decode_add_x_16_U48 ( .A(u_decode_add_x_16_n56), .B(
        u_decode_add_x_16_n58), .C(u_decode_add_x_16_n57), .Q(
        u_decode_add_x_16_n55) );
  OAI212 u_decode_add_x_16_U34 ( .A(u_decode_add_x_16_n48), .B(
        u_decode_add_x_16_n50), .C(u_decode_add_x_16_n49), .Q(
        u_decode_add_x_16_n47) );
  OAI212 u_decode_add_x_16_U20 ( .A(u_decode_add_x_16_n40), .B(
        u_decode_add_x_16_n42), .C(u_decode_add_x_16_n41), .Q(
        u_decode_add_x_16_n39) );
  OAI212 u_decode_add_x_16_U6 ( .A(u_decode_add_x_16_n32), .B(
        u_decode_add_x_16_n34), .C(u_decode_add_x_16_n33), .Q(
        u_decode_add_x_16_n31) );
  NAND22 add_x_1_U58 ( .A(mem_data_pc4[8]), .B(mem_data_pc4[9]), .Q(
        add_x_1_n49) );
  NAND22 add_x_1_U67 ( .A(mem_data_pc4[6]), .B(mem_data_pc4[7]), .Q(
        add_x_1_n56) );
  NOR21 add_x_1_U57 ( .A(add_x_1_n49), .B(add_x_1_n56), .Q(add_x_1_n48) );
  NAND22 add_x_1_U78 ( .A(mem_data_pc4[4]), .B(mem_data_pc4[5]), .Q(
        add_x_1_n65) );
  NAND22 add_x_1_U36 ( .A(mem_data_pc4[12]), .B(mem_data_pc4[13]), .Q(
        add_x_1_n31) );
  NAND22 add_x_1_U47 ( .A(mem_data_pc4[10]), .B(mem_data_pc4[11]), .Q(
        add_x_1_n40) );
  NAND22 add_x_1_U24 ( .A(mem_data_pc4[14]), .B(mem_data_pc4[15]), .Q(
        add_x_1_n21) );
  NOR21 add_x_1_U19 ( .A(mem_data_pc4[16]), .B(add_x_1_n21), .Q(add_x_1_n17)
         );
  NAND22 add_x_1_U18 ( .A(add_x_1_n30), .B(add_x_1_n17), .Q(add_x_1_n16) );
  ADD22 add_x_1_U3 ( .A(add_x_1_n3), .B(mem_data_pc4[29]), .CO(add_x_1_n2), 
        .S(u_mem_pc8[29]) );
  ADD22 add_x_1_U2 ( .A(add_x_1_n2), .B(mem_data_pc4[30]), .CO(add_x_1_n1), 
        .S(u_mem_pc8[30]) );
  OAI212 u_decode_add_x_16_U102 ( .A(u_decode_add_x_16_n89), .B(
        u_decode_add_x_16_n100), .C(u_decode_add_x_16_n90), .Q(
        u_decode_add_x_16_n88) );
  XOR21 u_decode_add_x_16_U111 ( .A(u_decode_add_x_16_n16), .B(
        u_decode_add_x_16_n100), .Q(u_decode_pcadd_o_addr_pcbranchE[14]) );
  NAND22 add_x_1_U45 ( .A(add_x_1_n46), .B(add_x_1_n39), .Q(add_x_1_n38) );
  XOR21 add_x_1_U39 ( .A(add_x_1_n37), .B(add_x_1_n38), .Q(u_mem_pc8[12]) );
  AOI211 u_decode_add_x_16_U86 ( .A(u_decode_add_x_16_n79), .B(
        u_decode_add_x_16_n92), .C(u_decode_add_x_16_n80), .Q(
        u_decode_add_x_16_n78) );
  AOI211 u_decode_add_x_16_U189 ( .A(u_decode_add_x_16_n154), .B(
        u_decode_add_x_16_n146), .C(u_decode_add_x_16_n147), .Q(
        u_decode_add_x_16_n145) );
  NOR21 add_x_4_U41 ( .A(add_x_4_n36), .B(add_x_4_n45), .Q(add_x_4_n35) );
  NOR21 add_x_1_U35 ( .A(add_x_1_n31), .B(add_x_1_n40), .Q(add_x_1_n30) );
  NAND22 u_decode_add_x_16_U15 ( .A(u_decode_add_x_16_n35), .B(
        u_decode_add_x_16_n38), .Q(u_decode_add_x_16_n3) );
  XOR21 add_x_1_U70 ( .A(add_x_1_n62), .B(add_x_1_n63), .Q(u_mem_pc8[6]) );
  NAND22 u_decode_add_x_16_U97 ( .A(u_decode_add_x_16_n84), .B(
        u_decode_add_x_16_n87), .Q(u_decode_add_x_16_n14) );
  ADD22 add_x_4_U5 ( .A(add_x_4_n5), .B(instruction_address[27]), .CO(
        add_x_4_n4), .S(u_fetch_jmux_i_addr_pc4_27_) );
  ADD22 add_x_4_U3 ( .A(add_x_4_n3), .B(instruction_address[29]), .CO(
        add_x_4_n2), .S(u_fetch_jmux_i_addr_pc4_29_) );
  ADD22 add_x_4_U2 ( .A(add_x_4_n2), .B(instruction_address[30]), .CO(
        add_x_4_n1), .S(u_fetch_jmux_i_addr_pc4_30_) );
  NAND22 add_x_4_U64 ( .A(instruction_address[8]), .B(instruction_address[9]), 
        .Q(add_x_4_n54) );
  NAND22 add_x_4_U73 ( .A(instruction_address[6]), .B(instruction_address[7]), 
        .Q(add_x_4_n61) );
  NOR21 u_decode_add_x_16_U79 ( .A(id_addr_pc4[18]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n72) );
  NOR21 u_decode_add_x_16_U163 ( .A(id_addr_pc4[9]), .B(if_addr_j[9]), .Q(
        u_decode_add_x_16_n129) );
  NOR21 u_decode_add_x_16_U194 ( .A(id_addr_pc4[5]), .B(if_addr_j[5]), .Q(
        u_decode_add_x_16_n148) );
  NOR21 u_decode_add_x_16_U146 ( .A(id_addr_pc4[11]), .B(if_addr_j[11]), .Q(
        u_decode_add_x_16_n118) );
  NOR21 u_decode_add_x_16_U128 ( .A(id_addr_pc4[13]), .B(if_addr_j[13]), .Q(
        u_decode_add_x_16_n106) );
  NOR21 u_decode_add_x_16_U109 ( .A(id_addr_pc4[15]), .B(if_addr_j[15]), .Q(
        u_decode_add_x_16_n93) );
  OAI212 u_decode_add_x_16_U121 ( .A(u_decode_add_x_16_n102), .B(
        u_decode_add_x_16_n123), .C(u_decode_add_x_16_n103), .Q(
        u_decode_add_x_16_n101) );
  OAI212 u_decode_add_x_16_U139 ( .A(u_decode_add_x_16_n114), .B(
        u_decode_add_x_16_n123), .C(u_decode_add_x_16_n115), .Q(
        u_decode_add_x_16_n113) );
  AOI211 u_decode_add_x_16_U172 ( .A(u_decode_add_x_16_n144), .B(
        u_decode_add_x_16_n135), .C(u_decode_add_x_16_n136), .Q(
        u_decode_add_x_16_n134) );
  DFC3 u_decode_pipe_con_Efamux_reg_0_ ( .D(u_decode_for_o_con_fa_0_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[0]) );
  DFC3 u_fetch_pipe_instr_reg_20_ ( .D(read_instruction[20]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[22]), .QN(n215) );
  DFC3 u_mem_pipe_addr_regdst_reg_3_ ( .D(mem_addr_regdst[3]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[3]) );
  NAND22 u_decode_add_x_16_U213 ( .A(if_addr_j[2]), .B(id_addr_pc4[2]), .Q(
        u_decode_add_x_16_n158) );
  NAND22 u_decode_add_x_16_U208 ( .A(if_addr_j[3]), .B(id_addr_pc4[3]), .Q(
        u_decode_add_x_16_n156) );
  NOR21 u_decode_add_x_16_U207 ( .A(id_addr_pc4[3]), .B(if_addr_j[3]), .Q(
        u_decode_add_x_16_n155) );
  NAND22 u_decode_add_x_16_U201 ( .A(if_addr_j[4]), .B(id_addr_pc4[4]), .Q(
        u_decode_add_x_16_n152) );
  NOR21 u_decode_add_x_16_U200 ( .A(id_addr_pc4[4]), .B(if_addr_j[4]), .Q(
        u_decode_add_x_16_n151) );
  NAND21 u_decode_add_x_16_U195 ( .A(if_addr_j[5]), .B(id_addr_pc4[5]), .Q(
        u_decode_add_x_16_n149) );
  NAND22 u_decode_add_x_16_U186 ( .A(if_addr_j[6]), .B(id_addr_pc4[6]), .Q(
        u_decode_add_x_16_n143) );
  NOR21 u_decode_add_x_16_U185 ( .A(id_addr_pc4[6]), .B(if_addr_j[6]), .Q(
        u_decode_add_x_16_n142) );
  NAND21 u_decode_add_x_16_U178 ( .A(if_addr_j[7]), .B(id_addr_pc4[7]), .Q(
        u_decode_add_x_16_n138) );
  NOR21 u_decode_add_x_16_U177 ( .A(id_addr_pc4[7]), .B(if_addr_j[7]), .Q(
        u_decode_add_x_16_n137) );
  NOR21 u_decode_add_x_16_U169 ( .A(id_addr_pc4[8]), .B(if_addr_j[8]), .Q(
        u_decode_add_x_16_n132) );
  NAND21 u_decode_add_x_16_U164 ( .A(if_addr_j[9]), .B(id_addr_pc4[9]), .Q(
        u_decode_add_x_16_n130) );
  NAND22 u_decode_add_x_16_U153 ( .A(if_addr_j[10]), .B(id_addr_pc4[10]), .Q(
        u_decode_add_x_16_n122) );
  NOR21 u_decode_add_x_16_U152 ( .A(id_addr_pc4[10]), .B(if_addr_j[10]), .Q(
        u_decode_add_x_16_n121) );
  NAND21 u_decode_add_x_16_U147 ( .A(if_addr_j[11]), .B(id_addr_pc4[11]), .Q(
        u_decode_add_x_16_n119) );
  NAND22 u_decode_add_x_16_U137 ( .A(if_addr_j[12]), .B(id_addr_pc4[12]), .Q(
        u_decode_add_x_16_n112) );
  NOR21 u_decode_add_x_16_U136 ( .A(id_addr_pc4[12]), .B(if_addr_j[12]), .Q(
        u_decode_add_x_16_n111) );
  NAND21 u_decode_add_x_16_U129 ( .A(if_addr_j[13]), .B(id_addr_pc4[13]), .Q(
        u_decode_add_x_16_n107) );
  NAND22 u_decode_add_x_16_U118 ( .A(if_addr_j[14]), .B(id_addr_pc4[14]), .Q(
        u_decode_add_x_16_n99) );
  NOR21 u_decode_add_x_16_U117 ( .A(id_addr_pc4[14]), .B(if_addr_j[14]), .Q(
        u_decode_add_x_16_n98) );
  NAND21 u_decode_add_x_16_U110 ( .A(if_addr_j[15]), .B(id_addr_pc4[15]), .Q(
        u_decode_add_x_16_n94) );
  NAND22 u_decode_add_x_16_U100 ( .A(if_addr_j[16]), .B(id_addr_pc4[16]), .Q(
        u_decode_add_x_16_n87) );
  NOR21 u_decode_add_x_16_U99 ( .A(id_addr_pc4[16]), .B(if_addr_j[16]), .Q(
        u_decode_add_x_16_n86) );
  NAND22 u_decode_add_x_16_U170 ( .A(if_addr_j[8]), .B(id_addr_pc4[8]), .Q(
        u_decode_add_x_16_n133) );
  NOR21 u_decode_add_x_16_U59 ( .A(id_addr_pc4[21]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n61) );
  NAND22 u_decode_add_x_16_U60 ( .A(if_addr_j[17]), .B(id_addr_pc4[21]), .Q(
        u_decode_add_x_16_n62) );
  NOR21 u_decode_add_x_16_U65 ( .A(id_addr_pc4[20]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n64) );
  OAI211 u_decode_add_x_16_U191 ( .A(u_decode_add_x_16_n152), .B(
        u_decode_add_x_16_n148), .C(u_decode_add_x_16_n149), .Q(
        u_decode_add_x_16_n147) );
  NAND22 u_decode_add_x_16_U66 ( .A(if_addr_j[17]), .B(id_addr_pc4[20]), .Q(
        u_decode_add_x_16_n65) );
  NAND21 u_decode_add_x_16_U92 ( .A(if_addr_j[17]), .B(id_addr_pc4[17]), .Q(
        u_decode_add_x_16_n82) );
  NOR21 u_decode_add_x_16_U73 ( .A(id_addr_pc4[19]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n69) );
  NAND22 u_decode_add_x_16_U74 ( .A(if_addr_j[17]), .B(id_addr_pc4[19]), .Q(
        u_decode_add_x_16_n70) );
  OAI211 u_decode_add_x_16_U174 ( .A(u_decode_add_x_16_n143), .B(
        u_decode_add_x_16_n137), .C(u_decode_add_x_16_n138), .Q(
        u_decode_add_x_16_n136) );
  NAND22 u_decode_add_x_16_U18 ( .A(if_addr_j[17]), .B(id_addr_pc4[27]), .Q(
        u_decode_add_x_16_n38) );
  NOR21 u_decode_add_x_16_U23 ( .A(id_addr_pc4[26]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n40) );
  NOR21 u_decode_add_x_16_U17 ( .A(id_addr_pc4[27]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n37) );
  NOR21 u_decode_add_x_16_U45 ( .A(id_addr_pc4[23]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n53) );
  NAND22 u_decode_add_x_16_U24 ( .A(if_addr_j[17]), .B(id_addr_pc4[26]), .Q(
        u_decode_add_x_16_n41) );
  NAND22 u_decode_add_x_16_U46 ( .A(if_addr_j[17]), .B(id_addr_pc4[23]), .Q(
        u_decode_add_x_16_n54) );
  NAND22 u_decode_add_x_16_U10 ( .A(if_addr_j[17]), .B(if_addr_j[28]), .Q(
        u_decode_add_x_16_n33) );
  NOR21 u_decode_add_x_16_U9 ( .A(if_addr_j[28]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n32) );
  NAND22 u_decode_add_x_16_U52 ( .A(if_addr_j[17]), .B(id_addr_pc4[22]), .Q(
        u_decode_add_x_16_n57) );
  NOR21 u_decode_add_x_16_U31 ( .A(id_addr_pc4[25]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n45) );
  NOR21 u_decode_add_x_16_U51 ( .A(id_addr_pc4[22]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n56) );
  NAND22 u_decode_add_x_16_U32 ( .A(if_addr_j[17]), .B(id_addr_pc4[25]), .Q(
        u_decode_add_x_16_n46) );
  NAND22 u_decode_add_x_16_U38 ( .A(if_addr_j[17]), .B(id_addr_pc4[24]), .Q(
        u_decode_add_x_16_n49) );
  OAI211 u_decode_add_x_16_U143 ( .A(u_decode_add_x_16_n122), .B(
        u_decode_add_x_16_n118), .C(u_decode_add_x_16_n119), .Q(
        u_decode_add_x_16_n117) );
  OAI211 u_decode_add_x_16_U106 ( .A(u_decode_add_x_16_n99), .B(
        u_decode_add_x_16_n93), .C(u_decode_add_x_16_n94), .Q(
        u_decode_add_x_16_n92) );
  NOR21 u_decode_add_x_16_U37 ( .A(id_addr_pc4[24]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n48) );
  NAND22 u_decode_add_x_16_U161 ( .A(u_decode_add_x_16_n178), .B(
        u_decode_add_x_16_n130), .Q(u_decode_add_x_16_n21) );
  NAND22 u_decode_add_x_16_U183 ( .A(u_decode_add_x_16_n181), .B(
        u_decode_add_x_16_n143), .Q(u_decode_add_x_16_n24) );
  NAND22 u_decode_add_x_16_U192 ( .A(u_decode_add_x_16_n182), .B(
        u_decode_add_x_16_n149), .Q(u_decode_add_x_16_n25) );
  NAND22 u_decode_add_x_16_U115 ( .A(u_decode_add_x_16_n96), .B(
        u_decode_add_x_16_n99), .Q(u_decode_add_x_16_n16) );
  NAND22 u_decode_add_x_16_U134 ( .A(u_decode_add_x_16_n175), .B(
        u_decode_add_x_16_n112), .Q(u_decode_add_x_16_n18) );
  NAND22 u_decode_add_x_16_U144 ( .A(u_decode_add_x_16_n176), .B(
        u_decode_add_x_16_n119), .Q(u_decode_add_x_16_n19) );
  XOR21 add_x_4_U81 ( .A(n235), .B(add_x_4_n73), .Q(u_fetch_jmux_i_addr_pc4_5_) );
  XOR21 add_x_4_U76 ( .A(n227), .B(add_x_4_n68), .Q(u_fetch_jmux_i_addr_pc4_6_) );
  NOR21 add_x_4_U77 ( .A(n227), .B(add_x_4_n68), .Q(add_x_4_n64) );
  NOR21 add_x_4_U72 ( .A(add_x_4_n61), .B(add_x_4_n68), .Q(add_x_4_n60) );
  NAND22 u_decode_add_x_16_U71 ( .A(u_decode_add_x_16_n67), .B(
        u_decode_add_x_16_n70), .Q(u_decode_add_x_16_n11) );
  OAI211 u_decode_add_x_16_U197 ( .A(u_decode_add_x_16_n151), .B(
        u_decode_add_x_16_n153), .C(u_decode_add_x_16_n152), .Q(
        u_decode_add_x_16_n150) );
  NAND22 u_decode_add_x_16_U57 ( .A(u_decode_add_x_16_n59), .B(
        u_decode_add_x_16_n62), .Q(u_decode_add_x_16_n9) );
  NOR21 add_x_1_U66 ( .A(add_x_1_n56), .B(add_x_1_n63), .Q(add_x_1_n55) );
  NOR21 add_x_1_U17 ( .A(add_x_1_n47), .B(add_x_1_n16), .Q(add_x_1_n15) );
  NAND22 add_x_4_U68 ( .A(add_x_4_n60), .B(instruction_address[8]), .Q(
        add_x_4_n57) );
  NAND22 add_x_4_U57 ( .A(add_x_4_n51), .B(instruction_address[10]), .Q(
        add_x_4_n48) );
  NAND22 add_x_4_U40 ( .A(add_x_4_n51), .B(add_x_4_n35), .Q(add_x_4_n34) );
  ADD22 add_x_4_U14 ( .A(add_x_4_n14), .B(instruction_address[18]), .CO(
        add_x_4_n13), .S(u_fetch_jmux_i_addr_pc4_18_) );
  ADD22 add_x_1_U15 ( .A(add_x_1_n15), .B(mem_data_pc4[17]), .CO(add_x_1_n14), 
        .S(u_mem_pc8[17]) );
  OAI211 u_decode_add_x_16_U84 ( .A(u_decode_add_x_16_n103), .B(
        u_decode_add_x_16_n77), .C(u_decode_add_x_16_n78), .Q(
        u_decode_add_x_16_n76) );
  AOI211 u_decode_add_x_16_U82 ( .A(u_decode_add_x_16_n124), .B(
        u_decode_add_x_16_n75), .C(u_decode_add_x_16_n76), .Q(
        u_decode_add_x_16_n74) );
  OAI211 u_decode_add_x_16_U149 ( .A(u_decode_add_x_16_n121), .B(
        u_decode_add_x_16_n123), .C(u_decode_add_x_16_n122), .Q(
        u_decode_add_x_16_n120) );
  OAI211 u_decode_add_x_16_U166 ( .A(u_decode_add_x_16_n132), .B(
        u_decode_add_x_16_n134), .C(u_decode_add_x_16_n133), .Q(
        u_decode_add_x_16_n131) );
  NOR21 add_x_4_U34 ( .A(n224), .B(add_x_4_n34), .Q(add_x_4_n29) );
  XOR21 add_x_4_U60 ( .A(n234), .B(add_x_4_n57), .Q(u_fetch_jmux_i_addr_pc4_9_) );
  XOR21 add_x_4_U50 ( .A(n233), .B(add_x_4_n48), .Q(
        u_fetch_jmux_i_addr_pc4_11_) );
  ADD22 add_x_4_U13 ( .A(add_x_4_n13), .B(instruction_address[19]), .CO(
        add_x_4_n12), .S(u_fetch_jmux_i_addr_pc4_19_) );
  NOR21 add_x_4_U46 ( .A(n226), .B(add_x_4_n43), .Q(add_x_4_n39) );
  XOR21 add_x_4_U45 ( .A(n226), .B(add_x_4_n43), .Q(
        u_fetch_jmux_i_addr_pc4_12_) );
  ADD22 add_x_1_U14 ( .A(add_x_1_n14), .B(mem_data_pc4[18]), .CO(add_x_1_n13), 
        .S(u_mem_pc8[18]) );
  ADD22 add_x_4_U12 ( .A(add_x_4_n12), .B(instruction_address[20]), .CO(
        add_x_4_n11), .S(u_fetch_jmux_i_addr_pc4_20_) );
  ADD22 add_x_1_U13 ( .A(add_x_1_n13), .B(mem_data_pc4[19]), .CO(add_x_1_n12), 
        .S(u_mem_pc8[19]) );
  AOI211 u_decode_add_x_16_U68 ( .A(u_decode_add_x_16_n71), .B(
        u_decode_add_x_16_n67), .C(u_decode_add_x_16_n68), .Q(
        u_decode_add_x_16_n66) );
  XOR21 add_x_4_U22 ( .A(n225), .B(add_x_4_n24), .Q(
        u_fetch_jmux_i_addr_pc4_16_) );
  NOR21 add_x_4_U23 ( .A(n225), .B(add_x_4_n24), .Q(add_x_4_n20) );
  ADD22 add_x_4_U11 ( .A(add_x_4_n11), .B(instruction_address[21]), .CO(
        add_x_4_n10), .S(u_fetch_jmux_i_addr_pc4_21_) );
  ADD22 add_x_1_U12 ( .A(add_x_1_n12), .B(mem_data_pc4[20]), .CO(add_x_1_n11), 
        .S(u_mem_pc8[20]) );
  ADD22 add_x_1_U11 ( .A(add_x_1_n11), .B(mem_data_pc4[21]), .CO(add_x_1_n10), 
        .S(u_mem_pc8[21]) );
  ADD22 add_x_4_U10 ( .A(add_x_4_n10), .B(instruction_address[22]), .CO(
        add_x_4_n9), .S(u_fetch_jmux_i_addr_pc4_22_) );
  ADD22 add_x_4_U9 ( .A(add_x_4_n9), .B(instruction_address[23]), .CO(
        add_x_4_n8), .S(u_fetch_jmux_i_addr_pc4_23_) );
  ADD22 add_x_1_U10 ( .A(add_x_1_n10), .B(mem_data_pc4[22]), .CO(add_x_1_n9), 
        .S(u_mem_pc8[22]) );
  AOI211 u_decode_add_x_16_U54 ( .A(u_decode_add_x_16_n63), .B(
        u_decode_add_x_16_n59), .C(u_decode_add_x_16_n60), .Q(
        u_decode_add_x_16_n58) );
  ADD22 add_x_1_U9 ( .A(add_x_1_n9), .B(mem_data_pc4[23]), .CO(add_x_1_n8), 
        .S(u_mem_pc8[23]) );
  ADD22 add_x_4_U8 ( .A(add_x_4_n8), .B(instruction_address[24]), .CO(
        add_x_4_n7), .S(u_fetch_jmux_i_addr_pc4_24_) );
  ADD22 add_x_4_U7 ( .A(add_x_4_n7), .B(instruction_address[25]), .CO(
        add_x_4_n6), .S(u_fetch_jmux_i_addr_pc4_25_) );
  ADD22 add_x_1_U8 ( .A(add_x_1_n8), .B(mem_data_pc4[24]), .CO(add_x_1_n7), 
        .S(u_mem_pc8[24]) );
  AOI211 u_decode_add_x_16_U40 ( .A(u_decode_add_x_16_n55), .B(
        u_decode_add_x_16_n51), .C(u_decode_add_x_16_n52), .Q(
        u_decode_add_x_16_n50) );
  ADD22 add_x_4_U6 ( .A(add_x_4_n6), .B(instruction_address[26]), .CO(
        add_x_4_n5), .S(u_fetch_jmux_i_addr_pc4_26_) );
  ADD22 add_x_1_U7 ( .A(add_x_1_n7), .B(mem_data_pc4[25]), .CO(add_x_1_n6), 
        .S(u_mem_pc8[25]) );
  ADD22 add_x_1_U6 ( .A(add_x_1_n6), .B(mem_data_pc4[26]), .CO(add_x_1_n5), 
        .S(u_mem_pc8[26]) );
  AOI211 u_decode_add_x_16_U26 ( .A(u_decode_add_x_16_n47), .B(
        u_decode_add_x_16_n43), .C(u_decode_add_x_16_n44), .Q(
        u_decode_add_x_16_n42) );
  ADD22 add_x_4_U4 ( .A(add_x_4_n4), .B(instruction_address[28]), .CO(
        add_x_4_n3), .S(u_fetch_jmux_i_addr_pc4_28_) );
  AOI211 u_decode_add_x_16_U12 ( .A(u_decode_add_x_16_n39), .B(
        u_decode_add_x_16_n35), .C(u_decode_add_x_16_n36), .Q(
        u_decode_add_x_16_n34) );
  ADD32 u_decode_add_x_16_U4 ( .A(if_addr_j[17]), .B(if_addr_j[29]), .CI(
        u_decode_add_x_16_n31), .CO(u_decode_add_x_16_n30), .S(
        u_decode_pcadd_o_addr_pcbranchE[29]) );
  ADD32 u_decode_add_x_16_U3 ( .A(if_addr_j[17]), .B(if_addr_j[30]), .CI(
        u_decode_add_x_16_n30), .CO(u_decode_add_x_16_n29), .S(
        u_decode_pcadd_o_addr_pcbranchE[30]) );
  NAND22 u_decode_add_x_16_U80 ( .A(if_addr_j[17]), .B(id_addr_pc4[18]), .Q(
        u_decode_add_x_16_n73) );
  NAND22 add_x_1_U34 ( .A(add_x_1_n46), .B(add_x_1_n30), .Q(add_x_1_n29) );
  OAI211 u_decode_add_x_16_U160 ( .A(u_decode_add_x_16_n133), .B(
        u_decode_add_x_16_n129), .C(u_decode_add_x_16_n130), .Q(
        u_decode_add_x_16_n128) );
  NAND21 add_x_4_U88 ( .A(add_x_4_n76), .B(instruction_address[4]), .Q(
        add_x_4_n73) );
  NAND21 u_decode_add_x_16_U43 ( .A(u_decode_add_x_16_n51), .B(
        u_decode_add_x_16_n54), .Q(u_decode_add_x_16_n7) );
  NAND21 u_decode_add_x_16_U29 ( .A(u_decode_add_x_16_n43), .B(
        u_decode_add_x_16_n46), .Q(u_decode_add_x_16_n5) );
  DFC3 u_fetch_pipe_instr_reg_15_ ( .D(read_instruction[15]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[17]), .QN(n207) );
  INV3 U204 ( .A(n264), .Q(n343) );
  CLKIN0 U205 ( .A(data_address[15]), .Q(n140) );
  NOR20 U206 ( .A(add_x_1_n29), .B(add_x_1_n27), .Q(n141) );
  XNR20 U207 ( .A(mem_data_pc4[15]), .B(n141), .Q(n142) );
  IMUX20 U208 ( .A(n140), .B(n142), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[15]) );
  CLKIN0 U209 ( .A(u_decode_add_x_16_n99), .Q(n143) );
  AOI210 U210 ( .A(u_decode_add_x_16_n101), .B(u_decode_add_x_16_n96), .C(n143), .Q(n144) );
  CLKIN0 U211 ( .A(u_decode_add_x_16_n94), .Q(n145) );
  NOR20 U212 ( .A(u_decode_add_x_16_n93), .B(n145), .Q(n146) );
  XNR20 U213 ( .A(n144), .B(n146), .Q(u_decode_pcadd_o_addr_pcbranchE[15]) );
  CLKIN0 U214 ( .A(data_address[13]), .Q(n147) );
  NOR20 U215 ( .A(add_x_1_n38), .B(add_x_1_n37), .Q(n148) );
  XNR20 U216 ( .A(mem_data_pc4[13]), .B(n148), .Q(n149) );
  IMUX20 U217 ( .A(n147), .B(n149), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[13]) );
  NAND20 U218 ( .A(add_x_1_n55), .B(mem_data_pc4[8]), .Q(n150) );
  XNR20 U219 ( .A(mem_data_pc4[9]), .B(n150), .Q(n151) );
  MUX21 U220 ( .A(data_address[9]), .B(n151), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[9]) );
  CLKIN0 U221 ( .A(u_decode_add_x_16_n73), .Q(n152) );
  NOR20 U222 ( .A(u_decode_add_x_16_n72), .B(n152), .Q(n153) );
  XNR20 U223 ( .A(u_decode_add_x_16_n74), .B(n153), .Q(
        u_decode_pcadd_o_addr_pcbranchE[18]) );
  CLKIN0 U224 ( .A(u_decode_add_x_16_n112), .Q(n154) );
  AOI210 U225 ( .A(u_decode_add_x_16_n113), .B(u_decode_add_x_16_n175), .C(
        n154), .Q(n155) );
  CLKIN0 U226 ( .A(u_decode_add_x_16_n107), .Q(n156) );
  NOR20 U227 ( .A(u_decode_add_x_16_n106), .B(n156), .Q(n157) );
  XNR20 U228 ( .A(n155), .B(n157), .Q(u_decode_pcadd_o_addr_pcbranchE[13]) );
  CLKIN0 U229 ( .A(u_decode_add_x_16_n133), .Q(n158) );
  NOR20 U230 ( .A(u_decode_add_x_16_n132), .B(n158), .Q(n159) );
  XNR20 U231 ( .A(u_decode_add_x_16_n134), .B(n159), .Q(
        u_decode_pcadd_o_addr_pcbranchE[8]) );
  CLKIN0 U232 ( .A(u_decode_add_x_16_n156), .Q(n160) );
  NOR20 U233 ( .A(u_decode_add_x_16_n155), .B(n160), .Q(n161) );
  XNR20 U234 ( .A(u_decode_add_x_16_n158), .B(n161), .Q(
        u_decode_pcadd_o_addr_pcbranchE[3]) );
  NAND20 U235 ( .A(add_x_1_n46), .B(mem_data_pc4[10]), .Q(n162) );
  XNR20 U236 ( .A(mem_data_pc4[11]), .B(n162), .Q(n163) );
  MUX21 U237 ( .A(data_address[11]), .B(n163), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[11]) );
  CLKIN0 U238 ( .A(data_address[8]), .Q(n164) );
  XNR20 U239 ( .A(add_x_1_n55), .B(mem_data_pc4[8]), .Q(n165) );
  IMUX20 U240 ( .A(n164), .B(n165), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[8]) );
  NAND20 U241 ( .A(add_x_1_n71), .B(mem_data_pc4[4]), .Q(n166) );
  XNR20 U242 ( .A(mem_data_pc4[5]), .B(n166), .Q(n167) );
  MUX21 U243 ( .A(data_address[5]), .B(n167), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[5]) );
  CLKIN0 U244 ( .A(data_address[3]), .Q(n168) );
  XNR20 U245 ( .A(mem_data_pc4[2]), .B(mem_data_pc4[3]), .Q(n169) );
  IMUX20 U246 ( .A(n168), .B(n169), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[3]) );
  XOR30 U247 ( .A(if_addr_j[17]), .B(if_addr_j[31]), .C(u_decode_add_x_16_n29), 
        .Q(u_decode_pcadd_o_addr_pcbranchE[31]) );
  CLKIN0 U248 ( .A(u_decode_add_x_16_n33), .Q(n170) );
  NOR20 U249 ( .A(u_decode_add_x_16_n32), .B(n170), .Q(n171) );
  XNR20 U250 ( .A(u_decode_add_x_16_n34), .B(n171), .Q(
        u_decode_pcadd_o_addr_pcbranchE[28]) );
  CLKIN0 U251 ( .A(u_decode_add_x_16_n41), .Q(n172) );
  NOR20 U252 ( .A(u_decode_add_x_16_n40), .B(n172), .Q(n173) );
  XNR20 U253 ( .A(u_decode_add_x_16_n42), .B(n173), .Q(
        u_decode_pcadd_o_addr_pcbranchE[26]) );
  CLKIN0 U254 ( .A(u_decode_add_x_16_n49), .Q(n174) );
  NOR20 U255 ( .A(u_decode_add_x_16_n48), .B(n174), .Q(n175) );
  XNR20 U256 ( .A(u_decode_add_x_16_n50), .B(n175), .Q(
        u_decode_pcadd_o_addr_pcbranchE[24]) );
  CLKIN0 U257 ( .A(u_decode_add_x_16_n57), .Q(n176) );
  NOR20 U258 ( .A(u_decode_add_x_16_n56), .B(n176), .Q(n177) );
  XNR20 U259 ( .A(u_decode_add_x_16_n58), .B(n177), .Q(
        u_decode_pcadd_o_addr_pcbranchE[22]) );
  CLKIN0 U260 ( .A(u_decode_add_x_16_n65), .Q(n178) );
  NOR20 U261 ( .A(u_decode_add_x_16_n64), .B(n178), .Q(n179) );
  XNR20 U262 ( .A(u_decode_add_x_16_n66), .B(n179), .Q(
        u_decode_pcadd_o_addr_pcbranchE[20]) );
  CLKIN0 U263 ( .A(u_decode_add_x_16_n87), .Q(n180) );
  AOI210 U264 ( .A(u_decode_add_x_16_n88), .B(u_decode_add_x_16_n84), .C(n180), 
        .Q(n181) );
  CLKIN0 U265 ( .A(u_decode_add_x_16_n82), .Q(n182) );
  NOR20 U266 ( .A(u_decode_add_x_16_n81), .B(n182), .Q(n183) );
  XNR20 U267 ( .A(n181), .B(n183), .Q(u_decode_pcadd_o_addr_pcbranchE[17]) );
  CLKIN0 U268 ( .A(u_decode_add_x_16_n122), .Q(n184) );
  NOR20 U269 ( .A(u_decode_add_x_16_n121), .B(n184), .Q(n185) );
  XNR20 U270 ( .A(u_decode_add_x_16_n123), .B(n185), .Q(
        u_decode_pcadd_o_addr_pcbranchE[10]) );
  CLKIN0 U271 ( .A(u_decode_add_x_16_n143), .Q(n186) );
  AOI210 U272 ( .A(u_decode_add_x_16_n144), .B(u_decode_add_x_16_n181), .C(
        n186), .Q(n187) );
  CLKIN0 U273 ( .A(u_decode_add_x_16_n138), .Q(n188) );
  NOR20 U274 ( .A(u_decode_add_x_16_n137), .B(n188), .Q(n189) );
  XNR20 U275 ( .A(n187), .B(n189), .Q(u_decode_pcadd_o_addr_pcbranchE[7]) );
  CLKIN0 U276 ( .A(u_decode_add_x_16_n152), .Q(n190) );
  NOR20 U277 ( .A(u_decode_add_x_16_n151), .B(n190), .Q(n191) );
  XNR20 U278 ( .A(u_decode_add_x_16_n153), .B(n191), .Q(
        u_decode_pcadd_o_addr_pcbranchE[4]) );
  OAI210 U279 ( .A(if_addr_j[2]), .B(id_addr_pc4[2]), .C(
        u_decode_add_x_16_n158), .Q(n192) );
  CLKIN0 U280 ( .A(n192), .Q(u_decode_pcadd_o_addr_pcbranchE[2]) );
  CLKIN0 U281 ( .A(add_x_1_n28), .Q(n193) );
  NOR20 U282 ( .A(add_x_1_n21), .B(n193), .Q(n194) );
  XNR20 U283 ( .A(mem_data_pc4[16]), .B(n194), .Q(n195) );
  MUX21 U284 ( .A(data_address[16]), .B(n195), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[16]) );
  CLKIN0 U285 ( .A(data_address[10]), .Q(n196) );
  XNR20 U286 ( .A(add_x_1_n46), .B(mem_data_pc4[10]), .Q(n197) );
  IMUX20 U287 ( .A(n196), .B(n197), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[10]) );
  CLKIN0 U288 ( .A(data_address[7]), .Q(n198) );
  NOR20 U289 ( .A(add_x_1_n63), .B(add_x_1_n62), .Q(n199) );
  XNR20 U290 ( .A(mem_data_pc4[7]), .B(n199), .Q(n200) );
  IMUX20 U291 ( .A(n198), .B(n200), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[7]) );
  CLKIN0 U292 ( .A(data_address[4]), .Q(n201) );
  XNR20 U293 ( .A(add_x_1_n71), .B(mem_data_pc4[4]), .Q(n202) );
  IMUX20 U294 ( .A(n201), .B(n202), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[4]) );
  CLKIN0 U295 ( .A(data_address[2]), .Q(n203) );
  IMUX20 U296 ( .A(n203), .B(mem_data_pc4[2]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[2]) );
  NOR24 U297 ( .A(n250), .B(n249), .Q(n349) );
  INV3 U298 ( .A(n252), .Q(n249) );
  AOI221 U299 ( .A(n349), .B(id_data_jr[9]), .C(n343), .D(if_addr_j[9]), .Q(
        n323) );
  AOI221 U300 ( .A(n349), .B(id_data_jr[13]), .C(n343), .D(if_addr_j[13]), .Q(
        n311) );
  AOI221 U301 ( .A(n349), .B(id_data_jr[4]), .C(n343), .D(if_addr_j[4]), .Q(
        n338) );
  AOI221 U302 ( .A(n349), .B(id_data_jr[7]), .C(n343), .D(if_addr_j[7]), .Q(
        n329) );
  AOI221 U303 ( .A(n349), .B(id_data_jr[15]), .C(n343), .D(if_addr_j[15]), .Q(
        n305) );
  AOI221 U304 ( .A(n349), .B(id_data_jr[8]), .C(n343), .D(if_addr_j[8]), .Q(
        n326) );
  AOI221 U305 ( .A(n349), .B(id_data_jr[16]), .C(n343), .D(if_addr_j[16]), .Q(
        n302) );
  AOI221 U306 ( .A(n349), .B(id_data_jr[3]), .C(n343), .D(if_addr_j[3]), .Q(
        n341) );
  AOI221 U307 ( .A(n349), .B(id_data_jr[14]), .C(n343), .D(if_addr_j[14]), .Q(
        n308) );
  AOI221 U308 ( .A(n349), .B(id_data_jr[11]), .C(n343), .D(if_addr_j[11]), .Q(
        n317) );
  AOI221 U309 ( .A(n349), .B(id_data_jr[12]), .C(n343), .D(if_addr_j[12]), .Q(
        n314) );
  MUX22 U310 ( .A(data_address[31]), .B(u_mem_pc8[31]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[31]) );
  CLKIN6 U311 ( .A(n253), .Q(n350) );
  NOR21 U312 ( .A(n347), .B(if_con_b), .Q(n252) );
  MUX22 U313 ( .A(data_address[29]), .B(u_mem_pc8[29]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[29]) );
  INV2 U314 ( .A(add_x_1_n64), .Q(add_x_1_n63) );
  INV2 U315 ( .A(add_x_4_n69), .Q(add_x_4_n68) );
  INV2 U316 ( .A(u_decode_add_x_16_n92), .Q(u_decode_add_x_16_n90) );
  INV2 U317 ( .A(n439), .Q(n440) );
  INV2 U318 ( .A(add_x_4_n77), .Q(add_x_4_n76) );
  INV2 U319 ( .A(add_x_1_n72), .Q(add_x_1_n71) );
  NOR21 U320 ( .A(add_x_4_n77), .B(add_x_4_n70), .Q(add_x_4_n69) );
  INV1 U321 ( .A(u_decode_add_x_16_n118), .Q(u_decode_add_x_16_n176) );
  NOR21 U322 ( .A(add_x_1_n72), .B(add_x_1_n65), .Q(add_x_1_n64) );
  INV2 U323 ( .A(u_fetch_jmux_i_addr_pc4_16_), .Q(n303) );
  INV2 U324 ( .A(u_fetch_jmux_i_addr_pc4_11_), .Q(n318) );
  INV2 U325 ( .A(u_fetch_jmux_i_addr_pc4_12_), .Q(n315) );
  INV2 U326 ( .A(u_fetch_jmux_i_addr_pc4_9_), .Q(n324) );
  INV2 U327 ( .A(u_fetch_jmux_i_addr_pc4_6_), .Q(n333) );
  INV2 U328 ( .A(u_fetch_jmux_i_addr_pc4_5_), .Q(n336) );
  NOR21 U329 ( .A(add_x_4_n52), .B(add_x_4_n15), .Q(add_x_4_n14) );
  AOI210 U330 ( .A(n438), .B(n439), .C(u_decode_control_o_con_aluop_1_), .Q(
        n437) );
  NAND22 U331 ( .A(add_x_1_n48), .B(add_x_1_n64), .Q(add_x_1_n47) );
  NAND22 U332 ( .A(add_x_4_n53), .B(add_x_4_n69), .Q(add_x_4_n52) );
  INV2 U333 ( .A(u_decode_add_x_16_n98), .Q(u_decode_add_x_16_n96) );
  INV3 U334 ( .A(mem_data_pc4[14]), .Q(add_x_1_n27) );
  NAND22 U335 ( .A(mem_data_pc4[2]), .B(mem_data_pc4[3]), .Q(add_x_1_n72) );
  INV3 U336 ( .A(mem_data_pc4[12]), .Q(add_x_1_n37) );
  OAI211 U337 ( .A(n243), .B(n257), .C(n256), .Q(n138) );
  OAI211 U338 ( .A(n243), .B(n261), .C(n260), .Q(n107) );
  OAI211 U339 ( .A(n241), .B(n352), .C(n351), .Q(n137) );
  OAI211 U340 ( .A(n240), .B(n352), .C(n348), .Q(n136) );
  OAI2111 U341 ( .A(instruction_address[2]), .B(n243), .C(n345), .D(n344), .Q(
        n135) );
  INV3 U342 ( .A(n244), .Q(n243) );
  INV3 U343 ( .A(n346), .Q(n244) );
  NAND33 U344 ( .A(n252), .B(n250), .C(n248), .Q(n346) );
  INV2 U345 ( .A(u_fetch_jmux_i_addr_pc4_31_), .Q(n257) );
  XOR21 U346 ( .A(mem_data_pc4[31]), .B(add_x_1_n1), .Q(u_mem_pc8[31]) );
  MUX22 U347 ( .A(data_address[30]), .B(u_mem_pc8[30]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[30]) );
  INV2 U348 ( .A(u_fetch_jmux_i_addr_pc4_30_), .Q(n261) );
  INV2 U349 ( .A(u_fetch_jmux_i_addr_pc4_28_), .Q(n267) );
  INV2 U350 ( .A(u_fetch_jmux_i_addr_pc4_27_), .Q(n270) );
  INV2 U351 ( .A(u_fetch_jmux_i_addr_pc4_26_), .Q(n273) );
  INV2 U352 ( .A(u_fetch_jmux_i_addr_pc4_25_), .Q(n276) );
  INV2 U353 ( .A(u_fetch_jmux_i_addr_pc4_24_), .Q(n279) );
  INV2 U354 ( .A(u_fetch_jmux_i_addr_pc4_23_), .Q(n282) );
  INV2 U355 ( .A(u_fetch_jmux_i_addr_pc4_22_), .Q(n285) );
  INV2 U356 ( .A(u_fetch_jmux_i_addr_pc4_17_), .Q(n300) );
  INV2 U357 ( .A(u_fetch_jmux_i_addr_pc4_21_), .Q(n288) );
  INV2 U358 ( .A(u_fetch_jmux_i_addr_pc4_13_), .Q(n312) );
  INV2 U359 ( .A(u_fetch_jmux_i_addr_pc4_14_), .Q(n309) );
  INV2 U360 ( .A(u_fetch_jmux_i_addr_pc4_20_), .Q(n291) );
  INV2 U361 ( .A(u_fetch_jmux_i_addr_pc4_15_), .Q(n306) );
  INV2 U362 ( .A(n401), .Q(n400) );
  AOI211 U363 ( .A(n353), .B(n354), .C(n207), .Q(u_decode_n1) );
  INV2 U364 ( .A(u_fetch_jmux_i_addr_pc4_19_), .Q(n294) );
  INV2 U365 ( .A(u_fetch_jmux_i_addr_pc4_7_), .Q(n330) );
  INV2 U366 ( .A(u_fetch_jmux_i_addr_pc4_10_), .Q(n321) );
  INV2 U367 ( .A(u_fetch_jmux_i_addr_pc4_8_), .Q(n327) );
  INV2 U368 ( .A(u_decode_control_o_con_aluop_4_), .Q(n354) );
  OAI211 U369 ( .A(n367), .B(n368), .C(n369), .Q(u_decode_for_o_con_fb[2]) );
  INV2 U370 ( .A(u_fetch_jmux_i_addr_pc4_18_), .Q(n297) );
  INV2 U371 ( .A(n368), .Q(n370) );
  INV2 U372 ( .A(n404), .Q(n402) );
  INV2 U373 ( .A(n437), .Q(u_decode_control_o_con_regwrite) );
  AOI211 U374 ( .A(n449), .B(n443), .C(n212), .Q(
        u_decode_control_o_con_aluop_4_) );
  NAND41 U375 ( .A(mem_read), .B(n374), .C(n373), .D(n375), .Q(n369) );
  INV3 U376 ( .A(add_x_1_n47), .Q(add_x_1_n46) );
  NAND31 U377 ( .A(for_FWmemread), .B(n394), .C(n395), .Q(n368) );
  INV3 U378 ( .A(add_x_4_n52), .Q(add_x_4_n51) );
  INV3 U379 ( .A(u_decode_add_x_16_n145), .Q(u_decode_add_x_16_n144) );
  INV1 U380 ( .A(u_decode_control_o_con_aluop_5_), .Q(n447) );
  OAI211 U381 ( .A(id_data_instr[28]), .B(n360), .C(n358), .Q(if_con_j[0]) );
  NAND21 U382 ( .A(ex_con_Wregwrite), .B(n425), .Q(n420) );
  INV2 U383 ( .A(u_fetch_jmux_i_addr_pc4_4_), .Q(n339) );
  INV2 U384 ( .A(u_decode_add_x_16_n116), .Q(u_decode_add_x_16_n114) );
  INV2 U385 ( .A(u_decode_add_x_16_n117), .Q(u_decode_add_x_16_n115) );
  INV2 U386 ( .A(u_decode_add_x_16_n91), .Q(u_decode_add_x_16_n89) );
  INV2 U387 ( .A(n413), .Q(n406) );
  NOR21 U388 ( .A(id_data_instr[27]), .B(n361), .Q(n360) );
  NAND41 U389 ( .A(for_FWmemread), .B(n430), .C(n431), .D(n413), .Q(n403) );
  NOR20 U390 ( .A(n441), .B(n359), .Q(u_decode_control_o_con_regdst) );
  OAI211 U391 ( .A(n212), .B(n443), .C(n444), .Q(
        u_decode_control_o_con_memread) );
  NOR21 U392 ( .A(n219), .B(n442), .Q(u_decode_control_o_con_memwrite) );
  INV3 U393 ( .A(u_decode_add_x_16_n154), .Q(u_decode_add_x_16_n153) );
  NAND22 U394 ( .A(n380), .B(n215), .Q(n373) );
  OAI212 U395 ( .A(id_data_instr[28]), .B(n363), .C(n358), .Q(if_con_ifstall)
         );
  NAND22 U396 ( .A(n445), .B(n208), .Q(n359) );
  INV2 U397 ( .A(add_x_4_n45), .Q(add_x_4_n44) );
  NAND41 U398 ( .A(mem_read), .B(n410), .C(n411), .D(n412), .Q(n409) );
  INV2 U399 ( .A(u_decode_add_x_16_n111), .Q(u_decode_add_x_16_n175) );
  INV3 U400 ( .A(add_x_4_n26), .Q(add_x_4_n25) );
  AOI311 U401 ( .A(if_addr_j[5]), .B(n362), .C(n218), .D(id_data_instr[26]), 
        .Q(n361) );
  NAND22 U402 ( .A(n432), .B(n213), .Q(n413) );
  INV2 U403 ( .A(u_fetch_jmux_i_addr_pc4_3_), .Q(n342) );
  INV1 U404 ( .A(u_decode_add_x_16_n148), .Q(u_decode_add_x_16_n182) );
  NAND21 U405 ( .A(id_data_instr[26]), .B(n448), .Q(n443) );
  INV2 U406 ( .A(u_decode_add_x_16_n129), .Q(u_decode_add_x_16_n178) );
  INV1 U407 ( .A(n358), .Q(n441) );
  INV2 U408 ( .A(add_x_1_n40), .Q(add_x_1_n39) );
  INV2 U409 ( .A(n448), .Q(n446) );
  INV3 U410 ( .A(u_decode_add_x_16_n86), .Q(u_decode_add_x_16_n84) );
  INV2 U411 ( .A(u_decode_add_x_16_n142), .Q(u_decode_add_x_16_n181) );
  MUX22 U412 ( .A(mem_data_alures[4]), .B(wb_data_memout[4]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[4]) );
  MUX22 U413 ( .A(mem_data_alures[5]), .B(wb_data_memout[5]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[5]) );
  MUX22 U414 ( .A(mem_data_alures[3]), .B(wb_data_memout[3]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[3]) );
  NAND22 U415 ( .A(instruction_address[3]), .B(instruction_address[2]), .Q(
        add_x_4_n77) );
  MUX22 U416 ( .A(mem_data_alures[1]), .B(wb_data_memout[1]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[1]) );
  MUX22 U417 ( .A(mem_data_alures[31]), .B(wb_data_memout[31]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[31]) );
  NOR31 U418 ( .A(id_data_instr[30]), .B(id_data_instr[29]), .C(
        id_data_instr[31]), .Q(n358) );
  NOR21 U419 ( .A(id_data_instr[27]), .B(n204), .Q(n363) );
  NOR21 U420 ( .A(id_data_instr[26]), .B(id_data_instr[27]), .Q(n445) );
  MUX22 U421 ( .A(mem_data_alures[16]), .B(wb_data_memout[16]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[16]) );
  INV2 U422 ( .A(mem_data_pc4[6]), .Q(add_x_1_n62) );
  MUX22 U423 ( .A(mem_data_alures[22]), .B(wb_data_memout[22]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[22]) );
  MUX22 U424 ( .A(mem_data_alures[25]), .B(wb_data_memout[25]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[25]) );
  MUX22 U425 ( .A(mem_data_alures[23]), .B(wb_data_memout[23]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[23]) );
  MUX22 U426 ( .A(mem_data_alures[29]), .B(wb_data_memout[29]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[29]) );
  MUX22 U427 ( .A(mem_data_alures[28]), .B(wb_data_memout[28]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[28]) );
  MUX22 U428 ( .A(mem_data_alures[0]), .B(wb_data_memout[0]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[0]) );
  MUX22 U429 ( .A(mem_data_alures[21]), .B(wb_data_memout[21]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[21]) );
  MUX22 U430 ( .A(mem_data_alures[6]), .B(wb_data_memout[6]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[6]) );
  MUX22 U431 ( .A(mem_data_alures[30]), .B(wb_data_memout[30]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[30]) );
  MUX22 U432 ( .A(mem_data_alures[26]), .B(wb_data_memout[26]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[26]) );
  MUX22 U433 ( .A(mem_data_alures[19]), .B(wb_data_memout[19]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[19]) );
  MUX22 U434 ( .A(mem_data_alures[2]), .B(wb_data_memout[2]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[2]) );
  MUX22 U435 ( .A(mem_data_alures[24]), .B(wb_data_memout[24]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[24]) );
  MUX22 U436 ( .A(mem_data_alures[27]), .B(wb_data_memout[27]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[27]) );
  MUX22 U437 ( .A(mem_data_alures[11]), .B(wb_data_memout[11]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[11]) );
  MUX22 U438 ( .A(mem_data_alures[20]), .B(wb_data_memout[20]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[20]) );
  MUX22 U439 ( .A(mem_data_alures[7]), .B(wb_data_memout[7]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[7]) );
  MUX22 U440 ( .A(mem_data_alures[8]), .B(wb_data_memout[8]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[8]) );
  MUX22 U441 ( .A(mem_data_alures[9]), .B(wb_data_memout[9]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[9]) );
  MUX22 U442 ( .A(mem_data_alures[10]), .B(wb_data_memout[10]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[10]) );
  MUX22 U443 ( .A(mem_data_alures[12]), .B(wb_data_memout[12]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[12]) );
  MUX22 U444 ( .A(mem_data_alures[13]), .B(wb_data_memout[13]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[13]) );
  MUX22 U445 ( .A(mem_data_alures[14]), .B(wb_data_memout[14]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[14]) );
  MUX22 U446 ( .A(mem_data_alures[15]), .B(wb_data_memout[15]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[15]) );
  MUX22 U447 ( .A(mem_data_alures[17]), .B(wb_data_memout[17]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[17]) );
  MUX22 U448 ( .A(mem_data_alures[18]), .B(wb_data_memout[18]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[18]) );
  NOR21 U449 ( .A(n205), .B(id_data_instr[30]), .Q(n355) );
  INV1 U450 ( .A(mem_con_Wregwrite), .Q(n393) );
  ADD22 U451 ( .A(add_x_1_n4), .B(mem_data_pc4[28]), .CO(add_x_1_n3), .S(
        u_mem_pc8[28]) );
  ADD22 U452 ( .A(add_x_1_n5), .B(mem_data_pc4[27]), .CO(add_x_1_n4), .S(
        u_mem_pc8[27]) );
  OAI210 U453 ( .A(n363), .B(n446), .C(n447), .Q(
        u_decode_control_o_con_aluop_2_) );
  INV3 U454 ( .A(u_decode_add_x_16_n124), .Q(u_decode_add_x_16_n123) );
  OAI210 U455 ( .A(n445), .B(n446), .C(n354), .Q(
        u_decode_control_o_con_aluop_3_) );
  NAND31 U456 ( .A(ex_con_Wregwrite), .B(n384), .C(n385), .Q(n371) );
  OAI2111 U457 ( .A(mem_addr_regdst[1]), .B(n414), .C(n415), .D(n416), .Q(n405) );
  OAI2111 U458 ( .A(for_o_addr_Erd[2]), .B(n209), .C(n422), .D(n423), .Q(n421)
         );
  AOI220 U459 ( .A(n350), .B(ex_data_pc4[0]), .C(n349), .D(id_data_jr[0]), .Q(
        n351) );
  INV3 U460 ( .A(if_con_ifstall), .Q(n347) );
  AOI220 U461 ( .A(instruction_address[16]), .B(n347), .C(n350), .D(
        if_addr_b[16]), .Q(n301) );
  NOR21 U462 ( .A(n247), .B(if_con_j[1]), .Q(n251) );
  NOR40 U463 ( .A(n406), .B(n407), .C(n408), .D(n409), .Q(n404) );
  BUF6 U464 ( .A(ex_data_immext[8]), .Q(n246) );
  BUF6 U465 ( .A(ex_data_immext[6]), .Q(n245) );
  NAND30 U466 ( .A(id_data_instr[28]), .B(n358), .C(n204), .Q(n366) );
  NAND20 U467 ( .A(n358), .B(n363), .Q(n365) );
  NOR30 U468 ( .A(n204), .B(n212), .C(id_data_instr[28]), .Q(n439) );
  AOI221 U469 ( .A(instruction_address[14]), .B(n347), .C(n350), .D(
        if_addr_b[14]), .Q(n307) );
  AOI221 U470 ( .A(instruction_address[15]), .B(n347), .C(n350), .D(
        if_addr_b[15]), .Q(n304) );
  AOI221 U471 ( .A(instruction_address[12]), .B(n347), .C(n350), .D(
        if_addr_b[12]), .Q(n313) );
  AOI221 U472 ( .A(instruction_address[13]), .B(n347), .C(n350), .D(
        if_addr_b[13]), .Q(n310) );
  NOR21 U473 ( .A(n440), .B(n441), .Q(u_decode_jbcon_o_con_aluPC4) );
  INV3 U474 ( .A(add_x_1_n29), .Q(add_x_1_n28) );
  NOR31 U475 ( .A(n370), .B(n367), .C(n371), .Q(u_decode_for_o_con_fb[1]) );
  AOI211 U476 ( .A(n368), .B(n372), .C(n367), .Q(u_decode_for_o_con_fb[0]) );
  NAND41 U477 ( .A(n381), .B(n371), .C(n382), .D(n383), .Q(n372) );
  IMUX20 U478 ( .A(if_addr_j[20]), .B(n214), .S(for_o_addr_Erd[2]), .Q(n385)
         );
  IMUX20 U479 ( .A(n216), .B(if_addr_j[18]), .S(for_o_addr_Erd[0]), .Q(n389)
         );
  IMUX20 U480 ( .A(n220), .B(if_addr_j[21]), .S(for_o_addr_Erd[3]), .Q(n388)
         );
  IMUX20 U481 ( .A(n206), .B(if_addr_j[19]), .S(for_o_addr_Erd[1]), .Q(n387)
         );
  NOR21 U482 ( .A(n400), .B(u_decode_for_o_con_fa_2_), .Q(
        u_decode_for_o_con_fa_1_) );
  NAND22 U483 ( .A(n402), .B(n403), .Q(u_decode_for_o_con_fa_2_) );
  AOI211 U484 ( .A(n403), .B(n405), .C(n404), .Q(u_decode_for_o_con_fa_0_) );
  IMUX20 U485 ( .A(if_addr_j[23]), .B(n211), .S(for_o_addr_Erd[0]), .Q(n422)
         );
  INV3 U486 ( .A(u_decode_add_x_16_n38), .Q(u_decode_add_x_16_n36) );
  INV3 U487 ( .A(u_decode_add_x_16_n46), .Q(u_decode_add_x_16_n44) );
  INV3 U488 ( .A(u_decode_add_x_16_n54), .Q(u_decode_add_x_16_n52) );
  INV3 U489 ( .A(u_decode_add_x_16_n62), .Q(u_decode_add_x_16_n60) );
  INV3 U490 ( .A(u_decode_add_x_16_n70), .Q(u_decode_add_x_16_n68) );
  OAI2111 U491 ( .A(n346), .B(n309), .C(n308), .D(n307), .Q(n123) );
  AOI221 U492 ( .A(n350), .B(ex_data_pc4[1]), .C(n349), .D(id_data_jr[1]), .Q(
        n348) );
  OAI2111 U493 ( .A(n346), .B(n306), .C(n305), .D(n304), .Q(n122) );
  OAI2111 U494 ( .A(n346), .B(n318), .C(n317), .D(n316), .Q(n126) );
  OAI2111 U495 ( .A(n346), .B(n315), .C(n314), .D(n313), .Q(n125) );
  OAI2111 U496 ( .A(n346), .B(n333), .C(n332), .D(n331), .Q(n131) );
  OAI2111 U497 ( .A(n346), .B(n312), .C(n311), .D(n310), .Q(n124) );
  OAI2111 U498 ( .A(n346), .B(n300), .C(n299), .D(n298), .Q(n120) );
  AOI221 U499 ( .A(instruction_address[17]), .B(n347), .C(n350), .D(
        if_addr_b[17]), .Q(n298) );
  OAI2111 U500 ( .A(n346), .B(n330), .C(n329), .D(n328), .Q(n130) );
  OAI2111 U501 ( .A(n346), .B(n327), .C(n326), .D(n325), .Q(n129) );
  OAI2111 U502 ( .A(n243), .B(n336), .C(n335), .D(n334), .Q(n132) );
  OAI2111 U503 ( .A(n243), .B(n288), .C(n287), .D(n286), .Q(n116) );
  OAI2111 U504 ( .A(n243), .B(n297), .C(n296), .D(n295), .Q(n119) );
  AOI211 U505 ( .A(n349), .B(id_data_jr[31]), .C(n255), .Q(n256) );
  AOI211 U506 ( .A(n349), .B(id_data_jr[30]), .C(n259), .Q(n260) );
  OAI2111 U507 ( .A(n346), .B(n324), .C(n323), .D(n322), .Q(n128) );
  OAI2111 U508 ( .A(n243), .B(n267), .C(n266), .D(n265), .Q(n109) );
  OAI2111 U509 ( .A(n264), .B(n238), .C(n263), .D(n262), .Q(n108) );
  OAI2111 U510 ( .A(n346), .B(n342), .C(n341), .D(n340), .Q(n134) );
  OAI2111 U511 ( .A(n346), .B(n321), .C(n320), .D(n319), .Q(n127) );
  OAI2111 U512 ( .A(n346), .B(n339), .C(n338), .D(n337), .Q(n133) );
  NOR21 U513 ( .A(n347), .B(n244), .Q(n352) );
  OAI2111 U514 ( .A(n243), .B(n294), .C(n293), .D(n292), .Q(n118) );
  OAI2111 U515 ( .A(n243), .B(n285), .C(n284), .D(n283), .Q(n115) );
  OAI2111 U516 ( .A(n243), .B(n291), .C(n290), .D(n289), .Q(n117) );
  OAI2111 U517 ( .A(n346), .B(n303), .C(n302), .D(n301), .Q(n121) );
  OAI2111 U518 ( .A(n243), .B(n279), .C(n278), .D(n277), .Q(n113) );
  OAI2111 U519 ( .A(n243), .B(n282), .C(n281), .D(n280), .Q(n114) );
  OAI2111 U520 ( .A(n243), .B(n276), .C(n275), .D(n274), .Q(n112) );
  OAI2111 U521 ( .A(n243), .B(n273), .C(n272), .D(n271), .Q(n111) );
  OAI2111 U522 ( .A(n243), .B(n270), .C(n269), .D(n268), .Q(n110) );
  NAND22 U523 ( .A(if_con_b), .B(if_con_ifstall), .Q(n253) );
  MUX21 U524 ( .A(data_address[12]), .B(u_mem_pc8[12]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[12]) );
  MUX21 U525 ( .A(data_address[21]), .B(u_mem_pc8[21]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[21]) );
  MUX21 U526 ( .A(data_address[20]), .B(u_mem_pc8[20]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[20]) );
  MUX21 U527 ( .A(data_address[19]), .B(u_mem_pc8[19]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[19]) );
  MUX21 U528 ( .A(data_address[18]), .B(u_mem_pc8[18]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[18]) );
  MUX21 U529 ( .A(data_address[14]), .B(u_mem_pc8[14]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[14]) );
  MUX21 U530 ( .A(data_address[0]), .B(u_mem_pc8[0]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[0]) );
  MUX21 U531 ( .A(data_address[17]), .B(u_mem_pc8[17]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[17]) );
  MUX21 U532 ( .A(data_address[1]), .B(u_mem_pc8[1]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[1]) );
  MUX21 U533 ( .A(data_address[6]), .B(u_mem_pc8[6]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[6]) );
  MUX21 U534 ( .A(data_address[22]), .B(u_mem_pc8[22]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[22]) );
  MUX21 U535 ( .A(data_address[23]), .B(u_mem_pc8[23]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[23]) );
  MUX21 U536 ( .A(data_address[24]), .B(u_mem_pc8[24]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[24]) );
  MUX21 U537 ( .A(data_address[25]), .B(u_mem_pc8[25]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[25]) );
  MUX21 U538 ( .A(data_address[26]), .B(u_mem_pc8[26]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[26]) );
  MUX21 U539 ( .A(data_address[27]), .B(u_mem_pc8[27]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[27]) );
  MUX21 U540 ( .A(data_address[28]), .B(u_mem_pc8[28]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[28]) );
  NAND22 U541 ( .A(n252), .B(n251), .Q(n264) );
  NAND22 U542 ( .A(n247), .B(if_con_j[1]), .Q(n250) );
  NAND22 U543 ( .A(n358), .B(n359), .Q(if_con_j[1]) );
  INV3 U544 ( .A(u_decode_add_x_16_n101), .Q(u_decode_add_x_16_n100) );
  INV3 U545 ( .A(n355), .Q(n442) );
  NAND22 U546 ( .A(n373), .B(n369), .Q(n367) );
  INV3 U547 ( .A(u_decode_add_x_16_n37), .Q(u_decode_add_x_16_n35) );
  INV3 U548 ( .A(u_decode_add_x_16_n45), .Q(u_decode_add_x_16_n43) );
  INV3 U549 ( .A(u_decode_add_x_16_n53), .Q(u_decode_add_x_16_n51) );
  INV3 U550 ( .A(u_decode_add_x_16_n61), .Q(u_decode_add_x_16_n59) );
  INV3 U551 ( .A(u_decode_add_x_16_n69), .Q(u_decode_add_x_16_n67) );
  AOI220 U552 ( .A(instruction_address[11]), .B(n347), .C(n350), .D(
        if_addr_b[11]), .Q(n316) );
  AOI220 U553 ( .A(instruction_address[6]), .B(n347), .C(n350), .D(
        if_addr_b[6]), .Q(n331) );
  AOI220 U554 ( .A(n349), .B(id_data_jr[6]), .C(n343), .D(if_addr_j[6]), .Q(
        n332) );
  AOI220 U555 ( .A(n349), .B(id_data_jr[17]), .C(n343), .D(if_addr_j[17]), .Q(
        n299) );
  AOI220 U556 ( .A(instruction_address[7]), .B(n347), .C(n350), .D(
        if_addr_b[7]), .Q(n328) );
  AOI220 U557 ( .A(instruction_address[8]), .B(n347), .C(n350), .D(
        if_addr_b[8]), .Q(n325) );
  AOI220 U558 ( .A(instruction_address[5]), .B(n347), .C(n350), .D(
        if_addr_b[5]), .Q(n334) );
  AOI220 U559 ( .A(n349), .B(id_data_jr[5]), .C(n343), .D(if_addr_j[5]), .Q(
        n335) );
  AOI220 U560 ( .A(instruction_address[21]), .B(n347), .C(n350), .D(
        if_addr_b[21]), .Q(n286) );
  AOI220 U561 ( .A(n349), .B(id_data_jr[21]), .C(n343), .D(if_addr_j[21]), .Q(
        n287) );
  AOI220 U562 ( .A(instruction_address[18]), .B(n347), .C(n350), .D(
        if_addr_b[18]), .Q(n295) );
  AOI220 U563 ( .A(n349), .B(id_data_jr[18]), .C(n343), .D(if_addr_j[18]), .Q(
        n296) );
  OAI210 U564 ( .A(n239), .B(n264), .C(n254), .Q(n255) );
  AOI220 U565 ( .A(instruction_address[31]), .B(n347), .C(n350), .D(
        if_addr_b[31]), .Q(n254) );
  OAI210 U566 ( .A(n237), .B(n264), .C(n258), .Q(n259) );
  AOI220 U567 ( .A(instruction_address[30]), .B(n347), .C(n350), .D(
        if_addr_b[30]), .Q(n258) );
  AOI220 U568 ( .A(instruction_address[9]), .B(n347), .C(n350), .D(
        if_addr_b[9]), .Q(n322) );
  AOI220 U569 ( .A(instruction_address[28]), .B(n347), .C(n350), .D(
        if_addr_b[28]), .Q(n265) );
  AOI220 U570 ( .A(n349), .B(id_data_jr[28]), .C(n343), .D(if_addr_j[28]), .Q(
        n266) );
  AOI220 U571 ( .A(instruction_address[29]), .B(n347), .C(n350), .D(
        if_addr_b[29]), .Q(n262) );
  AOI220 U572 ( .A(n349), .B(id_data_jr[29]), .C(n244), .D(
        u_fetch_jmux_i_addr_pc4_29_), .Q(n263) );
  AOI220 U573 ( .A(instruction_address[3]), .B(n347), .C(n350), .D(
        if_addr_b[3]), .Q(n340) );
  AOI220 U574 ( .A(instruction_address[10]), .B(n347), .C(n350), .D(
        if_addr_b[10]), .Q(n319) );
  AOI220 U575 ( .A(n349), .B(id_data_jr[10]), .C(n343), .D(if_addr_j[10]), .Q(
        n320) );
  AOI220 U576 ( .A(instruction_address[4]), .B(n347), .C(n350), .D(
        if_addr_b[4]), .Q(n337) );
  AOI220 U577 ( .A(instruction_address[2]), .B(n347), .C(n350), .D(
        if_addr_b[2]), .Q(n344) );
  AOI220 U578 ( .A(n349), .B(id_data_jr[2]), .C(n343), .D(if_addr_j[2]), .Q(
        n345) );
  AOI220 U579 ( .A(instruction_address[19]), .B(n347), .C(n350), .D(
        if_addr_b[19]), .Q(n292) );
  AOI220 U580 ( .A(n349), .B(id_data_jr[19]), .C(n343), .D(if_addr_j[19]), .Q(
        n293) );
  AOI220 U581 ( .A(instruction_address[22]), .B(n347), .C(n350), .D(
        if_addr_b[22]), .Q(n283) );
  AOI220 U582 ( .A(n349), .B(id_data_jr[22]), .C(n343), .D(if_addr_j[22]), .Q(
        n284) );
  AOI220 U583 ( .A(instruction_address[20]), .B(n347), .C(n350), .D(
        if_addr_b[20]), .Q(n289) );
  AOI220 U584 ( .A(n349), .B(id_data_jr[20]), .C(n343), .D(if_addr_j[20]), .Q(
        n290) );
  INV3 U585 ( .A(add_x_4_n34), .Q(add_x_4_n33) );
  AOI220 U586 ( .A(instruction_address[24]), .B(n347), .C(n350), .D(
        if_addr_b[24]), .Q(n277) );
  AOI220 U587 ( .A(n349), .B(id_data_jr[24]), .C(n343), .D(if_addr_j[24]), .Q(
        n278) );
  AOI220 U588 ( .A(instruction_address[23]), .B(n347), .C(n350), .D(
        if_addr_b[23]), .Q(n280) );
  AOI220 U589 ( .A(n349), .B(id_data_jr[23]), .C(n343), .D(if_addr_j[23]), .Q(
        n281) );
  AOI220 U590 ( .A(instruction_address[25]), .B(n347), .C(n350), .D(
        if_addr_b[25]), .Q(n274) );
  AOI220 U591 ( .A(n349), .B(id_data_jr[25]), .C(n343), .D(if_addr_j[25]), .Q(
        n275) );
  AOI220 U592 ( .A(instruction_address[26]), .B(n347), .C(n350), .D(
        if_addr_b[26]), .Q(n271) );
  AOI220 U593 ( .A(n349), .B(id_data_jr[26]), .C(n343), .D(if_addr_j[26]), .Q(
        n272) );
  AOI220 U594 ( .A(instruction_address[27]), .B(n347), .C(n350), .D(
        if_addr_b[27]), .Q(n268) );
  AOI220 U595 ( .A(n349), .B(id_data_jr[27]), .C(n343), .D(if_addr_j[27]), .Q(
        n269) );
  INV3 U596 ( .A(n251), .Q(n248) );
  INV3 U597 ( .A(if_con_j[0]), .Q(n247) );
  LOGIC0 U598 ( .Q(n242) );
  AOI310 U599 ( .A(n355), .B(n208), .C(n356), .D(
        u_decode_control_o_con_memtoreg), .Q(n353) );
  AOI210 U600 ( .A(n208), .B(id_data_instr[27]), .C(n357), .Q(u_decode_n6) );
  OAI2110 U601 ( .A(n208), .B(id_data_instr[27]), .C(n358), .D(
        id_data_instr[26]), .Q(n357) );
  NOR40 U602 ( .A(if_addr_j[2]), .B(if_addr_j[3]), .C(if_addr_j[4]), .D(
        if_addr_j[6]), .Q(n362) );
  OAI220 U603 ( .A(n364), .B(n365), .C(n212), .D(n366), .Q(
        u_decode_jbcon_o_con_bop[1]) );
  NOR20 U604 ( .A(if_addr_j[18]), .B(id_data_instr[28]), .Q(n364) );
  OAI310 U605 ( .A(if_addr_j[18]), .B(id_data_instr[28]), .C(n365), .D(n366), 
        .Q(u_decode_jbcon_o_con_bop[0]) );
  IMUX20 U606 ( .A(if_addr_j[20]), .B(n214), .S(for_addr_rtM[2]), .Q(n375) );
  NOR40 U607 ( .A(n376), .B(n377), .C(n378), .D(n379), .Q(n374) );
  IMUX20 U608 ( .A(n220), .B(if_addr_j[21]), .S(for_addr_rtM[3]), .Q(n379) );
  IMUX20 U609 ( .A(n206), .B(if_addr_j[19]), .S(for_addr_rtM[1]), .Q(n378) );
  IMUX20 U610 ( .A(n215), .B(if_addr_j[22]), .S(for_addr_rtM[4]), .Q(n377) );
  IMUX20 U611 ( .A(n216), .B(if_addr_j[18]), .S(for_addr_rtM[0]), .Q(n376) );
  NOR40 U612 ( .A(if_addr_j[19]), .B(if_addr_j[21]), .C(if_addr_j[18]), .D(
        if_addr_j[20]), .Q(n380) );
  IMUX20 U613 ( .A(if_addr_j[18]), .B(n216), .S(mem_addr_regdst[0]), .Q(n383)
         );
  IMUX20 U614 ( .A(if_addr_j[19]), .B(n206), .S(mem_addr_regdst[1]), .Q(n382)
         );
  NOR40 U615 ( .A(n386), .B(n387), .C(n388), .D(n389), .Q(n384) );
  IMUX20 U616 ( .A(n215), .B(if_addr_j[22]), .S(for_o_addr_Erd[4]), .Q(n386)
         );
  NOR40 U617 ( .A(n390), .B(n391), .C(n392), .D(n393), .Q(n381) );
  IMUX20 U618 ( .A(n220), .B(if_addr_j[21]), .S(mem_addr_regdst[3]), .Q(n392)
         );
  IMUX20 U619 ( .A(n214), .B(if_addr_j[20]), .S(mem_addr_regdst[2]), .Q(n391)
         );
  IMUX20 U620 ( .A(n215), .B(if_addr_j[22]), .S(mem_addr_regdst[4]), .Q(n390)
         );
  IMUX20 U621 ( .A(if_addr_j[22]), .B(n215), .S(for_addr_rtW[4]), .Q(n395) );
  NOR40 U622 ( .A(n396), .B(n397), .C(n398), .D(n399), .Q(n394) );
  IMUX20 U623 ( .A(n216), .B(if_addr_j[18]), .S(for_addr_rtW[0]), .Q(n399) );
  IMUX20 U624 ( .A(n206), .B(if_addr_j[19]), .S(for_addr_rtW[1]), .Q(n398) );
  IMUX20 U625 ( .A(n214), .B(if_addr_j[20]), .S(for_addr_rtW[2]), .Q(n397) );
  IMUX20 U626 ( .A(n220), .B(if_addr_j[21]), .S(for_addr_rtW[3]), .Q(n396) );
  IMUX20 U627 ( .A(if_addr_j[25]), .B(n209), .S(for_addr_rtM[2]), .Q(n412) );
  IMUX20 U628 ( .A(if_addr_j[26]), .B(n217), .S(for_addr_rtM[3]), .Q(n411) );
  IMUX20 U629 ( .A(if_addr_j[27]), .B(n213), .S(for_addr_rtM[4]), .Q(n410) );
  IMUX20 U630 ( .A(n211), .B(if_addr_j[23]), .S(for_addr_rtM[0]), .Q(n408) );
  IMUX20 U631 ( .A(n210), .B(if_addr_j[24]), .S(for_addr_rtM[1]), .Q(n407) );
  AOI2110 U632 ( .A(mem_addr_regdst[1]), .B(n210), .C(n401), .D(n417), .Q(n416) );
  IMUX20 U633 ( .A(n209), .B(if_addr_j[25]), .S(mem_addr_regdst[2]), .Q(n417)
         );
  NOR40 U634 ( .A(n418), .B(n419), .C(n420), .D(n421), .Q(n401) );
  OAI210 U635 ( .A(for_o_addr_Erd[2]), .B(n424), .C(n209), .Q(n423) );
  NOR40 U636 ( .A(for_o_addr_Erd[1]), .B(for_o_addr_Erd[3]), .C(
        for_o_addr_Erd[0]), .D(if_addr_j[27]), .Q(n424) );
  IMUX20 U637 ( .A(if_addr_j[27]), .B(n213), .S(for_o_addr_Erd[4]), .Q(n425)
         );
  IMUX20 U638 ( .A(n217), .B(if_addr_j[26]), .S(for_o_addr_Erd[3]), .Q(n419)
         );
  IMUX20 U639 ( .A(n210), .B(if_addr_j[24]), .S(for_o_addr_Erd[1]), .Q(n418)
         );
  NOR40 U640 ( .A(n426), .B(n427), .C(n428), .D(n393), .Q(n415) );
  IMUX20 U641 ( .A(n213), .B(if_addr_j[27]), .S(mem_addr_regdst[4]), .Q(n428)
         );
  IMUX20 U642 ( .A(n217), .B(if_addr_j[26]), .S(mem_addr_regdst[3]), .Q(n427)
         );
  IMUX20 U643 ( .A(n211), .B(if_addr_j[23]), .S(mem_addr_regdst[0]), .Q(n426)
         );
  NOR20 U644 ( .A(if_addr_j[24]), .B(n429), .Q(n414) );
  NOR40 U645 ( .A(mem_addr_regdst[0]), .B(mem_addr_regdst[4]), .C(
        mem_addr_regdst[2]), .D(mem_addr_regdst[3]), .Q(n429) );
  NOR40 U646 ( .A(if_addr_j[23]), .B(if_addr_j[25]), .C(if_addr_j[26]), .D(
        if_addr_j[24]), .Q(n432) );
  IMUX20 U647 ( .A(if_addr_j[26]), .B(n217), .S(for_addr_rtW[3]), .Q(n431) );
  NOR40 U648 ( .A(n433), .B(n434), .C(n435), .D(n436), .Q(n430) );
  IMUX20 U649 ( .A(n209), .B(if_addr_j[25]), .S(for_addr_rtW[2]), .Q(n436) );
  IMUX20 U650 ( .A(n213), .B(if_addr_j[27]), .S(for_addr_rtW[4]), .Q(n435) );
  IMUX20 U651 ( .A(n211), .B(if_addr_j[23]), .S(for_addr_rtW[0]), .Q(n434) );
  IMUX20 U652 ( .A(n210), .B(if_addr_j[24]), .S(for_addr_rtW[1]), .Q(n433) );
  AOI2110 U653 ( .A(n205), .B(n440), .C(id_data_instr[30]), .D(n219), .Q(
        u_decode_control_o_con_memtoreg) );
  NAND30 U654 ( .A(n438), .B(n439), .C(id_data_instr[31]), .Q(n444) );
  NOR20 U655 ( .A(id_data_instr[30]), .B(id_data_instr[29]), .Q(n438) );
  OAI310 U656 ( .A(id_data_instr[30]), .B(n440), .C(n219), .D(n442), .Q(
        u_decode_control_o_con_alusrc) );
  AOI2110 U657 ( .A(n205), .B(n359), .C(id_data_instr[30]), .D(
        id_data_instr[31]), .Q(u_decode_control_o_con_aluop_1_) );
  NOR40 U658 ( .A(id_data_instr[28]), .B(id_data_instr[31]), .C(n356), .D(n442), .Q(u_decode_control_o_con_aluop_5_) );
  NAND20 U659 ( .A(id_data_instr[26]), .B(id_data_instr[27]), .Q(n356) );
  NOR40 U660 ( .A(id_data_instr[30]), .B(id_data_instr[31]), .C(n205), .D(n208), .Q(n448) );
  NAND30 U661 ( .A(u_decode_control_o_con_aluop_0_), .B(n208), .C(n204), .Q(
        n449) );
  NOR20 U662 ( .A(id_data_instr[31]), .B(n442), .Q(
        u_decode_control_o_con_aluop_0_) );
endmodule

