module W_byte_extend