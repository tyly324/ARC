
module F_jumpmux ( i_addr_j, i_addr_jr, i_addr_pc4, i_con_jump, o_addr_jumpmux
 );
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [31:0] i_addr_pc4;
  input [1:0] i_con_jump;
  output [31:0] o_addr_jumpmux;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n23, n24,
         n45, n46, n67, n68, n1, n2, n3, n4, n5, n6, n19, n20, n21, n22, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n69, n70, n71,
         n72, n73, n74, n75, n76;

  BUF6 U1 ( .A(n75), .Q(n3) );
  NAND22 U2 ( .A(n73), .B(n72), .Q(o_addr_jumpmux[31]) );
  NAND22 U3 ( .A(i_addr_jr[28]), .B(n2), .Q(n64) );
  INV3 U4 ( .A(n19), .Q(n76) );
  AOI221 U5 ( .A(i_addr_j[23]), .B(n5), .C(i_addr_pc4[23]), .D(n4), .Q(n55) );
  BUF6 U6 ( .A(n76), .Q(n5) );
  NAND24 U7 ( .A(n17), .B(n18), .Q(o_addr_jumpmux[3]) );
  NAND23 U8 ( .A(n11), .B(n12), .Q(o_addr_jumpmux[6]) );
  NAND23 U9 ( .A(n67), .B(n68), .Q(o_addr_jumpmux[0]) );
  INV0 U10 ( .A(i_con_jump[0]), .Q(n20) );
  NAND21 U11 ( .A(i_con_jump[1]), .B(n20), .Q(n21) );
  AOI222 U12 ( .A(i_addr_pc4[3]), .B(n4), .C(i_addr_jr[3]), .D(n1), .Q(n17) );
  AOI222 U13 ( .A(i_addr_pc4[2]), .B(n3), .C(i_addr_jr[2]), .D(n1), .Q(n23) );
  BUF6 U14 ( .A(n74), .Q(n1) );
  AOI220 U15 ( .A(i_addr_j[10]), .B(n5), .C(i_addr_pc4[10]), .D(n3), .Q(n27)
         );
  AOI220 U16 ( .A(i_addr_j[12]), .B(n5), .C(i_addr_pc4[12]), .D(n3), .Q(n31)
         );
  AOI220 U17 ( .A(i_addr_j[13]), .B(n5), .C(i_addr_pc4[13]), .D(n3), .Q(n33)
         );
  AOI220 U18 ( .A(i_addr_j[14]), .B(n5), .C(i_addr_pc4[14]), .D(n3), .Q(n35)
         );
  AOI220 U19 ( .A(i_addr_j[17]), .B(n5), .C(i_addr_pc4[17]), .D(n3), .Q(n41)
         );
  AOI220 U20 ( .A(i_addr_j[18]), .B(n5), .C(i_addr_pc4[18]), .D(n3), .Q(n43)
         );
  AOI220 U21 ( .A(i_addr_j[21]), .B(n5), .C(i_addr_pc4[21]), .D(n3), .Q(n51)
         );
  AOI222 U22 ( .A(i_addr_j[31]), .B(n76), .C(i_addr_pc4[31]), .D(n4), .Q(n73)
         );
  BUF4 U23 ( .A(n74), .Q(n2) );
  CLKBU4 U24 ( .A(n75), .Q(n4) );
  NAND20 U25 ( .A(i_addr_j[1]), .B(n76), .Q(n46) );
  NAND20 U26 ( .A(i_addr_j[2]), .B(n76), .Q(n24) );
  NAND21 U27 ( .A(i_addr_j[7]), .B(n76), .Q(n10) );
  NAND21 U28 ( .A(i_addr_j[8]), .B(n76), .Q(n8) );
  NAND20 U29 ( .A(i_addr_j[6]), .B(n76), .Q(n12) );
  NAND20 U30 ( .A(i_addr_j[4]), .B(n76), .Q(n16) );
  NAND20 U31 ( .A(i_addr_j[3]), .B(n76), .Q(n18) );
  NAND20 U32 ( .A(i_addr_j[0]), .B(n76), .Q(n68) );
  NAND21 U33 ( .A(i_addr_j[5]), .B(n76), .Q(n14) );
  AOI221 U34 ( .A(i_addr_pc4[6]), .B(n4), .C(i_addr_jr[6]), .D(n1), .Q(n11) );
  AOI221 U35 ( .A(i_addr_pc4[7]), .B(n4), .C(i_addr_jr[7]), .D(n1), .Q(n9) );
  AOI221 U36 ( .A(i_addr_pc4[8]), .B(n4), .C(i_addr_jr[8]), .D(n1), .Q(n7) );
  AOI221 U37 ( .A(i_addr_pc4[4]), .B(n3), .C(i_addr_jr[4]), .D(n1), .Q(n15) );
  AOI221 U38 ( .A(i_addr_pc4[5]), .B(n3), .C(i_addr_jr[5]), .D(n1), .Q(n13) );
  INV3 U39 ( .A(n21), .Q(n74) );
  AOI221 U40 ( .A(i_addr_pc4[0]), .B(n3), .C(i_addr_jr[0]), .D(n1), .Q(n67) );
  AOI221 U41 ( .A(i_addr_pc4[1]), .B(n3), .C(i_addr_jr[1]), .D(n1), .Q(n45) );
  NAND22 U42 ( .A(n45), .B(n46), .Q(o_addr_jumpmux[1]) );
  NAND22 U43 ( .A(n23), .B(n24), .Q(o_addr_jumpmux[2]) );
  NAND22 U44 ( .A(n15), .B(n16), .Q(o_addr_jumpmux[4]) );
  NAND22 U45 ( .A(n13), .B(n14), .Q(o_addr_jumpmux[5]) );
  NAND22 U46 ( .A(n9), .B(n10), .Q(o_addr_jumpmux[7]) );
  NAND22 U47 ( .A(n7), .B(n8), .Q(o_addr_jumpmux[8]) );
  AOI221 U48 ( .A(i_addr_j[9]), .B(n5), .C(i_addr_pc4[9]), .D(n3), .Q(n25) );
  AOI221 U49 ( .A(i_addr_j[11]), .B(n5), .C(i_addr_pc4[11]), .D(n3), .Q(n29)
         );
  AOI221 U50 ( .A(i_addr_j[15]), .B(n5), .C(i_addr_pc4[15]), .D(n3), .Q(n37)
         );
  AOI221 U51 ( .A(i_addr_j[16]), .B(n5), .C(i_addr_pc4[16]), .D(n3), .Q(n39)
         );
  AOI221 U52 ( .A(i_addr_j[19]), .B(n5), .C(i_addr_pc4[19]), .D(n3), .Q(n47)
         );
  AOI221 U53 ( .A(i_addr_j[20]), .B(n5), .C(i_addr_pc4[20]), .D(n3), .Q(n49)
         );
  AOI221 U54 ( .A(i_addr_j[22]), .B(n5), .C(i_addr_pc4[22]), .D(n4), .Q(n53)
         );
  AOI221 U55 ( .A(i_addr_j[24]), .B(n5), .C(i_addr_pc4[24]), .D(n4), .Q(n57)
         );
  AOI221 U56 ( .A(i_addr_j[25]), .B(n5), .C(i_addr_pc4[25]), .D(n4), .Q(n59)
         );
  AOI221 U57 ( .A(i_addr_j[26]), .B(n5), .C(i_addr_pc4[26]), .D(n4), .Q(n61)
         );
  AOI221 U58 ( .A(i_addr_j[27]), .B(n76), .C(i_addr_pc4[27]), .D(n4), .Q(n63)
         );
  AOI221 U59 ( .A(i_addr_j[28]), .B(n76), .C(i_addr_pc4[28]), .D(n4), .Q(n65)
         );
  AOI221 U60 ( .A(i_addr_j[29]), .B(n76), .C(i_addr_pc4[29]), .D(n4), .Q(n69)
         );
  AOI221 U61 ( .A(i_addr_j[30]), .B(n76), .C(i_addr_pc4[30]), .D(n4), .Q(n71)
         );
  CLKIN3 U62 ( .A(i_con_jump[1]), .Q(n6) );
  NAND22 U63 ( .A(i_con_jump[0]), .B(n6), .Q(n19) );
  XNR21 U64 ( .A(i_con_jump[0]), .B(i_con_jump[1]), .Q(n75) );
  NAND22 U65 ( .A(i_addr_jr[9]), .B(n1), .Q(n22) );
  NAND22 U66 ( .A(n25), .B(n22), .Q(o_addr_jumpmux[9]) );
  NAND22 U67 ( .A(i_addr_jr[10]), .B(n1), .Q(n26) );
  NAND22 U68 ( .A(n27), .B(n26), .Q(o_addr_jumpmux[10]) );
  NAND22 U69 ( .A(i_addr_jr[11]), .B(n1), .Q(n28) );
  NAND22 U70 ( .A(n29), .B(n28), .Q(o_addr_jumpmux[11]) );
  NAND22 U71 ( .A(i_addr_jr[12]), .B(n1), .Q(n30) );
  NAND22 U72 ( .A(n31), .B(n30), .Q(o_addr_jumpmux[12]) );
  NAND22 U73 ( .A(i_addr_jr[13]), .B(n1), .Q(n32) );
  NAND22 U74 ( .A(n33), .B(n32), .Q(o_addr_jumpmux[13]) );
  NAND22 U75 ( .A(i_addr_jr[14]), .B(n1), .Q(n34) );
  NAND22 U76 ( .A(n35), .B(n34), .Q(o_addr_jumpmux[14]) );
  NAND22 U77 ( .A(i_addr_jr[15]), .B(n2), .Q(n36) );
  NAND22 U78 ( .A(n37), .B(n36), .Q(o_addr_jumpmux[15]) );
  NAND22 U79 ( .A(i_addr_jr[16]), .B(n2), .Q(n38) );
  NAND22 U80 ( .A(n39), .B(n38), .Q(o_addr_jumpmux[16]) );
  NAND22 U81 ( .A(i_addr_jr[17]), .B(n2), .Q(n40) );
  NAND22 U82 ( .A(n41), .B(n40), .Q(o_addr_jumpmux[17]) );
  NAND22 U83 ( .A(i_addr_jr[18]), .B(n2), .Q(n42) );
  NAND22 U84 ( .A(n43), .B(n42), .Q(o_addr_jumpmux[18]) );
  NAND22 U85 ( .A(i_addr_jr[19]), .B(n2), .Q(n44) );
  NAND22 U86 ( .A(n47), .B(n44), .Q(o_addr_jumpmux[19]) );
  NAND22 U87 ( .A(i_addr_jr[20]), .B(n2), .Q(n48) );
  NAND22 U88 ( .A(n49), .B(n48), .Q(o_addr_jumpmux[20]) );
  NAND22 U89 ( .A(i_addr_jr[21]), .B(n2), .Q(n50) );
  NAND22 U90 ( .A(n51), .B(n50), .Q(o_addr_jumpmux[21]) );
  NAND22 U91 ( .A(i_addr_jr[22]), .B(n2), .Q(n52) );
  NAND22 U92 ( .A(n53), .B(n52), .Q(o_addr_jumpmux[22]) );
  NAND22 U93 ( .A(i_addr_jr[23]), .B(n2), .Q(n54) );
  NAND22 U94 ( .A(n55), .B(n54), .Q(o_addr_jumpmux[23]) );
  NAND22 U95 ( .A(i_addr_jr[24]), .B(n2), .Q(n56) );
  NAND22 U96 ( .A(n57), .B(n56), .Q(o_addr_jumpmux[24]) );
  NAND22 U97 ( .A(i_addr_jr[25]), .B(n2), .Q(n58) );
  NAND22 U98 ( .A(n59), .B(n58), .Q(o_addr_jumpmux[25]) );
  NAND22 U99 ( .A(i_addr_jr[26]), .B(n2), .Q(n60) );
  NAND22 U100 ( .A(n61), .B(n60), .Q(o_addr_jumpmux[26]) );
  NAND22 U101 ( .A(i_addr_jr[27]), .B(n2), .Q(n62) );
  NAND22 U102 ( .A(n63), .B(n62), .Q(o_addr_jumpmux[27]) );
  NAND22 U103 ( .A(n65), .B(n64), .Q(o_addr_jumpmux[28]) );
  NAND22 U104 ( .A(i_addr_jr[29]), .B(n2), .Q(n66) );
  NAND22 U105 ( .A(n69), .B(n66), .Q(o_addr_jumpmux[29]) );
  NAND22 U106 ( .A(i_addr_jr[30]), .B(n2), .Q(n70) );
  NAND22 U107 ( .A(n71), .B(n70), .Q(o_addr_jumpmux[30]) );
  NAND22 U108 ( .A(i_addr_jr[31]), .B(n2), .Q(n72) );
endmodule


module F_branchmux ( i_addr_jumpmux, i_addr_b, i_con_ifbranch, o_addr_nextpc
 );
  input [31:0] i_addr_jumpmux;
  input [31:0] i_addr_b;
  output [31:0] o_addr_nextpc;
  input i_con_ifbranch;
  wire   n35, n36, n37, n38, n39, n40, n43, n54, n65, n1, n2, n3, n4;

  INV3 U1 ( .A(i_con_ifbranch), .Q(n3) );
  AOI222 U2 ( .A(i_addr_b[3]), .B(n1), .C(i_addr_jumpmux[3]), .D(n4), .Q(n40)
         );
  AOI222 U3 ( .A(i_addr_b[6]), .B(n2), .C(i_addr_jumpmux[6]), .D(n4), .Q(n37)
         );
  AOI222 U4 ( .A(i_addr_b[0]), .B(n1), .C(i_addr_jumpmux[0]), .D(n4), .Q(n65)
         );
  MUX24 U5 ( .A(i_addr_jumpmux[20]), .B(i_addr_b[20]), .S(n2), .Q(
        o_addr_nextpc[20]) );
  MUX24 U6 ( .A(i_addr_jumpmux[19]), .B(i_addr_b[19]), .S(n1), .Q(
        o_addr_nextpc[19]) );
  MUX24 U7 ( .A(i_addr_jumpmux[24]), .B(i_addr_b[24]), .S(n1), .Q(
        o_addr_nextpc[24]) );
  MUX24 U8 ( .A(i_addr_jumpmux[16]), .B(i_addr_b[16]), .S(n2), .Q(
        o_addr_nextpc[16]) );
  CLKIN6 U9 ( .A(n54), .Q(o_addr_nextpc[1]) );
  AOI222 U10 ( .A(i_addr_b[1]), .B(n1), .C(i_addr_jumpmux[1]), .D(n4), .Q(n54)
         );
  CLKIN3 U11 ( .A(n3), .Q(n1) );
  INV1 U12 ( .A(i_con_ifbranch), .Q(n4) );
  CLKIN3 U13 ( .A(n65), .Q(o_addr_nextpc[0]) );
  CLKIN3 U14 ( .A(n43), .Q(o_addr_nextpc[2]) );
  CLKIN3 U15 ( .A(n40), .Q(o_addr_nextpc[3]) );
  CLKIN3 U16 ( .A(n37), .Q(o_addr_nextpc[6]) );
  CLKIN3 U17 ( .A(n36), .Q(o_addr_nextpc[7]) );
  CLKIN3 U18 ( .A(n35), .Q(o_addr_nextpc[8]) );
  CLKIN3 U19 ( .A(n39), .Q(o_addr_nextpc[4]) );
  CLKIN3 U20 ( .A(n38), .Q(o_addr_nextpc[5]) );
  INV3 U21 ( .A(n3), .Q(n2) );
  AOI221 U22 ( .A(i_addr_b[2]), .B(n1), .C(i_addr_jumpmux[2]), .D(n4), .Q(n43)
         );
  AOI221 U23 ( .A(i_addr_b[4]), .B(n2), .C(i_addr_jumpmux[4]), .D(n4), .Q(n39)
         );
  AOI221 U24 ( .A(i_addr_b[5]), .B(n2), .C(i_addr_jumpmux[5]), .D(n4), .Q(n38)
         );
  AOI221 U25 ( .A(i_addr_b[7]), .B(n2), .C(i_addr_jumpmux[7]), .D(n3), .Q(n36)
         );
  AOI221 U26 ( .A(i_addr_b[8]), .B(n2), .C(i_addr_jumpmux[8]), .D(n3), .Q(n35)
         );
  MUX22 U27 ( .A(i_addr_jumpmux[9]), .B(i_addr_b[9]), .S(n2), .Q(
        o_addr_nextpc[9]) );
  MUX22 U28 ( .A(i_addr_jumpmux[10]), .B(i_addr_b[10]), .S(n2), .Q(
        o_addr_nextpc[10]) );
  MUX22 U29 ( .A(i_addr_jumpmux[11]), .B(i_addr_b[11]), .S(n2), .Q(
        o_addr_nextpc[11]) );
  MUX22 U30 ( .A(i_addr_jumpmux[12]), .B(i_addr_b[12]), .S(n2), .Q(
        o_addr_nextpc[12]) );
  MUX22 U31 ( .A(i_addr_jumpmux[13]), .B(i_addr_b[13]), .S(n2), .Q(
        o_addr_nextpc[13]) );
  MUX22 U32 ( .A(i_addr_jumpmux[14]), .B(i_addr_b[14]), .S(n2), .Q(
        o_addr_nextpc[14]) );
  MUX22 U33 ( .A(i_addr_jumpmux[15]), .B(i_addr_b[15]), .S(n2), .Q(
        o_addr_nextpc[15]) );
  MUX22 U34 ( .A(i_addr_jumpmux[17]), .B(i_addr_b[17]), .S(n2), .Q(
        o_addr_nextpc[17]) );
  MUX22 U35 ( .A(i_addr_jumpmux[18]), .B(i_addr_b[18]), .S(n2), .Q(
        o_addr_nextpc[18]) );
  MUX22 U36 ( .A(i_addr_jumpmux[21]), .B(i_addr_b[21]), .S(n2), .Q(
        o_addr_nextpc[21]) );
  MUX22 U37 ( .A(i_addr_jumpmux[22]), .B(i_addr_b[22]), .S(n1), .Q(
        o_addr_nextpc[22]) );
  MUX22 U38 ( .A(i_addr_jumpmux[23]), .B(i_addr_b[23]), .S(n1), .Q(
        o_addr_nextpc[23]) );
  MUX22 U39 ( .A(i_addr_jumpmux[25]), .B(i_addr_b[25]), .S(n1), .Q(
        o_addr_nextpc[25]) );
  MUX22 U40 ( .A(i_addr_jumpmux[26]), .B(i_addr_b[26]), .S(n1), .Q(
        o_addr_nextpc[26]) );
  MUX22 U41 ( .A(i_addr_jumpmux[27]), .B(i_addr_b[27]), .S(n1), .Q(
        o_addr_nextpc[27]) );
  MUX22 U42 ( .A(i_addr_jumpmux[28]), .B(i_addr_b[28]), .S(n1), .Q(
        o_addr_nextpc[28]) );
  MUX22 U43 ( .A(i_addr_jumpmux[29]), .B(i_addr_b[29]), .S(n1), .Q(
        o_addr_nextpc[29]) );
  MUX22 U44 ( .A(i_addr_jumpmux[30]), .B(i_addr_b[30]), .S(n1), .Q(
        o_addr_nextpc[30]) );
  MUX22 U45 ( .A(i_addr_jumpmux[31]), .B(i_addr_b[31]), .S(n1), .Q(
        o_addr_nextpc[31]) );
endmodule


module F_pc ( i_clk, i_rst_n, i_con_stall, i_addr_next_pc, o_addr_pc );
  input [31:0] i_addr_next_pc;
  output [31:0] o_addr_pc;
  input i_clk, i_rst_n, i_con_stall;
  wire   n1, n2;

  DFEC1 program_counter_reg_30_ ( .D(i_addr_next_pc[30]), .E(n2), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[30]) );
  DFEC1 program_counter_reg_28_ ( .D(i_addr_next_pc[28]), .E(n2), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[28]) );
  DFEC1 program_counter_reg_25_ ( .D(i_addr_next_pc[25]), .E(n1), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[25]) );
  DFEC1 program_counter_reg_15_ ( .D(i_addr_next_pc[15]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[15]) );
  DFEC1 program_counter_reg_23_ ( .D(i_addr_next_pc[23]), .E(n1), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[23]) );
  DFEC1 program_counter_reg_20_ ( .D(i_addr_next_pc[20]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[20]) );
  DFEC1 program_counter_reg_19_ ( .D(i_addr_next_pc[19]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[19]) );
  DFEC1 program_counter_reg_24_ ( .D(i_addr_next_pc[24]), .E(n1), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[24]) );
  DFEC1 program_counter_reg_13_ ( .D(i_addr_next_pc[13]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[13]) );
  DFEC1 program_counter_reg_6_ ( .D(i_addr_next_pc[6]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[6]) );
  DFEC1 program_counter_reg_10_ ( .D(i_addr_next_pc[10]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[10]) );
  DFEC1 program_counter_reg_16_ ( .D(i_addr_next_pc[16]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[16]) );
  DFEC1 program_counter_reg_11_ ( .D(i_addr_next_pc[11]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[11]) );
  DFEC1 program_counter_reg_9_ ( .D(i_addr_next_pc[9]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[9]) );
  DFEC1 program_counter_reg_12_ ( .D(i_addr_next_pc[12]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[12]) );
  DFEC1 program_counter_reg_3_ ( .D(i_addr_next_pc[3]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[3]) );
  DFEC1 program_counter_reg_21_ ( .D(i_addr_next_pc[21]), .E(n1), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[21]) );
  DFEC1 program_counter_reg_0_ ( .D(i_addr_next_pc[0]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[0]) );
  DFEC1 program_counter_reg_5_ ( .D(i_addr_next_pc[5]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[5]) );
  DFEC1 program_counter_reg_22_ ( .D(i_addr_next_pc[22]), .E(n1), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[22]) );
  DFEC1 program_counter_reg_17_ ( .D(i_addr_next_pc[17]), .E(n2), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[17]) );
  DFEC1 program_counter_reg_1_ ( .D(i_addr_next_pc[1]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[1]) );
  DFEC1 program_counter_reg_7_ ( .D(i_addr_next_pc[7]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[7]) );
  DFEC1 program_counter_reg_4_ ( .D(i_addr_next_pc[4]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[4]) );
  DFEC1 program_counter_reg_2_ ( .D(i_addr_next_pc[2]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[2]) );
  DFEC1 program_counter_reg_18_ ( .D(i_addr_next_pc[18]), .E(n2), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[18]) );
  DFEC1 program_counter_reg_27_ ( .D(i_addr_next_pc[27]), .E(n1), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[27]) );
  DFEC1 program_counter_reg_26_ ( .D(i_addr_next_pc[26]), .E(n1), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[26]) );
  DFEC1 program_counter_reg_14_ ( .D(i_addr_next_pc[14]), .E(n2), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[14]) );
  DFEC1 program_counter_reg_29_ ( .D(i_addr_next_pc[29]), .E(n2), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[29]) );
  DFEC1 program_counter_reg_31_ ( .D(i_addr_next_pc[31]), .E(n2), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[31]) );
  DFEC1 program_counter_reg_8_ ( .D(i_addr_next_pc[8]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[8]) );
  BUF2 U2 ( .A(i_con_stall), .Q(n1) );
  BUF2 U3 ( .A(i_con_stall), .Q(n2) );
endmodule


module F_add4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV6 U2 ( .A(n65), .Q(n46) );
  NOR22 U3 ( .A(n6), .B(n106), .Q(n104) );
  INV3 U4 ( .A(A[22]), .Q(n57) );
  NAND22 U5 ( .A(n44), .B(n46), .Q(n52) );
  NAND22 U6 ( .A(n67), .B(n46), .Q(n68) );
  NAND22 U7 ( .A(n18), .B(n23), .Q(n19) );
  NAND21 U8 ( .A(n2), .B(n3), .Q(n1) );
  NAND31 U9 ( .A(n94), .B(n3), .C(A[12]), .Q(n97) );
  XOR21 U10 ( .A(n70), .B(n78), .Q(SUM[17]) );
  NAND22 U11 ( .A(A[16]), .B(n46), .Q(n78) );
  NAND22 U12 ( .A(n74), .B(n46), .Q(n76) );
  NAND22 U13 ( .A(n60), .B(n46), .Q(n66) );
  NAND31 U14 ( .A(n46), .B(n49), .C(n44), .Q(n48) );
  CLKIN3 U15 ( .A(n96), .Q(n92) );
  INV3 U16 ( .A(A[2]), .Q(SUM[2]) );
  NOR22 U17 ( .A(n24), .B(n25), .Q(n23) );
  NAND22 U18 ( .A(A[19]), .B(A[16]), .Q(n69) );
  INV3 U19 ( .A(A[17]), .Q(n70) );
  NAND31 U20 ( .A(A[3]), .B(A[2]), .C(A[4]), .Q(n108) );
  NAND42 U21 ( .A(n79), .B(n80), .C(n81), .D(n82), .Q(n65) );
  XNR22 U22 ( .A(A[15]), .B(n89), .Q(SUM[15]) );
  NAND31 U23 ( .A(A[13]), .B(n94), .C(A[12]), .Q(n93) );
  XNR22 U24 ( .A(A[7]), .B(n7), .Q(SUM[7]) );
  NAND42 U25 ( .A(A[18]), .B(A[21]), .C(n53), .D(n54), .Q(n30) );
  XOR21 U26 ( .A(A[19]), .B(n72), .Q(SUM[19]) );
  NAND42 U27 ( .A(n31), .B(n32), .C(n33), .D(n34), .Q(n24) );
  INV1 U28 ( .A(n61), .Q(n60) );
  INV0 U29 ( .A(A[13]), .Q(n95) );
  NAND22 U30 ( .A(n44), .B(n46), .Q(n51) );
  XOR21 U31 ( .A(A[25]), .B(n50), .Q(SUM[25]) );
  XOR21 U32 ( .A(n27), .B(n48), .Q(SUM[26]) );
  XOR21 U33 ( .A(n62), .B(n66), .Q(SUM[21]) );
  XOR21 U34 ( .A(n71), .B(n76), .Q(SUM[18]) );
  XNR21 U35 ( .A(A[29]), .B(n22), .Q(SUM[29]) );
  XNR20 U36 ( .A(n11), .B(n12), .Q(SUM[5]) );
  CLKIN0 U37 ( .A(A[8]), .Q(n4) );
  CLKIN0 U38 ( .A(A[16]), .Q(n77) );
  CLKIN0 U39 ( .A(A[9]), .Q(n5) );
  XOR21 U40 ( .A(n23), .B(A[28]), .Q(SUM[28]) );
  CLKIN0 U41 ( .A(A[3]), .Q(n16) );
  XNR21 U42 ( .A(A[11]), .B(n103), .Q(SUM[11]) );
  INV3 U43 ( .A(n65), .Q(n75) );
  NAND20 U44 ( .A(n74), .B(n75), .Q(n73) );
  NOR20 U45 ( .A(n61), .B(n65), .Q(n64) );
  XOR21 U46 ( .A(n95), .B(n97), .Q(SUM[13]) );
  XOR21 U47 ( .A(n57), .B(n63), .Q(SUM[22]) );
  XOR21 U48 ( .A(n5), .B(n1), .Q(SUM[9]) );
  NAND30 U49 ( .A(A[6]), .B(A[5]), .C(A[7]), .Q(n109) );
  XOR20 U50 ( .A(n46), .B(A[16]), .Q(SUM[16]) );
  XNR20 U51 ( .A(A[12]), .B(n99), .Q(SUM[12]) );
  XNR21 U52 ( .A(A[27]), .B(n43), .Q(SUM[27]) );
  XOR20 U53 ( .A(n14), .B(A[4]), .Q(SUM[4]) );
  XNR20 U54 ( .A(A[8]), .B(n6), .Q(SUM[8]) );
  NAND20 U55 ( .A(A[4]), .B(A[3]), .Q(n36) );
  NAND20 U56 ( .A(A[2]), .B(A[8]), .Q(n35) );
  INV0 U57 ( .A(A[5]), .Q(n12) );
  NAND20 U58 ( .A(A[6]), .B(A[5]), .Q(n38) );
  NAND20 U59 ( .A(A[12]), .B(A[11]), .Q(n40) );
  NAND20 U60 ( .A(A[10]), .B(A[9]), .Q(n39) );
  NAND20 U61 ( .A(A[14]), .B(A[13]), .Q(n42) );
  CLKIN3 U62 ( .A(A[7]), .Q(n37) );
  NAND20 U63 ( .A(A[10]), .B(A[11]), .Q(n102) );
  NAND20 U64 ( .A(A[8]), .B(A[9]), .Q(n101) );
  NAND20 U65 ( .A(A[4]), .B(n14), .Q(n13) );
  CLKIN3 U66 ( .A(A[15]), .Q(n41) );
  XOR20 U67 ( .A(A[3]), .B(A[2]), .Q(SUM[3]) );
  INV0 U68 ( .A(A[10]), .Q(n105) );
  INV0 U69 ( .A(A[6]), .Q(n9) );
  INV0 U70 ( .A(A[14]), .Q(n91) );
  NOR21 U71 ( .A(n37), .B(n85), .Q(n81) );
  NOR21 U72 ( .A(n83), .B(n84), .Q(n82) );
  NOR21 U73 ( .A(n41), .B(n88), .Q(n79) );
  XNR21 U74 ( .A(n90), .B(n91), .Q(SUM[14]) );
  NAND22 U75 ( .A(n64), .B(A[21]), .Q(n63) );
  NOR21 U76 ( .A(n47), .B(n51), .Q(n50) );
  XNR21 U77 ( .A(n104), .B(n105), .Q(SUM[10]) );
  XNR21 U78 ( .A(n8), .B(n9), .Q(SUM[6]) );
  INV3 U79 ( .A(n30), .Q(n44) );
  INV3 U80 ( .A(n92), .Q(n3) );
  INV3 U81 ( .A(n107), .Q(n106) );
  NOR21 U82 ( .A(n5), .B(n4), .Q(n107) );
  NAND22 U83 ( .A(n44), .B(n26), .Q(n25) );
  INV3 U84 ( .A(n10), .Q(n8) );
  NAND22 U85 ( .A(n11), .B(A[5]), .Q(n10) );
  INV3 U86 ( .A(n98), .Q(n94) );
  NOR21 U87 ( .A(n70), .B(n77), .Q(n74) );
  NOR21 U88 ( .A(n47), .B(n29), .Q(n49) );
  NOR21 U89 ( .A(n57), .B(n62), .Q(n59) );
  INV3 U90 ( .A(n4), .Q(n2) );
  NOR21 U91 ( .A(n57), .B(n70), .Q(n53) );
  NOR21 U92 ( .A(n55), .B(n56), .Q(n54) );
  NAND22 U93 ( .A(n67), .B(A[20]), .Q(n61) );
  NAND22 U94 ( .A(n104), .B(A[10]), .Q(n103) );
  XNR21 U95 ( .A(A[24]), .B(n52), .Q(SUM[24]) );
  NOR21 U96 ( .A(n73), .B(n71), .Q(n72) );
  XNR21 U97 ( .A(A[20]), .B(n68), .Q(SUM[20]) );
  NAND22 U98 ( .A(n90), .B(A[14]), .Q(n89) );
  NAND31 U99 ( .A(n45), .B(n46), .C(n44), .Q(n43) );
  NOR31 U100 ( .A(n47), .B(n27), .C(n29), .Q(n45) );
  NOR31 U101 ( .A(n71), .B(n69), .C(n70), .Q(n67) );
  INV3 U102 ( .A(A[25]), .Q(n29) );
  XNR21 U103 ( .A(A[23]), .B(n58), .Q(SUM[23]) );
  NAND31 U104 ( .A(n59), .B(n60), .C(n46), .Q(n58) );
  XNR21 U105 ( .A(A[31]), .B(n17), .Q(SUM[31]) );
  NAND31 U106 ( .A(n23), .B(n18), .C(A[30]), .Q(n17) );
  NOR21 U107 ( .A(SUM[2]), .B(n16), .Q(n14) );
  NOR31 U108 ( .A(n29), .B(n27), .C(n28), .Q(n26) );
  NAND22 U109 ( .A(A[27]), .B(A[24]), .Q(n28) );
  NOR21 U110 ( .A(n108), .B(n109), .Q(n96) );
  INV3 U111 ( .A(A[18]), .Q(n71) );
  NOR21 U112 ( .A(n92), .B(n93), .Q(n90) );
  INV3 U113 ( .A(A[26]), .Q(n27) );
  NAND22 U114 ( .A(A[2]), .B(A[8]), .Q(n83) );
  NAND22 U115 ( .A(A[4]), .B(A[3]), .Q(n84) );
  NAND22 U116 ( .A(A[16]), .B(A[19]), .Q(n55) );
  NAND22 U117 ( .A(A[6]), .B(A[5]), .Q(n85) );
  NAND22 U118 ( .A(A[14]), .B(A[13]), .Q(n88) );
  NAND22 U119 ( .A(A[20]), .B(A[23]), .Q(n56) );
  NAND22 U120 ( .A(n94), .B(n3), .Q(n99) );
  NAND22 U121 ( .A(A[28]), .B(n23), .Q(n22) );
  XNR21 U122 ( .A(A[30]), .B(n19), .Q(SUM[30]) );
  NAND22 U123 ( .A(n8), .B(A[6]), .Q(n7) );
  NOR21 U124 ( .A(n41), .B(n42), .Q(n31) );
  INV3 U125 ( .A(n100), .Q(n98) );
  NOR21 U126 ( .A(n101), .B(n102), .Q(n100) );
  NOR21 U127 ( .A(n37), .B(n38), .Q(n33) );
  NOR21 U128 ( .A(n86), .B(n87), .Q(n80) );
  NAND22 U129 ( .A(A[12]), .B(A[11]), .Q(n87) );
  NAND22 U130 ( .A(A[10]), .B(A[9]), .Q(n86) );
  NOR21 U131 ( .A(n39), .B(n40), .Q(n32) );
  INV3 U132 ( .A(n13), .Q(n11) );
  NOR21 U133 ( .A(n35), .B(n36), .Q(n34) );
  INV3 U134 ( .A(A[24]), .Q(n47) );
  INV3 U135 ( .A(A[21]), .Q(n62) );
  NOR21 U136 ( .A(n20), .B(n21), .Q(n18) );
  INV3 U137 ( .A(A[29]), .Q(n21) );
  INV3 U138 ( .A(A[28]), .Q(n20) );
  CLKIN3 U139 ( .A(n3), .Q(n6) );
endmodule


module F_add4 ( i_addr_pc, o_addr_pcadd4 );
  input [31:0] i_addr_pc;
  output [31:0] o_addr_pcadd4;
  wire   n2, n1;

  F_add4_DW01_add_1 add_5 ( .A(i_addr_pc), .B({n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n2, n1, n1}), .CI(n1), .SUM(o_addr_pcadd4) );
  LOGIC0 U3 ( .Q(n1) );
  LOGIC1 U4 ( .Q(n2) );
endmodule


module fetch ( i_clk, i_nrst, i_addr_b, i_addr_j, i_addr_jr, i_con_b, i_con_j, 
        i_data_instr, i_con_ifstall, o_addr_pc, o_addr_pc4, o_data_instr );
  input [31:0] i_addr_b;
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [1:0] i_con_j;
  input [31:0] i_data_instr;
  output [31:0] o_addr_pc;
  output [31:0] o_addr_pc4;
  output [31:0] o_data_instr;
  input i_clk, i_nrst, i_con_b, i_con_ifstall;

  wire   [31:0] jmux_i_addr_pc4;
  wire   [31:0] bmux_i_addr_jumpmux;
  wire   [31:0] pc_i_addr_next_pc;

  DFC3 pipe_instr_reg_31_ ( .D(i_data_instr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[31]) );
  DFC3 pipe_instr_reg_30_ ( .D(i_data_instr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[30]) );
  DFC3 pipe_instr_reg_29_ ( .D(i_data_instr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[29]) );
  DFC3 pipe_instr_reg_28_ ( .D(i_data_instr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[28]) );
  DFC3 pipe_instr_reg_27_ ( .D(i_data_instr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[27]) );
  DFC3 pipe_instr_reg_26_ ( .D(i_data_instr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[26]) );
  DFC3 pipe_instr_reg_25_ ( .D(i_data_instr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[25]) );
  DFC3 pipe_instr_reg_24_ ( .D(i_data_instr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[24]) );
  DFC3 pipe_instr_reg_23_ ( .D(i_data_instr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[23]) );
  DFC3 pipe_instr_reg_22_ ( .D(i_data_instr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[22]) );
  DFC3 pipe_instr_reg_21_ ( .D(i_data_instr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[21]) );
  DFC3 pipe_instr_reg_20_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[20]) );
  DFC3 pipe_instr_reg_19_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[19]) );
  DFC3 pipe_instr_reg_18_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[18]) );
  DFC3 pipe_instr_reg_17_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[17]) );
  DFC3 pipe_instr_reg_16_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[16]) );
  DFC3 pipe_instr_reg_15_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[15]) );
  DFC3 pipe_instr_reg_14_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[14]) );
  DFC3 pipe_instr_reg_13_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[13]) );
  DFC3 pipe_instr_reg_12_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[12]) );
  DFC3 pipe_instr_reg_11_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[11]) );
  DFC3 pipe_instr_reg_10_ ( .D(i_data_instr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[10]) );
  DFC3 pipe_instr_reg_9_ ( .D(i_data_instr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[9]) );
  DFC3 pipe_instr_reg_8_ ( .D(i_data_instr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[8]) );
  DFC3 pipe_instr_reg_7_ ( .D(i_data_instr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[7]) );
  DFC3 pipe_instr_reg_6_ ( .D(i_data_instr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[6]) );
  DFC3 pipe_instr_reg_5_ ( .D(i_data_instr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[5]) );
  DFC3 pipe_instr_reg_4_ ( .D(i_data_instr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[4]) );
  DFC3 pipe_instr_reg_3_ ( .D(i_data_instr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[3]) );
  DFC3 pipe_instr_reg_2_ ( .D(i_data_instr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[2]) );
  DFC3 pipe_instr_reg_1_ ( .D(i_data_instr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[1]) );
  DFC3 pipe_instr_reg_0_ ( .D(i_data_instr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[0]) );
  DFC3 pipe_pc4_reg_29_ ( .D(jmux_i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(jmux_i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(jmux_i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(jmux_i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(jmux_i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_pc4_reg_22_ ( .D(jmux_i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(jmux_i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_pc4_reg_19_ ( .D(jmux_i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(jmux_i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(jmux_i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(jmux_i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(jmux_i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(jmux_i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(jmux_i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(jmux_i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(jmux_i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(jmux_i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(jmux_i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(jmux_i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(jmux_i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(jmux_i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(jmux_i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(jmux_i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(jmux_i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(jmux_i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(jmux_i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(jmux_i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  F_jumpmux u_jumpmux ( .i_addr_j(i_addr_j), .i_addr_jr(i_addr_jr), 
        .i_addr_pc4(jmux_i_addr_pc4), .i_con_jump(i_con_j), .o_addr_jumpmux(
        bmux_i_addr_jumpmux) );
  F_branchmux u_branchmux ( .i_addr_jumpmux(bmux_i_addr_jumpmux), .i_addr_b(
        i_addr_b), .i_con_ifbranch(i_con_b), .o_addr_nextpc(pc_i_addr_next_pc)
         );
  F_pc u_pc ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_con_stall(i_con_ifstall), 
        .i_addr_next_pc(pc_i_addr_next_pc), .o_addr_pc(o_addr_pc) );
  F_add4 u_add4 ( .i_addr_pc(o_addr_pc), .o_addr_pcadd4(jmux_i_addr_pc4) );
  DFC1 pipe_pc4_reg_31_ ( .D(jmux_i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC1 pipe_pc4_reg_30_ ( .D(jmux_i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC1 pipe_pc4_reg_23_ ( .D(jmux_i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC1 pipe_pc4_reg_20_ ( .D(jmux_i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC1 pipe_pc4_reg_24_ ( .D(jmux_i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
endmodule


module D_control ( o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite, 
        o_con_alusrc, o_con_regwrite, o_con_ifsign, o_con_loadsig, o_con_aluop, 
        i_con_instru );
  output [1:0] o_con_loadsig;
  output [5:0] o_con_aluop;
  input [5:0] i_con_instru;
  output o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite,
         o_con_alusrc, o_con_regwrite, o_con_ifsign;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n1, n2, n3, n5, n6, n7, n8, n9, n10, n12, n13, n14,
         n16, n17, n18, n19, n20, n52;

  OAI212 U24 ( .A(n2), .B(n10), .C(n17), .Q(o_con_aluop[2]) );
  NOR41 U2 ( .A(n36), .B(n5), .C(n6), .D(n7), .Q(n21) );
  NAND31 U3 ( .A(n38), .B(i_con_instru[0]), .C(n39), .Q(n28) );
  INV1 U4 ( .A(i_con_instru[4]), .Q(n1) );
  NAND22 U5 ( .A(n14), .B(n39), .Q(n40) );
  INV1 U6 ( .A(i_con_instru[5]), .Q(n9) );
  CLKIN1 U7 ( .A(i_con_instru[3]), .Q(n18) );
  CLKIN2 U8 ( .A(i_con_instru[2]), .Q(n19) );
  INV1 U9 ( .A(n46), .Q(n14) );
  AOI2110 U10 ( .A(n1), .B(n7), .C(o_con_loadsig[0]), .D(o_con_loadsig[1]), 
        .Q(n25) );
  NOR21 U11 ( .A(n9), .B(i_con_instru[3]), .Q(n38) );
  NOR20 U12 ( .A(n27), .B(i_con_instru[4]), .Q(o_con_loadsig[1]) );
  NAND30 U13 ( .A(n23), .B(n20), .C(n50), .Q(n34) );
  NOR20 U14 ( .A(n28), .B(i_con_instru[4]), .Q(o_con_loadsig[0]) );
  NAND21 U15 ( .A(n50), .B(n52), .Q(n46) );
  NAND20 U16 ( .A(n36), .B(n1), .Q(n43) );
  OAI210 U17 ( .A(n2), .B(n26), .C(n25), .Q(o_con_memread) );
  NAND30 U18 ( .A(n40), .B(n26), .C(n45), .Q(n49) );
  NAND30 U19 ( .A(n50), .B(n23), .C(i_con_instru[1]), .Q(n41) );
  NAND20 U20 ( .A(i_con_instru[5]), .B(i_con_instru[3]), .Q(n33) );
  NAND30 U21 ( .A(n50), .B(i_con_instru[0]), .C(n39), .Q(n44) );
  AOI310 U22 ( .A(n21), .B(n8), .C(n22), .D(n2), .Q(o_con_regwrite) );
  INV0 U23 ( .A(i_con_instru[1]), .Q(n20) );
  NAND30 U25 ( .A(n20), .B(n19), .C(n52), .Q(n24) );
  OAI2111 U26 ( .A(n2), .B(n8), .C(n43), .D(n17), .Q(o_con_aluop[1]) );
  INV3 U27 ( .A(o_con_aluop[5]), .Q(n17) );
  NAND22 U28 ( .A(n25), .B(n3), .Q(o_con_memtoreg) );
  INV3 U29 ( .A(o_con_memwrite), .Q(n3) );
  INV3 U30 ( .A(n43), .Q(o_con_aluop[4]) );
  INV3 U31 ( .A(n42), .Q(o_con_aluop[3]) );
  AOI211 U32 ( .A(n1), .B(n32), .C(o_con_aluop[4]), .Q(n42) );
  INV3 U33 ( .A(n27), .Q(n6) );
  INV3 U34 ( .A(n28), .Q(n5) );
  NAND31 U35 ( .A(n38), .B(n52), .C(n39), .Q(n27) );
  NOR40 U36 ( .A(n16), .B(n12), .C(n32), .D(n30), .Q(n31) );
  INV3 U37 ( .A(n40), .Q(n12) );
  INV3 U38 ( .A(n51), .Q(n13) );
  NAND31 U39 ( .A(n35), .B(n44), .C(n34), .Q(n51) );
  INV3 U40 ( .A(n47), .Q(n8) );
  NAND41 U41 ( .A(n13), .B(n48), .C(n45), .D(n40), .Q(n47) );
  NAND41 U42 ( .A(n52), .B(n20), .C(n19), .D(n9), .Q(n48) );
  AOI311 U43 ( .A(n13), .B(n41), .C(n10), .D(n2), .Q(o_con_aluop[0]) );
  NAND22 U44 ( .A(n44), .B(n45), .Q(n32) );
  NAND22 U45 ( .A(n14), .B(n19), .Q(n35) );
  NOR21 U46 ( .A(n41), .B(n2), .Q(o_con_aluop[5]) );
  INV3 U47 ( .A(n1), .Q(n2) );
  INV3 U48 ( .A(n41), .Q(n16) );
  INV3 U49 ( .A(n49), .Q(n10) );
  NOR31 U50 ( .A(n18), .B(n2), .C(n9), .Q(o_con_memwrite) );
  NAND41 U51 ( .A(i_con_instru[2]), .B(i_con_instru[1]), .C(n50), .D(
        i_con_instru[0]), .Q(n26) );
  NAND41 U52 ( .A(n21), .B(n33), .C(n34), .D(n35), .Q(n30) );
  OAI311 U53 ( .A(n46), .B(i_con_instru[2]), .C(n20), .D(n26), .Q(n36) );
  NOR21 U54 ( .A(n19), .B(i_con_instru[1]), .Q(n39) );
  NOR21 U55 ( .A(n18), .B(i_con_instru[5]), .Q(n50) );
  NOR21 U56 ( .A(n52), .B(i_con_instru[2]), .Q(n23) );
  INV3 U57 ( .A(i_con_instru[0]), .Q(n52) );
  AOI311 U58 ( .A(n23), .B(n18), .C(i_con_instru[1]), .D(n16), .Q(n22) );
  INV3 U59 ( .A(n29), .Q(o_con_ifsign) );
  NAND22 U60 ( .A(n1), .B(n30), .Q(n29) );
  INV3 U61 ( .A(n37), .Q(n7) );
  NAND31 U62 ( .A(i_con_instru[1]), .B(n23), .C(n38), .Q(n37) );
  NAND31 U63 ( .A(i_con_instru[2]), .B(i_con_instru[1]), .C(n14), .Q(n45) );
  NOR40 U64 ( .A(n24), .B(i_con_instru[3]), .C(i_con_instru[5]), .D(n2), .Q(
        o_con_regdst) );
  NOR21 U65 ( .A(n2), .B(n31), .Q(o_con_alusrc) );
endmodule


module D_jb_control ( o_con_jump, o_con_bop, o_con_aluPC4, o_con_ifstall, 
        i_con_instru, i_con_func, i_con_rt );
  output [1:0] o_con_jump;
  output [2:0] o_con_bop;
  input [5:0] i_con_instru;
  input [5:0] i_con_func;
  input i_con_rt;
  output o_con_aluPC4, o_con_ifstall;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n1, n3, n4,
         n5, n6;

  OAI2112 U4 ( .A(n9), .B(n8), .C(n10), .D(n7), .Q(o_con_jump[0]) );
  OAI222 U13 ( .A(n5), .B(n16), .C(n14), .D(n17), .Q(o_con_bop[1]) );
  CLKIN3 U3 ( .A(i_con_instru[2]), .Q(n4) );
  NOR42 U5 ( .A(n11), .B(i_con_func[2]), .C(i_con_func[5]), .D(i_con_func[4]), 
        .Q(n9) );
  NAND22 U6 ( .A(n12), .B(i_con_func[3]), .Q(n11) );
  NOR31 U7 ( .A(i_con_instru[3]), .B(i_con_instru[5]), .C(i_con_instru[4]), 
        .Q(n7) );
  NOR20 U8 ( .A(i_con_func[1]), .B(i_con_func[0]), .Q(n12) );
  CLKIN6 U9 ( .A(i_con_instru[1]), .Q(n5) );
  CLKIN3 U10 ( .A(i_con_instru[0]), .Q(n6) );
  NAND30 U11 ( .A(n7), .B(n6), .C(i_con_instru[2]), .Q(n16) );
  NAND20 U12 ( .A(i_con_instru[0]), .B(n5), .Q(n14) );
  NOR20 U14 ( .A(i_con_instru[2]), .B(i_con_rt), .Q(n18) );
  NOR30 U15 ( .A(n15), .B(n3), .C(n6), .Q(o_con_bop[2]) );
  XNR20 U16 ( .A(n5), .B(i_con_instru[2]), .Q(n15) );
  NAND31 U17 ( .A(n5), .B(n4), .C(n6), .Q(n8) );
  NAND22 U18 ( .A(n7), .B(n8), .Q(o_con_jump[1]) );
  INV3 U19 ( .A(n7), .Q(n3) );
  NAND22 U20 ( .A(n7), .B(n1), .Q(n17) );
  OAI311 U21 ( .A(n1), .B(n3), .C(n14), .D(n16), .Q(o_con_bop[0]) );
  INV3 U22 ( .A(n13), .Q(o_con_ifstall) );
  AOI211 U23 ( .A(n4), .B(n14), .C(n3), .Q(n13) );
  NAND22 U24 ( .A(i_con_instru[1]), .B(n4), .Q(n10) );
  NOR40 U25 ( .A(i_con_instru[2]), .B(n3), .C(n5), .D(n6), .Q(o_con_aluPC4) );
  INV3 U26 ( .A(n18), .Q(n1) );
endmodule


module D_pcadd_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309;

  INV3 U2 ( .A(n165), .Q(n127) );
  INV3 U3 ( .A(B[21]), .Q(n10) );
  AOI211 U4 ( .A(n110), .B(n65), .C(n111), .Q(n107) );
  OAI2111 U5 ( .A(n135), .B(n136), .C(n137), .D(n138), .Q(n132) );
  NOR21 U6 ( .A(B[8]), .B(A[8]), .Q(n269) );
  INV3 U7 ( .A(n9), .Q(n8) );
  NAND22 U8 ( .A(n122), .B(n123), .Q(n121) );
  NAND22 U9 ( .A(n17), .B(n18), .Q(n15) );
  NAND22 U10 ( .A(n226), .B(n224), .Q(n251) );
  NAND22 U11 ( .A(n139), .B(n137), .Q(n154) );
  NAND22 U12 ( .A(n28), .B(n30), .Q(n31) );
  NAND22 U13 ( .A(n173), .B(n174), .Q(n194) );
  XNR21 U14 ( .A(n57), .B(n4), .Q(SUM[30]) );
  NAND22 U15 ( .A(n307), .B(n308), .Q(n17) );
  CLKIN3 U16 ( .A(n17), .Q(n233) );
  MUX22 U17 ( .A(B[0]), .B(n309), .S(A[0]), .Q(SUM[0]) );
  NAND22 U18 ( .A(n8), .B(A[20]), .Q(n136) );
  NOR22 U19 ( .A(n142), .B(n143), .Q(n141) );
  AOI211 U20 ( .A(n81), .B(n65), .C(n79), .Q(n84) );
  XOR20 U21 ( .A(n83), .B(n84), .Q(SUM[28]) );
  INV1 U22 ( .A(B[18]), .Q(n6) );
  INV1 U23 ( .A(B[25]), .Q(n13) );
  NOR21 U24 ( .A(B[24]), .B(A[24]), .Q(n98) );
  NOR21 U25 ( .A(B[27]), .B(A[27]), .Q(n99) );
  NAND22 U26 ( .A(B[21]), .B(A[21]), .Q(n137) );
  NAND31 U27 ( .A(n90), .B(n96), .C(n97), .Q(n95) );
  NAND33 U28 ( .A(n131), .B(n139), .C(n141), .Q(n125) );
  AOI211 U29 ( .A(n115), .B(n65), .C(n109), .Q(n114) );
  AOI211 U30 ( .A(n76), .B(n65), .C(n61), .Q(n75) );
  INV0 U31 ( .A(n65), .Q(n119) );
  NAND26 U32 ( .A(n120), .B(n121), .Q(n65) );
  NAND23 U33 ( .A(n199), .B(n200), .Q(n123) );
  AOI211 U34 ( .A(n188), .B(n177), .C(n189), .Q(n187) );
  NOR42 U35 ( .A(n268), .B(n233), .C(n269), .D(n270), .Q(n206) );
  AOI212 U36 ( .A(n126), .B(n127), .C(n128), .Q(n120) );
  NAND21 U37 ( .A(B[25]), .B(A[25]), .Q(n93) );
  NAND33 U38 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  INV1 U39 ( .A(n124), .Q(n159) );
  CLKIN0 U40 ( .A(B[3]), .Q(n300) );
  CLKIN0 U41 ( .A(B[6]), .Q(n286) );
  INV3 U42 ( .A(n211), .Q(n40) );
  CLKIN3 U43 ( .A(n129), .Q(n128) );
  AOI2110 U44 ( .A(n286), .B(n287), .C(n288), .D(n36), .Q(n281) );
  INV3 U45 ( .A(n177), .Q(n175) );
  NOR20 U46 ( .A(A[23]), .B(B[23]), .Q(n140) );
  OAI2111 U47 ( .A(n40), .B(n235), .C(n209), .D(n204), .Q(n263) );
  AOI311 U48 ( .A(n130), .B(n131), .C(n132), .D(n133), .Q(n129) );
  NAND22 U49 ( .A(n17), .B(n16), .Q(n279) );
  XOR20 U50 ( .A(n34), .B(n38), .Q(SUM[5]) );
  NAND22 U51 ( .A(n250), .B(n226), .Q(n249) );
  AOI210 U52 ( .A(n233), .B(n231), .C(n214), .Q(n265) );
  XNR20 U53 ( .A(n31), .B(n27), .Q(SUM[6]) );
  INV0 U54 ( .A(n231), .Q(n277) );
  NAND22 U55 ( .A(B[9]), .B(A[9]), .Q(n18) );
  NAND22 U56 ( .A(n64), .B(n65), .Q(n58) );
  CLKIN3 U57 ( .A(B[14]), .Q(n247) );
  CLKIN0 U58 ( .A(B[26]), .Q(n14) );
  NOR21 U59 ( .A(B[4]), .B(A[4]), .Q(n291) );
  NAND22 U60 ( .A(B[4]), .B(A[4]), .Q(n288) );
  CLKIN2 U61 ( .A(A[3]), .Q(n299) );
  NOR24 U62 ( .A(B[12]), .B(A[12]), .Q(n237) );
  NOR23 U63 ( .A(n237), .B(n238), .Q(n236) );
  NAND21 U64 ( .A(B[14]), .B(A[14]), .Q(n225) );
  NOR21 U65 ( .A(B[7]), .B(A[7]), .Q(n292) );
  CLKIN3 U66 ( .A(B[20]), .Q(n9) );
  CLKIN3 U67 ( .A(B[19]), .Q(n7) );
  CLKIN2 U68 ( .A(B[23]), .Q(n12) );
  INV3 U69 ( .A(n204), .Q(n203) );
  NAND20 U70 ( .A(n256), .B(n206), .Q(n252) );
  NOR20 U71 ( .A(n134), .B(n12), .Q(n133) );
  NOR20 U72 ( .A(n169), .B(n7), .Q(n168) );
  NAND20 U73 ( .A(n193), .B(n174), .Q(n192) );
  XOR20 U74 ( .A(n147), .B(n149), .Q(SUM[22]) );
  NOR20 U75 ( .A(n277), .B(n234), .Q(n278) );
  XOR20 U76 ( .A(n243), .B(n245), .Q(SUM[14]) );
  INV0 U77 ( .A(n36), .Q(n35) );
  AOI310 U78 ( .A(n267), .B(n18), .C(n231), .D(n234), .Q(n266) );
  XNR20 U79 ( .A(n251), .B(n250), .Q(SUM[13]) );
  XNR20 U80 ( .A(n154), .B(n153), .Q(SUM[21]) );
  XNR20 U81 ( .A(n193), .B(n194), .Q(SUM[17]) );
  INV3 U82 ( .A(n96), .Q(n94) );
  INV2 U83 ( .A(n125), .Q(n126) );
  INV3 U84 ( .A(n139), .Q(n135) );
  INV0 U85 ( .A(n37), .Q(n28) );
  NAND20 U86 ( .A(B[29]), .B(A[29]), .Q(n59) );
  INV0 U87 ( .A(B[17]), .Q(n5) );
  NOR20 U88 ( .A(A[24]), .B(B[24]), .Q(n112) );
  NOR20 U89 ( .A(A[29]), .B(B[29]), .Q(n63) );
  NAND21 U90 ( .A(B[10]), .B(A[10]), .Q(n231) );
  NOR20 U91 ( .A(A[11]), .B(B[11]), .Q(n214) );
  NAND21 U92 ( .A(B[6]), .B(A[6]), .Q(n30) );
  CLKIN0 U93 ( .A(B[22]), .Q(n11) );
  NAND21 U94 ( .A(B[13]), .B(A[13]), .Q(n224) );
  NAND21 U95 ( .A(B[17]), .B(A[17]), .Q(n173) );
  NOR24 U96 ( .A(B[15]), .B(A[15]), .Q(n238) );
  NOR20 U97 ( .A(A[8]), .B(B[8]), .Q(n280) );
  NOR20 U98 ( .A(A[28]), .B(B[28]), .Q(n82) );
  NOR20 U99 ( .A(A[4]), .B(B[4]), .Q(n41) );
  NOR20 U100 ( .A(A[27]), .B(B[27]), .Q(n91) );
  NOR20 U101 ( .A(A[7]), .B(B[7]), .Q(n284) );
  NOR20 U102 ( .A(A[20]), .B(n8), .Q(n160) );
  NAND20 U103 ( .A(B[24]), .B(A[24]), .Q(n92) );
  NAND20 U104 ( .A(B[22]), .B(A[22]), .Q(n138) );
  XNR20 U105 ( .A(B[28]), .B(A[28]), .Q(n83) );
  XNR20 U106 ( .A(B[27]), .B(A[27]), .Q(n100) );
  AOI212 U107 ( .A(n102), .B(n90), .C(n88), .Q(n101) );
  XOR20 U108 ( .A(n74), .B(n75), .Q(SUM[29]) );
  XNR20 U109 ( .A(B[29]), .B(A[29]), .Q(n74) );
  XNR21 U110 ( .A(n2), .B(n146), .Q(SUM[23]) );
  XOR20 U111 ( .A(B[23]), .B(A[23]), .Q(n2) );
  XNR20 U112 ( .A(B[15]), .B(A[15]), .Q(n241) );
  XNR20 U113 ( .A(B[19]), .B(A[19]), .Q(n186) );
  XNR20 U114 ( .A(B[7]), .B(A[7]), .Q(n25) );
  XNR20 U115 ( .A(B[11]), .B(A[11]), .Q(n273) );
  INV0 U116 ( .A(n234), .Q(n276) );
  IMUX20 U117 ( .A(n19), .B(n20), .S(n21), .Q(SUM[8]) );
  XNR20 U118 ( .A(B[8]), .B(A[8]), .Q(n20) );
  NOR20 U119 ( .A(B[8]), .B(A[8]), .Q(n22) );
  XNR20 U120 ( .A(B[12]), .B(A[12]), .Q(n261) );
  AOI210 U121 ( .A(n206), .B(n263), .C(n255), .Q(n262) );
  IMUX20 U122 ( .A(n197), .B(n198), .S(n155), .Q(SUM[16]) );
  XNR20 U123 ( .A(n8), .B(A[20]), .Q(n163) );
  AOI210 U124 ( .A(n181), .B(n9), .C(n182), .Q(n162) );
  AOI210 U125 ( .A(n159), .B(n123), .C(n127), .Q(n164) );
  NAND20 U126 ( .A(B[7]), .B(A[7]), .Q(n209) );
  NAND20 U127 ( .A(B[18]), .B(A[18]), .Q(n172) );
  NOR20 U128 ( .A(A[19]), .B(B[19]), .Q(n176) );
  NAND20 U129 ( .A(B[11]), .B(A[11]), .Q(n230) );
  NAND20 U130 ( .A(B[28]), .B(A[28]), .Q(n78) );
  NAND20 U131 ( .A(B[27]), .B(A[27]), .Q(n85) );
  XNR20 U132 ( .A(B[30]), .B(A[30]), .Q(n4) );
  NAND20 U133 ( .A(A[5]), .B(B[5]), .Q(n285) );
  NAND20 U134 ( .A(B[24]), .B(A[24]), .Q(n145) );
  NAND20 U135 ( .A(B[26]), .B(A[26]), .Q(n106) );
  XNR20 U136 ( .A(B[31]), .B(A[31]), .Q(n54) );
  NAND20 U137 ( .A(B[30]), .B(A[30]), .Q(n55) );
  NAND20 U138 ( .A(B[8]), .B(A[8]), .Q(n267) );
  XNR20 U139 ( .A(B[24]), .B(A[24]), .Q(n118) );
  NAND20 U140 ( .A(A[12]), .B(B[12]), .Q(n223) );
  INV0 U141 ( .A(A[6]), .Q(n287) );
  NOR20 U142 ( .A(A[15]), .B(B[15]), .Q(n227) );
  INV0 U143 ( .A(B[15]), .Q(n221) );
  INV0 U144 ( .A(A[15]), .Q(n220) );
  NOR20 U145 ( .A(A[2]), .B(B[2]), .Q(n52) );
  NOR20 U146 ( .A(A[12]), .B(B[12]), .Q(n257) );
  NOR20 U147 ( .A(B[24]), .B(A[24]), .Q(n144) );
  NAND20 U148 ( .A(B[8]), .B(A[8]), .Q(n24) );
  NAND20 U149 ( .A(B[4]), .B(A[4]), .Q(n42) );
  NAND20 U150 ( .A(B[12]), .B(A[12]), .Q(n254) );
  NAND20 U151 ( .A(B[5]), .B(A[5]), .Q(n32) );
  XNR21 U152 ( .A(n47), .B(n3), .Q(SUM[3]) );
  XNR20 U153 ( .A(B[3]), .B(A[3]), .Q(n3) );
  IMUX20 U154 ( .A(n43), .B(n44), .S(n40), .Q(SUM[4]) );
  XNR20 U155 ( .A(B[4]), .B(A[4]), .Q(n44) );
  NOR20 U156 ( .A(B[4]), .B(A[4]), .Q(n45) );
  NAND20 U157 ( .A(B[2]), .B(A[2]), .Q(n48) );
  NOR20 U158 ( .A(B[12]), .B(A[12]), .Q(n271) );
  NOR30 U159 ( .A(n303), .B(n52), .C(n304), .Q(n302) );
  XOR21 U160 ( .A(n188), .B(n190), .Q(SUM[18]) );
  NOR21 U161 ( .A(n189), .B(n175), .Q(n190) );
  OAI2111 U162 ( .A(n21), .B(n252), .C(n253), .D(n254), .Q(n250) );
  NAND22 U163 ( .A(n255), .B(n256), .Q(n253) );
  INV3 U164 ( .A(n257), .Q(n256) );
  OAI2111 U165 ( .A(n155), .B(n156), .C(n157), .D(n136), .Q(n153) );
  NAND22 U166 ( .A(n127), .B(n158), .Q(n157) );
  NAND22 U167 ( .A(n158), .B(n159), .Q(n156) );
  INV3 U168 ( .A(n160), .Q(n158) );
  OAI2111 U169 ( .A(n170), .B(n171), .C(n172), .D(n173), .Q(n167) );
  INV3 U170 ( .A(n284), .Q(n283) );
  INV3 U171 ( .A(n140), .Q(n130) );
  AOI311 U172 ( .A(n206), .B(n210), .C(n211), .D(n212), .Q(n199) );
  AOI221 U173 ( .A(n201), .B(n202), .C(n203), .D(n202), .Q(n200) );
  NOR21 U174 ( .A(n208), .B(n235), .Q(n210) );
  NAND31 U175 ( .A(n294), .B(n295), .C(n293), .Q(n211) );
  INV3 U176 ( .A(n302), .Q(n294) );
  AOI211 U177 ( .A(n296), .B(n297), .C(n298), .Q(n295) );
  INV3 U178 ( .A(n305), .Q(n293) );
  OAI311 U179 ( .A(n213), .B(n214), .C(n208), .D(n215), .Q(n212) );
  AOI311 U180 ( .A(n216), .B(n217), .C(n218), .D(n219), .Q(n215) );
  NOR21 U181 ( .A(n228), .B(n229), .Q(n213) );
  NOR21 U182 ( .A(n220), .B(n221), .Q(n219) );
  NAND22 U183 ( .A(n81), .B(n80), .Q(n66) );
  NAND22 U184 ( .A(n279), .B(n18), .Q(n275) );
  NAND22 U185 ( .A(n192), .B(n173), .Q(n188) );
  NAND22 U186 ( .A(n152), .B(n137), .Q(n147) );
  NAND22 U187 ( .A(n153), .B(n139), .Q(n152) );
  NAND22 U188 ( .A(n206), .B(n207), .Q(n205) );
  NAND22 U189 ( .A(n224), .B(n249), .Q(n243) );
  NAND22 U190 ( .A(n107), .B(n108), .Q(n102) );
  NAND22 U191 ( .A(n109), .B(n96), .Q(n108) );
  INV3 U192 ( .A(n93), .Q(n111) );
  NAND22 U193 ( .A(n230), .B(n264), .Q(n255) );
  NAND22 U194 ( .A(n265), .B(n266), .Q(n264) );
  XOR21 U195 ( .A(n275), .B(n278), .Q(SUM[10]) );
  NOR21 U196 ( .A(n148), .B(n150), .Q(n149) );
  NOR21 U197 ( .A(n244), .B(n246), .Q(n245) );
  XOR21 U198 ( .A(n102), .B(n103), .Q(SUM[26]) );
  NOR21 U199 ( .A(n88), .B(n104), .Q(n103) );
  XNR21 U200 ( .A(n15), .B(n16), .Q(SUM[9]) );
  XOR21 U201 ( .A(n113), .B(n114), .Q(SUM[25]) );
  NAND22 U202 ( .A(n96), .B(n93), .Q(n113) );
  INV3 U203 ( .A(n112), .Q(n115) );
  NAND22 U204 ( .A(n32), .B(n33), .Q(n27) );
  NAND22 U205 ( .A(n34), .B(n35), .Q(n33) );
  NAND22 U206 ( .A(n230), .B(n231), .Q(n229) );
  AOI211 U207 ( .A(n166), .B(n167), .C(n168), .Q(n165) );
  NOR21 U208 ( .A(n175), .B(n176), .Q(n166) );
  NOR21 U209 ( .A(n66), .B(n63), .Q(n64) );
  NOR21 U210 ( .A(n124), .B(n125), .Q(n122) );
  NOR21 U211 ( .A(n299), .B(n300), .Q(n298) );
  XOR21 U212 ( .A(n50), .B(n67), .Q(SUM[2]) );
  NOR21 U213 ( .A(n68), .B(n52), .Q(n67) );
  NOR21 U214 ( .A(n36), .B(n39), .Q(n38) );
  INV3 U215 ( .A(n32), .Q(n39) );
  NOR21 U216 ( .A(n112), .B(n94), .Q(n110) );
  INV3 U217 ( .A(n63), .Q(n62) );
  XOR21 U218 ( .A(n71), .B(n183), .Q(SUM[1]) );
  NOR21 U219 ( .A(n184), .B(n73), .Q(n183) );
  NAND22 U220 ( .A(n69), .B(n70), .Q(n50) );
  NAND22 U221 ( .A(n71), .B(n72), .Q(n70) );
  INV3 U222 ( .A(n73), .Q(n72) );
  AOI211 U223 ( .A(n300), .B(n299), .C(n73), .Q(n296) );
  INV3 U224 ( .A(n52), .Q(n51) );
  NOR21 U225 ( .A(A[10]), .B(B[10]), .Q(n270) );
  NOR21 U226 ( .A(B[11]), .B(A[11]), .Q(n268) );
  NAND22 U227 ( .A(n85), .B(n86), .Q(n79) );
  OAI2111 U228 ( .A(n87), .B(n88), .C(n89), .D(n90), .Q(n86) );
  INV3 U229 ( .A(n91), .Q(n89) );
  NOR21 U230 ( .A(A[5]), .B(B[5]), .Q(n36) );
  OAI2111 U231 ( .A(n222), .B(n223), .C(n224), .D(n225), .Q(n218) );
  NAND31 U232 ( .A(n177), .B(n174), .C(n178), .Q(n124) );
  NOR21 U233 ( .A(n179), .B(n180), .Q(n178) );
  NOR21 U234 ( .A(B[16]), .B(A[16]), .Q(n179) );
  NOR21 U235 ( .A(B[19]), .B(A[19]), .Q(n180) );
  NOR21 U236 ( .A(B[23]), .B(A[23]), .Q(n143) );
  NOR21 U237 ( .A(n8), .B(A[20]), .Q(n142) );
  NAND22 U238 ( .A(n5), .B(n195), .Q(n174) );
  INV3 U239 ( .A(A[17]), .Q(n195) );
  NAND22 U240 ( .A(n61), .B(n62), .Q(n60) );
  NOR21 U241 ( .A(A[10]), .B(B[10]), .Q(n234) );
  INV3 U242 ( .A(B[9]), .Q(n307) );
  INV3 U243 ( .A(A[9]), .Q(n308) );
  NAND22 U244 ( .A(n258), .B(n259), .Q(n226) );
  INV3 U245 ( .A(A[13]), .Q(n259) );
  INV3 U246 ( .A(B[13]), .Q(n258) );
  NAND22 U247 ( .A(n10), .B(n161), .Q(n139) );
  INV3 U248 ( .A(A[21]), .Q(n161) );
  AOI2111 U249 ( .A(n232), .B(n18), .C(n233), .D(n234), .Q(n228) );
  NAND22 U250 ( .A(B[8]), .B(A[8]), .Q(n232) );
  NAND22 U251 ( .A(n14), .B(n105), .Q(n90) );
  INV3 U252 ( .A(A[26]), .Q(n105) );
  NAND22 U253 ( .A(n247), .B(n248), .Q(n217) );
  INV3 U254 ( .A(A[14]), .Q(n248) );
  NAND22 U255 ( .A(n11), .B(n151), .Q(n131) );
  INV3 U256 ( .A(A[22]), .Q(n151) );
  XOR21 U257 ( .A(n25), .B(n26), .Q(SUM[7]) );
  AOI211 U258 ( .A(n27), .B(n28), .C(n29), .Q(n26) );
  NAND22 U259 ( .A(B[16]), .B(A[16]), .Q(n171) );
  NOR21 U260 ( .A(A[6]), .B(B[6]), .Q(n37) );
  NOR21 U261 ( .A(A[3]), .B(B[3]), .Q(n304) );
  AOI211 U262 ( .A(n92), .B(n93), .C(n94), .Q(n87) );
  NAND22 U263 ( .A(n6), .B(n191), .Q(n177) );
  INV3 U264 ( .A(A[18]), .Q(n191) );
  NAND22 U265 ( .A(n196), .B(n171), .Q(n193) );
  NAND22 U266 ( .A(n289), .B(n290), .Q(n235) );
  NOR21 U267 ( .A(n291), .B(n292), .Q(n289) );
  NOR21 U268 ( .A(n36), .B(n37), .Q(n290) );
  NAND22 U269 ( .A(n77), .B(n78), .Q(n61) );
  NAND22 U270 ( .A(n79), .B(n80), .Q(n77) );
  NOR21 U271 ( .A(n304), .B(n306), .Q(n305) );
  NAND22 U272 ( .A(A[2]), .B(B[2]), .Q(n306) );
  XOR21 U273 ( .A(n273), .B(n274), .Q(SUM[11]) );
  AOI211 U274 ( .A(n275), .B(n276), .C(n277), .Q(n274) );
  XOR21 U275 ( .A(n241), .B(n242), .Q(SUM[15]) );
  AOI211 U276 ( .A(n243), .B(n217), .C(n244), .Q(n242) );
  XOR21 U277 ( .A(n100), .B(n101), .Q(SUM[27]) );
  AOI211 U278 ( .A(n147), .B(n131), .C(n148), .Q(n146) );
  XOR21 U279 ( .A(n186), .B(n187), .Q(SUM[19]) );
  NOR21 U280 ( .A(n98), .B(n99), .Q(n97) );
  IMUX21 U281 ( .A(n162), .B(n163), .S(n164), .Q(SUM[20]) );
  IMUX21 U282 ( .A(n117), .B(n118), .S(n119), .Q(SUM[24]) );
  NOR21 U283 ( .A(n144), .B(n109), .Q(n117) );
  XNR21 U284 ( .A(B[16]), .B(A[16]), .Q(n198) );
  NOR21 U285 ( .A(n239), .B(n240), .Q(n197) );
  NOR21 U286 ( .A(B[16]), .B(A[16]), .Q(n239) );
  XNR21 U287 ( .A(n53), .B(n54), .Q(SUM[31]) );
  NAND22 U288 ( .A(n55), .B(n56), .Q(n53) );
  INV3 U289 ( .A(n227), .Q(n216) );
  NAND22 U290 ( .A(n13), .B(n116), .Q(n96) );
  INV3 U291 ( .A(A[25]), .Q(n116) );
  NOR21 U292 ( .A(n22), .B(n23), .Q(n19) );
  NOR21 U293 ( .A(n45), .B(n46), .Q(n43) );
  IMUX21 U294 ( .A(n260), .B(n261), .S(n262), .Q(SUM[12]) );
  NOR21 U295 ( .A(n271), .B(n272), .Q(n260) );
  INV3 U296 ( .A(n82), .Q(n80) );
  INV3 U297 ( .A(A[23]), .Q(n134) );
  INV3 U298 ( .A(A[19]), .Q(n169) );
  NAND22 U299 ( .A(n48), .B(n49), .Q(n47) );
  NAND22 U300 ( .A(n50), .B(n51), .Q(n49) );
  NOR21 U301 ( .A(A[1]), .B(B[1]), .Q(n73) );
  INV3 U302 ( .A(A[20]), .Q(n181) );
  INV3 U303 ( .A(B[0]), .Q(n309) );
  NAND22 U304 ( .A(B[1]), .B(A[1]), .Q(n303) );
  NAND22 U305 ( .A(B[1]), .B(A[1]), .Q(n69) );
  NOR21 U306 ( .A(n52), .B(n301), .Q(n297) );
  NAND22 U307 ( .A(B[0]), .B(A[0]), .Q(n301) );
  INV3 U308 ( .A(n185), .Q(n71) );
  NAND22 U309 ( .A(B[0]), .B(A[0]), .Q(n185) );
  CLKIN3 U310 ( .A(n24), .Q(n23) );
  CLKIN3 U311 ( .A(n30), .Q(n29) );
  OAI212 U312 ( .A(n40), .B(n41), .C(n42), .Q(n34) );
  CLKIN3 U313 ( .A(n42), .Q(n46) );
  OAI212 U314 ( .A(A[30]), .B(B[30]), .C(n57), .Q(n56) );
  CLKIN3 U315 ( .A(n48), .Q(n68) );
  CLKIN3 U316 ( .A(n66), .Q(n76) );
  CLKIN3 U317 ( .A(n95), .Q(n81) );
  CLKIN3 U318 ( .A(n90), .Q(n104) );
  CLKIN3 U319 ( .A(n106), .Q(n88) );
  CLKIN3 U320 ( .A(n145), .Q(n109) );
  CLKIN3 U321 ( .A(n131), .Q(n150) );
  CLKIN3 U322 ( .A(n138), .Q(n148) );
  CLKIN3 U323 ( .A(n174), .Q(n170) );
  CLKIN3 U324 ( .A(n136), .Q(n182) );
  CLKIN3 U325 ( .A(n69), .Q(n184) );
  CLKIN3 U326 ( .A(n172), .Q(n189) );
  OAI212 U327 ( .A(A[16]), .B(B[16]), .C(n123), .Q(n196) );
  CLKIN3 U328 ( .A(n123), .Q(n155) );
  CLKIN3 U329 ( .A(n205), .Q(n202) );
  CLKIN3 U330 ( .A(n208), .Q(n207) );
  CLKIN3 U331 ( .A(n209), .Q(n201) );
  CLKIN3 U332 ( .A(n226), .Q(n222) );
  NAND33 U333 ( .A(n217), .B(n226), .C(n236), .Q(n208) );
  CLKIN3 U334 ( .A(n171), .Q(n240) );
  CLKIN3 U335 ( .A(n217), .Q(n246) );
  CLKIN3 U336 ( .A(n225), .Q(n244) );
  CLKIN3 U337 ( .A(n254), .Q(n272) );
  OAI212 U338 ( .A(n21), .B(n280), .C(n24), .Q(n16) );
  CLKIN3 U339 ( .A(n263), .Q(n21) );
  OAI212 U340 ( .A(n281), .B(n282), .C(n283), .Q(n204) );
  OAI212 U341 ( .A(n37), .B(n285), .C(n30), .Q(n282) );
endmodule


module D_pcadd ( i_addr_pcadd4E, i_data_immshiftl, o_addr_pcbranchE );
  input [31:0] i_addr_pcadd4E;
  input [31:0] i_data_immshiftl;
  output [31:0] o_addr_pcbranchE;
  wire   n1;

  D_pcadd_DW01_add_1 add_5 ( .A(i_addr_pcadd4E), .B(i_data_immshiftl), .CI(n1), 
        .SUM(o_addr_pcbranchE) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_addr_Rt, i_con_RegWr, 
        i_addr_Rd, i_data_Rd, o_data_Rs, o_data_Rt );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rt;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr;
  wire   n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985;
  wire   [1023:0] regs;

  DFEC1 regs_reg_31__31_ ( .D(n926), .E(n958), .C(i_clk), .RN(n928), .Q(
        regs[1023]) );
  DFEC1 regs_reg_31__30_ ( .D(n922), .E(n958), .C(i_clk), .RN(n928), .Q(
        regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(n918), .E(n958), .C(i_clk), .RN(n928), .Q(
        regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(n914), .E(n958), .C(i_clk), .RN(n928), .Q(
        regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(n910), .E(n958), .C(i_clk), .RN(n928), .Q(
        regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(n906), .E(n958), .C(i_clk), .RN(n928), .Q(
        regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(n902), .E(n958), .C(i_clk), .RN(n928), .Q(
        regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(n898), .E(n958), .C(i_clk), .RN(n928), .Q(
        regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(n894), .E(n958), .C(i_clk), .RN(n928), .Q(
        regs[1015]) );
  DFEC1 regs_reg_30__31_ ( .D(n926), .E(n959), .C(i_clk), .RN(n931), .Q(
        regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(n922), .E(n959), .C(i_clk), .RN(n931), .Q(
        regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(n918), .E(n959), .C(i_clk), .RN(n931), .Q(
        regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(n914), .E(n959), .C(i_clk), .RN(n931), .Q(
        regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(n910), .E(n959), .C(i_clk), .RN(n932), .Q(
        regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(n906), .E(n959), .C(i_clk), .RN(n932), .Q(
        regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(n902), .E(n959), .C(i_clk), .RN(n932), .Q(
        regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(n898), .E(n959), .C(i_clk), .RN(n932), .Q(
        regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(n894), .E(n959), .C(i_clk), .RN(n932), .Q(
        regs[983]) );
  DFEC1 regs_reg_29__31_ ( .D(n926), .E(n960), .C(i_clk), .RN(n935), .Q(
        regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(n922), .E(n960), .C(i_clk), .RN(n935), .Q(
        regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(n918), .E(n960), .C(i_clk), .RN(n935), .Q(
        regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(n914), .E(n960), .C(i_clk), .RN(n935), .Q(
        regs[956]) );
  DFEC1 regs_reg_29__27_ ( .D(n910), .E(n960), .C(i_clk), .RN(n935), .Q(
        regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(n906), .E(n960), .C(i_clk), .RN(n935), .Q(
        regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(n902), .E(n960), .C(i_clk), .RN(n935), .Q(
        regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(n898), .E(n960), .C(i_clk), .RN(n935), .Q(
        regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(n894), .E(n960), .C(i_clk), .RN(n936), .Q(
        regs[951]) );
  DFEC1 regs_reg_28__31_ ( .D(n926), .E(n961), .C(i_clk), .RN(n938), .Q(
        regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(n922), .E(n961), .C(i_clk), .RN(n938), .Q(
        regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(n918), .E(n961), .C(i_clk), .RN(n938), .Q(
        regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(n914), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(
        regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(n910), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(
        regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(n906), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(
        regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(n902), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(
        regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(n898), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(
        regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(n894), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(
        regs[919]) );
  DFEC1 regs_reg_27__31_ ( .D(n926), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(n922), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(n918), .E(n962), .C(i_clk), .RN(n940), .Q(
        regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(n914), .E(n962), .C(i_clk), .RN(n939), .Q(
        regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(n910), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(n906), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(n902), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(n898), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(n894), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[887]) );
  DFEC1 regs_reg_26__31_ ( .D(n926), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(n922), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(n918), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(n914), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(n910), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(n906), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(n902), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(n898), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(n894), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[855]) );
  DFEC1 regs_reg_25__31_ ( .D(n926), .E(n956), .C(i_clk), .RN(n935), .Q(
        regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(n922), .E(n956), .C(i_clk), .RN(n936), .Q(
        regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(n918), .E(n956), .C(i_clk), .RN(n928), .Q(
        regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(n914), .E(n956), .C(i_clk), .RN(n929), .Q(
        regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(n910), .E(n956), .C(i_clk), .RN(n930), .Q(
        regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(n906), .E(n956), .C(i_clk), .RN(n931), .Q(
        regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(n902), .E(n956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(n898), .E(n956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(n894), .E(n956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[823]) );
  DFEC1 regs_reg_24__31_ ( .D(n926), .E(n957), .C(i_clk), .RN(n944), .Q(
        regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(n922), .E(n957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(n918), .E(n957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(n914), .E(n957), .C(i_clk), .RN(n934), .Q(
        regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(n910), .E(n957), .C(i_clk), .RN(n927), .Q(
        regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(n906), .E(n957), .C(i_clk), .RN(n935), .Q(
        regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(n902), .E(n957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(n898), .E(n957), .C(i_clk), .RN(n947), .Q(
        regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(n894), .E(n957), .C(i_clk), .RN(n946), .Q(
        regs[791]) );
  DFEC1 regs_reg_23__31_ ( .D(n925), .E(n948), .C(i_clk), .RN(n944), .Q(
        regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(n921), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(n917), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(n913), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(n909), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(n905), .E(n948), .C(i_clk), .RN(n928), .Q(
        regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(n901), .E(n948), .C(i_clk), .RN(n929), .Q(
        regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(n897), .E(n948), .C(i_clk), .RN(n930), .Q(
        regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(n893), .E(n948), .C(i_clk), .RN(n931), .Q(
        regs[759]) );
  DFEC1 regs_reg_22__31_ ( .D(n925), .E(n949), .C(i_clk), .RN(n942), .Q(
        regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(n921), .E(n949), .C(i_clk), .RN(n928), .Q(
        regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(n917), .E(n949), .C(i_clk), .RN(n929), .Q(
        regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(n913), .E(n949), .C(i_clk), .RN(n930), .Q(
        regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(n909), .E(n949), .C(i_clk), .RN(n931), .Q(
        regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(n905), .E(n949), .C(i_clk), .RN(n932), .Q(
        regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(n901), .E(n949), .C(i_clk), .RN(n933), .Q(
        regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(n897), .E(n949), .C(i_clk), .RN(n934), .Q(
        regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(n893), .E(n949), .C(i_clk), .RN(n935), .Q(
        regs[727]) );
  DFEC1 regs_reg_21__31_ ( .D(n925), .E(n950), .C(i_clk), .RN(n933), .Q(
        regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(n921), .E(n950), .C(i_clk), .RN(n934), .Q(
        regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(n917), .E(n950), .C(i_clk), .RN(n935), .Q(
        regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(n913), .E(n950), .C(i_clk), .RN(n936), .Q(
        regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(n909), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(n905), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(n901), .E(n950), .C(i_clk), .RN(n942), .Q(
        regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(n897), .E(n950), .C(i_clk), .RN(n930), .Q(
        regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(n893), .E(n950), .C(i_clk), .RN(n942), .Q(
        regs[695]) );
  DFEC1 regs_reg_20__31_ ( .D(n925), .E(n951), .C(i_clk), .RN(n939), .Q(
        regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(n921), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(n917), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(n913), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(n909), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(n905), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(n901), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(n897), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(n893), .E(n951), .C(i_clk), .RN(n940), .Q(
        regs[663]) );
  DFEC1 regs_reg_19__31_ ( .D(n925), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(n921), .E(n952), .C(i_clk), .RN(n928), .Q(
        regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(n917), .E(n952), .C(i_clk), .RN(n929), .Q(
        regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(n913), .E(n952), .C(i_clk), .RN(n946), .Q(
        regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(n909), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(n905), .E(n952), .C(i_clk), .RN(n938), .Q(
        regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(n901), .E(n952), .C(i_clk), .RN(n934), .Q(
        regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(n897), .E(n952), .C(i_clk), .RN(n940), .Q(
        regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(n893), .E(n952), .C(i_clk), .RN(n941), .Q(
        regs[631]) );
  DFEC1 regs_reg_18__31_ ( .D(n925), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(n921), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(n917), .E(n953), .C(i_clk), .RN(n942), .Q(
        regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(n913), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(n909), .E(n953), .C(i_clk), .RN(n931), .Q(
        regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(n905), .E(n953), .C(i_clk), .RN(n932), .Q(
        regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(n901), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(n897), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(n893), .E(n953), .C(i_clk), .RN(n939), .Q(
        regs[599]) );
  DFEC1 regs_reg_17__31_ ( .D(n925), .E(n954), .C(i_clk), .RN(n939), .Q(
        regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(n921), .E(n954), .C(i_clk), .RN(n929), .Q(
        regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(n917), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(n913), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(n909), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(n905), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(n901), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(n897), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(n893), .E(n954), .C(i_clk), .RN(n943), .Q(
        regs[567]) );
  DFEC1 regs_reg_16__31_ ( .D(n925), .E(n955), .C(i_clk), .RN(n943), .Q(
        regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(n921), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(n917), .E(n955), .C(i_clk), .RN(n937), .Q(
        regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(n913), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(n909), .E(n955), .C(i_clk), .RN(n946), .Q(
        regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(n905), .E(n955), .C(i_clk), .RN(n945), .Q(
        regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(n901), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(n897), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(n893), .E(n955), .C(i_clk), .RN(n946), .Q(
        regs[535]) );
  DFEC1 regs_reg_15__31_ ( .D(n924), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(n920), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(n916), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(n912), .E(n965), .C(i_clk), .RN(n933), .Q(
        regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(n908), .E(n965), .C(i_clk), .RN(n947), .Q(
        regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(n904), .E(n965), .C(i_clk), .RN(n935), .Q(
        regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(n900), .E(n965), .C(i_clk), .RN(n936), .Q(
        regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(n896), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(n892), .E(n965), .C(i_clk), .RN(n945), .Q(
        regs[503]) );
  DFEC1 regs_reg_14__31_ ( .D(n924), .E(n966), .C(i_clk), .RN(n939), .Q(
        regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(n920), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(n916), .E(n966), .C(i_clk), .RN(n947), .Q(
        regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(n912), .E(n966), .C(i_clk), .RN(n947), .Q(
        regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(n908), .E(n966), .C(i_clk), .RN(n935), .Q(
        regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(n904), .E(n966), .C(i_clk), .RN(n944), .Q(
        regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(n900), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(n896), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(n892), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[471]) );
  DFEC1 regs_reg_13__31_ ( .D(n924), .E(n967), .C(i_clk), .RN(n941), .Q(
        regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(n920), .E(n967), .C(i_clk), .RN(n936), .Q(
        regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(n916), .E(n967), .C(i_clk), .RN(n946), .Q(
        regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(n912), .E(n967), .C(i_clk), .RN(n945), .Q(
        regs[444]) );
  DFEC1 regs_reg_13__27_ ( .D(n908), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(n904), .E(n967), .C(i_clk), .RN(n942), .Q(
        regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(n900), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(n896), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(n892), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[439]) );
  DFEC1 regs_reg_12__31_ ( .D(n924), .E(n968), .C(i_clk), .RN(n937), .Q(
        regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(n920), .E(n968), .C(i_clk), .RN(n934), .Q(
        regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(n916), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(n912), .E(n968), .C(i_clk), .RN(n945), .Q(
        regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(n908), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(n904), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(n900), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(n896), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(n892), .E(n968), .C(i_clk), .RN(n945), .Q(
        regs[407]) );
  DFEC1 regs_reg_11__31_ ( .D(n924), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(n920), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(n916), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(n912), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(n908), .E(n969), .C(i_clk), .RN(n938), .Q(
        regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(n904), .E(n969), .C(i_clk), .RN(n946), .Q(
        regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(n900), .E(n969), .C(i_clk), .RN(n931), .Q(
        regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(n896), .E(n969), .C(i_clk), .RN(n940), .Q(
        regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(n892), .E(n969), .C(i_clk), .RN(n933), .Q(
        regs[375]) );
  DFEC1 regs_reg_10__31_ ( .D(n924), .E(n970), .C(i_clk), .RN(n937), .Q(
        regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(n920), .E(n970), .C(i_clk), .RN(n947), .Q(
        regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(n916), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(n912), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(n908), .E(n970), .C(i_clk), .RN(n936), .Q(
        regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(n904), .E(n970), .C(i_clk), .RN(n927), .Q(
        regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(n900), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(n896), .E(n970), .C(i_clk), .RN(n947), .Q(
        regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(n892), .E(n970), .C(i_clk), .RN(n946), .Q(
        regs[343]) );
  DFEC1 regs_reg_9__31_ ( .D(n924), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(n920), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(n916), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(n912), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(n908), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(n904), .E(n971), .C(i_clk), .RN(n946), .Q(
        regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(n900), .E(n971), .C(i_clk), .RN(n945), .Q(
        regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(n896), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(n892), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[311]) );
  DFEC1 regs_reg_8__31_ ( .D(n924), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(n920), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(n916), .E(n972), .C(i_clk), .RN(n943), .Q(
        regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(n912), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(n908), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(n904), .E(n972), .C(i_clk), .RN(n946), .Q(
        regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(n900), .E(n972), .C(i_clk), .RN(n945), .Q(
        regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(n896), .E(n972), .C(i_clk), .RN(n944), .Q(
        regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(n892), .E(n972), .C(i_clk), .RN(n927), .Q(
        regs[279]) );
  DFEC1 regs_reg_7__31_ ( .D(n923), .E(n973), .C(i_clk), .RN(n943), .Q(
        regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(n919), .E(n973), .C(i_clk), .RN(n937), .Q(
        regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(n915), .E(n973), .C(i_clk), .RN(n935), .Q(
        regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(n911), .E(n973), .C(i_clk), .RN(n930), .Q(
        regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(n907), .E(n973), .C(i_clk), .RN(n927), .Q(
        regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(n903), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(n899), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(n895), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(n891), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[247]) );
  DFEC1 regs_reg_6__31_ ( .D(n923), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(n919), .E(n974), .C(i_clk), .RN(n947), .Q(
        regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(n915), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(n911), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(n907), .E(n974), .C(i_clk), .RN(n940), .Q(
        regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(n903), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(n899), .E(n974), .C(i_clk), .RN(n933), .Q(
        regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(n895), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(n891), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[215]) );
  DFEC1 regs_reg_5__31_ ( .D(n923), .E(n975), .C(i_clk), .RN(n939), .Q(
        regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(n919), .E(n975), .C(i_clk), .RN(n930), .Q(
        regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(n915), .E(n975), .C(i_clk), .RN(n928), .Q(
        regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(n911), .E(n975), .C(i_clk), .RN(n929), .Q(
        regs[188]) );
  DFEC1 regs_reg_5__27_ ( .D(n907), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(n903), .E(n975), .C(i_clk), .RN(n943), .Q(
        regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(n899), .E(n975), .C(i_clk), .RN(n943), .Q(
        regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(n895), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(n891), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[183]) );
  DFEC1 regs_reg_4__31_ ( .D(n923), .E(n976), .C(i_clk), .RN(n939), .Q(
        regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(n919), .E(n976), .C(i_clk), .RN(n942), .Q(
        regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(n915), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(n911), .E(n976), .C(i_clk), .RN(n928), .Q(
        regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(n907), .E(n976), .C(i_clk), .RN(n935), .Q(
        regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(n903), .E(n976), .C(i_clk), .RN(n946), .Q(
        regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(n899), .E(n976), .C(i_clk), .RN(n945), .Q(
        regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(n895), .E(n976), .C(i_clk), .RN(n944), .Q(
        regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(n891), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[151]) );
  DFEC1 regs_reg_3__31_ ( .D(n923), .E(n977), .C(i_clk), .RN(n944), .Q(
        regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(n919), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(n915), .E(n977), .C(i_clk), .RN(n945), .Q(
        regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(n911), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(n907), .E(n977), .C(i_clk), .RN(n927), .Q(
        regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(n903), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(n899), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(n895), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(n891), .E(n977), .C(i_clk), .RN(n943), .Q(
        regs[119]) );
  DFEC1 regs_reg_2__31_ ( .D(n923), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(n919), .E(n978), .C(i_clk), .RN(n929), .Q(
        regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(n915), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(n911), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(n907), .E(n978), .C(i_clk), .RN(n929), .Q(
        regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(n903), .E(n978), .C(i_clk), .RN(n942), .Q(
        regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(n899), .E(n978), .C(i_clk), .RN(n930), .Q(
        regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(n895), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(n891), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[87]) );
  DFEC1 regs_reg_1__31_ ( .D(n923), .E(n979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(n919), .E(n979), .C(i_clk), .RN(n927), .Q(
        regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(n915), .E(n979), .C(i_clk), .RN(n944), .Q(
        regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(n911), .E(n979), .C(i_clk), .RN(n946), .Q(
        regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(n907), .E(n979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(n903), .E(n979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(n899), .E(n979), .C(i_clk), .RN(n942), .Q(
        regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(n895), .E(n979), .C(i_clk), .RN(n927), .Q(
        regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(n891), .E(n979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[55]) );
  DFEC1 regs_reg_0__31_ ( .D(n923), .E(n980), .C(i_clk), .RN(n942), .Q(
        regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(n919), .E(n980), .C(i_clk), .RN(n942), .Q(
        regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(n915), .E(n980), .C(i_clk), .RN(n942), .Q(
        regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(n911), .E(n980), .C(i_clk), .RN(n942), .Q(
        regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(n907), .E(n980), .C(i_clk), .RN(n942), .Q(
        regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(n903), .E(n980), .C(i_clk), .RN(n942), .Q(
        regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(n899), .E(n980), .C(i_clk), .RN(n942), .Q(
        regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(n895), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(n891), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[23]) );
  DFEC1 regs_reg_31__22_ ( .D(i_data_Rd[22]), .E(n958), .C(i_clk), .RN(n929), 
        .Q(regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(i_data_Rd[21]), .E(n958), .C(i_clk), .RN(n929), 
        .Q(regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(n884), .E(n958), .C(i_clk), .RN(n929), .Q(
        regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n958), .C(i_clk), .RN(n929), 
        .Q(regs[1011]) );
  DFEC1 regs_reg_31__17_ ( .D(i_data_Rd[17]), .E(n958), .C(i_clk), .RN(n929), 
        .Q(regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(i_data_Rd[16]), .E(n958), .C(i_clk), .RN(n929), 
        .Q(regs[1008]) );
  DFEC1 regs_reg_30__22_ ( .D(i_data_Rd[22]), .E(n959), .C(i_clk), .RN(n932), 
        .Q(regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(i_data_Rd[21]), .E(n959), .C(i_clk), .RN(n932), 
        .Q(regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(n884), .E(n959), .C(i_clk), .RN(n932), .Q(
        regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n959), .C(i_clk), .RN(n932), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__17_ ( .D(i_data_Rd[17]), .E(n959), .C(i_clk), .RN(n933), 
        .Q(regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(i_data_Rd[16]), .E(n959), .C(i_clk), .RN(n933), 
        .Q(regs[976]) );
  DFEC1 regs_reg_29__22_ ( .D(i_data_Rd[22]), .E(n960), .C(i_clk), .RN(n936), 
        .Q(regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(i_data_Rd[21]), .E(n960), .C(i_clk), .RN(n936), 
        .Q(regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(n884), .E(n960), .C(i_clk), .RN(n936), .Q(
        regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n960), .C(i_clk), .RN(n936), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__17_ ( .D(i_data_Rd[17]), .E(n960), .C(i_clk), .RN(n936), 
        .Q(regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(i_data_Rd[16]), .E(n960), .C(i_clk), .RN(n936), 
        .Q(regs[944]) );
  DFEC1 regs_reg_28__22_ ( .D(i_data_Rd[22]), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(i_data_Rd[21]), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(n884), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(
        regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n961), .C(i_clk), .RN(n939), 
        .Q(regs[915]) );
  DFEC1 regs_reg_28__17_ ( .D(i_data_Rd[17]), .E(n961), .C(i_clk), .RN(n939), 
        .Q(regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(i_data_Rd[16]), .E(n961), .C(i_clk), .RN(n939), 
        .Q(regs[912]) );
  DFEC1 regs_reg_27__22_ ( .D(i_data_Rd[22]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(i_data_Rd[21]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(n884), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__17_ ( .D(i_data_Rd[17]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(i_data_Rd[16]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[880]) );
  DFEC1 regs_reg_26__22_ ( .D(i_data_Rd[22]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(i_data_Rd[21]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(n884), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__17_ ( .D(i_data_Rd[17]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(i_data_Rd[16]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[848]) );
  DFEC1 regs_reg_25__22_ ( .D(i_data_Rd[22]), .E(n956), .C(i_clk), .RN(i_rst_n), .Q(regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(i_data_Rd[21]), .E(n956), .C(i_clk), .RN(i_rst_n), .Q(regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(n884), .E(n956), .C(i_clk), .RN(n946), .Q(
        regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(i_data_Rd[19]), .E(n956), .C(i_clk), .RN(i_rst_n), .Q(regs[819]) );
  DFEC1 regs_reg_25__17_ ( .D(i_data_Rd[17]), .E(n956), .C(i_clk), .RN(i_rst_n), .Q(regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(i_data_Rd[16]), .E(n956), .C(i_clk), .RN(i_rst_n), .Q(regs[816]) );
  DFEC1 regs_reg_24__22_ ( .D(i_data_Rd[22]), .E(n957), .C(i_clk), .RN(n945), 
        .Q(regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(i_data_Rd[21]), .E(n957), .C(i_clk), .RN(n936), 
        .Q(regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(n884), .E(n957), .C(i_clk), .RN(n928), .Q(
        regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(i_data_Rd[19]), .E(n957), .C(i_clk), .RN(n929), 
        .Q(regs[787]) );
  DFEC1 regs_reg_24__17_ ( .D(i_data_Rd[17]), .E(n957), .C(i_clk), .RN(n930), 
        .Q(regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(i_data_Rd[16]), .E(n957), .C(i_clk), .RN(n931), 
        .Q(regs[784]) );
  DFEC1 regs_reg_23__22_ ( .D(n890), .E(n948), .C(i_clk), .RN(n932), .Q(
        regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(n887), .E(n948), .C(i_clk), .RN(n933), .Q(
        regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(i_data_Rd[20]), .E(n948), .C(i_clk), .RN(n934), 
        .Q(regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(n881), .E(n948), .C(i_clk), .RN(n935), .Q(
        regs[755]) );
  DFEC1 regs_reg_23__17_ ( .D(n874), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(n871), .E(n948), .C(i_clk), .RN(n941), .Q(
        regs[752]) );
  DFEC1 regs_reg_22__22_ ( .D(n890), .E(n949), .C(i_clk), .RN(n939), .Q(
        regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(n887), .E(n949), .C(i_clk), .RN(n940), .Q(
        regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(i_data_Rd[20]), .E(n949), .C(i_clk), .RN(n941), 
        .Q(regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(n881), .E(n949), .C(i_clk), .RN(n942), .Q(
        regs[723]) );
  DFEC1 regs_reg_22__17_ ( .D(n874), .E(n949), .C(i_clk), .RN(n928), .Q(
        regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(n871), .E(n949), .C(i_clk), .RN(n929), .Q(
        regs[720]) );
  DFEC1 regs_reg_21__22_ ( .D(n890), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(n887), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(i_data_Rd[20]), .E(n950), .C(i_clk), .RN(n927), 
        .Q(regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(n881), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[691]) );
  DFEC1 regs_reg_21__17_ ( .D(n874), .E(n950), .C(i_clk), .RN(n937), .Q(
        regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(n871), .E(n950), .C(i_clk), .RN(n947), .Q(
        regs[688]) );
  DFEC1 regs_reg_20__22_ ( .D(n890), .E(n951), .C(i_clk), .RN(n941), .Q(
        regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(n887), .E(n951), .C(i_clk), .RN(n942), .Q(
        regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(i_data_Rd[20]), .E(n951), .C(i_clk), .RN(n928), 
        .Q(regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(n881), .E(n951), .C(i_clk), .RN(n929), .Q(
        regs[659]) );
  DFEC1 regs_reg_20__17_ ( .D(n874), .E(n951), .C(i_clk), .RN(n930), .Q(
        regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(n871), .E(n951), .C(i_clk), .RN(n931), .Q(
        regs[656]) );
  DFEC1 regs_reg_19__22_ ( .D(n890), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(n887), .E(n952), .C(i_clk), .RN(n938), .Q(
        regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(i_data_Rd[20]), .E(n952), .C(i_clk), .RN(n940), 
        .Q(regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(n881), .E(n952), .C(i_clk), .RN(n940), .Q(
        regs[627]) );
  DFEC1 regs_reg_19__17_ ( .D(n874), .E(n952), .C(i_clk), .RN(n939), .Q(
        regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(n871), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[624]) );
  DFEC1 regs_reg_18__22_ ( .D(n890), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(n887), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(i_data_Rd[20]), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(n881), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[595]) );
  DFEC1 regs_reg_18__17_ ( .D(n874), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(n871), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[592]) );
  DFEC1 regs_reg_17__22_ ( .D(n890), .E(n954), .C(i_clk), .RN(n937), .Q(
        regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(n887), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(i_data_Rd[20]), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(n881), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[563]) );
  DFEC1 regs_reg_17__17_ ( .D(n874), .E(n954), .C(i_clk), .RN(n940), .Q(
        regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(n871), .E(n954), .C(i_clk), .RN(n941), .Q(
        regs[560]) );
  DFEC1 regs_reg_16__22_ ( .D(n890), .E(n955), .C(i_clk), .RN(n945), .Q(
        regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(n887), .E(n955), .C(i_clk), .RN(n928), .Q(
        regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(i_data_Rd[20]), .E(n955), .C(i_clk), .RN(n929), 
        .Q(regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(n881), .E(n955), .C(i_clk), .RN(n930), .Q(
        regs[531]) );
  DFEC1 regs_reg_16__17_ ( .D(n874), .E(n955), .C(i_clk), .RN(n931), .Q(
        regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(n871), .E(n955), .C(i_clk), .RN(n944), .Q(
        regs[528]) );
  DFEC1 regs_reg_15__22_ ( .D(n889), .E(n965), .C(i_clk), .RN(n934), .Q(
        regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(n886), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(n883), .E(n965), .C(i_clk), .RN(n939), .Q(
        regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(n880), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[499]) );
  DFEC1 regs_reg_15__17_ ( .D(n873), .E(n965), .C(i_clk), .RN(n946), .Q(
        regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(n870), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[496]) );
  DFEC1 regs_reg_14__22_ ( .D(n889), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(n886), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(n883), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(n880), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[467]) );
  DFEC1 regs_reg_14__17_ ( .D(n873), .E(n966), .C(i_clk), .RN(n927), .Q(
        regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(n870), .E(n966), .C(i_clk), .RN(n943), .Q(
        regs[464]) );
  DFEC1 regs_reg_13__22_ ( .D(n889), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(n886), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(n883), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(n880), .E(n967), .C(i_clk), .RN(n935), .Q(
        regs[435]) );
  DFEC1 regs_reg_13__17_ ( .D(n873), .E(n967), .C(i_clk), .RN(n941), .Q(
        regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(n870), .E(n967), .C(i_clk), .RN(n937), .Q(
        regs[432]) );
  DFEC1 regs_reg_12__22_ ( .D(n889), .E(n968), .C(i_clk), .RN(n932), .Q(
        regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(n886), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(n883), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(n880), .E(n968), .C(i_clk), .RN(n940), .Q(
        regs[403]) );
  DFEC1 regs_reg_12__17_ ( .D(n873), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(n870), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[400]) );
  DFEC1 regs_reg_11__22_ ( .D(n889), .E(n969), .C(i_clk), .RN(n936), .Q(
        regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(n886), .E(n969), .C(i_clk), .RN(n945), .Q(
        regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(n883), .E(n969), .C(i_clk), .RN(n935), .Q(
        regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(n880), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[371]) );
  DFEC1 regs_reg_11__17_ ( .D(n873), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(n870), .E(n969), .C(i_clk), .RN(n932), .Q(
        regs[368]) );
  DFEC1 regs_reg_10__22_ ( .D(n889), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(n886), .E(n970), .C(i_clk), .RN(n934), .Q(
        regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(n883), .E(n970), .C(i_clk), .RN(n946), .Q(
        regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(n880), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[339]) );
  DFEC1 regs_reg_10__17_ ( .D(n873), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(n870), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[336]) );
  DFEC1 regs_reg_9__22_ ( .D(n889), .E(n971), .C(i_clk), .RN(n947), .Q(
        regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(n886), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(n883), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(n880), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[307]) );
  DFEC1 regs_reg_9__17_ ( .D(n873), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(n870), .E(n971), .C(i_clk), .RN(n934), .Q(
        regs[304]) );
  DFEC1 regs_reg_8__22_ ( .D(n889), .E(n972), .C(i_clk), .RN(n947), .Q(
        regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(n886), .E(n972), .C(i_clk), .RN(n947), .Q(
        regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(n883), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(n880), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[275]) );
  DFEC1 regs_reg_8__17_ ( .D(n873), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(n870), .E(n972), .C(i_clk), .RN(n946), .Q(
        regs[272]) );
  DFEC1 regs_reg_7__22_ ( .D(n888), .E(n973), .C(i_clk), .RN(n934), .Q(
        regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(n885), .E(n973), .C(i_clk), .RN(n930), .Q(
        regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(n882), .E(n973), .C(i_clk), .RN(n944), .Q(
        regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(n879), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[243]) );
  DFEC1 regs_reg_7__17_ ( .D(n872), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(n869), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[240]) );
  DFEC1 regs_reg_6__22_ ( .D(n888), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(n885), .E(n974), .C(i_clk), .RN(n944), .Q(
        regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(n882), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(n879), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[211]) );
  DFEC1 regs_reg_6__17_ ( .D(n872), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(n869), .E(n974), .C(i_clk), .RN(n936), .Q(
        regs[208]) );
  DFEC1 regs_reg_5__22_ ( .D(n888), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(n885), .E(n975), .C(i_clk), .RN(n930), .Q(
        regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(n882), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(n879), .E(n975), .C(i_clk), .RN(n947), .Q(
        regs[179]) );
  DFEC1 regs_reg_5__17_ ( .D(n872), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(n869), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[176]) );
  DFEC1 regs_reg_4__22_ ( .D(n888), .E(n976), .C(i_clk), .RN(n946), .Q(
        regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(n885), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(n882), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(n879), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[147]) );
  DFEC1 regs_reg_4__17_ ( .D(n872), .E(n976), .C(i_clk), .RN(n932), .Q(
        regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(n869), .E(n976), .C(i_clk), .RN(n935), .Q(
        regs[144]) );
  DFEC1 regs_reg_3__22_ ( .D(n888), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(n885), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(n882), .E(n977), .C(i_clk), .RN(n945), .Q(
        regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(n879), .E(n977), .C(i_clk), .RN(n943), .Q(
        regs[115]) );
  DFEC1 regs_reg_3__17_ ( .D(n872), .E(n977), .C(i_clk), .RN(n946), .Q(
        regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(n869), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[112]) );
  DFEC1 regs_reg_2__22_ ( .D(n888), .E(n978), .C(i_clk), .RN(n938), .Q(
        regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(n885), .E(n978), .C(i_clk), .RN(n943), .Q(
        regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(n882), .E(n978), .C(i_clk), .RN(n941), .Q(
        regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(n879), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[83]) );
  DFEC1 regs_reg_2__17_ ( .D(n872), .E(n978), .C(i_clk), .RN(n927), .Q(
        regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(n869), .E(n978), .C(i_clk), .RN(n943), .Q(
        regs[80]) );
  DFEC1 regs_reg_1__22_ ( .D(n888), .E(n979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(n885), .E(n979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(n882), .E(n979), .C(i_clk), .RN(n928), .Q(
        regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(n879), .E(n979), .C(i_clk), .RN(n940), .Q(
        regs[51]) );
  DFEC1 regs_reg_1__17_ ( .D(n872), .E(n979), .C(i_clk), .RN(n940), .Q(
        regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(n869), .E(n979), .C(i_clk), .RN(n940), .Q(
        regs[48]) );
  DFEC1 regs_reg_0__22_ ( .D(n888), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(n885), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(n882), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(n879), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[19]) );
  DFEC1 regs_reg_0__17_ ( .D(n872), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(n869), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[16]) );
  DFEC1 regs_reg_31__18_ ( .D(n878), .E(n958), .C(i_clk), .RN(n929), .Q(
        regs[1010]) );
  DFEC1 regs_reg_30__18_ ( .D(n878), .E(n959), .C(i_clk), .RN(n933), .Q(
        regs[978]) );
  DFEC1 regs_reg_29__18_ ( .D(n878), .E(n960), .C(i_clk), .RN(n936), .Q(
        regs[946]) );
  DFEC1 regs_reg_28__18_ ( .D(n878), .E(n961), .C(i_clk), .RN(n939), .Q(
        regs[914]) );
  DFEC1 regs_reg_27__18_ ( .D(n878), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[882]) );
  DFEC1 regs_reg_26__18_ ( .D(n878), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[850]) );
  DFEC1 regs_reg_25__18_ ( .D(n878), .E(n956), .C(i_clk), .RN(n947), .Q(
        regs[818]) );
  DFEC1 regs_reg_24__18_ ( .D(n878), .E(n957), .C(i_clk), .RN(n932), .Q(
        regs[786]) );
  DFEC1 regs_reg_23__18_ ( .D(n877), .E(n948), .C(i_clk), .RN(n936), .Q(
        regs[754]) );
  DFEC1 regs_reg_22__18_ ( .D(n877), .E(n949), .C(i_clk), .RN(n930), .Q(
        regs[722]) );
  DFEC1 regs_reg_21__18_ ( .D(n877), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[690]) );
  DFEC1 regs_reg_20__18_ ( .D(n877), .E(n951), .C(i_clk), .RN(n932), .Q(
        regs[658]) );
  DFEC1 regs_reg_19__18_ ( .D(n877), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[626]) );
  DFEC1 regs_reg_18__18_ ( .D(n877), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[594]) );
  DFEC1 regs_reg_17__18_ ( .D(n877), .E(n954), .C(i_clk), .RN(n942), .Q(
        regs[562]) );
  DFEC1 regs_reg_16__18_ ( .D(n877), .E(n955), .C(i_clk), .RN(n932), .Q(
        regs[530]) );
  DFEC1 regs_reg_15__18_ ( .D(n876), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[498]) );
  DFEC1 regs_reg_14__18_ ( .D(n876), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[466]) );
  DFEC1 regs_reg_13__18_ ( .D(n876), .E(n967), .C(i_clk), .RN(n942), .Q(
        regs[434]) );
  DFEC1 regs_reg_12__18_ ( .D(n876), .E(n968), .C(i_clk), .RN(n934), .Q(
        regs[402]) );
  DFEC1 regs_reg_11__18_ ( .D(n876), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[370]) );
  DFEC1 regs_reg_10__18_ ( .D(n876), .E(n970), .C(i_clk), .RN(n947), .Q(
        regs[338]) );
  DFEC1 regs_reg_9__18_ ( .D(n876), .E(n971), .C(i_clk), .RN(n944), .Q(
        regs[306]) );
  DFEC1 regs_reg_8__18_ ( .D(n876), .E(n972), .C(i_clk), .RN(n945), .Q(
        regs[274]) );
  DFEC1 regs_reg_7__18_ ( .D(n875), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[242]) );
  DFEC1 regs_reg_6__18_ ( .D(n875), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[210]) );
  DFEC1 regs_reg_5__18_ ( .D(n875), .E(n975), .C(i_clk), .RN(n937), .Q(
        regs[178]) );
  DFEC1 regs_reg_4__18_ ( .D(n875), .E(n976), .C(i_clk), .RN(n928), .Q(
        regs[146]) );
  DFEC1 regs_reg_3__18_ ( .D(n875), .E(n977), .C(i_clk), .RN(n946), .Q(
        regs[114]) );
  DFEC1 regs_reg_2__18_ ( .D(n875), .E(n978), .C(i_clk), .RN(n943), .Q(
        regs[82]) );
  DFEC1 regs_reg_1__18_ ( .D(n875), .E(n979), .C(i_clk), .RN(n940), .Q(
        regs[50]) );
  DFEC1 regs_reg_0__18_ ( .D(n875), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[18]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n958), .C(i_clk), .RN(n930), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(i_data_Rd[5]), .E(n958), .C(i_clk), .RN(n930), 
        .Q(regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(i_data_Rd[4]), .E(n958), .C(i_clk), .RN(n931), 
        .Q(regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(i_data_Rd[3]), .E(n958), .C(i_clk), .RN(n931), 
        .Q(regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(i_data_Rd[2]), .E(n958), .C(i_clk), .RN(n931), 
        .Q(regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n958), .C(i_clk), .RN(n931), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(i_data_Rd[0]), .E(n958), .C(i_clk), .RN(n931), 
        .Q(regs[992]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n959), .C(i_clk), .RN(n934), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(i_data_Rd[5]), .E(n959), .C(i_clk), .RN(n934), 
        .Q(regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(i_data_Rd[4]), .E(n959), .C(i_clk), .RN(n934), 
        .Q(regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(i_data_Rd[3]), .E(n959), .C(i_clk), .RN(n934), 
        .Q(regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(i_data_Rd[2]), .E(n959), .C(i_clk), .RN(n934), 
        .Q(regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n959), .C(i_clk), .RN(n934), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(i_data_Rd[0]), .E(n959), .C(i_clk), .RN(n935), 
        .Q(regs[960]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n960), .C(i_clk), .RN(n937), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(i_data_Rd[5]), .E(n960), .C(i_clk), .RN(n938), 
        .Q(regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(i_data_Rd[4]), .E(n960), .C(i_clk), .RN(n938), 
        .Q(regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(i_data_Rd[3]), .E(n960), .C(i_clk), .RN(n938), 
        .Q(regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(i_data_Rd[2]), .E(n960), .C(i_clk), .RN(n938), 
        .Q(regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n960), .C(i_clk), .RN(n938), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(i_data_Rd[0]), .E(n960), .C(i_clk), .RN(n938), 
        .Q(regs[928]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n961), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(i_data_Rd[5]), .E(n961), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(i_data_Rd[4]), .E(n961), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(i_data_Rd[3]), .E(n961), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(i_data_Rd[2]), .E(n961), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n961), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(i_data_Rd[0]), .E(n961), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[896]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(i_data_Rd[5]), .E(n962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(i_data_Rd[4]), .E(n962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(i_data_Rd[3]), .E(n962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(i_data_Rd[2]), .E(n962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(i_data_Rd[1]), .E(n962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(i_data_Rd[0]), .E(n962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[864]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(i_data_Rd[5]), .E(n963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(i_data_Rd[4]), .E(n963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(i_data_Rd[3]), .E(n963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(i_data_Rd[2]), .E(n963), .C(i_clk), .RN(n932), 
        .Q(regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n963), .C(i_clk), .RN(n933), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(i_data_Rd[0]), .E(n963), .C(i_clk), .RN(n937), 
        .Q(regs[832]) );
  DFEC1 regs_reg_25__6_ ( .D(i_data_Rd[6]), .E(n956), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(i_data_Rd[5]), .E(n956), .C(i_clk), .RN(n928), 
        .Q(regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(i_data_Rd[4]), .E(n956), .C(i_clk), .RN(n929), 
        .Q(regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(i_data_Rd[3]), .E(n956), .C(i_clk), .RN(n940), 
        .Q(regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(i_data_Rd[2]), .E(n956), .C(i_clk), .RN(n941), 
        .Q(regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(i_data_Rd[1]), .E(n956), .C(i_clk), .RN(n942), 
        .Q(regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(i_data_Rd[0]), .E(n956), .C(i_clk), .RN(n939), 
        .Q(regs[800]) );
  DFEC1 regs_reg_24__6_ ( .D(i_data_Rd[6]), .E(n957), .C(i_clk), .RN(n928), 
        .Q(regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(i_data_Rd[5]), .E(n957), .C(i_clk), .RN(n929), 
        .Q(regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(i_data_Rd[4]), .E(n957), .C(i_clk), .RN(n930), 
        .Q(regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(i_data_Rd[3]), .E(n957), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(i_data_Rd[2]), .E(n957), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(i_data_Rd[1]), .E(n957), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(i_data_Rd[0]), .E(n957), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[768]) );
  DFEC1 regs_reg_23__6_ ( .D(n840), .E(n948), .C(i_clk), .RN(n943), .Q(
        regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(n837), .E(n948), .C(i_clk), .RN(n946), .Q(
        regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(n834), .E(n948), .C(i_clk), .RN(n945), .Q(
        regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(n831), .E(n948), .C(i_clk), .RN(n944), .Q(
        regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(n828), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(n825), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(n822), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[736]) );
  DFEC1 regs_reg_22__6_ ( .D(n840), .E(n949), .C(i_clk), .RN(i_rst_n), .Q(
        regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(n837), .E(n949), .C(i_clk), .RN(n947), .Q(
        regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(n834), .E(n949), .C(i_clk), .RN(n937), .Q(
        regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(n831), .E(n949), .C(i_clk), .RN(n938), .Q(
        regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(n828), .E(n949), .C(i_clk), .RN(i_rst_n), .Q(
        regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(n825), .E(n949), .C(i_clk), .RN(i_rst_n), .Q(
        regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(n822), .E(n949), .C(i_clk), .RN(i_rst_n), .Q(
        regs[704]) );
  DFEC1 regs_reg_21__6_ ( .D(n840), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(n837), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(n834), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(n831), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(n828), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(n825), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(n822), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[672]) );
  DFEC1 regs_reg_20__6_ ( .D(n840), .E(n951), .C(i_clk), .RN(n938), .Q(
        regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(n837), .E(n951), .C(i_clk), .RN(n930), .Q(
        regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(n834), .E(n951), .C(i_clk), .RN(n931), .Q(
        regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(n831), .E(n951), .C(i_clk), .RN(n932), .Q(
        regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(n828), .E(n951), .C(i_clk), .RN(n933), .Q(
        regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(n825), .E(n951), .C(i_clk), .RN(n934), .Q(
        regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(n822), .E(n951), .C(i_clk), .RN(n935), .Q(
        regs[640]) );
  DFEC1 regs_reg_19__6_ ( .D(n840), .E(n952), .C(i_clk), .RN(n943), .Q(
        regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(n837), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(n834), .E(n952), .C(i_clk), .RN(n946), .Q(
        regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(n831), .E(n952), .C(i_clk), .RN(n945), .Q(
        regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(n828), .E(n952), .C(i_clk), .RN(n944), .Q(
        regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(n825), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(n822), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[608]) );
  DFEC1 regs_reg_18__6_ ( .D(n840), .E(n953), .C(i_clk), .RN(n930), .Q(
        regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(n837), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(n834), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(n831), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(n828), .E(n953), .C(i_clk), .RN(n936), .Q(
        regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(n825), .E(n953), .C(i_clk), .RN(n941), .Q(
        regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(n822), .E(n953), .C(i_clk), .RN(n947), .Q(
        regs[576]) );
  DFEC1 regs_reg_17__6_ ( .D(n840), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(n837), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(n834), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(n831), .E(n954), .C(i_clk), .RN(n940), .Q(
        regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(n828), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(n825), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(n822), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[544]) );
  DFEC1 regs_reg_16__6_ ( .D(n840), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(n837), .E(n955), .C(i_clk), .RN(n947), .Q(
        regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(n834), .E(n955), .C(i_clk), .RN(n943), .Q(
        regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(n831), .E(n955), .C(i_clk), .RN(n947), .Q(
        regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(n828), .E(n955), .C(i_clk), .RN(n935), .Q(
        regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(n825), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(n822), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[512]) );
  DFEC1 regs_reg_15__6_ ( .D(n839), .E(n965), .C(i_clk), .RN(n928), .Q(
        regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(n836), .E(n965), .C(i_clk), .RN(n929), .Q(
        regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(n833), .E(n965), .C(i_clk), .RN(n930), .Q(
        regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(n830), .E(n965), .C(i_clk), .RN(n927), .Q(
        regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(n827), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(n824), .E(n965), .C(i_clk), .RN(n934), .Q(
        regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(n821), .E(n965), .C(i_clk), .RN(n936), .Q(
        regs[480]) );
  DFEC1 regs_reg_14__6_ ( .D(n839), .E(n966), .C(i_clk), .RN(n945), .Q(
        regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(n836), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(n833), .E(n966), .C(i_clk), .RN(n935), .Q(
        regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(n830), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(n827), .E(n966), .C(i_clk), .RN(n945), .Q(
        regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(n824), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(n821), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[448]) );
  DFEC1 regs_reg_13__6_ ( .D(n839), .E(n967), .C(i_clk), .RN(n932), .Q(
        regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(n836), .E(n967), .C(i_clk), .RN(n938), .Q(
        regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(n833), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(n830), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(n827), .E(n967), .C(i_clk), .RN(n938), .Q(
        regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(n824), .E(n967), .C(i_clk), .RN(n943), .Q(
        regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(n821), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[416]) );
  DFEC1 regs_reg_12__6_ ( .D(n839), .E(n968), .C(i_clk), .RN(n942), .Q(
        regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(n836), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(n833), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(n830), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(n827), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(n824), .E(n968), .C(i_clk), .RN(n944), .Q(
        regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(n821), .E(n968), .C(i_clk), .RN(n941), .Q(
        regs[384]) );
  DFEC1 regs_reg_11__6_ ( .D(n839), .E(n969), .C(i_clk), .RN(n943), .Q(
        regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(n836), .E(n969), .C(i_clk), .RN(n933), .Q(
        regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(n833), .E(n969), .C(i_clk), .RN(n938), .Q(
        regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(n830), .E(n969), .C(i_clk), .RN(n946), .Q(
        regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(n827), .E(n969), .C(i_clk), .RN(n938), .Q(
        regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(n824), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(n821), .E(n969), .C(i_clk), .RN(n937), .Q(
        regs[352]) );
  DFEC1 regs_reg_10__6_ ( .D(n839), .E(n970), .C(i_clk), .RN(n946), .Q(
        regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(n836), .E(n970), .C(i_clk), .RN(n941), .Q(
        regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(n833), .E(n970), .C(i_clk), .RN(n939), .Q(
        regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(n830), .E(n970), .C(i_clk), .RN(n937), .Q(
        regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(n827), .E(n970), .C(i_clk), .RN(n927), .Q(
        regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(n824), .E(n970), .C(i_clk), .RN(n944), .Q(
        regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(n821), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[320]) );
  DFEC1 regs_reg_9__6_ ( .D(n839), .E(n971), .C(i_clk), .RN(n931), .Q(
        regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(n836), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(n833), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(n830), .E(n971), .C(i_clk), .RN(n940), .Q(
        regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(n827), .E(n971), .C(i_clk), .RN(n933), .Q(
        regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(n824), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(n821), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[288]) );
  DFEC1 regs_reg_8__6_ ( .D(n839), .E(n972), .C(i_clk), .RN(n944), .Q(
        regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(n836), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(n833), .E(n972), .C(i_clk), .RN(n931), .Q(
        regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(n830), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(n827), .E(n972), .C(i_clk), .RN(n927), .Q(
        regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(n824), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(n821), .E(n972), .C(i_clk), .RN(n937), .Q(
        regs[256]) );
  DFEC1 regs_reg_7__6_ ( .D(n838), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(n835), .E(n973), .C(i_clk), .RN(n943), .Q(
        regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(n832), .E(n973), .C(i_clk), .RN(n933), .Q(
        regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(n829), .E(n973), .C(i_clk), .RN(n927), .Q(
        regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(n826), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(n823), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(n820), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[224]) );
  DFEC1 regs_reg_6__6_ ( .D(n838), .E(n974), .C(i_clk), .RN(n945), .Q(
        regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(n835), .E(n974), .C(i_clk), .RN(n941), .Q(
        regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(n832), .E(n974), .C(i_clk), .RN(n942), .Q(
        regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(n829), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(n826), .E(n974), .C(i_clk), .RN(n933), .Q(
        regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(n823), .E(n974), .C(i_clk), .RN(n940), .Q(
        regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(n820), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[192]) );
  DFEC1 regs_reg_5__6_ ( .D(n838), .E(n975), .C(i_clk), .RN(n931), .Q(
        regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(n835), .E(n975), .C(i_clk), .RN(n929), .Q(
        regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(n832), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(n829), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(n826), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(n823), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(n820), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[160]) );
  DFEC1 regs_reg_4__6_ ( .D(n838), .E(n976), .C(i_clk), .RN(n938), .Q(
        regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(n835), .E(n976), .C(i_clk), .RN(n927), .Q(
        regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(n832), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(n829), .E(n976), .C(i_clk), .RN(n939), .Q(
        regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(n826), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(n823), .E(n976), .C(i_clk), .RN(n942), .Q(
        regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(n820), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[128]) );
  DFEC1 regs_reg_3__6_ ( .D(n838), .E(n977), .C(i_clk), .RN(n931), .Q(
        regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(n835), .E(n977), .C(i_clk), .RN(n941), .Q(
        regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(n832), .E(n977), .C(i_clk), .RN(n939), .Q(
        regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(n829), .E(n977), .C(i_clk), .RN(n947), .Q(regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(n826), .E(n977), .C(i_clk), .RN(n947), .Q(regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(n823), .E(n977), .C(i_clk), .RN(n941), .Q(regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(n820), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[96]) );
  DFEC1 regs_reg_2__6_ ( .D(n838), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(n835), .E(n978), .C(i_clk), .RN(n937), .Q(regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(n832), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(n829), .E(n978), .C(i_clk), .RN(n936), .Q(regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(n826), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(n823), .E(n978), .C(i_clk), .RN(n934), .Q(regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(n820), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[64]) );
  DFEC1 regs_reg_1__6_ ( .D(n838), .E(n979), .C(i_clk), .RN(n941), .Q(regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(n835), .E(n979), .C(i_clk), .RN(n941), .Q(regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(n832), .E(n979), .C(i_clk), .RN(n941), .Q(regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(n829), .E(n979), .C(i_clk), .RN(n941), .Q(regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(n826), .E(n979), .C(i_clk), .RN(n941), .Q(regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(n823), .E(n979), .C(i_clk), .RN(n942), .Q(regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(n820), .E(n979), .C(i_clk), .RN(n942), .Q(regs[32]) );
  DFEC1 regs_reg_0__6_ ( .D(n838), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(n835), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(n832), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(n829), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(n826), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(n823), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(n820), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[0]) );
  DFEC1 regs_reg_31__9_ ( .D(i_data_Rd[9]), .E(n958), .C(i_clk), .RN(n930), 
        .Q(regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(i_data_Rd[8]), .E(n958), .C(i_clk), .RN(n930), 
        .Q(regs[1000]) );
  DFEC1 regs_reg_30__9_ ( .D(i_data_Rd[9]), .E(n959), .C(i_clk), .RN(n934), 
        .Q(regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(i_data_Rd[8]), .E(n959), .C(i_clk), .RN(n934), 
        .Q(regs[968]) );
  DFEC1 regs_reg_29__9_ ( .D(i_data_Rd[9]), .E(n960), .C(i_clk), .RN(n937), 
        .Q(regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(i_data_Rd[8]), .E(n960), .C(i_clk), .RN(n937), 
        .Q(regs[936]) );
  DFEC1 regs_reg_28__9_ ( .D(i_data_Rd[9]), .E(n961), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(i_data_Rd[8]), .E(n961), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[904]) );
  DFEC1 regs_reg_27__9_ ( .D(i_data_Rd[9]), .E(n962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(i_data_Rd[8]), .E(n962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[872]) );
  DFEC1 regs_reg_26__9_ ( .D(i_data_Rd[9]), .E(n963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(i_data_Rd[8]), .E(n963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[840]) );
  DFEC1 regs_reg_25__9_ ( .D(i_data_Rd[9]), .E(n956), .C(i_clk), .RN(n944), 
        .Q(regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(i_data_Rd[8]), .E(n956), .C(i_clk), .RN(n941), 
        .Q(regs[808]) );
  DFEC1 regs_reg_24__9_ ( .D(i_data_Rd[9]), .E(n957), .C(i_clk), .RN(n931), 
        .Q(regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(i_data_Rd[8]), .E(n957), .C(i_clk), .RN(n932), 
        .Q(regs[776]) );
  DFEC1 regs_reg_23__9_ ( .D(n850), .E(n948), .C(i_clk), .RN(n943), .Q(
        regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(n847), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[744]) );
  DFEC1 regs_reg_22__9_ ( .D(n850), .E(n949), .C(i_clk), .RN(i_rst_n), .Q(
        regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(n847), .E(n949), .C(i_clk), .RN(n944), .Q(
        regs[712]) );
  DFEC1 regs_reg_21__9_ ( .D(n850), .E(n950), .C(i_clk), .RN(n939), .Q(
        regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(n847), .E(n950), .C(i_clk), .RN(n940), .Q(
        regs[680]) );
  DFEC1 regs_reg_20__9_ ( .D(n850), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(n847), .E(n951), .C(i_clk), .RN(n939), .Q(
        regs[648]) );
  DFEC1 regs_reg_19__9_ ( .D(n850), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(n847), .E(n952), .C(i_clk), .RN(n928), .Q(
        regs[616]) );
  DFEC1 regs_reg_18__9_ ( .D(n850), .E(n953), .C(i_clk), .RN(n938), .Q(
        regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(n847), .E(n953), .C(i_clk), .RN(n936), .Q(
        regs[584]) );
  DFEC1 regs_reg_17__9_ ( .D(n850), .E(n954), .C(i_clk), .RN(n944), .Q(
        regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(n847), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[552]) );
  DFEC1 regs_reg_16__9_ ( .D(n850), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(n847), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[520]) );
  DFEC1 regs_reg_15__9_ ( .D(n849), .E(n965), .C(i_clk), .RN(n931), .Q(
        regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(n846), .E(n965), .C(i_clk), .RN(n932), .Q(
        regs[488]) );
  DFEC1 regs_reg_14__9_ ( .D(n849), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(n846), .E(n966), .C(i_clk), .RN(n933), .Q(
        regs[456]) );
  DFEC1 regs_reg_13__9_ ( .D(n849), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(n846), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[424]) );
  DFEC1 regs_reg_12__9_ ( .D(n849), .E(n968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(n846), .E(n968), .C(i_clk), .RN(n942), .Q(
        regs[392]) );
  DFEC1 regs_reg_11__9_ ( .D(n849), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(n846), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[360]) );
  DFEC1 regs_reg_10__9_ ( .D(n849), .E(n970), .C(i_clk), .RN(n941), .Q(
        regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(n846), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[328]) );
  DFEC1 regs_reg_9__9_ ( .D(n849), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(n846), .E(n971), .C(i_clk), .RN(n944), .Q(
        regs[296]) );
  DFEC1 regs_reg_8__9_ ( .D(n849), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(n846), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[264]) );
  DFEC1 regs_reg_7__9_ ( .D(n848), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(n845), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[232]) );
  DFEC1 regs_reg_6__9_ ( .D(n848), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(n845), .E(n974), .C(i_clk), .RN(n946), .Q(
        regs[200]) );
  DFEC1 regs_reg_5__9_ ( .D(n848), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(n845), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[168]) );
  DFEC1 regs_reg_4__9_ ( .D(n848), .E(n976), .C(i_clk), .RN(n940), .Q(
        regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(n845), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[136]) );
  DFEC1 regs_reg_3__9_ ( .D(n848), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(n845), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[104]) );
  DFEC1 regs_reg_2__9_ ( .D(n848), .E(n978), .C(i_clk), .RN(n938), .Q(regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(n845), .E(n978), .C(i_clk), .RN(n937), .Q(regs[72]) );
  DFEC1 regs_reg_1__9_ ( .D(n848), .E(n979), .C(i_clk), .RN(n941), .Q(regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(n845), .E(n979), .C(i_clk), .RN(n941), .Q(regs[40]) );
  DFEC1 regs_reg_0__9_ ( .D(n848), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(n845), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[8]) );
  DFEC1 regs_reg_31__15_ ( .D(i_data_Rd[15]), .E(n958), .C(i_clk), .RN(n929), 
        .Q(regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(i_data_Rd[14]), .E(n958), .C(i_clk), .RN(n929), 
        .Q(regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(i_data_Rd[13]), .E(n958), .C(i_clk), .RN(n930), 
        .Q(regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(i_data_Rd[12]), .E(n958), .C(i_clk), .RN(n930), 
        .Q(regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(i_data_Rd[11]), .E(n958), .C(i_clk), .RN(n930), 
        .Q(regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(n853), .E(n958), .C(i_clk), .RN(n930), .Q(
        regs[1002]) );
  DFEC1 regs_reg_30__15_ ( .D(i_data_Rd[15]), .E(n959), .C(i_clk), .RN(n933), 
        .Q(regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(i_data_Rd[14]), .E(n959), .C(i_clk), .RN(n933), 
        .Q(regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(i_data_Rd[13]), .E(n959), .C(i_clk), .RN(n933), 
        .Q(regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(i_data_Rd[12]), .E(n959), .C(i_clk), .RN(n933), 
        .Q(regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(i_data_Rd[11]), .E(n959), .C(i_clk), .RN(n933), 
        .Q(regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(n853), .E(n959), .C(i_clk), .RN(n933), .Q(
        regs[970]) );
  DFEC1 regs_reg_29__15_ ( .D(i_data_Rd[15]), .E(n960), .C(i_clk), .RN(n936), 
        .Q(regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(i_data_Rd[14]), .E(n960), .C(i_clk), .RN(n937), 
        .Q(regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(i_data_Rd[13]), .E(n960), .C(i_clk), .RN(n937), 
        .Q(regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(i_data_Rd[12]), .E(n960), .C(i_clk), .RN(n937), 
        .Q(regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(i_data_Rd[11]), .E(n960), .C(i_clk), .RN(n937), 
        .Q(regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(n853), .E(n960), .C(i_clk), .RN(n937), .Q(
        regs[938]) );
  DFEC1 regs_reg_28__15_ ( .D(i_data_Rd[15]), .E(n961), .C(i_clk), .RN(n939), 
        .Q(regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(i_data_Rd[14]), .E(n961), .C(i_clk), .RN(n939), 
        .Q(regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(i_data_Rd[13]), .E(n961), .C(i_clk), .RN(n939), 
        .Q(regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(i_data_Rd[12]), .E(n961), .C(i_clk), .RN(n939), 
        .Q(regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(i_data_Rd[11]), .E(n961), .C(i_clk), .RN(n939), 
        .Q(regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(n853), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(
        regs[906]) );
  DFEC1 regs_reg_27__15_ ( .D(i_data_Rd[15]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(i_data_Rd[14]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(i_data_Rd[13]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(i_data_Rd[12]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(i_data_Rd[11]), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(n853), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[874]) );
  DFEC1 regs_reg_26__15_ ( .D(i_data_Rd[15]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(i_data_Rd[14]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(i_data_Rd[13]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(i_data_Rd[12]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(i_data_Rd[11]), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(n853), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[842]) );
  DFEC1 regs_reg_25__15_ ( .D(i_data_Rd[15]), .E(n956), .C(i_clk), .RN(n934), 
        .Q(regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(i_data_Rd[14]), .E(n956), .C(i_clk), .RN(n935), 
        .Q(regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(i_data_Rd[13]), .E(n956), .C(i_clk), .RN(n936), 
        .Q(regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(i_data_Rd[12]), .E(n956), .C(i_clk), .RN(n928), 
        .Q(regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(i_data_Rd[11]), .E(n956), .C(i_clk), .RN(n929), 
        .Q(regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(n853), .E(n956), .C(i_clk), .RN(n930), .Q(
        regs[810]) );
  DFEC1 regs_reg_24__15_ ( .D(i_data_Rd[15]), .E(n957), .C(i_clk), .RN(n933), 
        .Q(regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(i_data_Rd[14]), .E(n957), .C(i_clk), .RN(n937), 
        .Q(regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(i_data_Rd[13]), .E(n957), .C(i_clk), .RN(n938), 
        .Q(regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(i_data_Rd[12]), .E(n957), .C(i_clk), .RN(n933), 
        .Q(regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(i_data_Rd[11]), .E(n957), .C(i_clk), .RN(n937), 
        .Q(regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(n853), .E(n957), .C(i_clk), .RN(n938), .Q(
        regs[778]) );
  DFEC1 regs_reg_23__15_ ( .D(n868), .E(n948), .C(i_clk), .RN(n941), .Q(
        regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(n865), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(n862), .E(n948), .C(i_clk), .RN(n939), .Q(
        regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(n859), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(n856), .E(n948), .C(i_clk), .RN(n944), .Q(
        regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(n852), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[746]) );
  DFEC1 regs_reg_22__15_ ( .D(n868), .E(n949), .C(i_clk), .RN(n931), .Q(
        regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(n865), .E(n949), .C(i_clk), .RN(n932), .Q(
        regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(n862), .E(n949), .C(i_clk), .RN(n934), .Q(
        regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(n859), .E(n949), .C(i_clk), .RN(n946), .Q(
        regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(n856), .E(n949), .C(i_clk), .RN(n945), .Q(
        regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(n852), .E(n949), .C(i_clk), .RN(n944), .Q(
        regs[714]) );
  DFEC1 regs_reg_21__15_ ( .D(n868), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(n865), .E(n950), .C(i_clk), .RN(n945), .Q(
        regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(n862), .E(n950), .C(i_clk), .RN(n936), .Q(
        regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(n859), .E(n950), .C(i_clk), .RN(n943), .Q(
        regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(n856), .E(n950), .C(i_clk), .RN(n946), .Q(
        regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(n852), .E(n950), .C(i_clk), .RN(n945), .Q(
        regs[682]) );
  DFEC1 regs_reg_20__15_ ( .D(n868), .E(n951), .C(i_clk), .RN(n933), .Q(
        regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(n865), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(n862), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(n859), .E(n951), .C(i_clk), .RN(n927), .Q(
        regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(n856), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(n852), .E(n951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[650]) );
  DFEC1 regs_reg_19__15_ ( .D(n868), .E(n952), .C(i_clk), .RN(n947), .Q(
        regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(n865), .E(n952), .C(i_clk), .RN(n927), .Q(
        regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(n862), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(n859), .E(n952), .C(i_clk), .RN(n928), .Q(
        regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(n856), .E(n952), .C(i_clk), .RN(n944), .Q(
        regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(n852), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[618]) );
  DFEC1 regs_reg_18__15_ ( .D(n868), .E(n953), .C(i_clk), .RN(n944), .Q(
        regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(n865), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(n862), .E(n953), .C(i_clk), .RN(n946), .Q(
        regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(n859), .E(n953), .C(i_clk), .RN(n945), .Q(
        regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(n856), .E(n953), .C(i_clk), .RN(n944), .Q(
        regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(n852), .E(n953), .C(i_clk), .RN(n947), .Q(
        regs[586]) );
  DFEC1 regs_reg_17__15_ ( .D(n868), .E(n954), .C(i_clk), .RN(n947), .Q(
        regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(n865), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(n862), .E(n954), .C(i_clk), .RN(n933), .Q(
        regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(n859), .E(n954), .C(i_clk), .RN(n943), .Q(
        regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(n856), .E(n954), .C(i_clk), .RN(n941), .Q(
        regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(n852), .E(n954), .C(i_clk), .RN(n927), .Q(
        regs[554]) );
  DFEC1 regs_reg_16__15_ ( .D(n868), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(n865), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(n862), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(n859), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(n856), .E(n955), .C(i_clk), .RN(n940), .Q(
        regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(n852), .E(n955), .C(i_clk), .RN(n938), .Q(
        regs[522]) );
  DFEC1 regs_reg_15__15_ ( .D(n867), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(n864), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(n861), .E(n965), .C(i_clk), .RN(i_rst_n), .Q(
        regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(n858), .E(n965), .C(i_clk), .RN(n933), .Q(
        regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(n855), .E(n965), .C(i_clk), .RN(n934), .Q(
        regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n965), .C(i_clk), .RN(n935), 
        .Q(regs[490]) );
  DFEC1 regs_reg_14__15_ ( .D(n867), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(n864), .E(n966), .C(i_clk), .RN(n943), .Q(
        regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(n861), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(n858), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(n855), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n966), .C(i_clk), .RN(i_rst_n), .Q(regs[458]) );
  DFEC1 regs_reg_13__15_ ( .D(n867), .E(n967), .C(i_clk), .RN(n942), .Q(
        regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(n864), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(n861), .E(n967), .C(i_clk), .RN(n937), .Q(
        regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(n858), .E(n967), .C(i_clk), .RN(n943), .Q(
        regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(n855), .E(n967), .C(i_clk), .RN(i_rst_n), .Q(
        regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n967), .C(i_clk), .RN(n938), 
        .Q(regs[426]) );
  DFEC1 regs_reg_12__15_ ( .D(n867), .E(n968), .C(i_clk), .RN(n935), .Q(
        regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(n864), .E(n968), .C(i_clk), .RN(n928), .Q(
        regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(n861), .E(n968), .C(i_clk), .RN(n929), .Q(
        regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(n858), .E(n968), .C(i_clk), .RN(n930), .Q(
        regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(n855), .E(n968), .C(i_clk), .RN(n931), .Q(
        regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n968), .C(i_clk), .RN(n932), 
        .Q(regs[394]) );
  DFEC1 regs_reg_11__15_ ( .D(n867), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(n864), .E(n969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(n861), .E(n969), .C(i_clk), .RN(n936), .Q(
        regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(n858), .E(n969), .C(i_clk), .RN(n927), .Q(
        regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(n855), .E(n969), .C(i_clk), .RN(n943), .Q(
        regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(i_data_Rd[10]), .E(n969), .C(i_clk), .RN(n937), 
        .Q(regs[362]) );
  DFEC1 regs_reg_10__15_ ( .D(n867), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(n864), .E(n970), .C(i_clk), .RN(n927), .Q(
        regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(n861), .E(n970), .C(i_clk), .RN(n938), .Q(
        regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(n858), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(n855), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n970), .C(i_clk), .RN(i_rst_n), .Q(regs[330]) );
  DFEC1 regs_reg_9__15_ ( .D(n867), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(n864), .E(n971), .C(i_clk), .RN(n947), .Q(
        regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(n861), .E(n971), .C(i_clk), .RN(n933), .Q(
        regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(n858), .E(n971), .C(i_clk), .RN(n927), .Q(
        regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(n855), .E(n971), .C(i_clk), .RN(n936), .Q(
        regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(i_data_Rd[10]), .E(n971), .C(i_clk), .RN(n927), 
        .Q(regs[298]) );
  DFEC1 regs_reg_8__15_ ( .D(n867), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(n864), .E(n972), .C(i_clk), .RN(n943), .Q(
        regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(n861), .E(n972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(n858), .E(n972), .C(i_clk), .RN(n935), .Q(
        regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(n855), .E(n972), .C(i_clk), .RN(n932), .Q(
        regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(i_data_Rd[10]), .E(n972), .C(i_clk), .RN(n947), 
        .Q(regs[266]) );
  DFEC1 regs_reg_7__15_ ( .D(n866), .E(n973), .C(i_clk), .RN(n927), .Q(
        regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(n863), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(n860), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(n857), .E(n973), .C(i_clk), .RN(n931), .Q(
        regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(n854), .E(n973), .C(i_clk), .RN(n932), .Q(
        regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(n851), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[234]) );
  DFEC1 regs_reg_6__15_ ( .D(n866), .E(n974), .C(i_clk), .RN(n939), .Q(
        regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(n863), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(n860), .E(n974), .C(i_clk), .RN(n947), .Q(
        regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(n857), .E(n974), .C(i_clk), .RN(n945), .Q(
        regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(n854), .E(n974), .C(i_clk), .RN(n944), .Q(
        regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(n851), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[202]) );
  DFEC1 regs_reg_5__15_ ( .D(n866), .E(n975), .C(i_clk), .RN(n942), .Q(
        regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(n863), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(n860), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(n857), .E(n975), .C(i_clk), .RN(n927), .Q(
        regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(n854), .E(n975), .C(i_clk), .RN(n945), .Q(
        regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(n851), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[170]) );
  DFEC1 regs_reg_4__15_ ( .D(n866), .E(n976), .C(i_clk), .RN(n940), .Q(
        regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(n863), .E(n976), .C(i_clk), .RN(n939), .Q(
        regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(n860), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(n857), .E(n976), .C(i_clk), .RN(n945), .Q(
        regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(n854), .E(n976), .C(i_clk), .RN(n943), .Q(
        regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(n851), .E(n976), .C(i_clk), .RN(n940), .Q(
        regs[138]) );
  DFEC1 regs_reg_3__15_ ( .D(n866), .E(n977), .C(i_clk), .RN(n929), .Q(
        regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(n863), .E(n977), .C(i_clk), .RN(n927), .Q(
        regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(n860), .E(n977), .C(i_clk), .RN(n947), .Q(
        regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(n857), .E(n977), .C(i_clk), .RN(n927), .Q(
        regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(n854), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(n851), .E(n977), .C(i_clk), .RN(n946), .Q(
        regs[106]) );
  DFEC1 regs_reg_2__15_ ( .D(n866), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(n863), .E(n978), .C(i_clk), .RN(n945), .Q(
        regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(n860), .E(n978), .C(i_clk), .RN(n927), .Q(
        regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(n857), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(n854), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(n851), .E(n978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[74]) );
  DFEC1 regs_reg_1__15_ ( .D(n866), .E(n979), .C(i_clk), .RN(n940), .Q(
        regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(n863), .E(n979), .C(i_clk), .RN(n940), .Q(
        regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(n860), .E(n979), .C(i_clk), .RN(n940), .Q(
        regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(n857), .E(n979), .C(i_clk), .RN(n940), .Q(
        regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(n854), .E(n979), .C(i_clk), .RN(n940), .Q(
        regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(n851), .E(n979), .C(i_clk), .RN(n941), .Q(
        regs[42]) );
  DFEC1 regs_reg_0__15_ ( .D(n866), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(n863), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(n860), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(n857), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(n854), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(n851), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[10]) );
  DFEC1 regs_reg_31__7_ ( .D(n844), .E(n958), .C(i_clk), .RN(n930), .Q(
        regs[999]) );
  DFEC1 regs_reg_30__7_ ( .D(n844), .E(n959), .C(i_clk), .RN(n934), .Q(
        regs[967]) );
  DFEC1 regs_reg_29__7_ ( .D(n844), .E(n960), .C(i_clk), .RN(n937), .Q(
        regs[935]) );
  DFEC1 regs_reg_28__7_ ( .D(n844), .E(n961), .C(i_clk), .RN(i_rst_n), .Q(
        regs[903]) );
  DFEC1 regs_reg_27__7_ ( .D(n844), .E(n962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[871]) );
  DFEC1 regs_reg_26__7_ ( .D(n844), .E(n963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[839]) );
  DFEC1 regs_reg_25__7_ ( .D(n844), .E(n956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[807]) );
  DFEC1 regs_reg_24__7_ ( .D(n844), .E(n957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[775]) );
  DFEC1 regs_reg_23__7_ ( .D(n843), .E(n948), .C(i_clk), .RN(i_rst_n), .Q(
        regs[743]) );
  DFEC1 regs_reg_22__7_ ( .D(n843), .E(n949), .C(i_clk), .RN(i_rst_n), .Q(
        regs[711]) );
  DFEC1 regs_reg_21__7_ ( .D(n843), .E(n950), .C(i_clk), .RN(i_rst_n), .Q(
        regs[679]) );
  DFEC1 regs_reg_20__7_ ( .D(n843), .E(n951), .C(i_clk), .RN(n943), .Q(
        regs[647]) );
  DFEC1 regs_reg_19__7_ ( .D(n843), .E(n952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[615]) );
  DFEC1 regs_reg_18__7_ ( .D(n843), .E(n953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[583]) );
  DFEC1 regs_reg_17__7_ ( .D(n843), .E(n954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[551]) );
  DFEC1 regs_reg_16__7_ ( .D(n843), .E(n955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[519]) );
  DFEC1 regs_reg_15__7_ ( .D(n842), .E(n965), .C(i_clk), .RN(n936), .Q(
        regs[487]) );
  DFEC1 regs_reg_14__7_ ( .D(n842), .E(n966), .C(i_clk), .RN(n931), .Q(
        regs[455]) );
  DFEC1 regs_reg_13__7_ ( .D(n842), .E(n967), .C(i_clk), .RN(n934), .Q(
        regs[423]) );
  DFEC1 regs_reg_12__7_ ( .D(n842), .E(n968), .C(i_clk), .RN(n934), .Q(
        regs[391]) );
  DFEC1 regs_reg_11__7_ ( .D(n842), .E(n969), .C(i_clk), .RN(n936), .Q(
        regs[359]) );
  DFEC1 regs_reg_10__7_ ( .D(n842), .E(n970), .C(i_clk), .RN(n932), .Q(
        regs[327]) );
  DFEC1 regs_reg_9__7_ ( .D(n842), .E(n971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[295]) );
  DFEC1 regs_reg_8__7_ ( .D(n842), .E(n972), .C(i_clk), .RN(n938), .Q(
        regs[263]) );
  DFEC1 regs_reg_7__7_ ( .D(n841), .E(n973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[231]) );
  DFEC1 regs_reg_6__7_ ( .D(n841), .E(n974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[199]) );
  DFEC1 regs_reg_5__7_ ( .D(n841), .E(n975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[167]) );
  DFEC1 regs_reg_4__7_ ( .D(n841), .E(n976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[135]) );
  DFEC1 regs_reg_3__7_ ( .D(n841), .E(n977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[103]) );
  DFEC1 regs_reg_2__7_ ( .D(n841), .E(n978), .C(i_clk), .RN(n944), .Q(regs[71]) );
  DFEC1 regs_reg_1__7_ ( .D(n841), .E(n979), .C(i_clk), .RN(n941), .Q(regs[39]) );
  DFEC1 regs_reg_0__7_ ( .D(n841), .E(n980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[7]) );
  IMUX40 U2 ( .A(n504), .B(n505), .C(n506), .D(n507), .S0(n765), .S1(n770), 
        .Q(n503) );
  IMUX40 U3 ( .A(n634), .B(n635), .C(n636), .D(n637), .S0(n766), .S1(n773), 
        .Q(n633) );
  CLKIN6 U4 ( .A(n816), .Q(n3) );
  CLKBU12 U5 ( .A(n819), .Q(n7) );
  INV8 U6 ( .A(n3), .Q(n4) );
  BUF6 U7 ( .A(n814), .Q(n811) );
  IMUX40 U8 ( .A(n444), .B(n445), .C(n446), .D(n447), .S0(n768), .S1(n771), 
        .Q(n443) );
  IMUX40 U9 ( .A(n599), .B(n600), .C(n601), .D(n602), .S0(n766), .S1(n772), 
        .Q(n598) );
  IMUX40 U10 ( .A(n604), .B(n605), .C(n606), .D(n607), .S0(n766), .S1(n772), 
        .Q(n603) );
  IMUX40 U11 ( .A(n644), .B(n645), .C(n646), .D(n647), .S0(n767), .S1(n773), 
        .Q(n643) );
  IMUX40 U12 ( .A(n674), .B(n675), .C(n676), .D(n677), .S0(n767), .S1(n770), 
        .Q(n673) );
  IMUX40 U13 ( .A(n684), .B(n685), .C(n686), .D(n687), .S0(n767), .S1(
        i_addr_Rs[2]), .Q(n683) );
  IMUX40 U14 ( .A(n689), .B(n690), .C(n691), .D(n692), .S0(n767), .S1(
        i_addr_Rs[2]), .Q(n688) );
  IMUX40 U15 ( .A(n699), .B(n700), .C(n701), .D(n702), .S0(n767), .S1(
        i_addr_Rs[2]), .Q(n698) );
  IMUX40 U16 ( .A(n694), .B(n695), .C(n696), .D(n697), .S0(n767), .S1(n769), 
        .Q(n693) );
  MUX22 U17 ( .A(n728), .B(n723), .S(n764), .Q(o_data_Rs[28]) );
  IMUX40 U18 ( .A(n729), .B(n730), .C(n731), .D(n732), .S0(n768), .S1(n773), 
        .Q(n728) );
  IMUX40 U19 ( .A(n724), .B(n725), .C(n726), .D(n727), .S0(n768), .S1(
        i_addr_Rs[2]), .Q(n723) );
  IMUX40 U20 ( .A(n734), .B(n735), .C(n736), .D(n737), .S0(n768), .S1(n773), 
        .Q(n733) );
  IMUX40 U21 ( .A(n749), .B(n750), .C(n751), .D(n752), .S0(n768), .S1(n769), 
        .Q(n748) );
  IMUX40 U22 ( .A(n744), .B(n745), .C(n746), .D(n747), .S0(n768), .S1(n772), 
        .Q(n743) );
  IMUX40 U23 ( .A(n759), .B(n760), .C(n761), .D(n762), .S0(n768), .S1(n771), 
        .Q(n758) );
  IMUX40 U24 ( .A(n754), .B(n755), .C(n756), .D(n757), .S0(n768), .S1(
        i_addr_Rs[2]), .Q(n753) );
  BUF4 U25 ( .A(n815), .Q(n807) );
  BUF2 U26 ( .A(i_addr_Rs[0]), .Q(n816) );
  IMUX41 U27 ( .A(n524), .B(n525), .C(n526), .D(n527), .S0(n767), .S1(n770), 
        .Q(n523) );
  IMUX41 U28 ( .A(n529), .B(n530), .C(n531), .D(n532), .S0(n766), .S1(n770), 
        .Q(n528) );
  CLKBU4 U29 ( .A(i_addr_Rs[0]), .Q(n815) );
  CLKBU4 U30 ( .A(i_addr_Rs[3]), .Q(n765) );
  CLKBU4 U31 ( .A(n814), .Q(n805) );
  CLKBU4 U32 ( .A(i_addr_Rs[0]), .Q(n814) );
  BUF8 U33 ( .A(n819), .Q(n813) );
  CLKBU15 U34 ( .A(n10), .Q(n2) );
  BUF2 U35 ( .A(i_addr_Rs[0]), .Q(n819) );
  BUF6 U36 ( .A(n809), .Q(n1) );
  CLKBU15 U37 ( .A(n10), .Q(n5) );
  BUF6 U38 ( .A(n809), .Q(n6) );
  BUF6 U39 ( .A(n817), .Q(n808) );
  CLKBU4 U40 ( .A(i_addr_Rs[0]), .Q(n817) );
  CLKBU4 U41 ( .A(i_addr_Rs[3]), .Q(n767) );
  BUF2 U42 ( .A(n815), .Q(n10) );
  IMUX41 U43 ( .A(n719), .B(n720), .C(n721), .D(n722), .S0(n768), .S1(
        i_addr_Rs[2]), .Q(n718) );
  CLKBU4 U44 ( .A(i_addr_Rs[3]), .Q(n768) );
  BUF6 U45 ( .A(n810), .Q(n8) );
  CLKBU4 U46 ( .A(i_addr_Rs[3]), .Q(n766) );
  IMUX41 U47 ( .A(n629), .B(n630), .C(n631), .D(n632), .S0(n766), .S1(n773), 
        .Q(n628) );
  IMUX41 U48 ( .A(n704), .B(n705), .C(n706), .D(n707), .S0(n768), .S1(
        i_addr_Rs[2]), .Q(n703) );
  CLKBU12 U49 ( .A(n818), .Q(n9) );
  IMUX41 U50 ( .A(n714), .B(n715), .C(n716), .D(n717), .S0(n768), .S1(
        i_addr_Rs[2]), .Q(n713) );
  IMUX41 U51 ( .A(n654), .B(n655), .C(n656), .D(n657), .S0(n767), .S1(n773), 
        .Q(n653) );
  IMUX41 U52 ( .A(n614), .B(n615), .C(n616), .D(n617), .S0(n766), .S1(n772), 
        .Q(n613) );
  IMUX41 U53 ( .A(n594), .B(n595), .C(n596), .D(n597), .S0(n766), .S1(n772), 
        .Q(n593) );
  IMUX41 U54 ( .A(n624), .B(n625), .C(n626), .D(n627), .S0(n766), .S1(n772), 
        .Q(n623) );
  BUF2 U55 ( .A(i_addr_Rs[4]), .Q(n764) );
  BUF2 U56 ( .A(n942), .Q(n939) );
  BUF2 U57 ( .A(n927), .Q(n938) );
  BUF2 U58 ( .A(n947), .Q(n937) );
  BUF2 U59 ( .A(n944), .Q(n936) );
  BUF2 U60 ( .A(n944), .Q(n935) );
  BUF2 U61 ( .A(n944), .Q(n934) );
  BUF2 U62 ( .A(n945), .Q(n933) );
  BUF2 U63 ( .A(n945), .Q(n932) );
  BUF2 U64 ( .A(n945), .Q(n931) );
  BUF2 U65 ( .A(n946), .Q(n930) );
  BUF2 U66 ( .A(n946), .Q(n929) );
  BUF2 U67 ( .A(n946), .Q(n928) );
  BUF2 U68 ( .A(n943), .Q(n942) );
  BUF2 U69 ( .A(n943), .Q(n941) );
  BUF2 U70 ( .A(n943), .Q(n940) );
  BUF2 U71 ( .A(n947), .Q(n944) );
  BUF2 U72 ( .A(n937), .Q(n945) );
  BUF2 U73 ( .A(n938), .Q(n946) );
  BUF2 U74 ( .A(n947), .Q(n943) );
  BUF2 U75 ( .A(n815), .Q(n806) );
  BUF2 U76 ( .A(n817), .Q(n809) );
  BUF2 U77 ( .A(n817), .Q(n810) );
  BUF2 U78 ( .A(n814), .Q(n812) );
  BUF2 U79 ( .A(n778), .Q(n780) );
  BUF2 U80 ( .A(n804), .Q(n781) );
  BUF2 U81 ( .A(n778), .Q(n782) );
  BUF2 U82 ( .A(n778), .Q(n783) );
  BUF2 U83 ( .A(n778), .Q(n784) );
  BUF2 U84 ( .A(n778), .Q(n785) );
  BUF2 U85 ( .A(n778), .Q(n786) );
  BUF2 U86 ( .A(n778), .Q(n787) );
  BUF2 U87 ( .A(n777), .Q(n788) );
  BUF2 U88 ( .A(n777), .Q(n789) );
  BUF2 U89 ( .A(n775), .Q(n790) );
  BUF2 U90 ( .A(n774), .Q(n791) );
  BUF2 U91 ( .A(n804), .Q(n792) );
  BUF2 U92 ( .A(n777), .Q(n793) );
  BUF2 U93 ( .A(n777), .Q(n794) );
  BUF2 U94 ( .A(n776), .Q(n795) );
  BUF2 U95 ( .A(n776), .Q(n796) );
  BUF2 U96 ( .A(n776), .Q(n797) );
  BUF2 U97 ( .A(n775), .Q(n798) );
  BUF2 U98 ( .A(n775), .Q(n799) );
  BUF2 U99 ( .A(n774), .Q(n800) );
  BUF2 U100 ( .A(n774), .Q(n801) );
  BUF2 U101 ( .A(n774), .Q(n802) );
  BUF2 U102 ( .A(i_data_Rd[0]), .Q(n820) );
  BUF2 U103 ( .A(i_data_Rd[1]), .Q(n823) );
  BUF2 U104 ( .A(i_data_Rd[2]), .Q(n826) );
  BUF2 U105 ( .A(i_data_Rd[3]), .Q(n829) );
  BUF2 U106 ( .A(i_data_Rd[4]), .Q(n832) );
  BUF2 U107 ( .A(i_data_Rd[5]), .Q(n835) );
  BUF2 U108 ( .A(i_data_Rd[6]), .Q(n838) );
  BUF2 U109 ( .A(i_data_Rd[7]), .Q(n841) );
  BUF2 U110 ( .A(i_data_Rd[10]), .Q(n851) );
  BUF2 U111 ( .A(i_data_Rd[11]), .Q(n854) );
  BUF2 U112 ( .A(i_data_Rd[12]), .Q(n857) );
  BUF2 U113 ( .A(i_data_Rd[13]), .Q(n860) );
  BUF2 U114 ( .A(i_data_Rd[14]), .Q(n863) );
  BUF2 U115 ( .A(i_data_Rd[15]), .Q(n866) );
  BUF2 U116 ( .A(i_data_Rd[16]), .Q(n869) );
  BUF2 U117 ( .A(i_data_Rd[17]), .Q(n872) );
  BUF2 U118 ( .A(i_data_Rd[19]), .Q(n879) );
  BUF2 U119 ( .A(i_data_Rd[20]), .Q(n882) );
  BUF2 U120 ( .A(i_data_Rd[21]), .Q(n885) );
  BUF2 U121 ( .A(i_data_Rd[22]), .Q(n888) );
  BUF2 U122 ( .A(i_data_Rd[23]), .Q(n891) );
  BUF2 U123 ( .A(i_data_Rd[24]), .Q(n895) );
  BUF2 U124 ( .A(i_data_Rd[25]), .Q(n899) );
  BUF2 U125 ( .A(i_data_Rd[26]), .Q(n903) );
  BUF2 U126 ( .A(i_data_Rd[27]), .Q(n907) );
  BUF2 U127 ( .A(i_data_Rd[28]), .Q(n911) );
  BUF2 U128 ( .A(i_data_Rd[29]), .Q(n915) );
  BUF2 U129 ( .A(i_data_Rd[30]), .Q(n919) );
  BUF2 U130 ( .A(i_data_Rd[31]), .Q(n923) );
  BUF2 U131 ( .A(i_data_Rd[0]), .Q(n821) );
  BUF2 U132 ( .A(i_data_Rd[1]), .Q(n824) );
  BUF2 U133 ( .A(i_data_Rd[2]), .Q(n827) );
  BUF2 U134 ( .A(i_data_Rd[3]), .Q(n830) );
  BUF2 U135 ( .A(i_data_Rd[4]), .Q(n833) );
  BUF2 U136 ( .A(i_data_Rd[5]), .Q(n836) );
  BUF2 U137 ( .A(i_data_Rd[6]), .Q(n839) );
  BUF2 U138 ( .A(i_data_Rd[7]), .Q(n842) );
  BUF2 U139 ( .A(i_data_Rd[11]), .Q(n855) );
  BUF2 U140 ( .A(i_data_Rd[12]), .Q(n858) );
  BUF2 U141 ( .A(i_data_Rd[13]), .Q(n861) );
  BUF2 U142 ( .A(i_data_Rd[14]), .Q(n864) );
  BUF2 U143 ( .A(i_data_Rd[15]), .Q(n867) );
  BUF2 U144 ( .A(i_data_Rd[16]), .Q(n870) );
  BUF2 U145 ( .A(i_data_Rd[17]), .Q(n873) );
  BUF2 U146 ( .A(i_data_Rd[19]), .Q(n880) );
  BUF2 U147 ( .A(i_data_Rd[20]), .Q(n883) );
  BUF2 U148 ( .A(i_data_Rd[21]), .Q(n886) );
  BUF2 U149 ( .A(i_data_Rd[22]), .Q(n889) );
  BUF2 U150 ( .A(i_data_Rd[23]), .Q(n892) );
  BUF2 U151 ( .A(i_data_Rd[24]), .Q(n896) );
  BUF2 U152 ( .A(i_data_Rd[25]), .Q(n900) );
  BUF2 U153 ( .A(i_data_Rd[26]), .Q(n904) );
  BUF2 U154 ( .A(i_data_Rd[27]), .Q(n908) );
  BUF2 U155 ( .A(i_data_Rd[28]), .Q(n912) );
  BUF2 U156 ( .A(i_data_Rd[29]), .Q(n916) );
  BUF2 U157 ( .A(i_data_Rd[30]), .Q(n920) );
  BUF2 U158 ( .A(i_data_Rd[31]), .Q(n924) );
  BUF2 U159 ( .A(i_data_Rd[0]), .Q(n822) );
  BUF2 U160 ( .A(i_data_Rd[1]), .Q(n825) );
  BUF2 U161 ( .A(i_data_Rd[2]), .Q(n828) );
  BUF2 U162 ( .A(i_data_Rd[3]), .Q(n831) );
  BUF2 U163 ( .A(i_data_Rd[4]), .Q(n834) );
  BUF2 U164 ( .A(i_data_Rd[5]), .Q(n837) );
  BUF2 U165 ( .A(i_data_Rd[6]), .Q(n840) );
  BUF2 U166 ( .A(i_data_Rd[7]), .Q(n843) );
  BUF2 U167 ( .A(i_data_Rd[10]), .Q(n852) );
  BUF2 U168 ( .A(i_data_Rd[11]), .Q(n856) );
  BUF2 U169 ( .A(i_data_Rd[12]), .Q(n859) );
  BUF2 U170 ( .A(i_data_Rd[13]), .Q(n862) );
  BUF2 U171 ( .A(i_data_Rd[14]), .Q(n865) );
  BUF2 U172 ( .A(i_data_Rd[15]), .Q(n868) );
  BUF2 U173 ( .A(i_data_Rd[16]), .Q(n871) );
  BUF2 U174 ( .A(i_data_Rd[17]), .Q(n874) );
  BUF2 U175 ( .A(i_data_Rd[19]), .Q(n881) );
  BUF2 U176 ( .A(i_data_Rd[21]), .Q(n887) );
  BUF2 U177 ( .A(i_data_Rd[22]), .Q(n890) );
  BUF2 U178 ( .A(i_data_Rd[23]), .Q(n893) );
  BUF2 U179 ( .A(i_data_Rd[24]), .Q(n897) );
  BUF2 U180 ( .A(i_data_Rd[25]), .Q(n901) );
  BUF2 U181 ( .A(i_data_Rd[26]), .Q(n905) );
  BUF2 U182 ( .A(i_data_Rd[27]), .Q(n909) );
  BUF2 U183 ( .A(i_data_Rd[28]), .Q(n913) );
  BUF2 U184 ( .A(i_data_Rd[29]), .Q(n917) );
  BUF2 U185 ( .A(i_data_Rd[30]), .Q(n921) );
  BUF2 U186 ( .A(i_data_Rd[31]), .Q(n925) );
  BUF2 U187 ( .A(i_data_Rd[7]), .Q(n844) );
  BUF2 U188 ( .A(i_data_Rd[10]), .Q(n853) );
  BUF2 U189 ( .A(i_data_Rd[20]), .Q(n884) );
  BUF2 U190 ( .A(i_data_Rd[23]), .Q(n894) );
  BUF2 U191 ( .A(i_data_Rd[24]), .Q(n898) );
  BUF2 U192 ( .A(i_data_Rd[25]), .Q(n902) );
  BUF2 U193 ( .A(i_data_Rd[26]), .Q(n906) );
  BUF2 U194 ( .A(i_data_Rd[27]), .Q(n910) );
  BUF2 U195 ( .A(i_data_Rd[28]), .Q(n914) );
  BUF2 U196 ( .A(i_data_Rd[29]), .Q(n918) );
  BUF2 U197 ( .A(i_data_Rd[30]), .Q(n922) );
  BUF2 U198 ( .A(i_data_Rd[31]), .Q(n926) );
  BUF2 U199 ( .A(i_data_Rd[18]), .Q(n875) );
  BUF2 U200 ( .A(i_data_Rd[18]), .Q(n876) );
  BUF2 U201 ( .A(i_data_Rd[18]), .Q(n877) );
  BUF2 U202 ( .A(i_data_Rd[18]), .Q(n878) );
  BUF2 U203 ( .A(n776), .Q(n779) );
  BUF2 U204 ( .A(n438), .Q(n417) );
  BUF2 U205 ( .A(n438), .Q(n418) );
  BUF2 U206 ( .A(n438), .Q(n419) );
  BUF2 U207 ( .A(i_addr_Rt[0]), .Q(n420) );
  BUF2 U208 ( .A(i_addr_Rt[0]), .Q(n421) );
  BUF2 U209 ( .A(i_addr_Rt[0]), .Q(n422) );
  BUF2 U210 ( .A(n439), .Q(n423) );
  BUF2 U211 ( .A(n439), .Q(n424) );
  BUF2 U212 ( .A(n439), .Q(n425) );
  BUF2 U213 ( .A(n440), .Q(n426) );
  BUF2 U214 ( .A(n440), .Q(n427) );
  BUF2 U215 ( .A(n440), .Q(n428) );
  BUF2 U216 ( .A(i_addr_Rt[0]), .Q(n429) );
  BUF2 U217 ( .A(i_addr_Rt[0]), .Q(n430) );
  BUF2 U218 ( .A(i_addr_Rt[0]), .Q(n431) );
  BUF2 U219 ( .A(n441), .Q(n432) );
  BUF2 U220 ( .A(n441), .Q(n433) );
  BUF2 U221 ( .A(n441), .Q(n434) );
  BUF2 U222 ( .A(n442), .Q(n435) );
  BUF2 U223 ( .A(n442), .Q(n436) );
  BUF2 U224 ( .A(n442), .Q(n437) );
  INV3 U225 ( .A(n51), .Q(n958) );
  NAND22 U226 ( .A(n52), .B(n42), .Q(n51) );
  BUF2 U227 ( .A(n415), .Q(n397) );
  BUF2 U228 ( .A(n394), .Q(n398) );
  BUF2 U229 ( .A(n393), .Q(n399) );
  BUF2 U230 ( .A(n395), .Q(n400) );
  BUF2 U231 ( .A(n395), .Q(n401) );
  BUF2 U232 ( .A(n395), .Q(n402) );
  BUF2 U233 ( .A(n394), .Q(n403) );
  BUF2 U234 ( .A(n394), .Q(n404) );
  BUF2 U235 ( .A(n394), .Q(n405) );
  BUF2 U236 ( .A(n393), .Q(n406) );
  BUF2 U237 ( .A(n393), .Q(n407) );
  BUF2 U238 ( .A(n393), .Q(n408) );
  BUF2 U239 ( .A(n392), .Q(n409) );
  BUF2 U240 ( .A(n392), .Q(n410) );
  BUF2 U241 ( .A(n392), .Q(n411) );
  BUF2 U242 ( .A(i_data_Rd[8]), .Q(n845) );
  BUF2 U243 ( .A(i_data_Rd[9]), .Q(n848) );
  BUF2 U244 ( .A(i_data_Rd[8]), .Q(n846) );
  BUF2 U245 ( .A(i_data_Rd[9]), .Q(n849) );
  BUF2 U246 ( .A(i_data_Rd[8]), .Q(n847) );
  BUF2 U247 ( .A(i_data_Rd[9]), .Q(n850) );
  BUF2 U248 ( .A(n927), .Q(n947) );
  BUF2 U249 ( .A(i_rst_n), .Q(n927) );
  BUF2 U250 ( .A(i_addr_Rs[0]), .Q(n818) );
  BUF2 U251 ( .A(i_addr_Rs[1]), .Q(n778) );
  BUF2 U252 ( .A(n804), .Q(n777) );
  BUF2 U253 ( .A(n803), .Q(n776) );
  BUF2 U254 ( .A(n803), .Q(n775) );
  BUF2 U255 ( .A(n803), .Q(n774) );
  NOR31 U256 ( .A(n964), .B(n981), .C(n985), .Q(n42) );
  NOR31 U257 ( .A(n983), .B(n984), .C(n982), .Q(n52) );
  INV3 U258 ( .A(n39), .Q(n956) );
  NAND22 U259 ( .A(n42), .B(n57), .Q(n39) );
  INV3 U260 ( .A(n82), .Q(n957) );
  NAND22 U261 ( .A(n55), .B(n42), .Q(n82) );
  INV3 U262 ( .A(n40), .Q(n963) );
  NAND22 U263 ( .A(n41), .B(n42), .Q(n40) );
  INV3 U264 ( .A(n43), .Q(n962) );
  NAND22 U265 ( .A(n44), .B(n42), .Q(n43) );
  INV3 U266 ( .A(n45), .Q(n961) );
  NAND22 U267 ( .A(n46), .B(n42), .Q(n45) );
  INV3 U268 ( .A(n47), .Q(n960) );
  NAND22 U269 ( .A(n48), .B(n42), .Q(n47) );
  INV3 U270 ( .A(n49), .Q(n959) );
  NAND22 U271 ( .A(n50), .B(n42), .Q(n49) );
  INV3 U272 ( .A(n53), .Q(n980) );
  NAND22 U273 ( .A(n54), .B(n55), .Q(n53) );
  INV3 U274 ( .A(n56), .Q(n979) );
  NAND22 U275 ( .A(n54), .B(n57), .Q(n56) );
  INV3 U276 ( .A(n58), .Q(n978) );
  NAND22 U277 ( .A(n54), .B(n41), .Q(n58) );
  INV3 U278 ( .A(n59), .Q(n977) );
  NAND22 U279 ( .A(n54), .B(n44), .Q(n59) );
  INV3 U280 ( .A(n60), .Q(n976) );
  NAND22 U281 ( .A(n54), .B(n46), .Q(n60) );
  INV3 U282 ( .A(n61), .Q(n975) );
  NAND22 U283 ( .A(n54), .B(n48), .Q(n61) );
  INV3 U284 ( .A(n62), .Q(n974) );
  NAND22 U285 ( .A(n54), .B(n50), .Q(n62) );
  INV3 U286 ( .A(n63), .Q(n973) );
  NAND22 U287 ( .A(n54), .B(n52), .Q(n63) );
  INV3 U288 ( .A(n64), .Q(n972) );
  NAND22 U289 ( .A(n65), .B(n55), .Q(n64) );
  INV3 U290 ( .A(n66), .Q(n971) );
  NAND22 U291 ( .A(n65), .B(n57), .Q(n66) );
  INV3 U292 ( .A(n67), .Q(n970) );
  NAND22 U293 ( .A(n65), .B(n41), .Q(n67) );
  INV3 U294 ( .A(n68), .Q(n969) );
  NAND22 U295 ( .A(n65), .B(n44), .Q(n68) );
  INV3 U296 ( .A(n69), .Q(n968) );
  NAND22 U297 ( .A(n65), .B(n46), .Q(n69) );
  INV3 U298 ( .A(n70), .Q(n967) );
  NAND22 U299 ( .A(n65), .B(n48), .Q(n70) );
  INV3 U300 ( .A(n71), .Q(n966) );
  NAND22 U301 ( .A(n65), .B(n50), .Q(n71) );
  INV3 U302 ( .A(n72), .Q(n965) );
  NAND22 U303 ( .A(n65), .B(n52), .Q(n72) );
  INV3 U304 ( .A(n73), .Q(n955) );
  NAND22 U305 ( .A(n74), .B(n55), .Q(n73) );
  INV3 U306 ( .A(n75), .Q(n954) );
  NAND22 U307 ( .A(n74), .B(n57), .Q(n75) );
  INV3 U308 ( .A(n76), .Q(n953) );
  NAND22 U309 ( .A(n74), .B(n41), .Q(n76) );
  INV3 U310 ( .A(n77), .Q(n952) );
  NAND22 U311 ( .A(n74), .B(n44), .Q(n77) );
  INV3 U312 ( .A(n78), .Q(n951) );
  NAND22 U313 ( .A(n74), .B(n46), .Q(n78) );
  INV3 U314 ( .A(n79), .Q(n950) );
  NAND22 U315 ( .A(n74), .B(n48), .Q(n79) );
  INV3 U316 ( .A(n80), .Q(n949) );
  NAND22 U317 ( .A(n74), .B(n50), .Q(n80) );
  INV3 U318 ( .A(n81), .Q(n948) );
  NAND22 U319 ( .A(n74), .B(n52), .Q(n81) );
  BUF2 U320 ( .A(n414), .Q(n412) );
  BUF2 U321 ( .A(n395), .Q(n413) );
  BUF2 U322 ( .A(i_addr_Rt[0]), .Q(n438) );
  BUF2 U323 ( .A(i_addr_Rt[0]), .Q(n439) );
  BUF2 U324 ( .A(i_addr_Rt[0]), .Q(n440) );
  BUF2 U325 ( .A(i_addr_Rt[0]), .Q(n441) );
  BUF2 U326 ( .A(i_addr_Rt[0]), .Q(n442) );
  BUF2 U327 ( .A(n414), .Q(n396) );
  BUF2 U328 ( .A(n416), .Q(n395) );
  BUF2 U329 ( .A(n416), .Q(n394) );
  BUF2 U330 ( .A(n416), .Q(n393) );
  BUF2 U331 ( .A(n415), .Q(n392) );
  BUF2 U332 ( .A(n415), .Q(n391) );
  BUF2 U333 ( .A(n415), .Q(n390) );
  IMUX40 U334 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n806), .S1(n780), .Q(n449) );
  IMUX40 U335 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n5), .S1(n780), .Q(n450) );
  IMUX40 U336 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n806), .S1(n780), .Q(n452) );
  IMUX40 U337 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(n805), .S1(n779), .Q(n447) );
  IMUX40 U338 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(n805), .S1(n779), .Q(n445) );
  IMUX40 U339 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(n805), .S1(n779), .Q(n444) );
  IMUX40 U340 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n808), .S1(n780), .Q(n457) );
  IMUX40 U341 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n808), .S1(n780), .Q(n455) );
  IMUX40 U342 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n5), .S1(n780), .Q(n454) );
  IMUX40 U343 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(n2), 
        .S1(n781), .Q(n459) );
  IMUX40 U344 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n807), .S1(n781), .Q(n460) );
  IMUX40 U345 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n2), .S1(n780), .Q(n462) );
  IMUX40 U346 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n806), .S1(n781), .Q(n467) );
  IMUX40 U347 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n806), .S1(n781), .Q(n465) );
  IMUX40 U348 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n5), .S1(n781), .Q(n464) );
  IMUX40 U349 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n807), .S1(n782), .Q(n469) );
  IMUX40 U350 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n807), .S1(n781), .Q(n470) );
  IMUX40 U351 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n806), .S1(n781), .Q(n472) );
  IMUX40 U352 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n807), .S1(n782), .Q(n477) );
  IMUX40 U353 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n807), .S1(n782), .Q(n475) );
  IMUX40 U354 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n5), .S1(n782), .Q(n474) );
  IMUX40 U355 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n806), .S1(n783), .Q(n479) );
  IMUX40 U356 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n808), .S1(n782), .Q(n482) );
  IMUX40 U357 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n5), .S1(n782), .Q(n480) );
  IMUX40 U358 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n807), .S1(n783), .Q(n487) );
  IMUX40 U359 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n5), .S1(n783), .Q(n485) );
  IMUX40 U360 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n5), .S1(n783), .Q(n484) );
  IMUX40 U361 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n806), .S1(n783), .Q(n489) );
  IMUX40 U362 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n5), .S1(n783), .Q(n490) );
  IMUX40 U363 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n2), .S1(n783), .Q(n492) );
  IMUX40 U364 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n7), .S1(n784), .Q(n497) );
  IMUX40 U365 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n7), .S1(n784), .Q(n495) );
  IMUX40 U366 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n4), .S1(n784), .Q(n494) );
  IMUX40 U367 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(n4), .S1(n784), .Q(n499) );
  IMUX40 U368 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n4), .S1(n784), .Q(n500) );
  IMUX40 U369 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n4), .S1(n784), .Q(n502) );
  IMUX40 U370 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n7), .S1(n784), .Q(n507) );
  IMUX40 U371 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n7), .S1(n785), .Q(n505) );
  IMUX40 U372 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n4), .S1(n785), .Q(n504) );
  IMUX40 U373 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n805), .S1(n785), .Q(n509) );
  IMUX40 U374 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n818), .S1(n785), .Q(n510) );
  IMUX40 U375 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n816), .S1(n785), .Q(n512) );
  IMUX40 U376 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n816), .S1(n785), .Q(n517) );
  IMUX40 U377 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n812), .S1(n785), .Q(n515) );
  IMUX40 U378 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n816), .S1(n786), .Q(n514) );
  IMUX40 U379 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n812), .S1(n786), .Q(n519) );
  IMUX40 U380 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n816), .S1(n786), .Q(n520) );
  IMUX40 U381 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n7), .S1(n786), .Q(n522) );
  IMUX40 U382 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n813), .S1(n786), .Q(n527) );
  IMUX40 U383 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n813), .S1(n786), .Q(n525) );
  IMUX40 U384 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n813), .S1(n787), .Q(n524) );
  IMUX40 U385 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n813), .S1(n787), .Q(n529) );
  IMUX40 U386 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n813), .S1(n787), .Q(n530) );
  IMUX40 U387 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n5), .S1(n787), .Q(n532) );
  IMUX40 U388 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n2), .S1(n787), .Q(n537) );
  IMUX40 U389 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n2), .S1(n787), .Q(n535) );
  IMUX40 U390 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n7), .S1(n787), .Q(n534) );
  IMUX40 U391 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n808), .S1(n788), .Q(n542) );
  IMUX40 U392 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n808), .S1(n786), .Q(n539) );
  IMUX40 U393 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n808), .S1(n790), .Q(n540) );
  IMUX40 U394 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n808), .S1(n793), .Q(n547) );
  IMUX40 U395 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n808), .S1(n795), .Q(n545) );
  IMUX40 U396 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n808), .S1(n779), .Q(n544) );
  IMUX40 U397 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n808), .S1(n791), .Q(n552) );
  IMUX40 U398 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n808), .S1(n788), .Q(n549) );
  IMUX40 U399 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n808), .S1(n788), .Q(n550) );
  IMUX40 U400 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n4), .S1(n788), .Q(n557) );
  IMUX40 U401 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n5), .S1(n788), .Q(n555) );
  IMUX40 U402 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n5), .S1(n788), .Q(n554) );
  IMUX40 U403 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n5), .S1(n788), .Q(n562) );
  IMUX40 U404 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n5), .S1(n789), .Q(n559) );
  IMUX40 U405 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n4), .S1(n788), .Q(n560) );
  IMUX40 U406 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n808), .S1(n789), .Q(n567) );
  IMUX40 U407 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n7), .S1(n789), .Q(n565) );
  IMUX40 U408 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n808), .S1(n789), .Q(n564) );
  IMUX40 U409 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n6), .S1(n789), .Q(n572) );
  IMUX40 U410 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n6), .S1(n790), .Q(n569) );
  IMUX40 U411 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n6), .S1(n789), .Q(n570) );
  IMUX40 U412 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n6), .S1(n790), .Q(n577) );
  IMUX40 U413 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n6), .S1(n790), .Q(n575) );
  IMUX40 U414 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n6), .S1(n790), .Q(n574) );
  IMUX40 U415 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n6), .S1(n790), .Q(n582) );
  IMUX40 U416 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n6), .S1(n790), .Q(n579) );
  IMUX40 U417 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n6), .S1(n790), .Q(n580) );
  IMUX40 U418 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n9), .S1(n791), .Q(n587) );
  IMUX40 U419 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n4), .S1(n791), .Q(n585) );
  IMUX40 U420 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n4), .S1(n791), .Q(n584) );
  IMUX40 U421 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n7), .S1(n791), .Q(n592) );
  IMUX40 U422 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n4), .S1(n791), .Q(n589) );
  IMUX40 U423 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n7), .S1(n791), .Q(n590) );
  IMUX40 U424 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n7), .S1(n791), .Q(n597) );
  IMUX40 U425 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n9), .S1(n792), .Q(n595) );
  IMUX40 U426 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n9), .S1(n792), .Q(n594) );
  IMUX40 U427 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n2), .S1(n792), .Q(n602) );
  IMUX40 U428 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n2), .S1(n792), .Q(n599) );
  IMUX40 U429 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n2), .S1(n792), .Q(n600) );
  IMUX40 U430 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n2), .S1(n792), .Q(n607) );
  IMUX40 U431 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n2), .S1(n792), .Q(n605) );
  IMUX40 U432 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n2), .S1(n793), .Q(n604) );
  IMUX40 U433 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n2), .S1(n793), .Q(n612) );
  IMUX40 U434 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n2), .S1(n793), .Q(n609) );
  IMUX40 U435 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n2), .S1(n793), .Q(n610) );
  IMUX40 U436 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n8), .S1(n793), .Q(n617) );
  IMUX40 U437 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n8), .S1(n793), .Q(n615) );
  IMUX40 U438 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n8), .S1(n794), .Q(n614) );
  IMUX40 U439 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n9), .S1(n794), .Q(n622) );
  IMUX40 U440 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n9), .S1(n794), .Q(n619) );
  IMUX40 U441 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n9), .S1(n794), .Q(n620) );
  IMUX40 U442 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n8), .S1(n794), .Q(n627) );
  IMUX40 U443 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n8), .S1(n794), .Q(n625) );
  IMUX40 U444 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n8), .S1(n794), .Q(n624) );
  IMUX40 U445 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n818), .S1(n792), .Q(n632) );
  IMUX40 U446 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n4), .S1(n792), .Q(n629) );
  IMUX40 U447 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n811), .S1(n792), .Q(n630) );
  IMUX40 U448 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n9), .S1(n792), .Q(n637) );
  IMUX40 U449 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n818), .S1(n779), .Q(n635) );
  IMUX40 U450 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n9), .S1(n792), .Q(n634) );
  IMUX40 U451 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n9), .S1(n792), .Q(n642) );
  IMUX40 U452 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n9), .S1(n795), .Q(n639) );
  IMUX40 U453 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n9), .S1(n795), .Q(n640) );
  IMUX40 U454 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n1), .S1(n795), .Q(n647) );
  IMUX40 U455 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n1), .S1(n795), .Q(n645) );
  IMUX40 U456 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n1), .S1(n795), .Q(n644) );
  IMUX40 U457 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n1), .S1(n795), .Q(n652) );
  IMUX40 U458 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n1), .S1(n796), .Q(n649) );
  IMUX40 U459 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n1), .S1(n795), .Q(n650) );
  IMUX40 U460 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n1), .S1(n796), .Q(n657) );
  IMUX40 U461 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n1), .S1(n796), .Q(n655) );
  IMUX40 U462 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n1), .S1(n796), .Q(n654) );
  IMUX40 U463 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n9), .S1(n796), .Q(n662) );
  IMUX40 U464 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n9), .S1(n797), .Q(n659) );
  IMUX40 U465 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n9), .S1(n796), .Q(n660) );
  IMUX40 U466 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n9), .S1(n797), .Q(n667) );
  IMUX40 U467 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n9), .S1(n797), .Q(n665) );
  IMUX40 U468 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n9), .S1(n797), .Q(n664) );
  IMUX40 U469 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n9), .S1(n797), .Q(n672) );
  IMUX40 U470 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n9), .S1(n797), .Q(n669) );
  IMUX40 U471 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n9), .S1(n797), .Q(n670) );
  IMUX40 U472 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n811), .S1(n798), .Q(n677) );
  IMUX40 U473 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n805), .S1(n798), .Q(n675) );
  IMUX40 U474 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n807), .S1(n798), .Q(n674) );
  IMUX40 U475 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n807), .S1(n798), .Q(n682) );
  IMUX40 U476 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n807), .S1(n798), .Q(n679) );
  IMUX40 U477 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n805), .S1(n798), .Q(n680) );
  IMUX40 U478 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n813), .S1(n798), .Q(n687) );
  IMUX40 U479 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n805), .S1(n800), .Q(n685) );
  IMUX40 U480 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n813), .S1(n780), .Q(n684) );
  IMUX40 U481 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n811), .S1(n794), .Q(n692) );
  IMUX40 U482 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n811), .S1(n783), .Q(n689) );
  IMUX40 U483 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n811), .S1(n784), .Q(n690) );
  IMUX40 U484 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n811), .S1(n799), .Q(n697) );
  IMUX40 U485 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n811), .S1(n798), .Q(n695) );
  IMUX40 U486 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n811), .S1(n799), .Q(n694) );
  IMUX40 U487 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n811), .S1(n799), .Q(n702) );
  IMUX40 U488 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n811), .S1(n799), .Q(n699) );
  IMUX40 U489 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n811), .S1(n799), .Q(n700) );
  IMUX40 U490 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n811), .S1(n799), .Q(n707) );
  IMUX40 U491 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n812), .S1(n799), .Q(n705) );
  IMUX40 U492 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n811), .S1(n800), .Q(n704) );
  IMUX40 U493 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n811), .S1(n800), .Q(n712) );
  IMUX40 U494 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n807), .S1(n800), .Q(n709) );
  IMUX40 U495 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n7), .S1(n800), .Q(n710) );
  IMUX40 U496 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n811), .S1(n800), .Q(n717) );
  IMUX40 U497 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n812), .S1(n800), .Q(n715) );
  IMUX40 U498 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n811), .S1(n800), .Q(n714) );
  IMUX40 U499 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n813), .S1(n801), .Q(n722) );
  IMUX40 U500 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n7), .S1(n801), .Q(n719) );
  IMUX40 U501 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n2), .S1(n801), .Q(n720) );
  IMUX40 U502 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n813), .S1(n801), .Q(n727) );
  IMUX40 U503 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n813), .S1(n801), .Q(n725) );
  IMUX40 U504 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n7), .S1(n801), .Q(n724) );
  IMUX40 U505 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n813), .S1(n801), .Q(n732) );
  IMUX40 U506 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n1), .S1(n802), .Q(n729) );
  IMUX40 U507 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n7), .S1(n802), .Q(n730) );
  IMUX40 U508 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n7), .S1(n802), .Q(n737) );
  IMUX40 U509 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n7), .S1(n802), .Q(n735) );
  IMUX40 U510 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n7), .S1(n802), .Q(n734) );
  IMUX40 U511 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n811), .S1(n802), .Q(n742) );
  IMUX40 U512 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n7), .S1(n781), .Q(n739) );
  IMUX40 U513 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n812), .S1(n802), .Q(n740) );
  IMUX40 U514 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n7), .S1(n787), .Q(n747) );
  IMUX40 U515 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n7), .S1(n781), .Q(n745) );
  IMUX40 U516 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n7), .S1(n782), .Q(n744) );
  IMUX40 U517 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n813), .S1(n780), .Q(n752) );
  IMUX40 U518 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n813), .S1(n785), .Q(n749) );
  IMUX40 U519 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n813), .S1(n778), .Q(n750) );
  IMUX40 U520 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n813), .S1(n782), .Q(n757) );
  IMUX40 U521 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n813), .S1(n784), .Q(n755) );
  IMUX40 U522 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n813), .S1(n787), .Q(n754) );
  IMUX40 U523 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n813), .S1(n779), .Q(n762) );
  IMUX40 U524 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n813), .S1(n781), .Q(n759) );
  IMUX40 U525 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n813), .S1(n781), .Q(n760) );
  IMUX40 U526 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n808), .S1(n780), .Q(n451) );
  IMUX40 U527 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(n805), .S1(n779), .Q(n446) );
  IMUX40 U528 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n808), .S1(n780), .Q(n456) );
  IMUX40 U529 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(i_addr_Rs[0]), .S1(n781), .Q(n466) );
  IMUX40 U530 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n5), .S1(n782), .Q(n476) );
  IMUX40 U531 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n807), .S1(n783), .Q(n486) );
  IMUX40 U532 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n7), .S1(n784), .Q(n496) );
  IMUX40 U533 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n7), .S1(n785), .Q(n506) );
  IMUX40 U534 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n805), .S1(n786), .Q(n516) );
  IMUX40 U535 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n813), .S1(n786), .Q(n526) );
  IMUX40 U536 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n2), .S1(n787), .Q(n536) );
  IMUX40 U537 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n808), .S1(n781), .Q(n546) );
  IMUX40 U538 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n4), .S1(n788), .Q(n556) );
  IMUX40 U539 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n7), .S1(n789), .Q(n566) );
  IMUX40 U540 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n6), .S1(n790), .Q(n576) );
  IMUX40 U541 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n4), .S1(n791), .Q(n586) );
  IMUX40 U542 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n7), .S1(n792), .Q(n596) );
  IMUX40 U543 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n2), .S1(n793), .Q(n606) );
  IMUX40 U544 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n8), .S1(n793), .Q(n616) );
  IMUX40 U545 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n8), .S1(n794), .Q(n626) );
  IMUX40 U546 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n7), .S1(n779), .Q(n636) );
  IMUX40 U547 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n1), .S1(n795), .Q(n646) );
  IMUX40 U548 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n1), .S1(n796), .Q(n656) );
  IMUX40 U549 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n9), .S1(n797), .Q(n666) );
  IMUX40 U550 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n811), .S1(n798), .Q(n676) );
  IMUX40 U551 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n807), .S1(n790), .Q(n686) );
  IMUX40 U552 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n811), .S1(n799), .Q(n696) );
  IMUX40 U553 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n811), .S1(n799), .Q(n706) );
  IMUX40 U554 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n811), .S1(n800), .Q(n716) );
  IMUX40 U555 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n813), .S1(n801), .Q(n726) );
  IMUX40 U556 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n7), .S1(n802), .Q(n736) );
  IMUX40 U557 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n7), .S1(n787), .Q(n746) );
  IMUX40 U558 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n813), .S1(n780), .Q(n756) );
  MUX22 U559 ( .A(n448), .B(n443), .S(n763), .Q(o_data_Rs[0]) );
  IMUX40 U560 ( .A(n449), .B(n450), .C(n451), .D(n452), .S0(n767), .S1(n769), 
        .Q(n448) );
  MUX22 U561 ( .A(n458), .B(n453), .S(n763), .Q(o_data_Rs[1]) );
  IMUX40 U562 ( .A(n459), .B(n460), .C(n461), .D(n462), .S0(n768), .S1(n769), 
        .Q(n458) );
  IMUX40 U563 ( .A(n454), .B(n455), .C(n456), .D(n457), .S0(n768), .S1(n769), 
        .Q(n453) );
  IMUX40 U564 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n808), .S1(n781), .Q(n461) );
  MUX22 U565 ( .A(n468), .B(n463), .S(n763), .Q(o_data_Rs[2]) );
  IMUX40 U566 ( .A(n469), .B(n470), .C(n471), .D(n472), .S0(n765), .S1(n769), 
        .Q(n468) );
  IMUX40 U567 ( .A(n464), .B(n465), .C(n466), .D(n467), .S0(n765), .S1(n769), 
        .Q(n463) );
  IMUX40 U568 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n5), .S1(n782), .Q(n471) );
  MUX22 U569 ( .A(n478), .B(n473), .S(n763), .Q(o_data_Rs[3]) );
  IMUX40 U570 ( .A(n479), .B(n480), .C(n481), .D(n482), .S0(n765), .S1(n769), 
        .Q(n478) );
  IMUX40 U571 ( .A(n474), .B(n475), .C(n476), .D(n477), .S0(n765), .S1(n769), 
        .Q(n473) );
  IMUX40 U572 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n808), .S1(n782), .Q(n481) );
  MUX22 U573 ( .A(n488), .B(n483), .S(n763), .Q(o_data_Rs[4]) );
  IMUX40 U574 ( .A(n489), .B(n490), .C(n491), .D(n492), .S0(n765), .S1(n769), 
        .Q(n488) );
  IMUX40 U575 ( .A(n484), .B(n485), .C(n486), .D(n487), .S0(n765), .S1(n769), 
        .Q(n483) );
  IMUX40 U576 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n5), .S1(n783), .Q(n491) );
  MUX22 U577 ( .A(n498), .B(n493), .S(n763), .Q(o_data_Rs[5]) );
  IMUX40 U578 ( .A(n499), .B(n500), .C(n501), .D(n502), .S0(n765), .S1(n770), 
        .Q(n498) );
  IMUX40 U579 ( .A(n494), .B(n495), .C(n496), .D(n497), .S0(n765), .S1(n770), 
        .Q(n493) );
  IMUX40 U580 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n7), .S1(n784), .Q(n501) );
  MUX22 U581 ( .A(n508), .B(n503), .S(n763), .Q(o_data_Rs[6]) );
  IMUX40 U582 ( .A(n509), .B(n510), .C(n511), .D(n512), .S0(n765), .S1(n770), 
        .Q(n508) );
  IMUX40 U583 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n805), .S1(n785), .Q(n511) );
  MUX22 U584 ( .A(n518), .B(n513), .S(n763), .Q(o_data_Rs[7]) );
  IMUX40 U585 ( .A(n519), .B(n520), .C(n521), .D(n522), .S0(n765), .S1(n770), 
        .Q(n518) );
  IMUX40 U586 ( .A(n514), .B(n515), .C(n516), .D(n517), .S0(n765), .S1(n770), 
        .Q(n513) );
  IMUX40 U587 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n810), .S1(n786), .Q(n521) );
  MUX22 U588 ( .A(n528), .B(n523), .S(n763), .Q(o_data_Rs[8]) );
  IMUX40 U589 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n813), .S1(n787), .Q(n531) );
  BUF2 U590 ( .A(i_addr_Rs[1]), .Q(n804) );
  BUF2 U591 ( .A(i_addr_Rs[1]), .Q(n803) );
  MUX22 U592 ( .A(n538), .B(n533), .S(n763), .Q(o_data_Rs[9]) );
  IMUX40 U593 ( .A(n539), .B(n540), .C(n541), .D(n542), .S0(i_addr_Rs[3]), 
        .S1(n771), .Q(n538) );
  IMUX40 U594 ( .A(n534), .B(n535), .C(n536), .D(n537), .S0(i_addr_Rs[3]), 
        .S1(n770), .Q(n533) );
  IMUX40 U595 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n808), .S1(n789), .Q(n541) );
  MUX22 U596 ( .A(n548), .B(n543), .S(i_addr_Rs[4]), .Q(o_data_Rs[10]) );
  IMUX40 U597 ( .A(n549), .B(n550), .C(n551), .D(n552), .S0(n765), .S1(n771), 
        .Q(n548) );
  IMUX40 U598 ( .A(n544), .B(n545), .C(n546), .D(n547), .S0(n767), .S1(n771), 
        .Q(n543) );
  IMUX40 U599 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n808), .S1(n788), .Q(n551) );
  MUX22 U600 ( .A(n558), .B(n553), .S(i_addr_Rs[4]), .Q(o_data_Rs[11]) );
  IMUX40 U601 ( .A(n559), .B(n560), .C(n561), .D(n562), .S0(n765), .S1(n771), 
        .Q(n558) );
  IMUX40 U602 ( .A(n554), .B(n555), .C(n556), .D(n557), .S0(n765), .S1(n771), 
        .Q(n553) );
  IMUX40 U603 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n808), .S1(n789), .Q(n561) );
  MUX22 U604 ( .A(n568), .B(n563), .S(i_addr_Rs[4]), .Q(o_data_Rs[12]) );
  IMUX40 U605 ( .A(n569), .B(n570), .C(n571), .D(n572), .S0(n767), .S1(n771), 
        .Q(n568) );
  IMUX40 U606 ( .A(n564), .B(n565), .C(n566), .D(n567), .S0(n766), .S1(n771), 
        .Q(n563) );
  IMUX40 U607 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n6), .S1(n789), .Q(n571) );
  MUX22 U608 ( .A(n578), .B(n573), .S(i_addr_Rs[4]), .Q(o_data_Rs[13]) );
  IMUX40 U609 ( .A(n579), .B(n580), .C(n581), .D(n582), .S0(n766), .S1(n771), 
        .Q(n578) );
  IMUX40 U610 ( .A(n574), .B(n575), .C(n576), .D(n577), .S0(n765), .S1(n771), 
        .Q(n573) );
  IMUX40 U611 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n6), .S1(n790), .Q(n581) );
  MUX22 U612 ( .A(n588), .B(n583), .S(i_addr_Rs[4]), .Q(o_data_Rs[14]) );
  IMUX40 U613 ( .A(n589), .B(n590), .C(n591), .D(n592), .S0(n766), .S1(n772), 
        .Q(n588) );
  IMUX40 U614 ( .A(n584), .B(n585), .C(n586), .D(n587), .S0(n766), .S1(n772), 
        .Q(n583) );
  IMUX40 U615 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n9), .S1(n791), .Q(n591) );
  MUX22 U616 ( .A(n598), .B(n593), .S(n763), .Q(o_data_Rs[15]) );
  IMUX40 U617 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n2), .S1(n792), .Q(n601) );
  MUX22 U618 ( .A(n608), .B(n603), .S(i_addr_Rs[4]), .Q(o_data_Rs[16]) );
  IMUX40 U619 ( .A(n609), .B(n610), .C(n611), .D(n612), .S0(n766), .S1(n772), 
        .Q(n608) );
  IMUX40 U620 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n2), .S1(n793), .Q(n611) );
  MUX22 U621 ( .A(n618), .B(n613), .S(n763), .Q(o_data_Rs[17]) );
  IMUX40 U622 ( .A(n619), .B(n620), .C(n621), .D(n622), .S0(n766), .S1(n772), 
        .Q(n618) );
  IMUX40 U623 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n9), .S1(n794), .Q(n621) );
  MUX22 U624 ( .A(n628), .B(n623), .S(n763), .Q(o_data_Rs[18]) );
  IMUX40 U625 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n8), .S1(n792), .Q(n631) );
  MUX22 U626 ( .A(n638), .B(n633), .S(n764), .Q(o_data_Rs[19]) );
  IMUX40 U627 ( .A(n639), .B(n640), .C(n641), .D(n642), .S0(n766), .S1(n773), 
        .Q(n638) );
  IMUX40 U628 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n9), .S1(n795), .Q(n641) );
  MUX22 U629 ( .A(n648), .B(n643), .S(n764), .Q(o_data_Rs[20]) );
  IMUX40 U630 ( .A(n649), .B(n650), .C(n651), .D(n652), .S0(n767), .S1(n773), 
        .Q(n648) );
  IMUX40 U631 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n1), .S1(n796), .Q(n651) );
  MUX22 U632 ( .A(n658), .B(n653), .S(n764), .Q(o_data_Rs[21]) );
  IMUX40 U633 ( .A(n659), .B(n660), .C(n661), .D(n662), .S0(n767), .S1(n773), 
        .Q(n658) );
  IMUX40 U634 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n9), .S1(n796), .Q(n661) );
  MUX22 U635 ( .A(n668), .B(n663), .S(n764), .Q(o_data_Rs[22]) );
  IMUX40 U636 ( .A(n669), .B(n670), .C(n671), .D(n672), .S0(n767), .S1(n773), 
        .Q(n668) );
  IMUX40 U637 ( .A(n664), .B(n665), .C(n666), .D(n667), .S0(n767), .S1(n773), 
        .Q(n663) );
  IMUX40 U638 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n9), .S1(n797), .Q(n671) );
  MUX22 U639 ( .A(n678), .B(n673), .S(n764), .Q(o_data_Rs[23]) );
  IMUX40 U640 ( .A(n679), .B(n680), .C(n681), .D(n682), .S0(n767), .S1(
        i_addr_Rs[2]), .Q(n678) );
  IMUX40 U641 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n805), .S1(n798), .Q(n681) );
  MUX22 U642 ( .A(n688), .B(n683), .S(n764), .Q(o_data_Rs[24]) );
  IMUX40 U643 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n811), .S1(n796), .Q(n691) );
  MUX22 U644 ( .A(n698), .B(n693), .S(n764), .Q(o_data_Rs[25]) );
  IMUX40 U645 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n811), .S1(n799), .Q(n701) );
  MUX22 U646 ( .A(n708), .B(n703), .S(n764), .Q(o_data_Rs[26]) );
  IMUX40 U647 ( .A(n709), .B(n710), .C(n711), .D(n712), .S0(n768), .S1(
        i_addr_Rs[2]), .Q(n708) );
  IMUX40 U648 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n807), .S1(n800), .Q(n711) );
  MUX22 U649 ( .A(n718), .B(n713), .S(n764), .Q(o_data_Rs[27]) );
  IMUX40 U650 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n6), .S1(n801), .Q(n721) );
  IMUX40 U651 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n2), .S1(n802), .Q(n731) );
  MUX22 U652 ( .A(n738), .B(n733), .S(n764), .Q(o_data_Rs[29]) );
  IMUX40 U653 ( .A(n739), .B(n740), .C(n741), .D(n742), .S0(n768), .S1(n772), 
        .Q(n738) );
  IMUX40 U654 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n812), .S1(n785), .Q(n741) );
  MUX22 U655 ( .A(n748), .B(n743), .S(n764), .Q(o_data_Rs[30]) );
  IMUX40 U656 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n813), .S1(n786), .Q(n751) );
  MUX22 U657 ( .A(n758), .B(n753), .S(n764), .Q(o_data_Rs[31]) );
  IMUX40 U658 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n813), .S1(n783), .Q(n761) );
  NOR31 U659 ( .A(n964), .B(i_addr_Rd[3]), .C(n985), .Q(n74) );
  NOR31 U660 ( .A(i_addr_Rd[3]), .B(i_addr_Rd[4]), .C(n985), .Q(n54) );
  NOR31 U661 ( .A(n981), .B(i_addr_Rd[4]), .C(n985), .Q(n65) );
  NOR31 U662 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(n984), .Q(n57) );
  NOR31 U663 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n982), .Q(n46) );
  NOR31 U664 ( .A(n984), .B(i_addr_Rd[1]), .C(n982), .Q(n48) );
  NOR31 U665 ( .A(n983), .B(i_addr_Rd[0]), .C(n982), .Q(n50) );
  NOR31 U666 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(i_addr_Rd[0]), .Q(n55)
         );
  NOR31 U667 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[2]), .C(n983), .Q(n41) );
  NOR31 U668 ( .A(n984), .B(i_addr_Rd[2]), .C(n983), .Q(n44) );
  IMUX40 U669 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n417), .S1(n396), .Q(n20) );
  IMUX40 U670 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n417), .S1(n396), .Q(n18) );
  IMUX40 U671 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n417), .S1(n396), .Q(n17) );
  IMUX40 U672 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(n421), .S1(n396), .Q(n15) );
  IMUX40 U673 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(n420), .S1(n396), .Q(n13) );
  IMUX40 U674 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(n422), .S1(n407), .Q(n12) );
  IMUX40 U675 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n417), .S1(n396), .Q(n25) );
  IMUX40 U676 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n417), .S1(n396), .Q(n23) );
  IMUX40 U677 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n417), .S1(n396), .Q(n22) );
  IMUX40 U678 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n417), .S1(n396), .Q(n30) );
  IMUX40 U679 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n417), .S1(n396), .Q(n28) );
  IMUX40 U680 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n418), .S1(n392), .Q(n35) );
  IMUX40 U681 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n418), .S1(n391), .Q(n33) );
  IMUX40 U682 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n418), .S1(n401), .Q(n32) );
  IMUX40 U683 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n418), .S1(n415), .Q(n84) );
  IMUX40 U684 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n418), .S1(n400), .Q(n38) );
  IMUX40 U685 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n418), .S1(n415), .Q(n89) );
  IMUX40 U686 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n418), .S1(n399), .Q(n87) );
  IMUX40 U687 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n418), .S1(i_addr_Rt[1]), .Q(n86) );
  IMUX40 U688 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n419), .S1(n416), .Q(n94) );
  IMUX40 U689 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n419), .S1(n415), .Q(n92) );
  IMUX40 U690 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n419), .S1(n414), .Q(n99) );
  IMUX40 U691 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n419), .S1(n390), .Q(n97) );
  IMUX40 U692 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n419), .S1(n401), .Q(n96) );
  IMUX40 U693 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n419), .S1(n404), .Q(n104) );
  IMUX40 U694 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n419), .S1(n400), .Q(n102) );
  IMUX40 U695 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n420), .S1(n398), .Q(n109) );
  IMUX40 U696 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n420), .S1(n413), .Q(n107) );
  IMUX40 U697 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n420), .S1(n406), .Q(n106) );
  IMUX40 U698 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n420), .S1(n414), .Q(n114) );
  IMUX40 U699 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n420), .S1(n405), .Q(n112) );
  IMUX40 U700 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n420), .S1(n412), .Q(n119) );
  IMUX40 U701 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n420), .S1(n397), .Q(n117) );
  IMUX40 U702 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n420), .S1(n397), .Q(n116) );
  IMUX40 U703 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n421), .S1(n397), .Q(n124) );
  IMUX40 U704 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n421), .S1(n397), .Q(n122) );
  IMUX40 U705 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n421), .S1(n397), .Q(n129) );
  IMUX40 U706 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n421), .S1(n397), .Q(n127) );
  IMUX40 U707 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n421), .S1(n398), .Q(n126) );
  IMUX40 U708 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n421), .S1(n398), .Q(n134) );
  IMUX40 U709 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n421), .S1(n398), .Q(n132) );
  IMUX40 U710 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n422), .S1(n398), .Q(n139) );
  IMUX40 U711 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n422), .S1(n398), .Q(n137) );
  IMUX40 U712 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n422), .S1(n399), .Q(n136) );
  IMUX40 U713 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n422), .S1(n399), .Q(n144) );
  IMUX40 U714 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n422), .S1(n399), .Q(n142) );
  IMUX40 U715 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n422), .S1(n399), .Q(n149) );
  IMUX40 U716 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n422), .S1(n399), .Q(n147) );
  IMUX40 U717 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n422), .S1(n399), .Q(n146) );
  IMUX40 U718 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n423), .S1(n400), .Q(n154) );
  IMUX40 U719 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n423), .S1(n400), .Q(n152) );
  IMUX40 U720 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n423), .S1(n400), .Q(n159) );
  IMUX40 U721 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n423), .S1(n400), .Q(n157) );
  IMUX40 U722 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n423), .S1(n400), .Q(n156) );
  IMUX40 U723 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n423), .S1(n400), .Q(n164) );
  IMUX40 U724 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n423), .S1(n401), .Q(n162) );
  IMUX40 U725 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n424), .S1(n401), .Q(n169) );
  IMUX40 U726 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n424), .S1(n401), .Q(n167) );
  IMUX40 U727 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n424), .S1(n401), .Q(n166) );
  IMUX40 U728 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n424), .S1(n401), .Q(n174) );
  IMUX40 U729 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n424), .S1(n401), .Q(n172) );
  IMUX40 U730 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n424), .S1(n402), .Q(n179) );
  IMUX40 U731 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n424), .S1(n402), .Q(n177) );
  IMUX40 U732 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n424), .S1(n402), .Q(n176) );
  IMUX40 U733 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n425), .S1(n402), .Q(n184) );
  IMUX40 U734 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n425), .S1(n402), .Q(n182) );
  IMUX40 U735 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n425), .S1(n403), .Q(n189) );
  IMUX40 U736 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n425), .S1(n403), .Q(n187) );
  IMUX40 U737 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n425), .S1(n403), .Q(n186) );
  IMUX40 U738 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n425), .S1(n403), .Q(n194) );
  IMUX40 U739 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n425), .S1(n403), .Q(n192) );
  IMUX40 U740 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n426), .S1(n404), .Q(n199) );
  IMUX40 U741 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n426), .S1(n404), .Q(n197) );
  IMUX40 U742 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n426), .S1(n404), .Q(n196) );
  IMUX40 U743 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n426), .S1(n404), .Q(n204) );
  IMUX40 U744 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n426), .S1(n404), .Q(n202) );
  IMUX40 U745 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n426), .S1(n404), .Q(n209) );
  IMUX40 U746 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n426), .S1(n405), .Q(n207) );
  IMUX40 U747 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n426), .S1(n405), .Q(n206) );
  IMUX40 U748 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n427), .S1(n405), .Q(n214) );
  IMUX40 U749 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n427), .S1(n405), .Q(n212) );
  IMUX40 U750 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n427), .S1(n405), .Q(n219) );
  IMUX40 U751 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n427), .S1(n405), .Q(n217) );
  IMUX40 U752 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n427), .S1(n406), .Q(n216) );
  IMUX40 U753 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n427), .S1(n406), .Q(n224) );
  IMUX40 U754 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n427), .S1(n406), .Q(n222) );
  IMUX40 U755 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n428), .S1(n406), .Q(n229) );
  IMUX40 U756 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n428), .S1(n406), .Q(n227) );
  IMUX40 U757 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n428), .S1(n407), .Q(n226) );
  IMUX40 U758 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n428), .S1(n407), .Q(n234) );
  IMUX40 U759 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n428), .S1(n407), .Q(n232) );
  IMUX40 U760 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n428), .S1(n407), .Q(n239) );
  IMUX40 U761 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n428), .S1(n407), .Q(n237) );
  IMUX40 U762 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n428), .S1(n407), .Q(n236) );
  IMUX40 U763 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n429), .S1(n408), .Q(n244) );
  IMUX40 U764 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n429), .S1(n408), .Q(n242) );
  IMUX40 U765 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n429), .S1(n408), .Q(n249) );
  IMUX40 U766 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n429), .S1(n408), .Q(n247) );
  IMUX40 U767 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n429), .S1(n408), .Q(n246) );
  IMUX40 U768 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n429), .S1(n408), .Q(n254) );
  IMUX40 U769 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n429), .S1(n409), .Q(n252) );
  IMUX40 U770 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n430), .S1(n409), .Q(n259) );
  IMUX40 U771 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n430), .S1(n409), .Q(n257) );
  IMUX40 U772 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n430), .S1(n409), .Q(n256) );
  IMUX40 U773 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n430), .S1(n409), .Q(n264) );
  IMUX40 U774 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n430), .S1(n409), .Q(n262) );
  IMUX40 U775 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n430), .S1(n410), .Q(n269) );
  IMUX40 U776 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n430), .S1(n410), .Q(n267) );
  IMUX40 U777 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n430), .S1(n410), .Q(n266) );
  IMUX40 U778 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n431), .S1(n410), .Q(n274) );
  IMUX40 U779 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n431), .S1(n410), .Q(n272) );
  IMUX40 U780 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n431), .S1(n411), .Q(n279) );
  IMUX40 U781 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n431), .S1(n411), .Q(n277) );
  IMUX40 U782 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n431), .S1(n411), .Q(n276) );
  IMUX40 U783 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n431), .S1(n411), .Q(n284) );
  IMUX40 U784 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n431), .S1(n411), .Q(n282) );
  IMUX40 U785 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n432), .S1(n391), .Q(n289) );
  IMUX40 U786 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n432), .S1(n391), .Q(n287) );
  IMUX40 U787 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n432), .S1(n391), .Q(n286) );
  IMUX40 U788 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n432), .S1(n391), .Q(n294) );
  IMUX40 U789 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n432), .S1(n391), .Q(n292) );
  IMUX40 U790 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n432), .S1(n391), .Q(n299) );
  IMUX40 U791 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n432), .S1(n394), .Q(n297) );
  IMUX40 U792 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n432), .S1(n409), .Q(n296) );
  IMUX40 U793 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n433), .S1(n391), .Q(n304) );
  IMUX40 U794 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n433), .S1(n396), .Q(n302) );
  IMUX40 U795 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n433), .S1(n395), .Q(n309) );
  IMUX40 U796 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n433), .S1(n393), .Q(n307) );
  IMUX40 U797 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n433), .S1(n391), .Q(n306) );
  IMUX40 U798 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n433), .S1(n392), .Q(n314) );
  IMUX40 U799 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n433), .S1(n415), .Q(n312) );
  IMUX40 U800 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n434), .S1(n390), .Q(n319) );
  IMUX40 U801 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n434), .S1(n391), .Q(n317) );
  IMUX40 U802 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n434), .S1(n390), .Q(n316) );
  IMUX40 U803 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n434), .S1(n390), .Q(n324) );
  IMUX40 U804 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n434), .S1(n390), .Q(n322) );
  IMUX40 U805 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n434), .S1(n390), .Q(n329) );
  IMUX40 U806 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n434), .S1(n390), .Q(n327) );
  IMUX40 U807 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n434), .S1(n390), .Q(n326) );
  IMUX40 U808 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n435), .S1(n391), .Q(n334) );
  IMUX40 U809 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n435), .S1(n393), .Q(n332) );
  IMUX40 U810 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n435), .S1(n395), .Q(n339) );
  IMUX40 U811 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n435), .S1(n392), .Q(n337) );
  IMUX40 U812 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n435), .S1(n416), .Q(n336) );
  IMUX40 U813 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n435), .S1(n394), .Q(n344) );
  IMUX40 U814 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n435), .S1(n394), .Q(n342) );
  IMUX40 U815 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n436), .S1(n396), .Q(n349) );
  IMUX40 U816 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n436), .S1(n397), .Q(n347) );
  IMUX40 U817 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n436), .S1(n390), .Q(n346) );
  IMUX40 U818 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n436), .S1(n414), .Q(n354) );
  IMUX40 U819 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n436), .S1(n393), .Q(n352) );
  IMUX40 U820 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n436), .S1(n412), .Q(n359) );
  IMUX40 U821 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n436), .S1(n412), .Q(n357) );
  IMUX40 U822 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n436), .S1(n412), .Q(n356) );
  IMUX40 U823 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n437), .S1(n412), .Q(n364) );
  IMUX40 U824 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n437), .S1(n412), .Q(n362) );
  IMUX40 U825 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n437), .S1(n413), .Q(n369) );
  IMUX40 U826 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n437), .S1(n413), .Q(n367) );
  IMUX40 U827 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n437), .S1(n413), .Q(n366) );
  IMUX40 U828 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n437), .S1(n413), .Q(n374) );
  IMUX40 U829 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n437), .S1(n413), .Q(n372) );
  IMUX40 U830 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n417), .S1(n396), .Q(n19) );
  IMUX40 U831 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(n422), .S1(n397), .Q(n14) );
  IMUX40 U832 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n417), .S1(n396), .Q(n24) );
  IMUX40 U833 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n417), .S1(n408), .Q(n29) );
  IMUX40 U834 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n418), .S1(n396), .Q(n34) );
  IMUX40 U835 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n418), .S1(n394), .Q(n83) );
  IMUX40 U836 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n418), .S1(n397), .Q(n88) );
  IMUX40 U837 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n419), .S1(n393), .Q(n93) );
  IMUX40 U838 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n419), .S1(n397), .Q(n98) );
  IMUX40 U839 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n419), .S1(n395), .Q(n103) );
  IMUX40 U840 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n420), .S1(n397), .Q(n108) );
  IMUX40 U841 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n420), .S1(n391), .Q(n113) );
  IMUX40 U842 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n420), .S1(n397), .Q(n118) );
  IMUX40 U843 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n421), .S1(n397), .Q(n123) );
  IMUX40 U844 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n421), .S1(n398), .Q(n128) );
  IMUX40 U845 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n421), .S1(n398), .Q(n133) );
  IMUX40 U846 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n422), .S1(n398), .Q(n138) );
  IMUX40 U847 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n422), .S1(n399), .Q(n143) );
  IMUX40 U848 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n422), .S1(n399), .Q(n148) );
  IMUX40 U849 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n423), .S1(n400), .Q(n153) );
  IMUX40 U850 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n423), .S1(n400), .Q(n158) );
  IMUX40 U851 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n423), .S1(n401), .Q(n163) );
  IMUX40 U852 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n424), .S1(n401), .Q(n168) );
  IMUX40 U853 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n424), .S1(n402), .Q(n173) );
  IMUX40 U854 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n424), .S1(n402), .Q(n178) );
  IMUX40 U855 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n425), .S1(n402), .Q(n183) );
  IMUX40 U856 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n425), .S1(n403), .Q(n188) );
  IMUX40 U857 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n425), .S1(n403), .Q(n193) );
  IMUX40 U858 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n426), .S1(n404), .Q(n198) );
  IMUX40 U859 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n426), .S1(n404), .Q(n203) );
  IMUX40 U860 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n426), .S1(n405), .Q(n208) );
  IMUX40 U861 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n427), .S1(n405), .Q(n213) );
  IMUX40 U862 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n427), .S1(n406), .Q(n218) );
  IMUX40 U863 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n427), .S1(n406), .Q(n223) );
  IMUX40 U864 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n428), .S1(n406), .Q(n228) );
  IMUX40 U865 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n428), .S1(n407), .Q(n233) );
  IMUX40 U866 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n428), .S1(n407), .Q(n238) );
  IMUX40 U867 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n429), .S1(n408), .Q(n243) );
  IMUX40 U868 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n429), .S1(n408), .Q(n248) );
  IMUX40 U869 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n429), .S1(n409), .Q(n253) );
  IMUX40 U870 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n430), .S1(n409), .Q(n258) );
  IMUX40 U871 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n430), .S1(n410), .Q(n263) );
  IMUX40 U872 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n430), .S1(n410), .Q(n268) );
  IMUX40 U873 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n431), .S1(n410), .Q(n273) );
  IMUX40 U874 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n431), .S1(n411), .Q(n278) );
  IMUX40 U875 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n431), .S1(n411), .Q(n283) );
  IMUX40 U876 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n432), .S1(n391), .Q(n288) );
  IMUX40 U877 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n432), .S1(n391), .Q(n293) );
  IMUX40 U878 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n432), .S1(n391), .Q(n298) );
  IMUX40 U879 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n433), .S1(n416), .Q(n303) );
  IMUX40 U880 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n433), .S1(n390), .Q(n308) );
  IMUX40 U881 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n433), .S1(n397), .Q(n313) );
  IMUX40 U882 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n434), .S1(n390), .Q(n318) );
  IMUX40 U883 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n434), .S1(n390), .Q(n323) );
  IMUX40 U884 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n434), .S1(n390), .Q(n328) );
  IMUX40 U885 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n435), .S1(n391), .Q(n333) );
  IMUX40 U886 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n435), .S1(n390), .Q(n338) );
  IMUX40 U887 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n435), .S1(n396), .Q(n343) );
  IMUX40 U888 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n436), .S1(n396), .Q(n348) );
  IMUX40 U889 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n436), .S1(n412), .Q(n353) );
  IMUX40 U890 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n436), .S1(n412), .Q(n358) );
  IMUX40 U891 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n437), .S1(n412), .Q(n363) );
  IMUX40 U892 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n437), .S1(n413), .Q(n368) );
  IMUX40 U893 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n437), .S1(n413), .Q(n373) );
  BUF2 U894 ( .A(i_addr_Rt[4]), .Q(n376) );
  BUF2 U895 ( .A(i_addr_Rt[3]), .Q(n378) );
  BUF2 U896 ( .A(i_addr_Rt[3]), .Q(n379) );
  BUF2 U897 ( .A(i_addr_Rt[3]), .Q(n380) );
  BUF2 U898 ( .A(i_addr_Rt[3]), .Q(n381) );
  BUF2 U899 ( .A(i_addr_Rt[3]), .Q(n382) );
  INV3 U900 ( .A(i_addr_Rd[0]), .Q(n984) );
  INV3 U901 ( .A(i_addr_Rd[1]), .Q(n983) );
  INV3 U902 ( .A(i_addr_Rd[2]), .Q(n982) );
  INV3 U903 ( .A(i_con_RegWr), .Q(n985) );
  BUF2 U904 ( .A(i_addr_Rt[4]), .Q(n375) );
  BUF2 U905 ( .A(i_addr_Rs[4]), .Q(n763) );
  BUF2 U906 ( .A(i_addr_Rt[2]), .Q(n383) );
  BUF2 U907 ( .A(i_addr_Rt[2]), .Q(n384) );
  BUF2 U908 ( .A(i_addr_Rt[2]), .Q(n385) );
  BUF2 U909 ( .A(i_addr_Rt[2]), .Q(n386) );
  BUF2 U910 ( .A(i_addr_Rt[2]), .Q(n387) );
  BUF2 U911 ( .A(i_addr_Rt[2]), .Q(n388) );
  BUF2 U912 ( .A(i_addr_Rt[2]), .Q(n389) );
  INV3 U913 ( .A(i_addr_Rd[4]), .Q(n964) );
  INV3 U914 ( .A(i_addr_Rd[3]), .Q(n981) );
  BUF2 U915 ( .A(i_addr_Rs[2]), .Q(n769) );
  BUF2 U916 ( .A(i_addr_Rs[2]), .Q(n770) );
  BUF2 U917 ( .A(i_addr_Rs[2]), .Q(n771) );
  BUF2 U918 ( .A(i_addr_Rs[2]), .Q(n772) );
  BUF2 U919 ( .A(i_addr_Rs[2]), .Q(n773) );
  BUF2 U920 ( .A(i_addr_Rt[3]), .Q(n377) );
  BUF2 U921 ( .A(i_addr_Rt[1]), .Q(n416) );
  BUF2 U922 ( .A(i_addr_Rt[1]), .Q(n415) );
  BUF2 U923 ( .A(i_addr_Rt[1]), .Q(n414) );
  MUX22 U924 ( .A(n16), .B(n11), .S(n375), .Q(o_data_Rt[0]) );
  IMUX40 U925 ( .A(n12), .B(n13), .C(n14), .D(n15), .S0(n377), .S1(
        i_addr_Rt[2]), .Q(n11) );
  IMUX40 U926 ( .A(n17), .B(n18), .C(n19), .D(n20), .S0(n377), .S1(n383), .Q(
        n16) );
  MUX22 U927 ( .A(n26), .B(n21), .S(n375), .Q(o_data_Rt[1]) );
  IMUX40 U928 ( .A(n27), .B(n28), .C(n29), .D(n30), .S0(n377), .S1(n383), .Q(
        n26) );
  IMUX40 U929 ( .A(n22), .B(n23), .C(n24), .D(n25), .S0(n377), .S1(n383), .Q(
        n21) );
  IMUX40 U930 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n417), .S1(n402), .Q(n27) );
  MUX22 U931 ( .A(n36), .B(n31), .S(n375), .Q(o_data_Rt[2]) );
  IMUX40 U932 ( .A(n37), .B(n38), .C(n83), .D(n84), .S0(n378), .S1(n383), .Q(
        n36) );
  IMUX40 U933 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(n378), .S1(n383), .Q(
        n31) );
  IMUX40 U934 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n418), .S1(i_addr_Rt[1]), .Q(n37) );
  MUX22 U935 ( .A(n90), .B(n85), .S(n375), .Q(o_data_Rt[3]) );
  IMUX40 U936 ( .A(n91), .B(n92), .C(n93), .D(n94), .S0(n378), .S1(n383), .Q(
        n90) );
  IMUX40 U937 ( .A(n86), .B(n87), .C(n88), .D(n89), .S0(n378), .S1(n383), .Q(
        n85) );
  IMUX40 U938 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n419), .S1(n402), .Q(n91) );
  MUX22 U939 ( .A(n100), .B(n95), .S(n375), .Q(o_data_Rt[4]) );
  IMUX40 U940 ( .A(n101), .B(n102), .C(n103), .D(n104), .S0(n378), .S1(n383), 
        .Q(n100) );
  IMUX40 U941 ( .A(n96), .B(n97), .C(n98), .D(n99), .S0(n378), .S1(n383), .Q(
        n95) );
  IMUX40 U942 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n419), .S1(n403), .Q(n101) );
  MUX22 U943 ( .A(n110), .B(n105), .S(n375), .Q(o_data_Rt[5]) );
  IMUX40 U944 ( .A(n111), .B(n112), .C(n113), .D(n114), .S0(n378), .S1(n384), 
        .Q(n110) );
  IMUX40 U945 ( .A(n106), .B(n107), .C(n108), .D(n109), .S0(n378), .S1(n384), 
        .Q(n105) );
  IMUX40 U946 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n420), .S1(n414), .Q(n111) );
  MUX22 U947 ( .A(n120), .B(n115), .S(n376), .Q(o_data_Rt[6]) );
  IMUX40 U948 ( .A(n121), .B(n122), .C(n123), .D(n124), .S0(n378), .S1(n384), 
        .Q(n120) );
  IMUX40 U949 ( .A(n116), .B(n117), .C(n118), .D(n119), .S0(n378), .S1(n384), 
        .Q(n115) );
  IMUX40 U950 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n421), .S1(n397), .Q(n121) );
  MUX22 U951 ( .A(n130), .B(n125), .S(n376), .Q(o_data_Rt[7]) );
  IMUX40 U952 ( .A(n131), .B(n132), .C(n133), .D(n134), .S0(n378), .S1(n384), 
        .Q(n130) );
  IMUX40 U953 ( .A(n126), .B(n127), .C(n128), .D(n129), .S0(n378), .S1(n384), 
        .Q(n125) );
  IMUX40 U954 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n421), .S1(n398), .Q(n131) );
  MUX22 U955 ( .A(n140), .B(n135), .S(n376), .Q(o_data_Rt[8]) );
  IMUX40 U956 ( .A(n141), .B(n142), .C(n143), .D(n144), .S0(n379), .S1(n384), 
        .Q(n140) );
  IMUX40 U957 ( .A(n136), .B(n137), .C(n138), .D(n139), .S0(n379), .S1(n384), 
        .Q(n135) );
  IMUX40 U958 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n422), .S1(n399), .Q(n141) );
  MUX22 U959 ( .A(n150), .B(n145), .S(n376), .Q(o_data_Rt[9]) );
  IMUX40 U960 ( .A(n151), .B(n152), .C(n153), .D(n154), .S0(n379), .S1(n385), 
        .Q(n150) );
  IMUX40 U961 ( .A(n146), .B(n147), .C(n148), .D(n149), .S0(n379), .S1(n384), 
        .Q(n145) );
  IMUX40 U962 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n423), .S1(n400), .Q(n151) );
  MUX22 U963 ( .A(n160), .B(n155), .S(n376), .Q(o_data_Rt[10]) );
  IMUX40 U964 ( .A(n161), .B(n162), .C(n163), .D(n164), .S0(n379), .S1(n385), 
        .Q(n160) );
  IMUX40 U965 ( .A(n156), .B(n157), .C(n158), .D(n159), .S0(n379), .S1(n385), 
        .Q(n155) );
  IMUX40 U966 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n423), .S1(n401), .Q(n161) );
  MUX22 U967 ( .A(n170), .B(n165), .S(n376), .Q(o_data_Rt[11]) );
  IMUX40 U968 ( .A(n171), .B(n172), .C(n173), .D(n174), .S0(n379), .S1(n385), 
        .Q(n170) );
  IMUX40 U969 ( .A(n166), .B(n167), .C(n168), .D(n169), .S0(n379), .S1(n385), 
        .Q(n165) );
  IMUX40 U970 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n424), .S1(n402), .Q(n171) );
  MUX22 U971 ( .A(n180), .B(n175), .S(n376), .Q(o_data_Rt[12]) );
  IMUX40 U972 ( .A(n181), .B(n182), .C(n183), .D(n184), .S0(n379), .S1(n385), 
        .Q(n180) );
  IMUX40 U973 ( .A(n176), .B(n177), .C(n178), .D(n179), .S0(n379), .S1(n385), 
        .Q(n175) );
  IMUX40 U974 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n425), .S1(n403), .Q(n181) );
  MUX22 U975 ( .A(n190), .B(n185), .S(n376), .Q(o_data_Rt[13]) );
  IMUX40 U976 ( .A(n191), .B(n192), .C(n193), .D(n194), .S0(n379), .S1(n385), 
        .Q(n190) );
  IMUX40 U977 ( .A(n186), .B(n187), .C(n188), .D(n189), .S0(n379), .S1(n385), 
        .Q(n185) );
  IMUX40 U978 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n425), .S1(n403), .Q(n191) );
  MUX22 U979 ( .A(n200), .B(n195), .S(n376), .Q(o_data_Rt[14]) );
  IMUX40 U980 ( .A(n201), .B(n202), .C(n203), .D(n204), .S0(n380), .S1(n386), 
        .Q(n200) );
  IMUX40 U981 ( .A(n196), .B(n197), .C(n198), .D(n199), .S0(n380), .S1(n386), 
        .Q(n195) );
  IMUX40 U982 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n426), .S1(n404), .Q(n201) );
  MUX22 U983 ( .A(n210), .B(n205), .S(n376), .Q(o_data_Rt[15]) );
  IMUX40 U984 ( .A(n211), .B(n212), .C(n213), .D(n214), .S0(n380), .S1(n386), 
        .Q(n210) );
  IMUX40 U985 ( .A(n206), .B(n207), .C(n208), .D(n209), .S0(n380), .S1(n386), 
        .Q(n205) );
  IMUX40 U986 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n427), .S1(n405), .Q(n211) );
  MUX22 U987 ( .A(n220), .B(n215), .S(n376), .Q(o_data_Rt[16]) );
  IMUX40 U988 ( .A(n221), .B(n222), .C(n223), .D(n224), .S0(n380), .S1(n386), 
        .Q(n220) );
  IMUX40 U989 ( .A(n216), .B(n217), .C(n218), .D(n219), .S0(n380), .S1(n386), 
        .Q(n215) );
  IMUX40 U990 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n427), .S1(n406), .Q(n221) );
  MUX22 U991 ( .A(n230), .B(n225), .S(n376), .Q(o_data_Rt[17]) );
  IMUX40 U992 ( .A(n231), .B(n232), .C(n233), .D(n234), .S0(n380), .S1(n386), 
        .Q(n230) );
  IMUX40 U993 ( .A(n226), .B(n227), .C(n228), .D(n229), .S0(n380), .S1(n386), 
        .Q(n225) );
  IMUX40 U994 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n428), .S1(n407), .Q(n231) );
  MUX22 U995 ( .A(n240), .B(n235), .S(n376), .Q(o_data_Rt[18]) );
  IMUX40 U996 ( .A(n241), .B(n242), .C(n243), .D(n244), .S0(n380), .S1(n387), 
        .Q(n240) );
  IMUX40 U997 ( .A(n236), .B(n237), .C(n238), .D(n239), .S0(n380), .S1(n386), 
        .Q(n235) );
  IMUX40 U998 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n429), .S1(n408), .Q(n241) );
  MUX22 U999 ( .A(n250), .B(n245), .S(n375), .Q(o_data_Rt[19]) );
  IMUX40 U1000 ( .A(n251), .B(n252), .C(n253), .D(n254), .S0(n380), .S1(n387), 
        .Q(n250) );
  IMUX40 U1001 ( .A(n246), .B(n247), .C(n248), .D(n249), .S0(n380), .S1(n387), 
        .Q(n245) );
  IMUX40 U1002 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n429), .S1(n409), .Q(n251) );
  MUX22 U1003 ( .A(n260), .B(n255), .S(n375), .Q(o_data_Rt[20]) );
  IMUX40 U1004 ( .A(n261), .B(n262), .C(n263), .D(n264), .S0(n381), .S1(n387), 
        .Q(n260) );
  IMUX40 U1005 ( .A(n256), .B(n257), .C(n258), .D(n259), .S0(n381), .S1(n387), 
        .Q(n255) );
  IMUX40 U1006 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n430), .S1(n410), .Q(n261) );
  MUX22 U1007 ( .A(n270), .B(n265), .S(n375), .Q(o_data_Rt[21]) );
  IMUX40 U1008 ( .A(n271), .B(n272), .C(n273), .D(n274), .S0(n381), .S1(n387), 
        .Q(n270) );
  IMUX40 U1009 ( .A(n266), .B(n267), .C(n268), .D(n269), .S0(n381), .S1(n387), 
        .Q(n265) );
  IMUX40 U1010 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n431), .S1(n411), .Q(n271) );
  MUX22 U1011 ( .A(n280), .B(n275), .S(n375), .Q(o_data_Rt[22]) );
  IMUX40 U1012 ( .A(n281), .B(n282), .C(n283), .D(n284), .S0(n381), .S1(n387), 
        .Q(n280) );
  IMUX40 U1013 ( .A(n276), .B(n277), .C(n278), .D(n279), .S0(n381), .S1(n387), 
        .Q(n275) );
  IMUX40 U1014 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n431), .S1(n411), .Q(n281) );
  MUX22 U1015 ( .A(n290), .B(n285), .S(n375), .Q(o_data_Rt[23]) );
  IMUX40 U1016 ( .A(n291), .B(n292), .C(n293), .D(n294), .S0(n381), .S1(n388), 
        .Q(n290) );
  IMUX40 U1017 ( .A(n286), .B(n287), .C(n288), .D(n289), .S0(n381), .S1(n388), 
        .Q(n285) );
  IMUX40 U1018 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n432), .S1(n391), .Q(n291) );
  MUX22 U1019 ( .A(n300), .B(n295), .S(n375), .Q(o_data_Rt[24]) );
  IMUX40 U1020 ( .A(n301), .B(n302), .C(n303), .D(n304), .S0(n381), .S1(n388), 
        .Q(n300) );
  IMUX40 U1021 ( .A(n296), .B(n297), .C(n298), .D(n299), .S0(n381), .S1(n388), 
        .Q(n295) );
  IMUX40 U1022 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n433), .S1(n410), .Q(n301) );
  MUX22 U1023 ( .A(n310), .B(n305), .S(n375), .Q(o_data_Rt[25]) );
  IMUX40 U1024 ( .A(n311), .B(n312), .C(n313), .D(n314), .S0(n381), .S1(n388), 
        .Q(n310) );
  IMUX40 U1025 ( .A(n306), .B(n307), .C(n308), .D(n309), .S0(n381), .S1(n388), 
        .Q(n305) );
  IMUX40 U1026 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n433), .S1(n414), .Q(n311) );
  MUX22 U1027 ( .A(n320), .B(n315), .S(i_addr_Rt[4]), .Q(o_data_Rt[26]) );
  IMUX40 U1028 ( .A(n321), .B(n322), .C(n323), .D(n324), .S0(n382), .S1(n388), 
        .Q(n320) );
  IMUX40 U1029 ( .A(n316), .B(n317), .C(n318), .D(n319), .S0(n382), .S1(n388), 
        .Q(n315) );
  IMUX40 U1030 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n434), .S1(n390), .Q(n321) );
  MUX22 U1031 ( .A(n330), .B(n325), .S(i_addr_Rt[4]), .Q(o_data_Rt[27]) );
  IMUX40 U1032 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(n382), .S1(n389), 
        .Q(n330) );
  IMUX40 U1033 ( .A(n326), .B(n327), .C(n328), .D(n329), .S0(n382), .S1(n388), 
        .Q(n325) );
  IMUX40 U1034 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n435), .S1(n390), .Q(n331) );
  MUX22 U1035 ( .A(n340), .B(n335), .S(i_addr_Rt[4]), .Q(o_data_Rt[28]) );
  IMUX40 U1036 ( .A(n341), .B(n342), .C(n343), .D(n344), .S0(n382), .S1(n389), 
        .Q(n340) );
  IMUX40 U1037 ( .A(n336), .B(n337), .C(n338), .D(n339), .S0(n382), .S1(n389), 
        .Q(n335) );
  IMUX40 U1038 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n435), .S1(n397), .Q(n341) );
  MUX22 U1039 ( .A(n350), .B(n345), .S(i_addr_Rt[4]), .Q(o_data_Rt[29]) );
  IMUX40 U1040 ( .A(n351), .B(n352), .C(n353), .D(n354), .S0(n382), .S1(n389), 
        .Q(n350) );
  IMUX40 U1041 ( .A(n346), .B(n347), .C(n348), .D(n349), .S0(n382), .S1(n389), 
        .Q(n345) );
  IMUX40 U1042 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n436), .S1(n412), .Q(n351) );
  MUX22 U1043 ( .A(n360), .B(n355), .S(i_addr_Rt[4]), .Q(o_data_Rt[30]) );
  IMUX40 U1044 ( .A(n361), .B(n362), .C(n363), .D(n364), .S0(n382), .S1(n389), 
        .Q(n360) );
  IMUX40 U1045 ( .A(n356), .B(n357), .C(n358), .D(n359), .S0(n382), .S1(n389), 
        .Q(n355) );
  IMUX40 U1046 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n437), .S1(n413), .Q(n361) );
  MUX22 U1047 ( .A(n370), .B(n365), .S(i_addr_Rt[4]), .Q(o_data_Rt[31]) );
  IMUX40 U1048 ( .A(n371), .B(n372), .C(n373), .D(n374), .S0(n382), .S1(n389), 
        .Q(n370) );
  IMUX40 U1049 ( .A(n366), .B(n367), .C(n368), .D(n369), .S0(n382), .S1(n389), 
        .Q(n365) );
  IMUX40 U1050 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n437), .S1(n413), .Q(n371) );
endmodule


module D_shiftleft ( i_data_immE, o_data_immshiftl );
  input [15:0] i_data_immE;
  output [31:0] o_data_immshiftl;
  wire   n1;
  assign o_data_immshiftl[0] = o_data_immshiftl[1];
  assign o_data_immshiftl[31] = o_data_immshiftl[21];
  assign o_data_immshiftl[24] = o_data_immshiftl[21];
  assign o_data_immshiftl[27] = o_data_immshiftl[21];
  assign o_data_immshiftl[28] = o_data_immshiftl[19];
  assign o_data_immshiftl[25] = o_data_immshiftl[19];
  assign o_data_immshiftl[18] = o_data_immshiftl[19];
  assign o_data_immshiftl[30] = o_data_immshiftl[19];
  assign o_data_immshiftl[20] = o_data_immshiftl[19];
  assign o_data_immshiftl[29] = o_data_immshiftl[19];
  assign o_data_immshiftl[17] = o_data_immshiftl[19];
  assign o_data_immshiftl[26] = o_data_immshiftl[19];
  assign o_data_immshiftl[22] = o_data_immshiftl[19];
  assign o_data_immshiftl[23] = o_data_immshiftl[19];
  assign o_data_immshiftl[16] = i_data_immE[14];
  assign o_data_immshiftl[15] = i_data_immE[13];
  assign o_data_immshiftl[14] = i_data_immE[12];
  assign o_data_immshiftl[13] = i_data_immE[11];
  assign o_data_immshiftl[12] = i_data_immE[10];
  assign o_data_immshiftl[11] = i_data_immE[9];
  assign o_data_immshiftl[10] = i_data_immE[8];
  assign o_data_immshiftl[9] = i_data_immE[7];
  assign o_data_immshiftl[8] = i_data_immE[6];
  assign o_data_immshiftl[7] = i_data_immE[5];
  assign o_data_immshiftl[6] = i_data_immE[4];
  assign o_data_immshiftl[5] = i_data_immE[3];
  assign o_data_immshiftl[4] = i_data_immE[2];
  assign o_data_immshiftl[3] = i_data_immE[1];
  assign o_data_immshiftl[2] = i_data_immE[0];

  INV8 U2 ( .A(n1), .Q(o_data_immshiftl[19]) );
  INV3 U3 ( .A(i_data_immE[15]), .Q(n1) );
  CLKIN3 U4 ( .A(n1), .Q(o_data_immshiftl[21]) );
  LOGIC0 U5 ( .Q(o_data_immshiftl[1]) );
endmodule


module D_sign_extend ( i_data_immD, i_con_signext, o_data_immD );
  input [15:0] i_data_immD;
  output [31:0] o_data_immD;
  input i_con_signext;
  wire   n2;
  assign o_data_immD[15] = i_data_immD[15];
  assign o_data_immD[14] = i_data_immD[14];
  assign o_data_immD[13] = i_data_immD[13];
  assign o_data_immD[12] = i_data_immD[12];
  assign o_data_immD[11] = i_data_immD[11];
  assign o_data_immD[10] = i_data_immD[10];
  assign o_data_immD[9] = i_data_immD[9];
  assign o_data_immD[8] = i_data_immD[8];
  assign o_data_immD[7] = i_data_immD[7];
  assign o_data_immD[6] = i_data_immD[6];
  assign o_data_immD[5] = i_data_immD[5];
  assign o_data_immD[4] = i_data_immD[4];
  assign o_data_immD[3] = i_data_immD[3];
  assign o_data_immD[2] = i_data_immD[2];
  assign o_data_immD[1] = i_data_immD[1];
  assign o_data_immD[0] = i_data_immD[0];
  assign o_data_immD[16] = o_data_immD[31];
  assign o_data_immD[17] = o_data_immD[31];
  assign o_data_immD[18] = o_data_immD[31];
  assign o_data_immD[19] = o_data_immD[31];
  assign o_data_immD[20] = o_data_immD[31];
  assign o_data_immD[21] = o_data_immD[31];
  assign o_data_immD[22] = o_data_immD[31];
  assign o_data_immD[23] = o_data_immD[31];
  assign o_data_immD[24] = o_data_immD[31];
  assign o_data_immD[25] = o_data_immD[31];
  assign o_data_immD[26] = o_data_immD[31];
  assign o_data_immD[27] = o_data_immD[31];
  assign o_data_immD[28] = o_data_immD[31];
  assign o_data_immD[29] = o_data_immD[31];
  assign o_data_immD[30] = o_data_immD[31];

  INV6 U2 ( .A(n2), .Q(o_data_immD[31]) );
  NAND22 U3 ( .A(i_con_signext), .B(i_data_immD[15]), .Q(n2) );
endmodule


module D_jump_ext ( i_addr_j, i_PC4_j, o_addr_j );
  input [25:0] i_addr_j;
  input [3:0] i_PC4_j;
  output [31:0] o_addr_j;

  assign o_addr_j[0] = o_addr_j[1];
  assign o_addr_j[31] = i_PC4_j[3];
  assign o_addr_j[30] = i_PC4_j[2];
  assign o_addr_j[29] = i_PC4_j[1];
  assign o_addr_j[28] = i_PC4_j[0];
  assign o_addr_j[27] = i_addr_j[25];
  assign o_addr_j[26] = i_addr_j[24];
  assign o_addr_j[25] = i_addr_j[23];
  assign o_addr_j[24] = i_addr_j[22];
  assign o_addr_j[23] = i_addr_j[21];
  assign o_addr_j[22] = i_addr_j[20];
  assign o_addr_j[21] = i_addr_j[19];
  assign o_addr_j[20] = i_addr_j[18];
  assign o_addr_j[19] = i_addr_j[17];
  assign o_addr_j[18] = i_addr_j[16];
  assign o_addr_j[17] = i_addr_j[15];
  assign o_addr_j[16] = i_addr_j[14];
  assign o_addr_j[15] = i_addr_j[13];
  assign o_addr_j[14] = i_addr_j[12];
  assign o_addr_j[13] = i_addr_j[11];
  assign o_addr_j[12] = i_addr_j[10];
  assign o_addr_j[11] = i_addr_j[9];
  assign o_addr_j[10] = i_addr_j[8];
  assign o_addr_j[9] = i_addr_j[7];
  assign o_addr_j[8] = i_addr_j[6];
  assign o_addr_j[7] = i_addr_j[5];
  assign o_addr_j[6] = i_addr_j[4];
  assign o_addr_j[5] = i_addr_j[3];
  assign o_addr_j[4] = i_addr_j[2];
  assign o_addr_j[3] = i_addr_j[1];
  assign o_addr_j[2] = i_addr_j[0];

  LOGIC0 U2 ( .Q(o_addr_j[1]) );
endmodule


module E_forward ( i_addr_rs, i_addr_rt, i_addr_rdM, i_addr_rdW, i_addr_rtM, 
        i_addr_rtW, i_con_regwriteM, i_con_regwriteW, i_con_memreadM, 
        i_con_memreadW, o_con_fa, o_con_fb, o_con_cmpalu, o_con_cmpmem );
  input [4:0] i_addr_rs;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rdM;
  input [4:0] i_addr_rdW;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  output [2:0] o_con_fa;
  output [2:0] o_con_fb;
  input i_con_regwriteM, i_con_regwriteW, i_con_memreadM, i_con_memreadW;
  output o_con_cmpalu, o_con_cmpmem;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87;

  XOR21 U1 ( .A(n3), .B(i_addr_rdM[1]), .Q(n1) );
  INV3 U2 ( .A(n29), .Q(n40) );
  XNR20 U3 ( .A(i_addr_rs[0]), .B(i_addr_rdM[0]), .Q(n86) );
  NOR31 U4 ( .A(n41), .B(o_con_fa[2]), .C(n40), .Q(o_con_fa[1]) );
  XNR21 U5 ( .A(i_addr_rs[2]), .B(i_addr_rdM[2]), .Q(n87) );
  NAND41 U6 ( .A(n73), .B(n74), .C(n75), .D(n76), .Q(n44) );
  NOR30 U7 ( .A(n19), .B(n40), .C(n18), .Q(o_con_cmpalu) );
  OAI310 U8 ( .A(i_addr_rdM[1]), .B(i_addr_rdM[0]), .C(n27), .D(
        i_con_regwriteM), .Q(n41) );
  INV2 U9 ( .A(i_addr_rs[3]), .Q(n6) );
  INV1 U10 ( .A(i_addr_rs[1]), .Q(n4) );
  XNR20 U11 ( .A(n2), .B(i_addr_rdW[0]), .Q(n32) );
  NOR40 U12 ( .A(i_addr_rs[4]), .B(i_addr_rs[3]), .C(i_addr_rs[2]), .D(n8), 
        .Q(n19) );
  NOR40 U13 ( .A(n17), .B(n16), .C(n15), .D(n1), .Q(n29) );
  INV3 U14 ( .A(i_addr_rs[0]), .Q(n2) );
  INV3 U15 ( .A(n4), .Q(n3) );
  NAND41 U16 ( .A(n14), .B(n13), .C(n12), .D(n11), .Q(n26) );
  NAND41 U17 ( .A(n25), .B(n24), .C(n23), .D(n22), .Q(n39) );
  NOR40 U18 ( .A(n10), .B(n9), .C(n42), .D(n19), .Q(n11) );
  NOR40 U19 ( .A(n21), .B(n20), .C(n62), .D(n19), .Q(n22) );
  INV3 U20 ( .A(n59), .Q(n27) );
  AOI211 U21 ( .A(n30), .B(n29), .C(n28), .Q(n36) );
  IMUX21 U22 ( .A(n60), .B(i_addr_rs[4]), .S(i_addr_rdW[4]), .Q(n28) );
  AOI211 U23 ( .A(n70), .B(i_con_memreadM), .C(n43), .Q(n49) );
  NAND41 U24 ( .A(i_con_regwriteW), .B(n37), .C(n36), .D(n35), .Q(n38) );
  NOR40 U25 ( .A(n34), .B(n33), .C(n32), .D(n31), .Q(n35) );
  INV3 U26 ( .A(i_addr_rs[2]), .Q(n5) );
  INV3 U27 ( .A(i_addr_rs[4]), .Q(n7) );
  NOR31 U28 ( .A(i_addr_rt[0]), .B(i_addr_rt[1]), .C(n71), .Q(n43) );
  INV3 U29 ( .A(n44), .Q(n70) );
  CLKIN3 U30 ( .A(i_con_memreadM), .Q(n42) );
  CLKIN3 U31 ( .A(i_con_memreadW), .Q(n62) );
  CLKIN3 U32 ( .A(i_addr_rtM[1]), .Q(n79) );
  CLKIN3 U33 ( .A(i_addr_rtW[1]), .Q(n63) );
  XNR21 U34 ( .A(i_addr_rtM[4]), .B(i_addr_rs[4]), .Q(n14) );
  XNR21 U35 ( .A(i_addr_rtM[3]), .B(i_addr_rs[3]), .Q(n13) );
  XNR21 U36 ( .A(i_addr_rtM[2]), .B(i_addr_rs[2]), .Q(n12) );
  XNR21 U37 ( .A(n79), .B(n3), .Q(n10) );
  XNR21 U38 ( .A(n2), .B(i_addr_rtM[0]), .Q(n9) );
  NAND22 U39 ( .A(n2), .B(n4), .Q(n8) );
  CLKIN3 U40 ( .A(n26), .Q(o_con_cmpmem) );
  XNR21 U41 ( .A(n7), .B(i_addr_rdM[4]), .Q(n17) );
  XNR21 U42 ( .A(n6), .B(i_addr_rdM[3]), .Q(n16) );
  NAND22 U43 ( .A(n87), .B(n86), .Q(n15) );
  CLKIN3 U44 ( .A(i_con_regwriteM), .Q(n18) );
  XNR21 U45 ( .A(i_addr_rtW[4]), .B(i_addr_rs[4]), .Q(n25) );
  XNR21 U46 ( .A(i_addr_rtW[3]), .B(i_addr_rs[3]), .Q(n24) );
  XNR21 U47 ( .A(i_addr_rtW[2]), .B(i_addr_rs[2]), .Q(n23) );
  XNR21 U48 ( .A(n63), .B(n3), .Q(n21) );
  XNR21 U49 ( .A(n2), .B(i_addr_rtW[0]), .Q(n20) );
  NAND22 U50 ( .A(n39), .B(n26), .Q(o_con_fa[2]) );
  CLKIN3 U51 ( .A(o_con_fa[2]), .Q(n37) );
  CLKIN3 U52 ( .A(n41), .Q(n30) );
  XNR21 U53 ( .A(n5), .B(i_addr_rdW[2]), .Q(n34) );
  XNR21 U54 ( .A(n4), .B(i_addr_rdW[1]), .Q(n33) );
  XNR21 U55 ( .A(n6), .B(i_addr_rdW[3]), .Q(n31) );
  OAI212 U56 ( .A(o_con_cmpmem), .B(n39), .C(n38), .Q(o_con_fa[0]) );
  OAI310 U57 ( .A(n42), .B(n43), .C(n44), .D(n45), .Q(o_con_fb[2]) );
  OAI210 U58 ( .A(n46), .B(n47), .C(n45), .Q(o_con_fb[0]) );
  NAND30 U59 ( .A(n48), .B(n49), .C(i_con_memreadW), .Q(n45) );
  CLKIN0 U60 ( .A(n50), .Q(n48) );
  NAND40 U61 ( .A(n51), .B(n52), .C(n53), .D(n54), .Q(n47) );
  XNR20 U62 ( .A(i_addr_rt[1]), .B(i_addr_rdW[1]), .Q(n54) );
  XNR20 U63 ( .A(i_addr_rt[2]), .B(i_addr_rdW[2]), .Q(n53) );
  XNR20 U64 ( .A(i_addr_rt[3]), .B(i_addr_rdW[3]), .Q(n52) );
  XNR20 U65 ( .A(i_addr_rt[4]), .B(i_addr_rdW[4]), .Q(n51) );
  NAND40 U66 ( .A(n55), .B(i_con_regwriteW), .C(n56), .D(n57), .Q(n46) );
  CLKIN0 U67 ( .A(n58), .Q(n56) );
  XNR20 U68 ( .A(i_addr_rt[0]), .B(i_addr_rdW[0]), .Q(n55) );
  NOR30 U69 ( .A(i_addr_rdM[2]), .B(i_addr_rdM[4]), .C(i_addr_rdM[3]), .Q(n59)
         );
  NOR20 U70 ( .A(n61), .B(i_addr_rs[4]), .Q(n60) );
  NOR40 U71 ( .A(i_addr_rdW[3]), .B(i_addr_rdW[2]), .C(i_addr_rdW[1]), .D(
        i_addr_rdW[0]), .Q(n61) );
  NOR20 U72 ( .A(n58), .B(n57), .Q(o_con_fb[1]) );
  NAND40 U73 ( .A(n64), .B(i_con_regwriteM), .C(n65), .D(n66), .Q(n57) );
  NOR30 U74 ( .A(n67), .B(n68), .C(n69), .Q(n66) );
  XOR20 U75 ( .A(i_addr_rdM[2]), .B(i_addr_rt[2]), .Q(n69) );
  XOR20 U76 ( .A(i_addr_rdM[4]), .B(i_addr_rt[4]), .Q(n68) );
  XOR20 U77 ( .A(i_addr_rdM[3]), .B(i_addr_rt[3]), .Q(n67) );
  XNR20 U78 ( .A(i_addr_rt[0]), .B(i_addr_rdM[0]), .Q(n65) );
  XNR20 U79 ( .A(i_addr_rt[1]), .B(i_addr_rdM[1]), .Q(n64) );
  OAI210 U80 ( .A(n50), .B(n62), .C(n49), .Q(n58) );
  CLKIN0 U81 ( .A(n72), .Q(n71) );
  NOR30 U82 ( .A(i_addr_rt[2]), .B(i_addr_rt[4]), .C(i_addr_rt[3]), .Q(n72) );
  XNR20 U83 ( .A(i_addr_rt[0]), .B(i_addr_rtM[0]), .Q(n76) );
  NOR20 U84 ( .A(n77), .B(n78), .Q(n75) );
  XOR20 U85 ( .A(i_addr_rtM[3]), .B(i_addr_rt[3]), .Q(n78) );
  XNR20 U86 ( .A(n79), .B(i_addr_rt[1]), .Q(n77) );
  XNR20 U87 ( .A(i_addr_rt[2]), .B(i_addr_rtM[2]), .Q(n74) );
  XNR20 U88 ( .A(i_addr_rt[4]), .B(i_addr_rtM[4]), .Q(n73) );
  NAND40 U89 ( .A(n80), .B(n81), .C(n82), .D(n83), .Q(n50) );
  XNR20 U90 ( .A(i_addr_rt[0]), .B(i_addr_rtW[0]), .Q(n83) );
  NOR20 U91 ( .A(n84), .B(n85), .Q(n82) );
  XOR20 U92 ( .A(i_addr_rtW[3]), .B(i_addr_rt[3]), .Q(n85) );
  XNR20 U93 ( .A(n63), .B(i_addr_rt[1]), .Q(n84) );
  XNR20 U94 ( .A(i_addr_rt[2]), .B(i_addr_rtW[2]), .Q(n81) );
  XNR20 U95 ( .A(i_addr_rt[4]), .B(i_addr_rtW[4]), .Q(n80) );
endmodule


module decode ( i_clk, i_nrst, i_addr_pc4, i_data_instr, i_con_Wregwrite, 
        i_data_Wregwrite, i_addr_Wregwrite, i_addr_Erd, i_addr_Mrd, 
        i_con_Eregwrite, i_con_Mregwrite, i_addr_rtM, i_addr_rtW, 
        i_con_memreadM, i_con_memreadW, o_data_rs, o_data_rt, o_addr_rd, 
        o_addr_rt, o_data_jr, o_con_jump, o_addr_pc4, o_addr_branch, 
        o_addr_jump, o_con_Ealuop, o_con_Ealusrc, o_con_Eregdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Wloadmux, o_con_Walupc8, 
        o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall, o_con_Ebop, 
        o_data_signext, o_con_Efamux, o_con_Efbmux, o_data_Fmemout );
  input [31:0] i_addr_pc4;
  input [31:0] i_data_instr;
  input [31:0] i_data_Wregwrite;
  input [4:0] i_addr_Wregwrite;
  input [4:0] i_addr_Erd;
  input [4:0] i_addr_Mrd;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  output [31:0] o_data_rs;
  output [31:0] o_data_rt;
  output [4:0] o_addr_rd;
  output [4:0] o_addr_rt;
  output [31:0] o_data_jr;
  output [1:0] o_con_jump;
  output [31:0] o_addr_pc4;
  output [31:0] o_addr_branch;
  output [31:0] o_addr_jump;
  output [5:0] o_con_Ealuop;
  output [1:0] o_con_Wloadmux;
  output [2:0] o_con_Ebop;
  output [31:0] o_data_signext;
  output [2:0] o_con_Efamux;
  output [2:0] o_con_Efbmux;
  output [31:0] o_data_Fmemout;
  input i_clk, i_nrst, i_con_Wregwrite, i_con_Eregwrite, i_con_Mregwrite,
         i_con_memreadM, i_con_memreadW;
  output o_con_Ealusrc, o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite,
         o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall;
  wire   control_o_con_alusrc, control_o_con_regdst, jbcon_o_con_aluPC4,
         control_o_con_memread, control_o_con_memwrite, control_o_con_memtoreg,
         control_o_con_regwrite, signext_i_con_signext, n1, n2,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4;
  wire   [31:0] regbank_o_data_Rt;
  wire   [5:0] control_o_con_aluop;
  wire   [1:0] control_o_con_loadsig;
  wire   [31:0] signext_o_data_immD;
  wire   [2:0] for_o_con_fa;
  wire   [2:0] for_o_con_fb;
  wire   [31:0] pcadd_o_addr_pcbranchE;
  wire   [2:0] jbcon_o_con_bop;
  wire   [31:2] pcadd_i_data_immshiftl;
  assign o_addr_jump[1] = o_addr_jump[0];

  DFC3 pipe_bop_reg_2_ ( .D(jbcon_o_con_bop[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[2]) );
  DFC3 pipe_bop_reg_1_ ( .D(jbcon_o_con_bop[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[1]) );
  DFC3 pipe_bop_reg_0_ ( .D(jbcon_o_con_bop[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[0]) );
  DFC3 pipe_addr_rd_reg_3_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[3]) );
  DFC3 pipe_addr_rd_reg_1_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[1]) );
  DFC3 pipe_addr_rt_reg_4_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(n1), .C(i_clk), .RN(i_nrst), .Q(o_addr_rt[0])
         );
  DFC3 pipe_addr_pc4_reg_31_ ( .D(i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_addr_pc4_reg_30_ ( .D(i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_addr_pc4_reg_29_ ( .D(i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_addr_pc4_reg_28_ ( .D(i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_addr_pc4_reg_27_ ( .D(i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_addr_pc4_reg_26_ ( .D(i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_addr_pc4_reg_25_ ( .D(i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_addr_pc4_reg_24_ ( .D(i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_addr_pc4_reg_23_ ( .D(i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_addr_pc4_reg_22_ ( .D(i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_addr_pc4_reg_21_ ( .D(i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_addr_pc4_reg_20_ ( .D(i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_addr_pc4_reg_19_ ( .D(i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_addr_pc4_reg_18_ ( .D(i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_addr_pc4_reg_17_ ( .D(i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_addr_pc4_reg_16_ ( .D(i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_addr_pc4_reg_14_ ( .D(i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_addr_pc4_reg_12_ ( .D(i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_addr_pc4_reg_8_ ( .D(i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_addr_pc4_reg_7_ ( .D(i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_addr_pc4_reg_4_ ( .D(i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_addr_pc4_reg_1_ ( .D(i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_addr_pc4_reg_0_ ( .D(i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  DFC3 pipe_con_Ealuop_reg_5_ ( .D(control_o_con_aluop[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[5]) );
  DFC3 pipe_con_Ealuop_reg_4_ ( .D(control_o_con_aluop[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[4]) );
  DFC3 pipe_con_Ealuop_reg_3_ ( .D(control_o_con_aluop[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[3]) );
  DFC3 pipe_con_Ealuop_reg_2_ ( .D(control_o_con_aluop[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[2]) );
  DFC3 pipe_con_Ealuop_reg_1_ ( .D(control_o_con_aluop[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[1]) );
  DFC3 pipe_con_Ealuop_reg_0_ ( .D(control_o_con_aluop[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[0]) );
  DFC3 pipe_con_Ealusrc_reg ( .D(control_o_con_alusrc), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Ealusrc) );
  DFC3 pipe_con_Eregdst_reg ( .D(control_o_con_regdst), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Eregdst) );
  DFC3 pipe_con_EaluPC4_reg ( .D(jbcon_o_con_aluPC4), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Walupc8) );
  DFC3 pipe_con_Mmemread_reg ( .D(control_o_con_memread), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(control_o_con_memwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wloadmux_reg_1_ ( .D(control_o_con_loadsig[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_con_Wloadmux[1]) );
  DFC3 pipe_con_Wloadmux_reg_0_ ( .D(control_o_con_loadsig[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_con_Wloadmux[0]) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(control_o_con_memtoreg), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(control_o_con_regwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wregwrite) );
  DFC3 pipe_signext_o_data_immD_reg_21_ ( .D(signext_o_data_immD[21]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[21]) );
  DFC3 pipe_signext_o_data_immD_reg_20_ ( .D(signext_o_data_immD[20]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[20]) );
  DFC3 pipe_signext_o_data_immD_reg_19_ ( .D(signext_o_data_immD[19]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[19]) );
  DFC3 pipe_signext_o_data_immD_reg_18_ ( .D(signext_o_data_immD[18]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[18]) );
  DFC3 pipe_signext_o_data_immD_reg_17_ ( .D(signext_o_data_immD[17]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[17]) );
  DFC3 pipe_signext_o_data_immD_reg_16_ ( .D(signext_o_data_immD[16]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[16]) );
  DFC3 pipe_signext_o_data_immD_reg_15_ ( .D(signext_o_data_immD[15]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[15]) );
  DFC3 pipe_signext_o_data_immD_reg_14_ ( .D(signext_o_data_immD[14]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[14]) );
  DFC3 pipe_signext_o_data_immD_reg_12_ ( .D(signext_o_data_immD[12]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[12]) );
  DFC3 pipe_signext_o_data_immD_reg_11_ ( .D(signext_o_data_immD[11]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[11]) );
  DFC3 pipe_signext_o_data_immD_reg_10_ ( .D(signext_o_data_immD[10]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[10]) );
  DFC3 pipe_signext_o_data_immD_reg_9_ ( .D(signext_o_data_immD[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[9]) );
  DFC3 pipe_signext_o_data_immD_reg_8_ ( .D(signext_o_data_immD[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[8]) );
  DFC3 pipe_signext_o_data_immD_reg_7_ ( .D(signext_o_data_immD[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[7]) );
  DFC3 pipe_signext_o_data_immD_reg_6_ ( .D(signext_o_data_immD[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[6]) );
  DFC3 pipe_signext_o_data_immD_reg_5_ ( .D(signext_o_data_immD[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[5]) );
  DFC3 pipe_signext_o_data_immD_reg_4_ ( .D(signext_o_data_immD[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[4]) );
  DFC3 pipe_signext_o_data_immD_reg_3_ ( .D(signext_o_data_immD[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[3]) );
  DFC3 pipe_signext_o_data_immD_reg_2_ ( .D(signext_o_data_immD[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[2]) );
  DFC3 pipe_signext_o_data_immD_reg_1_ ( .D(signext_o_data_immD[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[1]) );
  DFC3 pipe_signext_o_data_immD_reg_0_ ( .D(signext_o_data_immD[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[0]) );
  DFC3 pipe_con_Efbmux_reg_2_ ( .D(for_o_con_fb[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[2]) );
  DFC3 pipe_addr_branch_reg_30_ ( .D(pcadd_o_addr_pcbranchE[30]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[30]) );
  DFC3 pipe_addr_branch_reg_29_ ( .D(pcadd_o_addr_pcbranchE[29]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[29]) );
  DFC3 pipe_addr_branch_reg_18_ ( .D(pcadd_o_addr_pcbranchE[18]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[18]) );
  DFC3 pipe_addr_branch_reg_17_ ( .D(pcadd_o_addr_pcbranchE[17]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[17]) );
  DFC3 pipe_addr_branch_reg_16_ ( .D(pcadd_o_addr_pcbranchE[16]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[16]) );
  DFC3 pipe_addr_branch_reg_6_ ( .D(pcadd_o_addr_pcbranchE[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[6]) );
  DFC3 pipe_addr_branch_reg_5_ ( .D(pcadd_o_addr_pcbranchE[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[5]) );
  DFC3 pipe_addr_branch_reg_4_ ( .D(pcadd_o_addr_pcbranchE[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[4]) );
  DFC3 pipe_addr_branch_reg_3_ ( .D(pcadd_o_addr_pcbranchE[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[3]) );
  DFC3 pipe_addr_branch_reg_2_ ( .D(pcadd_o_addr_pcbranchE[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[2]) );
  DFC3 pipe_addr_branch_reg_1_ ( .D(pcadd_o_addr_pcbranchE[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[1]) );
  DFC3 pipe_addr_branch_reg_0_ ( .D(pcadd_o_addr_pcbranchE[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[0]) );
  D_control u_control ( .o_con_regdst(control_o_con_regdst), .o_con_memread(
        control_o_con_memread), .o_con_memtoreg(control_o_con_memtoreg), 
        .o_con_memwrite(control_o_con_memwrite), .o_con_alusrc(
        control_o_con_alusrc), .o_con_regwrite(control_o_con_regwrite), 
        .o_con_ifsign(signext_i_con_signext), .o_con_loadsig(
        control_o_con_loadsig), .o_con_aluop(control_o_con_aluop), 
        .i_con_instru(i_data_instr[31:26]) );
  D_jb_control u_jb_control ( .o_con_jump(o_con_jump), .o_con_bop(
        jbcon_o_con_bop), .o_con_aluPC4(jbcon_o_con_aluPC4), .o_con_ifstall(
        o_con_ifstall), .i_con_instru(i_data_instr[31:26]), .i_con_func(
        i_data_instr[5:0]), .i_con_rt(o_addr_jump[0]) );
  D_pcadd u_pcadd ( .i_addr_pcadd4E(i_addr_pc4), .i_data_immshiftl({
        pcadd_i_data_immshiftl, o_addr_jump[0], o_addr_jump[0]}), 
        .o_addr_pcbranchE(pcadd_o_addr_pcbranchE) );
  D_register_bank u_regbank ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_addr_Rs({
        i_data_instr[25:22], n2}), .i_addr_Rt({i_data_instr[20:17], n1}), 
        .i_con_RegWr(i_con_Wregwrite), .i_addr_Rd(i_addr_Wregwrite), 
        .i_data_Rd(i_data_Wregwrite), .o_data_Rs(o_data_jr), .o_data_Rt(
        regbank_o_data_Rt) );
  D_shiftleft u_sl ( .i_data_immE(i_data_instr[15:0]), .o_data_immshiftl({
        pcadd_i_data_immshiftl, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}) );
  D_sign_extend u_signext ( .i_data_immD(i_data_instr[15:0]), .i_con_signext(
        signext_i_con_signext), .o_data_immD(signext_o_data_immD) );
  D_jump_ext u_jump_ext ( .i_addr_j({i_data_instr[25:22], n2, 
        i_data_instr[20:17], n1, i_data_instr[15:0]}), .i_PC4_j(
        i_addr_pc4[31:28]), .o_addr_j({o_addr_jump[31:2], 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4}) );
  E_forward u_forward ( .i_addr_rs({i_data_instr[25:22], n2}), .i_addr_rt({
        i_data_instr[20:17], n1}), .i_addr_rdM(i_addr_Erd), .i_addr_rdW(
        i_addr_Mrd), .i_addr_rtM(i_addr_rtM), .i_addr_rtW(i_addr_rtW), 
        .i_con_regwriteM(i_con_Eregwrite), .i_con_regwriteW(i_con_Mregwrite), 
        .i_con_memreadM(i_con_memreadM), .i_con_memreadW(i_con_memreadW), 
        .o_con_fa(for_o_con_fa), .o_con_fb(for_o_con_fb) );
  DFC1 pipe_signext_o_data_immD_reg_24_ ( .D(signext_o_data_immD[24]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[24]) );
  DFC1 pipe_signext_o_data_immD_reg_13_ ( .D(signext_o_data_immD[13]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[13]) );
  DFC1 pipe_data_rs_reg_31_ ( .D(o_data_jr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[31]) );
  DFC1 pipe_data_rs_reg_30_ ( .D(o_data_jr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[30]) );
  DFC1 pipe_data_rs_reg_29_ ( .D(o_data_jr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[29]) );
  DFC1 pipe_data_rs_reg_28_ ( .D(o_data_jr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[28]) );
  DFC1 pipe_data_rs_reg_27_ ( .D(o_data_jr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[27]) );
  DFC1 pipe_data_rs_reg_26_ ( .D(o_data_jr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[26]) );
  DFC1 pipe_data_rs_reg_25_ ( .D(o_data_jr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[25]) );
  DFC1 pipe_data_rs_reg_24_ ( .D(o_data_jr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[24]) );
  DFC1 pipe_data_rs_reg_23_ ( .D(o_data_jr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[23]) );
  DFC1 pipe_data_rs_reg_22_ ( .D(o_data_jr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[22]) );
  DFC1 pipe_data_rs_reg_21_ ( .D(o_data_jr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[21]) );
  DFC1 pipe_data_rs_reg_20_ ( .D(o_data_jr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[20]) );
  DFC1 pipe_data_rs_reg_19_ ( .D(o_data_jr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[19]) );
  DFC1 pipe_data_rs_reg_18_ ( .D(o_data_jr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[18]) );
  DFC1 pipe_data_rs_reg_17_ ( .D(o_data_jr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[17]) );
  DFC1 pipe_data_rs_reg_16_ ( .D(o_data_jr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[16]) );
  DFC1 pipe_data_rs_reg_15_ ( .D(o_data_jr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[15]) );
  DFC1 pipe_data_rs_reg_14_ ( .D(o_data_jr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[14]) );
  DFC1 pipe_data_rs_reg_13_ ( .D(o_data_jr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[13]) );
  DFC1 pipe_data_rs_reg_12_ ( .D(o_data_jr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[12]) );
  DFC1 pipe_data_rs_reg_11_ ( .D(o_data_jr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[11]) );
  DFC1 pipe_data_rs_reg_10_ ( .D(o_data_jr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[10]) );
  DFC1 pipe_data_rs_reg_9_ ( .D(o_data_jr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[9]) );
  DFC1 pipe_data_rs_reg_8_ ( .D(o_data_jr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[8]) );
  DFC1 pipe_data_rs_reg_7_ ( .D(o_data_jr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[7]) );
  DFC1 pipe_data_rs_reg_6_ ( .D(o_data_jr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[6]) );
  DFC1 pipe_data_rs_reg_5_ ( .D(o_data_jr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[5]) );
  DFC1 pipe_data_rs_reg_4_ ( .D(o_data_jr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[4]) );
  DFC1 pipe_data_rs_reg_3_ ( .D(o_data_jr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[3]) );
  DFC1 pipe_data_rs_reg_2_ ( .D(o_data_jr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[2]) );
  DFC1 pipe_data_rs_reg_1_ ( .D(o_data_jr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[1]) );
  DFC1 pipe_data_rs_reg_0_ ( .D(o_data_jr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[0]) );
  DFC1 pipe_data_rt_reg_31_ ( .D(regbank_o_data_Rt[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[31]) );
  DFC1 pipe_data_rt_reg_30_ ( .D(regbank_o_data_Rt[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC1 pipe_data_rt_reg_29_ ( .D(regbank_o_data_Rt[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[29]) );
  DFC1 pipe_data_rt_reg_28_ ( .D(regbank_o_data_Rt[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28]) );
  DFC1 pipe_data_rt_reg_27_ ( .D(regbank_o_data_Rt[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27]) );
  DFC1 pipe_data_rt_reg_26_ ( .D(regbank_o_data_Rt[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26]) );
  DFC1 pipe_data_rt_reg_25_ ( .D(regbank_o_data_Rt[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25]) );
  DFC1 pipe_data_rt_reg_24_ ( .D(regbank_o_data_Rt[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24]) );
  DFC1 pipe_data_rt_reg_23_ ( .D(regbank_o_data_Rt[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23]) );
  DFC1 pipe_data_rt_reg_22_ ( .D(regbank_o_data_Rt[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC1 pipe_data_rt_reg_21_ ( .D(regbank_o_data_Rt[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21]) );
  DFC1 pipe_data_rt_reg_20_ ( .D(regbank_o_data_Rt[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20]) );
  DFC1 pipe_data_rt_reg_19_ ( .D(regbank_o_data_Rt[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19]) );
  DFC1 pipe_data_rt_reg_18_ ( .D(regbank_o_data_Rt[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18]) );
  DFC1 pipe_data_rt_reg_17_ ( .D(regbank_o_data_Rt[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17]) );
  DFC1 pipe_data_rt_reg_16_ ( .D(regbank_o_data_Rt[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC1 pipe_data_rt_reg_15_ ( .D(regbank_o_data_Rt[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15]) );
  DFC1 pipe_data_rt_reg_14_ ( .D(regbank_o_data_Rt[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14]) );
  DFC1 pipe_data_rt_reg_13_ ( .D(regbank_o_data_Rt[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC1 pipe_data_rt_reg_12_ ( .D(regbank_o_data_Rt[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12]) );
  DFC1 pipe_data_rt_reg_11_ ( .D(regbank_o_data_Rt[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11]) );
  DFC1 pipe_data_rt_reg_10_ ( .D(regbank_o_data_Rt[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC1 pipe_data_rt_reg_9_ ( .D(regbank_o_data_Rt[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[9]) );
  DFC1 pipe_data_rt_reg_8_ ( .D(regbank_o_data_Rt[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[8]) );
  DFC1 pipe_data_rt_reg_7_ ( .D(regbank_o_data_Rt[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[7]) );
  DFC1 pipe_data_rt_reg_6_ ( .D(regbank_o_data_Rt[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[6]) );
  DFC1 pipe_data_rt_reg_5_ ( .D(regbank_o_data_Rt[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[5]) );
  DFC1 pipe_data_rt_reg_4_ ( .D(regbank_o_data_Rt[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[4]) );
  DFC1 pipe_data_rt_reg_3_ ( .D(regbank_o_data_Rt[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[3]) );
  DFC1 pipe_data_rt_reg_2_ ( .D(regbank_o_data_Rt[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[2]) );
  DFC1 pipe_data_rt_reg_1_ ( .D(regbank_o_data_Rt[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[1]) );
  DFC1 pipe_data_rt_reg_0_ ( .D(regbank_o_data_Rt[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[0]) );
  DFC1 pipe_memout_reg_31_ ( .D(i_data_Wregwrite[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[31]) );
  DFC1 pipe_memout_reg_30_ ( .D(i_data_Wregwrite[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[30]) );
  DFC1 pipe_memout_reg_29_ ( .D(i_data_Wregwrite[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[29]) );
  DFC1 pipe_memout_reg_28_ ( .D(i_data_Wregwrite[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[28]) );
  DFC1 pipe_memout_reg_27_ ( .D(i_data_Wregwrite[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[27]) );
  DFC1 pipe_memout_reg_26_ ( .D(i_data_Wregwrite[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[26]) );
  DFC1 pipe_memout_reg_25_ ( .D(i_data_Wregwrite[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[25]) );
  DFC1 pipe_memout_reg_24_ ( .D(i_data_Wregwrite[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[24]) );
  DFC1 pipe_memout_reg_23_ ( .D(i_data_Wregwrite[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[23]) );
  DFC1 pipe_memout_reg_22_ ( .D(i_data_Wregwrite[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[22]) );
  DFC1 pipe_memout_reg_21_ ( .D(i_data_Wregwrite[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[21]) );
  DFC1 pipe_memout_reg_20_ ( .D(i_data_Wregwrite[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[20]) );
  DFC1 pipe_memout_reg_19_ ( .D(i_data_Wregwrite[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[19]) );
  DFC1 pipe_memout_reg_18_ ( .D(i_data_Wregwrite[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[18]) );
  DFC1 pipe_memout_reg_17_ ( .D(i_data_Wregwrite[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[17]) );
  DFC1 pipe_memout_reg_16_ ( .D(i_data_Wregwrite[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[16]) );
  DFC1 pipe_memout_reg_15_ ( .D(i_data_Wregwrite[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[15]) );
  DFC1 pipe_memout_reg_14_ ( .D(i_data_Wregwrite[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[14]) );
  DFC1 pipe_memout_reg_13_ ( .D(i_data_Wregwrite[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[13]) );
  DFC1 pipe_memout_reg_12_ ( .D(i_data_Wregwrite[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[12]) );
  DFC1 pipe_memout_reg_11_ ( .D(i_data_Wregwrite[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[11]) );
  DFC1 pipe_memout_reg_10_ ( .D(i_data_Wregwrite[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[10]) );
  DFC1 pipe_memout_reg_9_ ( .D(i_data_Wregwrite[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[9]) );
  DFC1 pipe_memout_reg_8_ ( .D(i_data_Wregwrite[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[8]) );
  DFC1 pipe_memout_reg_7_ ( .D(i_data_Wregwrite[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[7]) );
  DFC1 pipe_memout_reg_6_ ( .D(i_data_Wregwrite[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[6]) );
  DFC1 pipe_memout_reg_5_ ( .D(i_data_Wregwrite[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[5]) );
  DFC1 pipe_memout_reg_4_ ( .D(i_data_Wregwrite[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[4]) );
  DFC1 pipe_memout_reg_3_ ( .D(i_data_Wregwrite[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[3]) );
  DFC1 pipe_memout_reg_2_ ( .D(i_data_Wregwrite[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[2]) );
  DFC1 pipe_memout_reg_1_ ( .D(i_data_Wregwrite[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[1]) );
  DFC1 pipe_memout_reg_0_ ( .D(i_data_Wregwrite[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[0]) );
  DFC1 pipe_con_Efamux_reg_2_ ( .D(for_o_con_fa[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[2]) );
  DFC1 pipe_con_Efamux_reg_0_ ( .D(for_o_con_fa[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[0]) );
  DFC1 pipe_con_Efbmux_reg_0_ ( .D(for_o_con_fb[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[0]) );
  DFC1 pipe_con_Efamux_reg_1_ ( .D(for_o_con_fa[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[1]) );
  DFC1 pipe_con_Efbmux_reg_1_ ( .D(for_o_con_fb[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[1]) );
  DFC1 pipe_addr_branch_reg_31_ ( .D(pcadd_o_addr_pcbranchE[31]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[31]) );
  DFC1 pipe_addr_branch_reg_28_ ( .D(pcadd_o_addr_pcbranchE[28]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[28]) );
  DFC1 pipe_addr_branch_reg_27_ ( .D(pcadd_o_addr_pcbranchE[27]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[27]) );
  DFC1 pipe_addr_branch_reg_26_ ( .D(pcadd_o_addr_pcbranchE[26]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[26]) );
  DFC1 pipe_addr_branch_reg_25_ ( .D(pcadd_o_addr_pcbranchE[25]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[25]) );
  DFC1 pipe_addr_branch_reg_24_ ( .D(pcadd_o_addr_pcbranchE[24]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[24]) );
  DFC1 pipe_addr_branch_reg_22_ ( .D(pcadd_o_addr_pcbranchE[22]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[22]) );
  DFC1 pipe_addr_branch_reg_19_ ( .D(pcadd_o_addr_pcbranchE[19]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[19]) );
  DFC1 pipe_addr_branch_reg_15_ ( .D(pcadd_o_addr_pcbranchE[15]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[15]) );
  DFC1 pipe_signext_o_data_immD_reg_30_ ( .D(signext_o_data_immD[30]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[30]) );
  DFC1 pipe_signext_o_data_immD_reg_29_ ( .D(signext_o_data_immD[29]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[29]) );
  DFC1 pipe_signext_o_data_immD_reg_31_ ( .D(signext_o_data_immD[31]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[31]) );
  DFC1 pipe_signext_o_data_immD_reg_23_ ( .D(signext_o_data_immD[23]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[23]) );
  DFC1 pipe_signext_o_data_immD_reg_26_ ( .D(signext_o_data_immD[26]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[26]) );
  DFC1 pipe_signext_o_data_immD_reg_22_ ( .D(signext_o_data_immD[22]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[22]) );
  DFC1 pipe_signext_o_data_immD_reg_28_ ( .D(signext_o_data_immD[28]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[28]) );
  DFC1 pipe_signext_o_data_immD_reg_27_ ( .D(signext_o_data_immD[27]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[27]) );
  DFC1 pipe_signext_o_data_immD_reg_25_ ( .D(signext_o_data_immD[25]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[25]) );
  DFC1 pipe_addr_branch_reg_8_ ( .D(pcadd_o_addr_pcbranchE[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[8]) );
  DFC1 pipe_addr_branch_reg_7_ ( .D(pcadd_o_addr_pcbranchE[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[7]) );
  DFC1 pipe_addr_branch_reg_21_ ( .D(pcadd_o_addr_pcbranchE[21]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[21]) );
  DFC1 pipe_addr_branch_reg_20_ ( .D(pcadd_o_addr_pcbranchE[20]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[20]) );
  DFC1 pipe_addr_branch_reg_14_ ( .D(pcadd_o_addr_pcbranchE[14]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[14]) );
  DFC1 pipe_addr_branch_reg_13_ ( .D(pcadd_o_addr_pcbranchE[13]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[13]) );
  DFC1 pipe_addr_branch_reg_12_ ( .D(pcadd_o_addr_pcbranchE[12]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[12]) );
  DFC1 pipe_addr_branch_reg_11_ ( .D(pcadd_o_addr_pcbranchE[11]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[11]) );
  DFC1 pipe_addr_branch_reg_10_ ( .D(pcadd_o_addr_pcbranchE[10]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[10]) );
  DFC1 pipe_addr_branch_reg_9_ ( .D(pcadd_o_addr_pcbranchE[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[9]) );
  DFC1 pipe_addr_pc4_reg_15_ ( .D(i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC1 pipe_addr_pc4_reg_13_ ( .D(i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC1 pipe_addr_pc4_reg_11_ ( .D(i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC1 pipe_addr_pc4_reg_10_ ( .D(i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC1 pipe_addr_pc4_reg_9_ ( .D(i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC1 pipe_addr_pc4_reg_6_ ( .D(i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC1 pipe_addr_pc4_reg_5_ ( .D(i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC1 pipe_addr_pc4_reg_3_ ( .D(i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC1 pipe_addr_pc4_reg_2_ ( .D(i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC1 pipe_addr_rd_reg_4_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[4]) );
  DFC1 pipe_addr_rd_reg_2_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[2]) );
  DFC1 pipe_addr_rd_reg_0_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[0]) );
  DFC1 pipe_addr_branch_reg_23_ ( .D(pcadd_o_addr_pcbranchE[23]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[23]) );
  BUF15 U3 ( .A(i_data_instr[21]), .Q(n2) );
  BUF12 U4 ( .A(i_data_instr[16]), .Q(n1) );
  LOGIC0 U5 ( .Q(o_addr_jump[0]) );
endmodule


module E_alu_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378;

  NOR23 U2 ( .A(n189), .B(n190), .Q(n179) );
  BUF2 U3 ( .A(n277), .Q(n19) );
  IMUX21 U4 ( .A(n275), .B(n276), .S(n19), .Q(SUM[16]) );
  INV4 U5 ( .A(n191), .Q(n190) );
  CLKIN6 U6 ( .A(n208), .Q(n205) );
  NOR24 U7 ( .A(B[26]), .B(A[26]), .Q(n1) );
  INV12 U8 ( .A(n1), .Q(n151) );
  BUF2 U9 ( .A(B[15]), .Q(n2) );
  CLKIN6 U10 ( .A(n245), .Q(n249) );
  NAND22 U11 ( .A(n3), .B(n4), .Q(n5) );
  NAND22 U12 ( .A(n5), .B(n245), .Q(n244) );
  INV3 U13 ( .A(A[19]), .Q(n3) );
  INV2 U14 ( .A(B[19]), .Q(n4) );
  INV12 U15 ( .A(n297), .Q(n294) );
  CLKIN3 U16 ( .A(B[12]), .Q(n49) );
  NAND26 U17 ( .A(n262), .B(n263), .Q(n245) );
  NAND23 U18 ( .A(B[2]), .B(A[2]), .Q(n91) );
  NAND23 U19 ( .A(B[1]), .B(A[1]), .Q(n365) );
  NOR24 U20 ( .A(B[24]), .B(A[24]), .Q(n212) );
  NAND22 U21 ( .A(B[0]), .B(A[0]), .Q(n257) );
  NOR22 U22 ( .A(B[4]), .B(A[4]), .Q(n87) );
  OAI2112 U23 ( .A(n67), .B(n348), .C(n349), .D(n63), .Q(n39) );
  NOR23 U24 ( .A(n184), .B(n185), .Q(n180) );
  BUF8 U25 ( .A(B[11]), .Q(n18) );
  NOR24 U26 ( .A(n108), .B(n115), .Q(n105) );
  NOR22 U27 ( .A(A[30]), .B(B[30]), .Q(n108) );
  NOR22 U28 ( .A(n250), .B(n251), .Q(n246) );
  NOR21 U29 ( .A(A[24]), .B(B[24]), .Q(n167) );
  INV3 U30 ( .A(n10), .Q(n152) );
  INV3 U31 ( .A(n108), .Q(n104) );
  NOR22 U32 ( .A(n95), .B(n257), .Q(n359) );
  NOR22 U33 ( .A(n364), .B(n91), .Q(n363) );
  NAND26 U34 ( .A(n300), .B(n301), .Q(n295) );
  NAND24 U35 ( .A(n120), .B(n121), .Q(n115) );
  NOR23 U36 ( .A(n212), .B(n154), .Q(n153) );
  INV6 U37 ( .A(n163), .Q(n183) );
  INV3 U38 ( .A(n216), .Q(n42) );
  INV3 U39 ( .A(n172), .Q(n9) );
  NAND21 U40 ( .A(B[15]), .B(A[15]), .Q(n286) );
  CLKIN10 U41 ( .A(n112), .Q(n169) );
  NAND26 U42 ( .A(n142), .B(n141), .Q(n138) );
  NAND24 U43 ( .A(n144), .B(n143), .Q(n142) );
  XOR22 U44 ( .A(n6), .B(n96), .Q(SUM[31]) );
  XOR20 U45 ( .A(B[31]), .B(A[31]), .Q(n6) );
  NAND22 U46 ( .A(B[6]), .B(A[6]), .Q(n75) );
  INV3 U47 ( .A(n188), .Q(n184) );
  CLKIN8 U48 ( .A(n99), .Q(n277) );
  XNR22 U49 ( .A(n7), .B(n213), .Q(SUM[23]) );
  XNR20 U50 ( .A(B[23]), .B(A[23]), .Q(n7) );
  CLKIN3 U51 ( .A(n192), .Q(n189) );
  XNR22 U52 ( .A(n8), .B(n258), .Q(SUM[19]) );
  XNR20 U53 ( .A(B[19]), .B(A[19]), .Q(n8) );
  CLKIN4 U54 ( .A(n132), .Q(n15) );
  INV6 U55 ( .A(n133), .Q(n31) );
  BUF2 U56 ( .A(n290), .Q(n40) );
  NOR22 U57 ( .A(A[14]), .B(B[14]), .Q(n290) );
  NAND24 U58 ( .A(n160), .B(n161), .Q(n157) );
  NAND23 U59 ( .A(n99), .B(n162), .Q(n161) );
  NAND26 U60 ( .A(n295), .B(n188), .Q(n279) );
  NAND26 U61 ( .A(n191), .B(n192), .Q(n280) );
  NOR22 U62 ( .A(n223), .B(n205), .Q(n222) );
  NAND24 U63 ( .A(n366), .B(n367), .Q(n305) );
  INV3 U64 ( .A(n49), .Q(n14) );
  BUF2 U65 ( .A(n298), .Q(n24) );
  NAND21 U66 ( .A(n24), .B(n327), .Q(n322) );
  XNR22 U67 ( .A(n9), .B(n173), .Q(SUM[25]) );
  NOR24 U68 ( .A(B[25]), .B(A[25]), .Q(n10) );
  NOR23 U69 ( .A(n112), .B(n113), .Q(n106) );
  NAND23 U70 ( .A(n48), .B(n109), .Q(n119) );
  NAND21 U71 ( .A(n325), .B(n301), .Q(n323) );
  INV12 U72 ( .A(n169), .Q(n11) );
  NAND26 U73 ( .A(n193), .B(n194), .Q(n112) );
  NAND28 U74 ( .A(n332), .B(n333), .Q(n301) );
  INV2 U75 ( .A(n62), .Q(n12) );
  INV1 U76 ( .A(n64), .Q(n62) );
  CLKIN3 U77 ( .A(n283), .Q(n282) );
  BUF2 U78 ( .A(n150), .Q(n13) );
  NOR22 U79 ( .A(A[13]), .B(B[13]), .Q(n289) );
  NAND26 U80 ( .A(n374), .B(n375), .Q(n73) );
  BUF4 U81 ( .A(n115), .Q(n48) );
  NAND21 U82 ( .A(n231), .B(n226), .Q(n227) );
  INV6 U83 ( .A(n288), .Q(n285) );
  NOR22 U84 ( .A(n51), .B(n291), .Q(n284) );
  NAND26 U85 ( .A(n103), .B(n104), .Q(n101) );
  NAND24 U86 ( .A(n131), .B(n15), .Q(n16) );
  NAND22 U87 ( .A(n132), .B(n41), .Q(n17) );
  NAND24 U88 ( .A(n16), .B(n17), .Q(SUM[29]) );
  NOR22 U89 ( .A(A[11]), .B(B[11]), .Q(n303) );
  NAND23 U90 ( .A(n86), .B(n304), .Q(n353) );
  CLKIN3 U91 ( .A(n86), .Q(n81) );
  NAND23 U92 ( .A(B[8]), .B(A[8]), .Q(n336) );
  NAND22 U93 ( .A(B[21]), .B(A[21]), .Q(n203) );
  BUF2 U94 ( .A(n75), .Q(n20) );
  INV6 U95 ( .A(B[22]), .Q(n218) );
  NOR31 U96 ( .A(n163), .B(n164), .C(n165), .Q(n162) );
  INV6 U97 ( .A(n102), .Q(n114) );
  INV12 U98 ( .A(n207), .Q(n206) );
  NAND23 U99 ( .A(B[17]), .B(A[17]), .Q(n243) );
  INV6 U100 ( .A(n75), .Q(n25) );
  AOI211 U101 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  XOR22 U102 ( .A(n70), .B(n71), .Q(SUM[7]) );
  CLKIN3 U103 ( .A(n370), .Q(n296) );
  NAND21 U104 ( .A(B[7]), .B(A[7]), .Q(n370) );
  XOR20 U105 ( .A(n79), .B(n80), .Q(SUM[5]) );
  INV6 U106 ( .A(n29), .Q(n30) );
  INV6 U107 ( .A(n305), .Q(n304) );
  NOR23 U108 ( .A(n87), .B(n369), .Q(n366) );
  NOR23 U109 ( .A(n186), .B(n187), .Q(n185) );
  NAND23 U110 ( .A(B[9]), .B(A[9]), .Q(n63) );
  INV4 U111 ( .A(n79), .Q(n78) );
  OAI221 U112 ( .A(A[9]), .B(B[9]), .C(A[10]), .D(B[10]), .Q(n340) );
  NOR22 U113 ( .A(A[9]), .B(B[9]), .Q(n64) );
  NOR20 U114 ( .A(A[15]), .B(B[15]), .Q(n283) );
  XOR22 U115 ( .A(n320), .B(n321), .Q(SUM[13]) );
  NAND21 U116 ( .A(n99), .B(n103), .Q(n122) );
  NAND28 U117 ( .A(n265), .B(n264), .Q(n259) );
  INV6 U118 ( .A(n59), .Q(n67) );
  NAND22 U119 ( .A(n221), .B(n220), .Q(n21) );
  NAND24 U120 ( .A(n220), .B(n221), .Q(n215) );
  CLKIN6 U121 ( .A(n226), .Q(n224) );
  CLKIN3 U122 ( .A(n301), .Q(n186) );
  CLKIN6 U123 ( .A(n346), .Q(n338) );
  NAND24 U124 ( .A(n359), .B(n358), .Q(n355) );
  NAND24 U125 ( .A(n114), .B(n104), .Q(n113) );
  NOR22 U126 ( .A(A[28]), .B(B[28]), .Q(n134) );
  NOR20 U127 ( .A(A[8]), .B(B[8]), .Q(n61) );
  NAND23 U128 ( .A(n99), .B(n266), .Q(n265) );
  XOR22 U129 ( .A(n116), .B(n117), .Q(SUM[30]) );
  NAND24 U130 ( .A(n299), .B(n302), .Q(n187) );
  INV2 U131 ( .A(n203), .Q(n225) );
  INV6 U132 ( .A(n259), .Q(n22) );
  INV6 U133 ( .A(n187), .Q(n300) );
  NOR24 U134 ( .A(n248), .B(n249), .Q(n247) );
  NAND28 U135 ( .A(n182), .B(n183), .Q(n124) );
  NAND28 U136 ( .A(n294), .B(n296), .Q(n188) );
  NAND20 U137 ( .A(n73), .B(n20), .Q(n76) );
  INV0 U138 ( .A(n20), .Q(n74) );
  XOR22 U139 ( .A(n343), .B(n344), .Q(SUM[11]) );
  AOI212 U140 ( .A(n39), .B(n345), .C(n338), .Q(n344) );
  NOR24 U141 ( .A(n77), .B(n368), .Q(n367) );
  CLKIN6 U142 ( .A(n73), .Q(n368) );
  NAND22 U143 ( .A(B[5]), .B(A[5]), .Q(n372) );
  BUF2 U144 ( .A(n14), .Q(n23) );
  NOR23 U145 ( .A(A[5]), .B(B[5]), .Q(n77) );
  INV0 U146 ( .A(n289), .Q(n314) );
  NOR33 U147 ( .A(n107), .B(n106), .C(n105), .Q(n97) );
  NOR33 U148 ( .A(n365), .B(n95), .C(n364), .Q(n362) );
  NOR24 U149 ( .A(n362), .B(n363), .Q(n354) );
  CLKIN3 U150 ( .A(B[6]), .Q(n374) );
  NAND22 U151 ( .A(B[14]), .B(A[14]), .Q(n287) );
  AOI312 U152 ( .A(n313), .B(n314), .C(n315), .D(n316), .Q(n312) );
  INV3 U153 ( .A(n315), .Q(n321) );
  NAND22 U154 ( .A(B[22]), .B(A[22]), .Q(n198) );
  NOR20 U155 ( .A(n268), .B(n248), .Q(n272) );
  NOR20 U156 ( .A(n267), .B(n248), .Q(n266) );
  INV12 U157 ( .A(n165), .Q(n182) );
  NAND28 U158 ( .A(n246), .B(n247), .Q(n165) );
  NOR24 U159 ( .A(n101), .B(n102), .Q(n100) );
  NAND21 U160 ( .A(n99), .B(n100), .Q(n98) );
  AOI210 U161 ( .A(n24), .B(n59), .C(n331), .Q(n330) );
  NAND24 U162 ( .A(n200), .B(n201), .Q(n195) );
  INV6 U163 ( .A(n215), .Q(n214) );
  NAND28 U164 ( .A(n52), .B(n121), .Q(n102) );
  NOR21 U165 ( .A(A[29]), .B(B[29]), .Q(n123) );
  INV3 U166 ( .A(n131), .Q(n41) );
  XOR22 U167 ( .A(n317), .B(n318), .Q(SUM[14]) );
  INV6 U168 ( .A(n124), .Q(n103) );
  NOR22 U169 ( .A(B[16]), .B(A[16]), .Q(n250) );
  NAND22 U170 ( .A(A[24]), .B(B[24]), .Q(n145) );
  NAND24 U171 ( .A(n99), .B(n222), .Q(n221) );
  NOR33 U172 ( .A(n25), .B(n26), .C(n27), .Q(n28) );
  NOR24 U173 ( .A(n373), .B(n28), .Q(n293) );
  CLKIN6 U174 ( .A(n371), .Q(n26) );
  CLKIN6 U175 ( .A(n372), .Q(n27) );
  OAI2112 U176 ( .A(A[5]), .B(B[5]), .C(B[4]), .D(A[4]), .Q(n371) );
  NAND22 U177 ( .A(n55), .B(n73), .Q(n373) );
  NAND24 U178 ( .A(n208), .B(n207), .Q(n29) );
  NAND28 U179 ( .A(n209), .B(n30), .Q(n163) );
  NAND28 U180 ( .A(n218), .B(n219), .Q(n207) );
  NAND28 U181 ( .A(n229), .B(n230), .Q(n208) );
  NOR24 U182 ( .A(n210), .B(n211), .Q(n209) );
  NAND24 U183 ( .A(n31), .B(n175), .Q(n32) );
  NAND22 U184 ( .A(n133), .B(n176), .Q(n33) );
  NAND24 U185 ( .A(n32), .B(n33), .Q(n34) );
  CLKIN6 U186 ( .A(n34), .Q(SUM[24]) );
  NAND28 U187 ( .A(n177), .B(n11), .Q(n133) );
  NAND22 U188 ( .A(n198), .B(n196), .Q(n35) );
  NAND33 U189 ( .A(n195), .B(n197), .C(n36), .Q(n194) );
  INV4 U190 ( .A(n35), .Q(n36) );
  NAND21 U191 ( .A(B[19]), .B(A[19]), .Q(n196) );
  NOR24 U192 ( .A(n37), .B(n277), .Q(n38) );
  NOR24 U193 ( .A(n38), .B(n239), .Q(n238) );
  INV1 U194 ( .A(n182), .Q(n37) );
  IMUX22 U195 ( .A(n236), .B(n237), .S(n238), .Q(SUM[20]) );
  OAI2112 U196 ( .A(A[17]), .B(B[17]), .C(B[16]), .D(A[16]), .Q(n242) );
  NAND34 U197 ( .A(n354), .B(n355), .C(n356), .Q(n86) );
  NAND28 U198 ( .A(n293), .B(n294), .Q(n191) );
  NOR24 U199 ( .A(n119), .B(n118), .Q(n117) );
  AOI212 U200 ( .A(n122), .B(n11), .C(n102), .Q(n118) );
  AOI312 U201 ( .A(n163), .B(n198), .C(n195), .D(n199), .Q(n193) );
  XNR22 U202 ( .A(n42), .B(n21), .Q(SUM[22]) );
  NAND22 U203 ( .A(B[23]), .B(A[23]), .Q(n202) );
  NOR24 U204 ( .A(A[17]), .B(B[17]), .Q(n248) );
  NAND20 U205 ( .A(n99), .B(n234), .Q(n231) );
  NAND28 U206 ( .A(n298), .B(n299), .Q(n297) );
  CLKIN6 U207 ( .A(n178), .Q(n177) );
  OAI2112 U208 ( .A(n145), .B(n10), .C(n146), .D(n147), .Q(n144) );
  NAND22 U209 ( .A(B[25]), .B(A[25]), .Q(n146) );
  NOR24 U210 ( .A(A[3]), .B(B[3]), .Q(n364) );
  CLKIN3 U211 ( .A(B[3]), .Q(n360) );
  NOR21 U212 ( .A(B[20]), .B(A[20]), .Q(n210) );
  NAND24 U213 ( .A(B[18]), .B(A[18]), .Q(n241) );
  AOI212 U214 ( .A(n148), .B(n149), .C(n1), .Q(n143) );
  XNR21 U215 ( .A(n347), .B(n39), .Q(SUM[10]) );
  XNR21 U216 ( .A(n76), .B(n72), .Q(SUM[6]) );
  AOI212 U217 ( .A(n72), .B(n73), .C(n74), .Q(n71) );
  CLKIN2 U218 ( .A(n350), .Q(n349) );
  NOR20 U219 ( .A(n303), .B(n326), .Q(n325) );
  NOR20 U220 ( .A(n126), .B(n95), .Q(n125) );
  XOR21 U221 ( .A(n157), .B(n159), .Q(SUM[26]) );
  INV3 U222 ( .A(n123), .Q(n121) );
  NAND22 U223 ( .A(B[10]), .B(A[10]), .Q(n346) );
  XOR22 U224 ( .A(n311), .B(n312), .Q(SUM[15]) );
  NOR24 U225 ( .A(A[2]), .B(B[2]), .Q(n95) );
  INV3 U226 ( .A(n228), .Q(n43) );
  NOR20 U227 ( .A(n225), .B(n205), .Q(n228) );
  NAND24 U228 ( .A(n182), .B(n233), .Q(n223) );
  NOR20 U229 ( .A(n248), .B(n270), .Q(n269) );
  NOR22 U230 ( .A(n268), .B(n269), .Q(n264) );
  CLKIN0 U231 ( .A(n267), .Q(n274) );
  NOR20 U232 ( .A(n261), .B(n249), .Q(n260) );
  NOR22 U233 ( .A(B[23]), .B(A[23]), .Q(n211) );
  OAI2112 U234 ( .A(n67), .B(n322), .C(n323), .D(n324), .Q(n315) );
  NAND21 U235 ( .A(n314), .B(n46), .Q(n320) );
  XNR22 U236 ( .A(n43), .B(n227), .Q(SUM[21]) );
  CLKIN3 U237 ( .A(n351), .Q(n348) );
  INV0 U238 ( .A(n130), .Q(n129) );
  NOR20 U239 ( .A(n186), .B(n303), .Q(n331) );
  CLKIN6 U240 ( .A(n303), .Q(n302) );
  INV1 U241 ( .A(n326), .Q(n327) );
  INV0 U242 ( .A(n61), .Q(n58) );
  INV0 U243 ( .A(B[30]), .Q(n111) );
  NOR20 U244 ( .A(A[16]), .B(B[16]), .Q(n267) );
  XOR22 U245 ( .A(n259), .B(n260), .Q(SUM[18]) );
  INV6 U246 ( .A(B[21]), .Q(n229) );
  NOR21 U247 ( .A(n158), .B(n1), .Q(n159) );
  XOR21 U248 ( .A(n93), .B(n125), .Q(SUM[2]) );
  INV3 U249 ( .A(n166), .Q(n164) );
  NOR21 U250 ( .A(n167), .B(n10), .Q(n166) );
  NAND22 U251 ( .A(n128), .B(n129), .Q(n127) );
  NOR21 U252 ( .A(n296), .B(n293), .Q(n352) );
  NAND22 U253 ( .A(n273), .B(n270), .Q(n271) );
  XOR21 U254 ( .A(n128), .B(n255), .Q(SUM[1]) );
  NAND22 U255 ( .A(n313), .B(n287), .Q(n317) );
  NAND26 U256 ( .A(n232), .B(n233), .Q(n226) );
  INV3 U257 ( .A(n167), .Q(n168) );
  NAND20 U258 ( .A(n196), .B(n197), .Q(n239) );
  NAND21 U259 ( .A(B[16]), .B(A[16]), .Q(n270) );
  INV3 U260 ( .A(A[28]), .Q(n136) );
  INV0 U261 ( .A(B[28]), .Q(n137) );
  NAND22 U262 ( .A(B[20]), .B(A[20]), .Q(n204) );
  NAND20 U263 ( .A(B[24]), .B(A[24]), .Q(n171) );
  NAND21 U264 ( .A(B[3]), .B(A[3]), .Q(n356) );
  NAND20 U265 ( .A(B[29]), .B(A[29]), .Q(n109) );
  XNR22 U266 ( .A(n44), .B(n140), .Q(SUM[28]) );
  XOR20 U267 ( .A(B[28]), .B(A[28]), .Q(n44) );
  XNR20 U268 ( .A(B[29]), .B(A[29]), .Q(n131) );
  AOI211 U269 ( .A(n308), .B(n309), .C(n310), .Q(n275) );
  INV3 U270 ( .A(A[16]), .Q(n308) );
  INV0 U271 ( .A(B[16]), .Q(n309) );
  NOR20 U272 ( .A(A[23]), .B(B[23]), .Q(n199) );
  IMUX21 U273 ( .A(n84), .B(n85), .S(n45), .Q(SUM[4]) );
  NOR21 U274 ( .A(n87), .B(n88), .Q(n84) );
  XNR20 U275 ( .A(B[16]), .B(A[16]), .Q(n276) );
  INV3 U276 ( .A(A[3]), .Q(n361) );
  INV3 U277 ( .A(A[21]), .Q(n230) );
  IMUX20 U278 ( .A(n65), .B(n66), .S(n67), .Q(SUM[8]) );
  AOI211 U279 ( .A(n68), .B(n69), .C(n60), .Q(n65) );
  INV3 U280 ( .A(A[8]), .Q(n68) );
  IMUX21 U281 ( .A(n328), .B(n329), .S(n330), .Q(SUM[12]) );
  NOR21 U282 ( .A(n341), .B(n342), .Q(n328) );
  AOI211 U283 ( .A(n252), .B(n253), .C(n254), .Q(n236) );
  INV3 U284 ( .A(A[27]), .Q(n149) );
  INV3 U285 ( .A(n235), .Q(n233) );
  NOR20 U286 ( .A(A[20]), .B(B[20]), .Q(n235) );
  XOR21 U287 ( .A(n89), .B(n90), .Q(SUM[3]) );
  NAND22 U288 ( .A(n93), .B(n94), .Q(n92) );
  INV3 U289 ( .A(A[22]), .Q(n219) );
  XNR20 U290 ( .A(B[30]), .B(A[30]), .Q(n116) );
  INV3 U291 ( .A(A[6]), .Q(n375) );
  XNR20 U292 ( .A(B[24]), .B(A[24]), .Q(n175) );
  NOR21 U293 ( .A(n212), .B(n174), .Q(n176) );
  INV3 U294 ( .A(n257), .Q(n128) );
  INV3 U295 ( .A(A[18]), .Q(n263) );
  INV0 U296 ( .A(B[0]), .Q(n376) );
  INV3 U297 ( .A(n378), .Q(n377) );
  INV3 U298 ( .A(A[20]), .Q(n252) );
  INV3 U299 ( .A(A[30]), .Q(n110) );
  INV3 U300 ( .A(A[0]), .Q(n357) );
  INV3 U301 ( .A(n40), .Q(n313) );
  OAI210 U302 ( .A(n40), .B(n46), .C(n287), .Q(n316) );
  INV3 U303 ( .A(n337), .Q(n345) );
  XNR20 U304 ( .A(B[27]), .B(A[27]), .Q(n155) );
  NAND21 U305 ( .A(B[27]), .B(A[27]), .Q(n141) );
  INV1 U306 ( .A(B[27]), .Q(n148) );
  NOR22 U307 ( .A(B[27]), .B(A[27]), .Q(n154) );
  NAND21 U308 ( .A(n99), .B(n274), .Q(n273) );
  NAND34 U309 ( .A(n196), .B(n204), .C(n197), .Q(n232) );
  NAND20 U310 ( .A(n14), .B(A[12]), .Q(n324) );
  NOR20 U311 ( .A(A[12]), .B(n14), .Q(n326) );
  NAND20 U312 ( .A(B[4]), .B(A[4]), .Q(n83) );
  NOR20 U313 ( .A(n23), .B(A[12]), .Q(n341) );
  BUF2 U314 ( .A(n81), .Q(n45) );
  NAND24 U315 ( .A(n336), .B(n63), .Q(n335) );
  NOR20 U316 ( .A(n77), .B(n27), .Q(n80) );
  NOR22 U317 ( .A(A[1]), .B(B[1]), .Q(n130) );
  NOR20 U318 ( .A(n256), .B(n130), .Q(n255) );
  BUF2 U319 ( .A(n292), .Q(n46) );
  NAND22 U320 ( .A(B[13]), .B(A[13]), .Q(n292) );
  CLKIN0 U321 ( .A(n135), .Q(n47) );
  INV6 U322 ( .A(n138), .Q(n135) );
  NAND24 U323 ( .A(n97), .B(n98), .Q(n96) );
  NAND26 U324 ( .A(n281), .B(n282), .Q(n192) );
  NOR21 U325 ( .A(n217), .B(n206), .Q(n216) );
  NAND33 U326 ( .A(n151), .B(n152), .C(n153), .Q(n150) );
  NAND20 U327 ( .A(n152), .B(n146), .Q(n172) );
  XNR20 U328 ( .A(n18), .B(A[11]), .Q(n343) );
  CLKIN0 U329 ( .A(n95), .Q(n94) );
  NAND22 U330 ( .A(n91), .B(n92), .Q(n89) );
  NOR22 U331 ( .A(n49), .B(n50), .Q(n51) );
  INV3 U332 ( .A(A[12]), .Q(n50) );
  NAND20 U333 ( .A(n62), .B(n63), .Q(n56) );
  NOR21 U334 ( .A(n12), .B(n336), .Q(n350) );
  NOR21 U335 ( .A(n12), .B(n61), .Q(n351) );
  XOR21 U336 ( .A(n56), .B(n57), .Q(SUM[9]) );
  XOR20 U337 ( .A(B[3]), .B(A[3]), .Q(n90) );
  NOR24 U338 ( .A(n150), .B(n134), .Q(n52) );
  INV4 U339 ( .A(n13), .Q(n139) );
  CLKIN0 U340 ( .A(B[8]), .Q(n69) );
  NAND22 U341 ( .A(n365), .B(n127), .Q(n93) );
  INV6 U342 ( .A(n240), .Q(n197) );
  NAND22 U343 ( .A(n53), .B(n54), .Q(n55) );
  INV3 U344 ( .A(A[7]), .Q(n53) );
  INV2 U345 ( .A(B[7]), .Q(n54) );
  NOR22 U346 ( .A(A[10]), .B(B[10]), .Q(n337) );
  NAND20 U347 ( .A(n345), .B(n346), .Q(n347) );
  NOR24 U348 ( .A(n337), .B(n64), .Q(n334) );
  NAND42 U349 ( .A(n299), .B(n298), .C(n304), .D(n86), .Q(n181) );
  NOR21 U350 ( .A(B[19]), .B(A[19]), .Q(n251) );
  XNR20 U351 ( .A(n2), .B(A[15]), .Q(n311) );
  XNR20 U352 ( .A(B[7]), .B(A[7]), .Q(n70) );
  NOR21 U353 ( .A(B[7]), .B(A[7]), .Q(n369) );
  NOR20 U354 ( .A(A[4]), .B(B[4]), .Q(n82) );
  OAI222 U355 ( .A(B[14]), .B(A[14]), .C(B[13]), .D(A[13]), .Q(n307) );
  XNR20 U356 ( .A(B[4]), .B(A[4]), .Q(n85) );
  CLKIN0 U357 ( .A(B[20]), .Q(n253) );
  XNR20 U358 ( .A(B[20]), .B(A[20]), .Q(n237) );
  NOR21 U359 ( .A(B[0]), .B(n357), .Q(n378) );
  XNR20 U360 ( .A(B[8]), .B(A[8]), .Q(n66) );
  XNR20 U361 ( .A(n23), .B(A[12]), .Q(n329) );
  NAND28 U362 ( .A(n181), .B(n278), .Q(n99) );
  CLKIN3 U363 ( .A(n336), .Q(n60) );
  OAI212 U364 ( .A(n77), .B(n78), .C(n372), .Q(n72) );
  OAI212 U365 ( .A(n81), .B(n82), .C(n83), .Q(n79) );
  CLKIN3 U366 ( .A(n83), .Q(n88) );
  OAI222 U367 ( .A(n108), .B(n109), .C(n110), .D(n111), .Q(n107) );
  CLKIN3 U368 ( .A(n91), .Q(n126) );
  AOI212 U369 ( .A(n133), .B(n52), .C(n120), .Q(n132) );
  OAI222 U370 ( .A(n134), .B(n135), .C(n136), .D(n137), .Q(n120) );
  AOI212 U371 ( .A(n133), .B(n139), .C(n47), .Q(n140) );
  XOR22 U372 ( .A(n155), .B(n156), .Q(SUM[27]) );
  AOI212 U373 ( .A(n157), .B(n151), .C(n158), .Q(n156) );
  CLKIN3 U374 ( .A(n147), .Q(n158) );
  NAND24 U375 ( .A(B[26]), .B(A[26]), .Q(n147) );
  AOI312 U376 ( .A(n168), .B(n152), .C(n169), .D(n170), .Q(n160) );
  OAI212 U377 ( .A(n10), .B(n171), .C(n146), .Q(n170) );
  AOI212 U378 ( .A(n133), .B(n168), .C(n174), .Q(n173) );
  AOI312 U379 ( .A(n179), .B(n181), .C(n180), .D(n124), .Q(n178) );
  NAND33 U380 ( .A(n202), .B(n203), .C(n204), .Q(n201) );
  OAI212 U381 ( .A(n205), .B(n206), .C(n202), .Q(n200) );
  CLKIN3 U382 ( .A(n171), .Q(n174) );
  OAI212 U383 ( .A(n206), .B(n214), .C(n198), .Q(n213) );
  CLKIN3 U384 ( .A(n198), .Q(n217) );
  AOI212 U385 ( .A(n224), .B(n208), .C(n225), .Q(n220) );
  CLKIN3 U386 ( .A(n223), .Q(n234) );
  AOI312 U387 ( .A(n241), .B(n243), .C(n242), .D(n244), .Q(n240) );
  CLKIN3 U388 ( .A(n204), .Q(n254) );
  CLKIN3 U389 ( .A(n365), .Q(n256) );
  OAI212 U390 ( .A(n249), .B(n22), .C(n241), .Q(n258) );
  CLKIN6 U391 ( .A(B[18]), .Q(n262) );
  CLKIN3 U392 ( .A(n241), .Q(n261) );
  XOR22 U393 ( .A(n271), .B(n272), .Q(SUM[17]) );
  CLKIN3 U394 ( .A(n243), .Q(n268) );
  NOR24 U395 ( .A(n279), .B(n280), .Q(n278) );
  OAI2112 U396 ( .A(n284), .B(n285), .C(n286), .D(n287), .Q(n281) );
  NOR24 U397 ( .A(n289), .B(n290), .Q(n288) );
  CLKIN6 U398 ( .A(n292), .Q(n291) );
  NOR24 U399 ( .A(n307), .B(n306), .Q(n299) );
  OAI222 U400 ( .A(B[15]), .B(A[15]), .C(B[12]), .D(A[12]), .Q(n306) );
  CLKIN3 U401 ( .A(n270), .Q(n310) );
  AOI212 U402 ( .A(n315), .B(n314), .C(n319), .Q(n318) );
  CLKIN3 U403 ( .A(n46), .Q(n319) );
  NAND24 U404 ( .A(n334), .B(n335), .Q(n333) );
  AOI212 U405 ( .A(n18), .B(A[11]), .C(n338), .Q(n332) );
  NOR24 U406 ( .A(n339), .B(n340), .Q(n298) );
  OAI222 U407 ( .A(B[8]), .B(A[8]), .C(B[11]), .D(A[11]), .Q(n339) );
  CLKIN3 U408 ( .A(n324), .Q(n342) );
  NAND24 U409 ( .A(n352), .B(n353), .Q(n59) );
  AOI212 U410 ( .A(n360), .B(n361), .C(n130), .Q(n358) );
  OAI212 U411 ( .A(A[0]), .B(n376), .C(n377), .Q(SUM[0]) );
endmodule


module E_alu_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255;

  CLKIN6 U1 ( .A(B[23]), .Q(n255) );
  NAND33 U2 ( .A(n221), .B(n222), .C(n223), .Q(n143) );
  NOR24 U3 ( .A(n143), .B(n144), .Q(n7) );
  CLKIN3 U4 ( .A(n149), .Q(n3) );
  NAND26 U5 ( .A(A[17]), .B(n252), .Q(n54) );
  INV3 U6 ( .A(n38), .Q(n56) );
  NOR20 U7 ( .A(n69), .B(n130), .Q(n126) );
  INV6 U8 ( .A(n33), .Q(n2) );
  NOR24 U9 ( .A(B[3]), .B(n206), .Q(n205) );
  NOR24 U10 ( .A(B[25]), .B(n133), .Q(n132) );
  NOR23 U11 ( .A(B[24]), .B(n134), .Q(n248) );
  NOR24 U12 ( .A(n246), .B(n247), .Q(n135) );
  NAND32 U13 ( .A(n54), .B(n80), .C(n66), .Q(n157) );
  NAND22 U14 ( .A(n66), .B(n54), .Q(n251) );
  NOR22 U15 ( .A(n40), .B(n41), .Q(n227) );
  NOR24 U16 ( .A(n41), .B(n42), .Q(n45) );
  NOR23 U17 ( .A(n156), .B(n157), .Q(n148) );
  NAND31 U18 ( .A(n81), .B(n158), .C(n83), .Q(n156) );
  AOI2111 U19 ( .A(n105), .B(n33), .C(n106), .D(n107), .Q(n8) );
  INV2 U20 ( .A(B[22]), .Q(n253) );
  NAND23 U21 ( .A(A[16]), .B(n57), .Q(n80) );
  NOR22 U22 ( .A(n205), .B(n217), .Q(n216) );
  NOR21 U23 ( .A(A[2]), .B(n219), .Q(n218) );
  CLKIN6 U24 ( .A(B[9]), .Q(n100) );
  INV6 U25 ( .A(n66), .Q(n42) );
  INV6 U26 ( .A(n80), .Q(n40) );
  INV3 U27 ( .A(n148), .Q(n1) );
  NAND31 U28 ( .A(n150), .B(n151), .C(n20), .Q(n24) );
  NOR21 U29 ( .A(n240), .B(n241), .Q(n239) );
  NOR22 U30 ( .A(n242), .B(n243), .Q(n238) );
  NOR21 U31 ( .A(n200), .B(n201), .Q(n182) );
  INV12 U32 ( .A(n110), .Q(n33) );
  AOI221 U33 ( .A(n125), .B(n60), .C(n126), .D(n127), .Q(n114) );
  INV1 U34 ( .A(B[15]), .Q(n231) );
  NAND34 U35 ( .A(n31), .B(n30), .C(n6), .Q(n27) );
  NOR23 U36 ( .A(n248), .B(n132), .Q(n131) );
  NAND22 U37 ( .A(n159), .B(n33), .Q(n146) );
  NOR24 U38 ( .A(n27), .B(n26), .Q(n9) );
  NAND31 U39 ( .A(n75), .B(n33), .C(n76), .Q(n74) );
  INV6 U40 ( .A(n67), .Q(n243) );
  NAND21 U41 ( .A(n66), .B(n67), .Q(n120) );
  NAND24 U42 ( .A(A[21]), .B(n244), .Q(n67) );
  NOR22 U43 ( .A(n160), .B(n161), .Q(n159) );
  NOR23 U44 ( .A(n4), .B(n24), .Q(n147) );
  NAND22 U45 ( .A(n224), .B(n33), .Q(n223) );
  OAI311 U46 ( .A(n181), .B(n182), .C(n183), .D(n184), .Q(n145) );
  INV0 U47 ( .A(B[12]), .Q(n167) );
  NAND30 U48 ( .A(n78), .B(n38), .C(B[7]), .Q(n155) );
  CLKIN1 U49 ( .A(B[10]), .Q(n192) );
  NAND20 U50 ( .A(B[11]), .B(n38), .Q(n44) );
  INV4 U51 ( .A(B[11]), .Q(n187) );
  OAI220 U52 ( .A(n108), .B(n109), .C(n110), .D(n111), .Q(n107) );
  NAND28 U53 ( .A(A[22]), .B(n253), .Q(n66) );
  OAI2111 U54 ( .A(n173), .B(n174), .C(n38), .D(n66), .Q(n160) );
  INV1 U55 ( .A(n172), .Q(n142) );
  NAND22 U56 ( .A(n131), .B(B[20]), .Q(n70) );
  INV2 U57 ( .A(B[2]), .Q(n219) );
  INV6 U58 ( .A(B[17]), .Q(n252) );
  INV3 U59 ( .A(n54), .Q(n41) );
  NAND31 U60 ( .A(n78), .B(n38), .C(B[8]), .Q(n77) );
  NOR22 U61 ( .A(n155), .B(n37), .Q(n149) );
  INV2 U62 ( .A(B[8]), .Q(n165) );
  NOR22 U63 ( .A(B[27]), .B(n136), .Q(n247) );
  INV1 U64 ( .A(B[20]), .Q(n245) );
  NOR20 U65 ( .A(B[5]), .B(n178), .Q(n176) );
  NAND42 U66 ( .A(n71), .B(n73), .C(n72), .D(n74), .Q(n26) );
  INV6 U67 ( .A(n135), .Q(n69) );
  INV4 U68 ( .A(n162), .Q(n78) );
  INV8 U69 ( .A(n166), .Q(n37) );
  INV1 U70 ( .A(B[5]), .Q(n177) );
  NAND21 U71 ( .A(B[31]), .B(n152), .Q(n20) );
  INV1 U72 ( .A(B[14]), .Q(n230) );
  NOR33 U73 ( .A(n1), .B(n2), .C(n3), .Q(n4) );
  NOR22 U74 ( .A(B[26]), .B(n137), .Q(n246) );
  NAND41 U75 ( .A(n93), .B(n94), .C(n95), .D(n33), .Q(n72) );
  AOI311 U76 ( .A(n47), .B(n48), .C(n33), .D(n49), .Q(n30) );
  NOR21 U77 ( .A(n69), .B(n70), .Q(n62) );
  NOR20 U78 ( .A(B[7]), .B(n158), .Q(n189) );
  NOR22 U79 ( .A(A[30]), .B(n19), .Q(n154) );
  INV1 U80 ( .A(B[30]), .Q(n19) );
  INV4 U81 ( .A(n5), .Q(n6) );
  AOI221 U82 ( .A(n32), .B(n33), .C(n34), .D(n33), .Q(n31) );
  NAND43 U83 ( .A(n237), .B(n135), .C(n238), .D(n239), .Q(n110) );
  NAND22 U84 ( .A(n28), .B(n29), .Q(n5) );
  NOR31 U85 ( .A(n251), .B(n40), .C(n91), .Q(n84) );
  NAND22 U86 ( .A(n81), .B(n99), .Q(n98) );
  NOR21 U87 ( .A(n50), .B(n51), .Q(n49) );
  INV3 U88 ( .A(n218), .Q(n217) );
  NOR21 U89 ( .A(n42), .B(n53), .Q(n48) );
  CLKIN6 U90 ( .A(n69), .Q(n60) );
  NOR20 U91 ( .A(n56), .B(n69), .Q(n117) );
  NAND20 U92 ( .A(n232), .B(n33), .Q(n222) );
  NOR20 U93 ( .A(n123), .B(n124), .Q(n116) );
  NOR20 U94 ( .A(n69), .B(n87), .Q(n86) );
  NOR21 U95 ( .A(n185), .B(n186), .Q(n184) );
  NAND20 U96 ( .A(n66), .B(n235), .Q(n234) );
  NAND20 U97 ( .A(n236), .B(n33), .Q(n221) );
  NAND20 U98 ( .A(n121), .B(n122), .Q(n119) );
  NOR21 U99 ( .A(n79), .B(n157), .Q(n75) );
  NAND20 U100 ( .A(n54), .B(n55), .Q(n53) );
  NAND20 U101 ( .A(A[30]), .B(n19), .Q(n18) );
  INV2 U102 ( .A(n88), .Q(n87) );
  NAND22 U103 ( .A(n131), .B(n60), .Q(n50) );
  NOR22 U104 ( .A(n248), .B(n132), .Q(n237) );
  INV3 U105 ( .A(B[16]), .Q(n57) );
  NOR20 U106 ( .A(n56), .B(n57), .Q(n47) );
  NAND22 U107 ( .A(n131), .B(B[21]), .Q(n130) );
  INV3 U108 ( .A(B[19]), .Q(n124) );
  NOR21 U109 ( .A(n101), .B(n102), .Q(n71) );
  NAND22 U110 ( .A(n58), .B(n59), .Q(n29) );
  NAND22 U111 ( .A(n62), .B(n63), .Q(n28) );
  NAND20 U112 ( .A(B[22]), .B(n131), .Q(n109) );
  NAND22 U113 ( .A(n113), .B(n60), .Q(n108) );
  NAND30 U114 ( .A(n80), .B(n81), .C(n54), .Q(n186) );
  NAND31 U115 ( .A(n11), .B(n12), .C(n13), .Q(n10) );
  NOR31 U116 ( .A(n35), .B(n36), .C(n37), .Q(n34) );
  NOR31 U117 ( .A(n43), .B(n44), .C(n37), .Q(n32) );
  NAND22 U118 ( .A(n45), .B(n39), .Q(n35) );
  NOR31 U119 ( .A(n96), .B(n97), .C(n98), .Q(n95) );
  NAND20 U120 ( .A(n54), .B(n80), .Q(n96) );
  NOR21 U121 ( .A(n225), .B(n226), .Q(n224) );
  NAND22 U122 ( .A(n227), .B(n228), .Q(n225) );
  NAND22 U123 ( .A(n202), .B(n203), .Q(n201) );
  INV3 U124 ( .A(n204), .Q(n203) );
  NOR21 U125 ( .A(A[0]), .B(n205), .Q(n202) );
  NOR21 U126 ( .A(B[18]), .B(n235), .Q(n240) );
  NAND22 U127 ( .A(n208), .B(n209), .Q(n200) );
  INV3 U128 ( .A(n210), .Q(n209) );
  INV0 U129 ( .A(B[0]), .Q(n210) );
  NOR21 U130 ( .A(n189), .B(n190), .Q(n188) );
  NAND22 U131 ( .A(n171), .B(n172), .Q(n168) );
  NOR21 U132 ( .A(n142), .B(n229), .Q(n228) );
  NAND22 U133 ( .A(n171), .B(n170), .Q(n229) );
  NAND22 U134 ( .A(n93), .B(n78), .Q(n161) );
  NOR21 U135 ( .A(n14), .B(n15), .Q(n13) );
  NOR21 U136 ( .A(n17), .B(n18), .Q(n14) );
  NOR21 U137 ( .A(n16), .B(n17), .Q(n15) );
  NAND22 U138 ( .A(n114), .B(n115), .Q(n106) );
  NAND31 U139 ( .A(n116), .B(n117), .C(n118), .Q(n115) );
  NOR21 U140 ( .A(n119), .B(n120), .Q(n118) );
  NOR31 U141 ( .A(n249), .B(n250), .C(n251), .Q(n236) );
  NAND20 U142 ( .A(n80), .B(n254), .Q(n250) );
  INV3 U143 ( .A(n131), .Q(n123) );
  NOR21 U144 ( .A(n233), .B(n234), .Q(n232) );
  NAND20 U145 ( .A(B[18]), .B(n38), .Q(n233) );
  NAND41 U146 ( .A(n213), .B(n180), .C(n214), .D(n215), .Q(n181) );
  INV3 U147 ( .A(n220), .Q(n213) );
  INV3 U148 ( .A(n216), .Q(n215) );
  NAND22 U149 ( .A(A[11]), .B(n187), .Q(n81) );
  INV3 U150 ( .A(A[8]), .Q(n82) );
  NOR21 U151 ( .A(A[24]), .B(n61), .Q(n58) );
  INV0 U152 ( .A(B[24]), .Q(n61) );
  NOR21 U153 ( .A(A[5]), .B(n177), .Q(n220) );
  NOR21 U154 ( .A(A[12]), .B(n40), .Q(n39) );
  INV3 U155 ( .A(A[5]), .Q(n178) );
  NOR21 U156 ( .A(A[27]), .B(n104), .Q(n101) );
  NAND22 U157 ( .A(n163), .B(n164), .Q(n162) );
  NAND22 U158 ( .A(A[9]), .B(n100), .Q(n163) );
  NAND22 U159 ( .A(A[8]), .B(n165), .Q(n164) );
  NAND22 U160 ( .A(A[20]), .B(n245), .Q(n121) );
  INV3 U161 ( .A(B[21]), .Q(n244) );
  NOR21 U162 ( .A(A[28]), .B(n103), .Q(n102) );
  INV0 U163 ( .A(B[28]), .Q(n103) );
  NOR20 U164 ( .A(A[22]), .B(n56), .Q(n113) );
  NAND22 U165 ( .A(A[15]), .B(n231), .Q(n172) );
  NAND20 U166 ( .A(B[29]), .B(n153), .Q(n151) );
  INV3 U167 ( .A(n154), .Q(n150) );
  INV3 U168 ( .A(A[29]), .Q(n153) );
  NAND22 U169 ( .A(A[14]), .B(n230), .Q(n171) );
  NOR21 U170 ( .A(A[25]), .B(n138), .Q(n125) );
  INV0 U171 ( .A(B[25]), .Q(n138) );
  INV3 U172 ( .A(A[31]), .Q(n152) );
  NAND22 U173 ( .A(n45), .B(n46), .Q(n43) );
  INV3 U174 ( .A(A[16]), .Q(n55) );
  NAND22 U175 ( .A(n81), .B(n92), .Q(n91) );
  INV3 U176 ( .A(A[10]), .Q(n92) );
  NOR21 U177 ( .A(n64), .B(n65), .Q(n63) );
  NAND20 U178 ( .A(n67), .B(n68), .Q(n64) );
  NAND20 U179 ( .A(n38), .B(n66), .Q(n65) );
  INV3 U180 ( .A(A[20]), .Q(n68) );
  NAND22 U181 ( .A(n21), .B(n22), .Q(n12) );
  NOR20 U182 ( .A(B[29]), .B(n153), .Q(n21) );
  NAND22 U183 ( .A(n23), .B(n22), .Q(n11) );
  NOR20 U184 ( .A(B[28]), .B(n25), .Q(n23) );
  INV3 U185 ( .A(A[28]), .Q(n25) );
  NOR21 U186 ( .A(n139), .B(n140), .Q(n105) );
  NAND30 U187 ( .A(B[14]), .B(n66), .C(n38), .Q(n140) );
  NAND22 U188 ( .A(n227), .B(n141), .Q(n139) );
  NOR21 U189 ( .A(A[14]), .B(n142), .Q(n141) );
  NOR21 U190 ( .A(n56), .B(n128), .Q(n127) );
  NAND20 U191 ( .A(n66), .B(n129), .Q(n128) );
  INV3 U192 ( .A(A[21]), .Q(n129) );
  NOR21 U193 ( .A(A[26]), .B(n89), .Q(n88) );
  INV0 U194 ( .A(B[26]), .Q(n89) );
  NAND20 U195 ( .A(B[23]), .B(n52), .Q(n51) );
  INV3 U196 ( .A(A[23]), .Q(n52) );
  INV3 U197 ( .A(n196), .Q(n195) );
  NOR21 U198 ( .A(A[3]), .B(n197), .Q(n196) );
  INV3 U199 ( .A(A[24]), .Q(n134) );
  INV3 U200 ( .A(A[3]), .Q(n206) );
  INV3 U201 ( .A(A[26]), .Q(n137) );
  INV3 U202 ( .A(A[0]), .Q(n207) );
  INV3 U203 ( .A(A[27]), .Q(n136) );
  INV3 U204 ( .A(A[18]), .Q(n235) );
  INV3 U205 ( .A(A[13]), .Q(n170) );
  INV3 U206 ( .A(A[9]), .Q(n99) );
  INV3 U207 ( .A(A[19]), .Q(n122) );
  INV3 U208 ( .A(A[4]), .Q(n179) );
  INV3 U209 ( .A(A[7]), .Q(n158) );
  INV3 U210 ( .A(A[15]), .Q(n254) );
  INV3 U211 ( .A(A[1]), .Q(n199) );
  INV3 U212 ( .A(A[2]), .Q(n198) );
  INV3 U213 ( .A(A[25]), .Q(n133) );
  INV3 U214 ( .A(A[6]), .Q(n191) );
  INV3 U215 ( .A(A[17]), .Q(n112) );
  NOR21 U216 ( .A(n77), .B(n37), .Q(n76) );
  INV0 U217 ( .A(B[27]), .Q(n104) );
  NAND20 U218 ( .A(B[12]), .B(n38), .Q(n36) );
  NAND20 U219 ( .A(B[4]), .B(n179), .Q(n214) );
  NOR31 U220 ( .A(n100), .B(n42), .C(n56), .Q(n94) );
  NAND40 U221 ( .A(n66), .B(n112), .C(B[17]), .D(n38), .Q(n111) );
  NAND30 U222 ( .A(B[13]), .B(n66), .C(n38), .Q(n226) );
  NOR20 U223 ( .A(B[13]), .B(n170), .Q(n169) );
  NAND20 U224 ( .A(B[10]), .B(n38), .Q(n90) );
  NOR21 U225 ( .A(n90), .B(n37), .Q(n85) );
  NAND31 U226 ( .A(n81), .B(n82), .C(n83), .Q(n79) );
  NAND22 U227 ( .A(n83), .B(n188), .Q(n185) );
  AOI311 U228 ( .A(n84), .B(n85), .C(n33), .D(n86), .Q(n73) );
  NAND22 U229 ( .A(A[10]), .B(n192), .Q(n83) );
  NOR20 U230 ( .A(B[2]), .B(n198), .Q(n204) );
  INV0 U231 ( .A(B[3]), .Q(n197) );
  NOR20 U232 ( .A(B[1]), .B(n199), .Q(n212) );
  CLKIN0 U233 ( .A(B[1]), .Q(n194) );
  NOR21 U234 ( .A(n211), .B(n212), .Q(n208) );
  OAI311 U235 ( .A(n193), .B(n205), .C(n194), .D(n195), .Q(n183) );
  NAND20 U236 ( .A(B[6]), .B(n191), .Q(n180) );
  NOR20 U237 ( .A(B[6]), .B(n191), .Q(n190) );
  XNR21 U238 ( .A(B[31]), .B(A[31]), .Q(n16) );
  NOR21 U239 ( .A(B[19]), .B(n122), .Q(n241) );
  OAI210 U240 ( .A(B[2]), .B(n198), .C(n199), .Q(n193) );
  NAND20 U241 ( .A(B[15]), .B(n38), .Q(n249) );
  NOR20 U242 ( .A(B[4]), .B(n179), .Q(n175) );
  NOR21 U243 ( .A(A[11]), .B(n40), .Q(n46) );
  NOR21 U244 ( .A(B[0]), .B(n207), .Q(n211) );
  NAND28 U245 ( .A(A[23]), .B(n255), .Q(n38) );
  AOI312 U246 ( .A(n7), .B(n8), .C(n9), .D(n10), .Q(LT_LE) );
  CLKIN3 U247 ( .A(n20), .Q(n17) );
  CLKIN3 U248 ( .A(n24), .Q(n22) );
  CLKIN3 U249 ( .A(n50), .Q(n59) );
  CLKIN3 U250 ( .A(n83), .Q(n97) );
  OAI212 U251 ( .A(n145), .B(n146), .C(n147), .Q(n144) );
  CLKIN3 U252 ( .A(n37), .Q(n93) );
  AOI2112 U253 ( .A(A[12]), .B(n167), .C(n168), .D(n169), .Q(n166) );
  OAI222 U254 ( .A(n175), .B(n176), .C(A[5]), .D(n177), .Q(n174) );
  CLKIN3 U255 ( .A(n180), .Q(n173) );
  CLKIN3 U256 ( .A(n121), .Q(n242) );
endmodule


module E_alu_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283;

  NAND22 U3 ( .A(n272), .B(n273), .Q(n42) );
  NAND24 U4 ( .A(n264), .B(n265), .Q(n120) );
  AOI222 U5 ( .A(n100), .B(n41), .C(n96), .D(n42), .Q(n271) );
  CLKIN3 U6 ( .A(SH[1]), .Q(n15) );
  NAND22 U7 ( .A(n196), .B(n197), .Q(n29) );
  NAND23 U8 ( .A(n137), .B(n138), .Q(n63) );
  NAND23 U9 ( .A(n227), .B(n228), .Q(n56) );
  AOI211 U10 ( .A(n18), .B(n117), .C(n200), .Q(n182) );
  CLKIN3 U11 ( .A(SH[0]), .Q(n14) );
  NOR20 U12 ( .A(SH[1]), .B(SH[0]), .Q(n6) );
  NAND34 U13 ( .A(n161), .B(n162), .C(n160), .Q(n159) );
  AOI220 U14 ( .A(A[21]), .B(n7), .C(A[22]), .D(n191), .Q(n197) );
  BUF2 U15 ( .A(n5), .Q(n7) );
  INV6 U16 ( .A(n283), .Q(n192) );
  INV6 U17 ( .A(n209), .Q(n193) );
  BUF2 U18 ( .A(n5), .Q(n8) );
  NAND41 U19 ( .A(n92), .B(n93), .C(n94), .D(n95), .Q(n91) );
  INV3 U20 ( .A(n117), .Q(n115) );
  BUF2 U21 ( .A(n190), .Q(n11) );
  NAND23 U22 ( .A(n223), .B(n224), .Q(n104) );
  INV3 U23 ( .A(n237), .Q(n139) );
  NAND23 U24 ( .A(n194), .B(n195), .Q(n116) );
  NAND24 U25 ( .A(n101), .B(n56), .Q(n94) );
  INV3 U26 ( .A(n254), .Q(n30) );
  INV3 U27 ( .A(n245), .Q(n28) );
  INV3 U28 ( .A(n248), .Q(n26) );
  NAND23 U29 ( .A(n243), .B(n244), .Q(n108) );
  NOR24 U30 ( .A(n18), .B(n153), .Q(B[18]) );
  AOI221 U31 ( .A(A[24]), .B(n192), .C(A[25]), .D(n193), .Q(n243) );
  NOR24 U32 ( .A(n18), .B(n150), .Q(B[19]) );
  AOI220 U33 ( .A(A[12]), .B(n8), .C(A[13]), .D(n191), .Q(n273) );
  INV3 U34 ( .A(SH[4]), .Q(n19) );
  AOI222 U35 ( .A(n100), .B(n116), .C(n96), .D(n159), .Q(n158) );
  AOI221 U36 ( .A(A[18]), .B(n8), .C(A[19]), .D(n191), .Q(n247) );
  INV8 U37 ( .A(n282), .Q(n191) );
  NAND24 U38 ( .A(n144), .B(n145), .Q(n143) );
  AOI221 U39 ( .A(A[20]), .B(n9), .C(A[21]), .D(n191), .Q(n267) );
  AOI221 U40 ( .A(n101), .B(n43), .C(n102), .D(n44), .Q(n260) );
  NAND21 U41 ( .A(n26), .B(n108), .Q(n180) );
  AOI220 U42 ( .A(n26), .B(n70), .C(n28), .D(n108), .Q(n242) );
  AOI221 U43 ( .A(n13), .B(n70), .C(n102), .D(n108), .Q(n154) );
  AOI222 U44 ( .A(n101), .B(n106), .C(n102), .D(n104), .Q(n134) );
  AOI221 U45 ( .A(A[25]), .B(n192), .C(A[26]), .D(n193), .Q(n225) );
  NAND21 U46 ( .A(n35), .B(n60), .Q(n57) );
  NAND21 U47 ( .A(n35), .B(n36), .Q(n32) );
  NAND21 U48 ( .A(n35), .B(n41), .Q(n89) );
  INV6 U49 ( .A(n251), .Q(n35) );
  AOI221 U50 ( .A(A[17]), .B(n11), .C(A[18]), .D(n191), .Q(n205) );
  NOR24 U51 ( .A(n18), .B(n133), .Q(B[23]) );
  AOI221 U52 ( .A(A[30]), .B(n192), .C(A[31]), .D(n193), .Q(n262) );
  INV3 U53 ( .A(n40), .Q(n129) );
  INV6 U54 ( .A(n112), .Q(n153) );
  AOI221 U55 ( .A(A[24]), .B(n7), .C(A[25]), .D(n191), .Q(n265) );
  NOR21 U56 ( .A(SH[1]), .B(SH[0]), .Q(n5) );
  NAND20 U57 ( .A(n26), .B(n29), .Q(n185) );
  NAND23 U58 ( .A(n141), .B(n142), .Q(n140) );
  AOI220 U59 ( .A(n28), .B(n29), .C(n30), .D(n31), .Q(n24) );
  AOI222 U60 ( .A(n12), .B(n29), .C(n102), .D(n116), .Q(n141) );
  NOR21 U61 ( .A(n18), .B(n156), .Q(B[17]) );
  AOI221 U62 ( .A(A[25]), .B(n8), .C(A[26]), .D(n191), .Q(n195) );
  NAND21 U63 ( .A(n42), .B(n26), .Q(n88) );
  NAND24 U64 ( .A(n134), .B(n135), .Q(n49) );
  NOR22 U65 ( .A(n18), .B(n129), .Q(B[24]) );
  NAND22 U66 ( .A(A[29]), .B(n7), .Q(n162) );
  AOI221 U67 ( .A(n101), .B(n44), .C(n102), .D(n120), .Q(n144) );
  NAND21 U68 ( .A(n100), .B(n159), .Q(n142) );
  NAND24 U69 ( .A(n93), .B(n94), .Q(n151) );
  NAND22 U70 ( .A(n102), .B(n106), .Q(n93) );
  AOI222 U71 ( .A(n100), .B(n110), .C(n96), .D(n139), .Q(n155) );
  AOI222 U72 ( .A(A[28]), .B(n9), .C(A[29]), .D(n191), .Q(n263) );
  INV3 U73 ( .A(n125), .Q(n20) );
  OAI211 U74 ( .A(n126), .B(n127), .C(n128), .Q(n125) );
  NAND24 U75 ( .A(n225), .B(n226), .Q(n106) );
  NAND22 U76 ( .A(A[31]), .B(n192), .Q(n160) );
  INV2 U77 ( .A(n63), .Q(n136) );
  NAND21 U78 ( .A(SH[1]), .B(SH[0]), .Q(n209) );
  OAI220 U79 ( .A(n12), .B(n222), .C(n104), .D(n222), .Q(n221) );
  NOR20 U80 ( .A(n173), .B(n127), .Q(n222) );
  NAND22 U81 ( .A(A[31]), .B(n8), .Q(n173) );
  NAND20 U82 ( .A(n28), .B(n104), .Q(n169) );
  NOR24 U83 ( .A(n126), .B(n208), .Q(n117) );
  AOI2112 U84 ( .A(n96), .B(n97), .C(n151), .D(n152), .Q(n150) );
  AOI220 U85 ( .A(A[21]), .B(n192), .C(A[22]), .D(n193), .Q(n227) );
  BUF6 U86 ( .A(n6), .Q(n9) );
  NAND21 U87 ( .A(n12), .B(n116), .Q(n128) );
  NAND21 U88 ( .A(n26), .B(n106), .Q(n170) );
  AOI221 U89 ( .A(A[23]), .B(n10), .C(A[24]), .D(n191), .Q(n226) );
  AOI221 U90 ( .A(n100), .B(n120), .C(n96), .D(n132), .Q(n261) );
  AOI221 U91 ( .A(A[29]), .B(n192), .C(A[30]), .D(n193), .Q(n223) );
  NAND21 U92 ( .A(A[30]), .B(n191), .Q(n161) );
  AOI221 U93 ( .A(A[22]), .B(n9), .C(A[23]), .D(n191), .Q(n244) );
  NAND26 U94 ( .A(n238), .B(n239), .Q(n110) );
  AOI221 U95 ( .A(A[28]), .B(n192), .C(A[29]), .D(n193), .Q(n238) );
  NAND21 U96 ( .A(n18), .B(n49), .Q(n48) );
  NAND24 U97 ( .A(n262), .B(n263), .Q(n132) );
  NAND21 U98 ( .A(SH[1]), .B(n14), .Q(n283) );
  NOR23 U99 ( .A(n18), .B(n83), .Q(B[20]) );
  AOI221 U100 ( .A(A[22]), .B(n192), .C(A[23]), .D(n193), .Q(n266) );
  NAND21 U101 ( .A(n30), .B(n59), .Q(n58) );
  AOI221 U102 ( .A(n12), .B(n27), .C(n102), .D(n29), .Q(n157) );
  AOI220 U103 ( .A(n96), .B(n69), .C(n100), .D(n74), .Q(n114) );
  NAND20 U104 ( .A(n30), .B(n73), .Q(n72) );
  CLKIN2 U105 ( .A(n32), .Q(n22) );
  AOI220 U106 ( .A(n102), .B(n73), .C(n101), .D(n64), .Q(n113) );
  NAND21 U107 ( .A(n26), .B(n69), .Q(n68) );
  NAND21 U108 ( .A(n102), .B(n19), .Q(n251) );
  NAND22 U109 ( .A(n30), .B(n36), .Q(n187) );
  NOR21 U110 ( .A(n18), .B(n20), .Q(B[25]) );
  CLKIN2 U111 ( .A(n181), .Q(n177) );
  AOI220 U112 ( .A(n30), .B(n60), .C(n35), .D(n55), .Q(n214) );
  NAND21 U113 ( .A(n96), .B(n19), .Q(n245) );
  NAND21 U114 ( .A(n100), .B(n19), .Q(n248) );
  AOI2111 U115 ( .A(n30), .B(n45), .C(n85), .D(n86), .Q(n84) );
  MUX22 U116 ( .A(n111), .B(n112), .S(n18), .Q(B[2]) );
  INV2 U117 ( .A(n101), .Q(n208) );
  CLKIN3 U118 ( .A(n172), .Q(n105) );
  INV6 U119 ( .A(n159), .Q(n126) );
  NAND20 U120 ( .A(n18), .B(n40), .Q(n39) );
  NAND20 U121 ( .A(n18), .B(n124), .Q(n234) );
  NAND20 U122 ( .A(SH[3]), .B(SH[2]), .Q(n274) );
  AOI220 U123 ( .A(n30), .B(n42), .C(n35), .D(n43), .Q(n210) );
  AOI220 U124 ( .A(n26), .B(n43), .C(n28), .D(n44), .Q(n37) );
  CLKIN3 U125 ( .A(n221), .Q(n122) );
  NAND20 U126 ( .A(n12), .B(n110), .Q(n235) );
  NOR20 U127 ( .A(SH[1]), .B(SH[0]), .Q(n190) );
  CLKIN3 U128 ( .A(n171), .Q(n167) );
  NAND21 U129 ( .A(n30), .B(n55), .Q(n171) );
  NAND24 U130 ( .A(n157), .B(n158), .Q(n147) );
  NAND24 U131 ( .A(n154), .B(n155), .Q(n112) );
  AOI222 U132 ( .A(n13), .B(n108), .C(n102), .D(n110), .Q(n137) );
  NAND20 U133 ( .A(n30), .B(n69), .Q(n181) );
  AOI220 U134 ( .A(n12), .B(n50), .C(n102), .D(n59), .Q(n98) );
  CLKIN3 U135 ( .A(n213), .Q(n119) );
  NAND20 U136 ( .A(n13), .B(n132), .Q(n213) );
  AOI220 U137 ( .A(n35), .B(n70), .C(n18), .D(n109), .Q(n175) );
  NAND20 U138 ( .A(n28), .B(n43), .Q(n87) );
  NAND20 U139 ( .A(n12), .B(n139), .Q(n176) );
  NAND20 U140 ( .A(n30), .B(n33), .Q(n82) );
  NAND20 U141 ( .A(n26), .B(n36), .Q(n79) );
  NAND20 U142 ( .A(n28), .B(n27), .Q(n80) );
  NAND20 U143 ( .A(n28), .B(n70), .Q(n67) );
  NAND20 U144 ( .A(n28), .B(n116), .Q(n186) );
  INV2 U145 ( .A(n184), .Q(n183) );
  NAND20 U146 ( .A(n35), .B(n27), .Q(n201) );
  MUX21 U147 ( .A(n259), .B(n164), .S(n18), .Q(B[0]) );
  NAND20 U148 ( .A(SH[3]), .B(n16), .Q(n277) );
  AOI220 U149 ( .A(A[19]), .B(n9), .C(A[20]), .D(n191), .Q(n228) );
  NAND21 U150 ( .A(SH[2]), .B(n17), .Q(n127) );
  NAND21 U151 ( .A(SH[0]), .B(n15), .Q(n282) );
  CLKIN3 U152 ( .A(n121), .Q(B[27]) );
  NAND20 U153 ( .A(n119), .B(n19), .Q(n118) );
  CLKIN3 U154 ( .A(n103), .Q(B[31]) );
  AOI220 U155 ( .A(n30), .B(n41), .C(n35), .D(n42), .Q(n38) );
  MUX21 U156 ( .A(n146), .B(n147), .S(n18), .Q(B[1]) );
  NAND22 U157 ( .A(n18), .B(n122), .Q(n216) );
  NAND22 U158 ( .A(n18), .B(n119), .Q(n212) );
  NAND22 U159 ( .A(n47), .B(n48), .Q(B[7]) );
  NOR21 U160 ( .A(n51), .B(n52), .Q(n47) );
  NAND22 U161 ( .A(n57), .B(n58), .Q(n51) );
  NAND22 U162 ( .A(n233), .B(n234), .Q(B[10]) );
  INV3 U163 ( .A(n240), .Q(n233) );
  NAND22 U164 ( .A(n241), .B(n242), .Q(n240) );
  BUF2 U165 ( .A(n190), .Q(n10) );
  NOR21 U166 ( .A(SH[3]), .B(SH[2]), .Q(n12) );
  NOR21 U167 ( .A(SH[3]), .B(SH[2]), .Q(n13) );
  NOR21 U168 ( .A(SH[3]), .B(SH[2]), .Q(n101) );
  AOI220 U169 ( .A(A[23]), .B(n192), .C(A[24]), .D(n193), .Q(n196) );
  NAND22 U170 ( .A(n113), .B(n114), .Q(n111) );
  INV3 U171 ( .A(n127), .Q(n102) );
  NAND22 U172 ( .A(n100), .B(n132), .Q(n145) );
  INV3 U173 ( .A(n274), .Q(n96) );
  NAND22 U174 ( .A(n100), .B(n104), .Q(n95) );
  NAND22 U175 ( .A(n130), .B(n131), .Q(n40) );
  NAND22 U176 ( .A(n120), .B(n13), .Q(n130) );
  NAND22 U177 ( .A(n102), .B(n132), .Q(n131) );
  NAND22 U178 ( .A(n235), .B(n236), .Q(n124) );
  NAND22 U179 ( .A(n102), .B(n139), .Q(n236) );
  NAND22 U180 ( .A(n260), .B(n261), .Q(n164) );
  CLKIN3 U181 ( .A(n95), .Q(n152) );
  NOR21 U182 ( .A(n18), .B(n136), .Q(B[22]) );
  NAND22 U183 ( .A(n100), .B(n97), .Q(n135) );
  NAND22 U184 ( .A(n148), .B(n149), .Q(n146) );
  AOI221 U185 ( .A(n102), .B(n33), .C(n13), .D(n34), .Q(n148) );
  NAND22 U186 ( .A(n100), .B(n139), .Q(n138) );
  NAND22 U187 ( .A(n98), .B(n99), .Q(n90) );
  AOI221 U188 ( .A(n100), .B(n60), .C(n96), .D(n55), .Q(n99) );
  NAND22 U189 ( .A(n217), .B(n218), .Q(n50) );
  NAND22 U190 ( .A(n81), .B(n82), .Q(n77) );
  NAND22 U191 ( .A(n71), .B(n72), .Q(n65) );
  NAND22 U192 ( .A(n24), .B(n25), .Q(n23) );
  NAND22 U193 ( .A(n26), .B(n27), .Q(n25) );
  NAND22 U194 ( .A(n79), .B(n80), .Q(n78) );
  NAND22 U195 ( .A(n53), .B(n54), .Q(n52) );
  NAND22 U196 ( .A(n28), .B(n56), .Q(n53) );
  NAND22 U197 ( .A(n26), .B(n55), .Q(n54) );
  NAND22 U198 ( .A(n67), .B(n68), .Q(n66) );
  NAND22 U199 ( .A(n179), .B(n180), .Q(n178) );
  NAND22 U200 ( .A(n28), .B(n110), .Q(n179) );
  INV3 U201 ( .A(n173), .Q(n97) );
  NOR21 U202 ( .A(n18), .B(n163), .Q(B[16]) );
  NAND22 U203 ( .A(n87), .B(n88), .Q(n86) );
  NOR21 U204 ( .A(n167), .B(n168), .Q(n166) );
  NAND22 U205 ( .A(n169), .B(n170), .Q(n168) );
  NOR21 U206 ( .A(n18), .B(n123), .Q(B[26]) );
  NAND22 U207 ( .A(n174), .B(n175), .Q(B[14]) );
  NOR21 U208 ( .A(n177), .B(n178), .Q(n174) );
  INV3 U209 ( .A(n176), .Q(n109) );
  INV3 U210 ( .A(n89), .Q(n85) );
  INV3 U211 ( .A(n201), .Q(n200) );
  NAND22 U212 ( .A(n270), .B(n271), .Q(n259) );
  AOI221 U213 ( .A(n13), .B(n46), .C(n102), .D(n45), .Q(n270) );
  NAND31 U214 ( .A(n185), .B(n186), .C(n187), .Q(n184) );
  NAND22 U215 ( .A(n204), .B(n205), .Q(n27) );
  INV3 U216 ( .A(n19), .Q(n18) );
  NAND22 U217 ( .A(n188), .B(n189), .Q(n36) );
  NAND22 U218 ( .A(n229), .B(n230), .Q(n55) );
  NAND22 U219 ( .A(n268), .B(n269), .Q(n43) );
  NAND22 U220 ( .A(n246), .B(n247), .Q(n70) );
  NAND22 U221 ( .A(n249), .B(n250), .Q(n69) );
  NAND22 U222 ( .A(n266), .B(n267), .Q(n44) );
  NAND22 U223 ( .A(n252), .B(n253), .Q(n74) );
  NAND22 U224 ( .A(n231), .B(n232), .Q(n60) );
  NAND31 U225 ( .A(n215), .B(n216), .C(n214), .Q(B[11]) );
  NOR21 U226 ( .A(n18), .B(n115), .Q(B[29]) );
  INV3 U227 ( .A(n277), .Q(n100) );
  NAND22 U228 ( .A(n206), .B(n207), .Q(n33) );
  NAND22 U229 ( .A(n255), .B(n256), .Q(n73) );
  NAND22 U230 ( .A(n275), .B(n276), .Q(n41) );
  NAND22 U231 ( .A(n202), .B(n203), .Q(n31) );
  NAND22 U232 ( .A(n12), .B(n19), .Q(n254) );
  NAND22 U233 ( .A(n219), .B(n220), .Q(n59) );
  NAND22 U234 ( .A(n165), .B(n166), .Q(B[15]) );
  NOR21 U235 ( .A(n18), .B(n75), .Q(B[21]) );
  INV3 U236 ( .A(n107), .Q(B[30]) );
  NAND22 U237 ( .A(n109), .B(n19), .Q(n107) );
  NAND22 U238 ( .A(n122), .B(n19), .Q(n121) );
  INV3 U239 ( .A(n118), .Q(B[28]) );
  NAND22 U240 ( .A(n105), .B(n19), .Q(n103) );
  MUX22 U241 ( .A(n90), .B(n91), .S(n18), .Q(B[3]) );
  NOR21 U242 ( .A(n22), .B(n23), .Q(n21) );
  NOR21 U243 ( .A(n77), .B(n78), .Q(n76) );
  NAND31 U244 ( .A(n211), .B(n212), .C(n210), .Q(B[12]) );
  AOI220 U245 ( .A(n26), .B(n44), .C(n28), .D(n120), .Q(n211) );
  NAND31 U246 ( .A(n38), .B(n39), .C(n37), .Q(B[8]) );
  NAND22 U247 ( .A(n61), .B(n62), .Q(B[6]) );
  NOR21 U248 ( .A(n65), .B(n66), .Q(n61) );
  OAI212 U249 ( .A(n75), .B(n19), .C(n76), .Q(B[5]) );
  AOI221 U250 ( .A(A[26]), .B(n9), .C(A[27]), .D(n191), .Q(n239) );
  AOI220 U251 ( .A(A[27]), .B(n192), .C(A[28]), .D(n193), .Q(n194) );
  AOI220 U252 ( .A(A[26]), .B(n192), .C(A[27]), .D(n193), .Q(n264) );
  AOI221 U253 ( .A(A[27]), .B(n7), .C(A[28]), .D(n191), .Q(n224) );
  INV1 U254 ( .A(SH[3]), .Q(n17) );
  AOI220 U255 ( .A(A[5]), .B(n9), .C(A[6]), .D(n191), .Q(n207) );
  NAND22 U256 ( .A(n278), .B(n279), .Q(n45) );
  NAND22 U257 ( .A(n257), .B(n258), .Q(n64) );
  AOI220 U258 ( .A(A[16]), .B(n9), .C(n191), .D(A[17]), .Q(n269) );
  AOI220 U259 ( .A(A[16]), .B(n192), .C(A[17]), .D(n193), .Q(n249) );
  AOI220 U260 ( .A(n192), .B(A[17]), .C(A[18]), .D(n193), .Q(n229) );
  NAND22 U261 ( .A(n35), .B(n31), .Q(n81) );
  AOI221 U262 ( .A(n96), .B(n36), .C(n100), .D(n31), .Q(n149) );
  NAND22 U263 ( .A(n35), .B(n74), .Q(n71) );
  AOI220 U264 ( .A(n30), .B(n74), .C(n35), .D(n69), .Q(n241) );
  AOI220 U265 ( .A(A[10]), .B(n7), .C(A[11]), .D(n191), .Q(n253) );
  AOI220 U266 ( .A(n35), .B(n56), .C(n18), .D(n105), .Q(n165) );
  AOI220 U267 ( .A(n26), .B(n56), .C(n28), .D(n106), .Q(n215) );
  NAND22 U268 ( .A(n280), .B(n281), .Q(n46) );
  NAND22 U269 ( .A(n198), .B(n199), .Q(n34) );
  AOI220 U270 ( .A(A[5]), .B(n192), .C(A[6]), .D(n193), .Q(n217) );
  AOI221 U271 ( .A(A[30]), .B(n9), .C(A[31]), .D(n191), .Q(n237) );
  AOI220 U272 ( .A(A[10]), .B(n192), .C(A[11]), .D(n193), .Q(n275) );
  NAND22 U273 ( .A(n96), .B(n97), .Q(n92) );
  NAND21 U274 ( .A(n13), .B(n97), .Q(n172) );
  AOI220 U275 ( .A(n192), .B(A[18]), .C(A[19]), .D(n193), .Q(n268) );
  NAND21 U276 ( .A(n18), .B(n63), .Q(n62) );
  AOI220 U277 ( .A(A[1]), .B(n11), .C(A[2]), .D(n191), .Q(n199) );
  AOI220 U278 ( .A(A[2]), .B(n192), .C(A[3]), .D(n193), .Q(n280) );
  AOI220 U279 ( .A(A[2]), .B(n10), .C(A[3]), .D(n191), .Q(n258) );
  INV3 U280 ( .A(SH[2]), .Q(n16) );
  AOI220 U281 ( .A(A[14]), .B(n192), .C(A[15]), .D(n193), .Q(n272) );
  AOI220 U282 ( .A(A[14]), .B(n8), .C(A[15]), .D(n191), .Q(n250) );
  AOI220 U283 ( .A(A[15]), .B(n11), .C(A[16]), .D(n191), .Q(n230) );
  AOI220 U284 ( .A(A[15]), .B(n192), .C(A[16]), .D(n193), .Q(n188) );
  AOI220 U285 ( .A(A[6]), .B(n192), .C(A[7]), .D(n193), .Q(n278) );
  AOI220 U286 ( .A(A[6]), .B(n11), .C(A[7]), .D(n191), .Q(n256) );
  AOI220 U287 ( .A(A[3]), .B(n192), .C(A[4]), .D(n193), .Q(n198) );
  AOI220 U288 ( .A(A[4]), .B(n8), .C(A[5]), .D(n191), .Q(n279) );
  AOI220 U289 ( .A(A[4]), .B(n192), .C(A[5]), .D(n193), .Q(n257) );
  AOI220 U290 ( .A(A[3]), .B(n9), .C(A[4]), .D(n191), .Q(n218) );
  AOI220 U291 ( .A(A[9]), .B(n192), .C(A[10]), .D(n193), .Q(n219) );
  AOI220 U292 ( .A(A[9]), .B(n10), .C(A[10]), .D(n191), .Q(n203) );
  AOI220 U293 ( .A(A[13]), .B(n192), .C(A[14]), .D(n193), .Q(n231) );
  AOI220 U294 ( .A(A[13]), .B(n10), .C(A[14]), .D(n191), .Q(n189) );
  AOI220 U295 ( .A(A[20]), .B(n192), .C(A[21]), .D(n193), .Q(n246) );
  AOI220 U296 ( .A(A[19]), .B(n192), .C(A[20]), .D(n193), .Q(n204) );
  AOI220 U297 ( .A(n11), .B(A[0]), .C(A[1]), .D(n191), .Q(n281) );
  AOI220 U298 ( .A(A[7]), .B(n9), .C(A[8]), .D(n191), .Q(n220) );
  AOI220 U299 ( .A(A[7]), .B(n192), .C(A[8]), .D(n193), .Q(n206) );
  AOI220 U300 ( .A(A[8]), .B(n192), .C(A[9]), .D(n193), .Q(n255) );
  AOI220 U301 ( .A(A[8]), .B(n7), .C(A[9]), .D(n191), .Q(n276) );
  AOI220 U302 ( .A(A[11]), .B(n192), .C(A[12]), .D(n193), .Q(n202) );
  AOI220 U303 ( .A(A[12]), .B(n192), .C(A[13]), .D(n193), .Q(n252) );
  AOI220 U304 ( .A(A[11]), .B(n10), .C(A[12]), .D(n191), .Q(n232) );
  OAI212 U305 ( .A(n20), .B(n19), .C(n21), .Q(B[9]) );
  OAI212 U306 ( .A(n83), .B(n19), .C(n84), .Q(B[4]) );
  CLKIN3 U307 ( .A(n124), .Q(n123) );
  CLKIN3 U308 ( .A(n49), .Q(n133) );
  CLKIN3 U309 ( .A(n140), .Q(n75) );
  CLKIN3 U310 ( .A(n143), .Q(n83) );
  CLKIN3 U311 ( .A(n147), .Q(n156) );
  CLKIN3 U312 ( .A(n164), .Q(n163) );
  NAND22 U313 ( .A(n182), .B(n183), .Q(B[13]) );
endmodule


module E_alu_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n_Logic0_, ML_int_1__31_, ML_int_1__30_, ML_int_1__29_, ML_int_1__28_,
         ML_int_1__27_, ML_int_1__26_, ML_int_1__25_, ML_int_1__24_,
         ML_int_1__23_, ML_int_1__22_, ML_int_1__21_, ML_int_1__20_,
         ML_int_1__19_, ML_int_1__18_, ML_int_1__17_, ML_int_1__16_,
         ML_int_1__15_, ML_int_1__14_, ML_int_1__13_, ML_int_1__12_,
         ML_int_1__11_, ML_int_1__10_, ML_int_1__9_, ML_int_1__8_,
         ML_int_1__7_, ML_int_1__6_, ML_int_1__5_, ML_int_1__4_, ML_int_1__3_,
         ML_int_1__2_, ML_int_1__1_, ML_int_1__0_, ML_int_2__31_,
         ML_int_2__30_, ML_int_2__29_, ML_int_2__28_, ML_int_2__27_,
         ML_int_2__26_, ML_int_2__25_, ML_int_2__24_, ML_int_2__23_,
         ML_int_2__22_, ML_int_2__21_, ML_int_2__20_, ML_int_2__19_,
         ML_int_2__18_, ML_int_2__17_, ML_int_2__16_, ML_int_2__15_,
         ML_int_2__14_, ML_int_2__13_, ML_int_2__12_, ML_int_2__11_,
         ML_int_2__10_, ML_int_2__9_, ML_int_2__8_, ML_int_2__7_, ML_int_2__6_,
         ML_int_2__5_, ML_int_2__4_, ML_int_2__3_, ML_int_2__2_, ML_int_2__1_,
         ML_int_2__0_, ML_int_3__31_, ML_int_3__30_, ML_int_3__29_,
         ML_int_3__28_, ML_int_3__27_, ML_int_3__26_, ML_int_3__25_,
         ML_int_3__24_, ML_int_3__23_, ML_int_3__22_, ML_int_3__21_,
         ML_int_3__20_, ML_int_3__19_, ML_int_3__18_, ML_int_3__17_,
         ML_int_3__16_, ML_int_3__15_, ML_int_3__14_, ML_int_3__13_,
         ML_int_3__12_, ML_int_3__11_, ML_int_3__10_, ML_int_3__9_,
         ML_int_3__8_, ML_int_3__7_, ML_int_3__6_, ML_int_3__5_, ML_int_3__4_,
         ML_int_3__3_, ML_int_3__2_, ML_int_3__1_, ML_int_3__0_, ML_int_4__31_,
         ML_int_4__30_, ML_int_4__29_, ML_int_4__28_, ML_int_4__27_,
         ML_int_4__26_, ML_int_4__25_, ML_int_4__24_, ML_int_4__23_,
         ML_int_4__22_, ML_int_4__21_, ML_int_4__20_, ML_int_4__19_,
         ML_int_4__18_, ML_int_4__17_, ML_int_4__16_, ML_int_4__15_,
         ML_int_4__14_, ML_int_4__13_, ML_int_4__12_, ML_int_4__11_,
         ML_int_4__10_, ML_int_4__9_, ML_int_4__8_, ML_int_4__7_, ML_int_4__6_,
         ML_int_4__5_, ML_int_4__4_, ML_int_4__3_, ML_int_4__2_, ML_int_4__1_,
         ML_int_4__0_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61;

  MUX26 M1_4_18 ( .A(ML_int_4__18_), .B(ML_int_4__2_), .S(n61), .Q(B[18]) );
  MUX26 M1_3_14 ( .A(ML_int_3__14_), .B(ML_int_3__6_), .S(n55), .Q(
        ML_int_4__14_) );
  MUX26 M1_3_12 ( .A(ML_int_3__12_), .B(ML_int_3__4_), .S(n55), .Q(
        ML_int_4__12_) );
  MUX22 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n39), .Q(ML_int_1__15_) );
  MUX22 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n41), .Q(ML_int_1__22_) );
  MUX22 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n41), .Q(ML_int_1__31_) );
  MUX22 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n37), .Q(ML_int_1__9_) );
  MUX22 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n41), .Q(ML_int_1__21_) );
  MUX22 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n39), .Q(ML_int_1__19_) );
  MUX22 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n40), .Q(ML_int_1__26_) );
  MUX22 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n38), .Q(ML_int_1__10_) );
  MUX22 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n40), .Q(ML_int_1__27_) );
  MUX22 M1_4_22 ( .A(ML_int_4__22_), .B(ML_int_4__6_), .S(n60), .Q(B[22]) );
  MUX22 M1_2_24 ( .A(ML_int_2__24_), .B(ML_int_2__20_), .S(n51), .Q(
        ML_int_3__24_) );
  MUX22 M1_4_23 ( .A(ML_int_4__23_), .B(ML_int_4__7_), .S(n60), .Q(B[23]) );
  MUX22 M1_3_28 ( .A(ML_int_3__28_), .B(ML_int_3__20_), .S(n58), .Q(
        ML_int_4__28_) );
  MUX21 M1_3_16 ( .A(ML_int_3__16_), .B(ML_int_3__8_), .S(n56), .Q(
        ML_int_4__16_) );
  MUX22 M1_4_21 ( .A(ML_int_4__21_), .B(ML_int_4__5_), .S(n60), .Q(B[21]) );
  MUX22 M1_3_31 ( .A(ML_int_3__31_), .B(ML_int_3__23_), .S(n59), .Q(
        ML_int_4__31_) );
  MUX22 M1_3_25 ( .A(ML_int_3__25_), .B(ML_int_3__17_), .S(n58), .Q(
        ML_int_4__25_) );
  MUX22 M1_2_29 ( .A(ML_int_2__29_), .B(ML_int_2__25_), .S(n52), .Q(
        ML_int_3__29_) );
  MUX22 M1_3_29 ( .A(ML_int_3__29_), .B(ML_int_3__21_), .S(n58), .Q(
        ML_int_4__29_) );
  MUX22 M1_3_20 ( .A(ML_int_3__20_), .B(ML_int_3__12_), .S(n57), .Q(
        ML_int_4__20_) );
  MUX22 M1_2_6 ( .A(ML_int_2__6_), .B(ML_int_2__2_), .S(n49), .Q(ML_int_3__6_)
         );
  MUX22 M1_2_4 ( .A(ML_int_2__4_), .B(ML_int_2__0_), .S(n48), .Q(ML_int_3__4_)
         );
  MUX22 M1_2_5 ( .A(ML_int_2__5_), .B(ML_int_2__1_), .S(n49), .Q(ML_int_3__5_)
         );
  MUX22 M1_2_19 ( .A(ML_int_2__19_), .B(ML_int_2__15_), .S(n52), .Q(
        ML_int_3__19_) );
  MUX22 M1_2_22 ( .A(ML_int_2__22_), .B(ML_int_2__18_), .S(n51), .Q(
        ML_int_3__22_) );
  MUX22 M1_1_19 ( .A(ML_int_1__19_), .B(ML_int_1__17_), .S(n45), .Q(
        ML_int_2__19_) );
  MUX22 M1_1_26 ( .A(ML_int_1__26_), .B(ML_int_1__24_), .S(n47), .Q(
        ML_int_2__26_) );
  MUX22 M1_2_16 ( .A(ML_int_2__16_), .B(ML_int_2__12_), .S(n52), .Q(
        ML_int_3__16_) );
  MUX22 M1_1_15 ( .A(ML_int_1__15_), .B(ML_int_1__13_), .S(n45), .Q(
        ML_int_2__15_) );
  MUX22 M1_1_22 ( .A(ML_int_1__22_), .B(ML_int_1__20_), .S(n46), .Q(
        ML_int_2__22_) );
  MUX22 M1_4_29 ( .A(ML_int_4__29_), .B(ML_int_4__13_), .S(n60), .Q(B[29]) );
  MUX22 M1_1_2 ( .A(ML_int_1__2_), .B(ML_int_1__0_), .S(n42), .Q(ML_int_2__2_)
         );
  MUX22 M1_4_20 ( .A(ML_int_4__20_), .B(ML_int_4__4_), .S(n60), .Q(B[20]) );
  MUX22 M1_3_19 ( .A(ML_int_3__19_), .B(ML_int_3__11_), .S(n56), .Q(
        ML_int_4__19_) );
  MUX22 M1_4_19 ( .A(ML_int_4__19_), .B(ML_int_4__3_), .S(n60), .Q(B[19]) );
  MUX22 M1_3_26 ( .A(ML_int_3__26_), .B(ML_int_3__18_), .S(n58), .Q(
        ML_int_4__26_) );
  MUX21 M1_1_28 ( .A(ML_int_1__28_), .B(ML_int_1__26_), .S(n47), .Q(
        ML_int_2__28_) );
  MUX21 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n41), .Q(ML_int_1__30_) );
  MUX21 M1_2_25 ( .A(ML_int_2__25_), .B(ML_int_2__21_), .S(n50), .Q(
        ML_int_3__25_) );
  MUX22 M1_2_8 ( .A(ML_int_2__8_), .B(ML_int_2__4_), .S(n49), .Q(ML_int_3__8_)
         );
  MUX22 M1_2_20 ( .A(ML_int_2__20_), .B(ML_int_2__16_), .S(n51), .Q(
        ML_int_3__20_) );
  MUX22 M1_2_28 ( .A(ML_int_2__28_), .B(ML_int_2__24_), .S(n49), .Q(
        ML_int_3__28_) );
  MUX21 M1_1_30 ( .A(ML_int_1__30_), .B(ML_int_1__28_), .S(n45), .Q(
        ML_int_2__30_) );
  MUX21 M1_2_31 ( .A(ML_int_2__31_), .B(ML_int_2__27_), .S(n52), .Q(
        ML_int_3__31_) );
  MUX22 M1_2_27 ( .A(ML_int_2__27_), .B(ML_int_2__23_), .S(n51), .Q(
        ML_int_3__27_) );
  MUX22 M1_3_27 ( .A(ML_int_3__27_), .B(ML_int_3__19_), .S(n58), .Q(
        ML_int_4__27_) );
  MUX21 M1_3_21 ( .A(ML_int_3__21_), .B(ML_int_3__13_), .S(n57), .Q(
        ML_int_4__21_) );
  MUX22 M1_2_26 ( .A(ML_int_2__26_), .B(ML_int_2__22_), .S(n52), .Q(
        ML_int_3__26_) );
  MUX24 M1_3_17 ( .A(ML_int_3__17_), .B(ML_int_3__9_), .S(n56), .Q(
        ML_int_4__17_) );
  MUX22 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n38), .Q(ML_int_1__11_) );
  MUX26 M1_2_7 ( .A(ML_int_2__7_), .B(ML_int_2__3_), .S(n49), .Q(ML_int_3__7_)
         );
  MUX22 M1_2_23 ( .A(ML_int_2__23_), .B(ML_int_2__19_), .S(n51), .Q(
        ML_int_3__23_) );
  MUX24 M1_1_12 ( .A(ML_int_1__12_), .B(ML_int_1__10_), .S(n44), .Q(
        ML_int_2__12_) );
  MUX24 M1_2_12 ( .A(ML_int_2__12_), .B(ML_int_2__8_), .S(n50), .Q(
        ML_int_3__12_) );
  MUX24 M1_2_15 ( .A(ML_int_2__15_), .B(ML_int_2__11_), .S(n52), .Q(
        ML_int_3__15_) );
  MUX22 M1_3_23 ( .A(ML_int_3__23_), .B(ML_int_3__15_), .S(n57), .Q(
        ML_int_4__23_) );
  MUX22 M1_3_15 ( .A(ML_int_3__15_), .B(ML_int_3__7_), .S(n56), .Q(
        ML_int_4__15_) );
  MUX24 M1_1_7 ( .A(ML_int_1__7_), .B(ML_int_1__5_), .S(n43), .Q(ML_int_2__7_)
         );
  MUX26 M1_1_5 ( .A(ML_int_1__5_), .B(ML_int_1__3_), .S(n43), .Q(ML_int_2__5_)
         );
  MUX22 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n38), .Q(ML_int_1__12_) );
  MUX24 M1_1_27 ( .A(ML_int_1__27_), .B(ML_int_1__25_), .S(n47), .Q(
        ML_int_2__27_) );
  MUX22 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n40), .Q(ML_int_1__25_) );
  MUX24 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n39), .Q(ML_int_1__17_) );
  MUX24 M1_1_17 ( .A(ML_int_1__17_), .B(ML_int_1__15_), .S(n45), .Q(
        ML_int_2__17_) );
  MUX24 M1_1_25 ( .A(ML_int_1__25_), .B(ML_int_1__23_), .S(n47), .Q(
        ML_int_2__25_) );
  MUX26 M1_1_23 ( .A(ML_int_1__23_), .B(ML_int_1__21_), .S(n46), .Q(
        ML_int_2__23_) );
  MUX22 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n36), .Q(ML_int_1__4_) );
  MUX22 M1_4_25 ( .A(ML_int_4__25_), .B(ML_int_4__9_), .S(n60), .Q(B[25]) );
  MUX24 M1_3_10 ( .A(ML_int_3__10_), .B(ML_int_3__2_), .S(n55), .Q(
        ML_int_4__10_) );
  MUX22 M1_2_30 ( .A(ML_int_2__30_), .B(ML_int_2__26_), .S(n52), .Q(
        ML_int_3__30_) );
  MUX24 M1_3_13 ( .A(ML_int_3__13_), .B(ML_int_3__5_), .S(n55), .Q(
        ML_int_4__13_) );
  MUX22 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n37), .Q(ML_int_1__8_) );
  MUX22 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n37), .Q(ML_int_1__6_) );
  MUX21 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n38), .Q(ML_int_1__13_) );
  MUX24 M1_4_30 ( .A(ML_int_4__30_), .B(ML_int_4__14_), .S(n60), .Q(B[30]) );
  MUX22 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n39), .Q(ML_int_1__16_) );
  MUX22 M1_1_9 ( .A(ML_int_1__9_), .B(ML_int_1__7_), .S(n43), .Q(ML_int_2__9_)
         );
  MUX24 M1_2_13 ( .A(ML_int_2__13_), .B(ML_int_2__9_), .S(n50), .Q(
        ML_int_3__13_) );
  MUX22 M1_1_13 ( .A(ML_int_1__13_), .B(ML_int_1__11_), .S(n44), .Q(
        ML_int_2__13_) );
  MUX24 M1_3_8 ( .A(ML_int_3__8_), .B(ML_int_3__0_), .S(n54), .Q(ML_int_4__8_)
         );
  MUX22 M1_4_17 ( .A(ML_int_4__17_), .B(ML_int_4__1_), .S(n61), .Q(B[17]) );
  MUX24 M1_1_8 ( .A(ML_int_1__8_), .B(ML_int_1__6_), .S(n43), .Q(ML_int_2__8_)
         );
  MUX22 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n37), .Q(ML_int_1__7_) );
  MUX24 M1_4_27 ( .A(ML_int_4__27_), .B(ML_int_4__11_), .S(n60), .Q(B[27]) );
  MUX24 M1_4_26 ( .A(ML_int_4__26_), .B(ML_int_4__10_), .S(n60), .Q(B[26]) );
  MUX24 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n41), .Q(ML_int_1__24_) );
  MUX22 M1_1_21 ( .A(ML_int_1__21_), .B(ML_int_1__19_), .S(n46), .Q(
        ML_int_2__21_) );
  MUX24 M1_2_21 ( .A(ML_int_2__21_), .B(ML_int_2__17_), .S(n51), .Q(
        ML_int_3__21_) );
  MUX24 M1_2_14 ( .A(ML_int_2__14_), .B(ML_int_2__10_), .S(n50), .Q(
        ML_int_3__14_) );
  MUX26 M1_1_14 ( .A(ML_int_1__14_), .B(ML_int_1__12_), .S(n44), .Q(
        ML_int_2__14_) );
  MUX24 M1_1_11 ( .A(ML_int_1__11_), .B(ML_int_1__9_), .S(n44), .Q(
        ML_int_2__11_) );
  MUX24 M1_3_11 ( .A(ML_int_3__11_), .B(ML_int_3__3_), .S(n55), .Q(
        ML_int_4__11_) );
  MUX22 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n38), .Q(ML_int_1__14_) );
  MUX24 M1_1_16 ( .A(ML_int_1__16_), .B(ML_int_1__14_), .S(n45), .Q(
        ML_int_2__16_) );
  MUX22 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n41), .Q(ML_int_1__20_) );
  MUX26 M1_1_20 ( .A(ML_int_1__20_), .B(ML_int_1__18_), .S(n46), .Q(
        ML_int_2__20_) );
  MUX26 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n39), .Q(ML_int_1__18_) );
  MUX24 M1_2_18 ( .A(ML_int_2__18_), .B(ML_int_2__14_), .S(n51), .Q(
        ML_int_3__18_) );
  MUX22 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n36), .Q(ML_int_1__3_) );
  MUX22 M1_2_17 ( .A(ML_int_2__17_), .B(ML_int_2__13_), .S(n52), .Q(
        ML_int_3__17_) );
  MUX22 M1_2_9 ( .A(ML_int_2__9_), .B(ML_int_2__5_), .S(n49), .Q(ML_int_3__9_)
         );
  MUX22 M1_2_11 ( .A(ML_int_2__11_), .B(ML_int_2__7_), .S(n50), .Q(
        ML_int_3__11_) );
  MUX22 M1_1_3 ( .A(ML_int_1__3_), .B(ML_int_1__1_), .S(n42), .Q(ML_int_2__3_)
         );
  MUX22 M1_1_4 ( .A(ML_int_1__4_), .B(ML_int_1__2_), .S(n42), .Q(ML_int_2__4_)
         );
  MUX21 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n36), .Q(ML_int_1__2_) );
  MUX21 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n36), .Q(ML_int_1__1_) );
  MUX24 M1_4_24 ( .A(ML_int_4__24_), .B(ML_int_4__8_), .S(n60), .Q(B[24]) );
  MUX24 M1_4_31 ( .A(ML_int_4__31_), .B(ML_int_4__15_), .S(n60), .Q(B[31]) );
  MUX24 M1_3_18 ( .A(ML_int_3__18_), .B(ML_int_3__10_), .S(n56), .Q(
        ML_int_4__18_) );
  MUX24 M1_1_6 ( .A(ML_int_1__6_), .B(ML_int_1__4_), .S(n43), .Q(ML_int_2__6_)
         );
  MUX24 M1_1_10 ( .A(ML_int_1__10_), .B(ML_int_1__8_), .S(n44), .Q(
        ML_int_2__10_) );
  MUX24 M1_2_10 ( .A(ML_int_2__10_), .B(ML_int_2__6_), .S(n50), .Q(
        ML_int_3__10_) );
  MUX22 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n40), .Q(ML_int_1__28_) );
  MUX22 M1_3_30 ( .A(ML_int_3__30_), .B(ML_int_3__22_), .S(n59), .Q(
        ML_int_4__30_) );
  MUX24 M1_3_22 ( .A(ML_int_3__22_), .B(ML_int_3__14_), .S(n57), .Q(
        ML_int_4__22_) );
  MUX22 M1_1_18 ( .A(ML_int_1__18_), .B(ML_int_1__16_), .S(n45), .Q(
        ML_int_2__18_) );
  MUX22 M1_4_16 ( .A(ML_int_4__16_), .B(ML_int_4__0_), .S(n61), .Q(B[16]) );
  MUX22 M1_1_31 ( .A(ML_int_1__31_), .B(ML_int_1__29_), .S(n47), .Q(
        ML_int_2__31_) );
  MUX22 M1_1_24 ( .A(ML_int_1__24_), .B(ML_int_1__22_), .S(n46), .Q(
        ML_int_2__24_) );
  MUX22 M1_3_24 ( .A(ML_int_3__24_), .B(ML_int_3__16_), .S(n57), .Q(
        ML_int_4__24_) );
  MUX22 M1_3_9 ( .A(ML_int_3__9_), .B(ML_int_3__1_), .S(n54), .Q(ML_int_4__9_)
         );
  MUX22 M1_1_29 ( .A(ML_int_1__29_), .B(ML_int_1__27_), .S(n47), .Q(
        ML_int_2__29_) );
  MUX22 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n40), .Q(ML_int_1__23_) );
  MUX22 M1_4_28 ( .A(ML_int_4__28_), .B(ML_int_4__12_), .S(n60), .Q(B[28]) );
  MUX22 M0_1_1 ( .A(ML_int_1__1_), .B(n_Logic0_), .S(n42), .Q(ML_int_2__1_) );
  NOR24 U3 ( .A(n48), .B(n1), .Q(ML_int_3__3_) );
  CLKIN6 U4 ( .A(ML_int_2__3_), .Q(n1) );
  INV1 U5 ( .A(ML_int_4__4_), .Q(n18) );
  NOR23 U6 ( .A(n53), .B(n26), .Q(ML_int_4__4_) );
  NAND22 U7 ( .A(n5), .B(n6), .Q(ML_int_1__29_) );
  NAND21 U8 ( .A(A[28]), .B(n40), .Q(n6) );
  NAND22 U9 ( .A(A[29]), .B(n4), .Q(n5) );
  NAND23 U10 ( .A(n2), .B(n3), .Q(ML_int_1__5_) );
  NOR23 U11 ( .A(n61), .B(n11), .Q(B[11]) );
  BUF2 U12 ( .A(SH[0]), .Q(n40) );
  INV3 U13 ( .A(ML_int_1__0_), .Q(n34) );
  INV3 U14 ( .A(ML_int_4__9_), .Q(n13) );
  NOR23 U15 ( .A(n61), .B(n8), .Q(B[14]) );
  NAND22 U16 ( .A(A[5]), .B(n4), .Q(n2) );
  NOR22 U17 ( .A(n54), .B(n23), .Q(ML_int_4__7_) );
  INV3 U18 ( .A(ML_int_3__7_), .Q(n23) );
  INV2 U19 ( .A(ML_int_4__7_), .Q(n15) );
  CLKIN4 U20 ( .A(ML_int_2__2_), .Q(n31) );
  INV2 U21 ( .A(A[0]), .Q(n35) );
  NOR23 U22 ( .A(n53), .B(n28), .Q(ML_int_4__2_) );
  CLKIN3 U23 ( .A(ML_int_3__2_), .Q(n28) );
  NOR22 U24 ( .A(n53), .B(n30), .Q(ML_int_4__0_) );
  CLKIN6 U25 ( .A(ML_int_4__0_), .Q(n22) );
  NOR23 U26 ( .A(n48), .B(n33), .Q(ML_int_3__0_) );
  CLKIN3 U27 ( .A(ML_int_4__13_), .Q(n9) );
  NOR22 U28 ( .A(n61), .B(n7), .Q(B[15]) );
  CLKIN2 U29 ( .A(ML_int_4__15_), .Q(n7) );
  NAND21 U30 ( .A(A[4]), .B(n37), .Q(n3) );
  INV3 U31 ( .A(n40), .Q(n4) );
  NOR22 U32 ( .A(n36), .B(n35), .Q(ML_int_1__0_) );
  NOR24 U33 ( .A(n42), .B(n34), .Q(ML_int_2__0_) );
  CLKIN0 U34 ( .A(ML_int_4__10_), .Q(n12) );
  CLKIN1 U35 ( .A(ML_int_4__6_), .Q(n16) );
  INV2 U36 ( .A(ML_int_2__0_), .Q(n33) );
  INV1 U37 ( .A(ML_int_3__0_), .Q(n30) );
  CLKIN0 U38 ( .A(ML_int_4__2_), .Q(n20) );
  INV3 U39 ( .A(ML_int_4__14_), .Q(n8) );
  CLKIN0 U40 ( .A(ML_int_4__12_), .Q(n10) );
  INV1 U41 ( .A(ML_int_4__1_), .Q(n21) );
  NOR23 U42 ( .A(n48), .B(n32), .Q(ML_int_3__1_) );
  CLKIN2 U43 ( .A(ML_int_2__1_), .Q(n32) );
  NOR24 U44 ( .A(n48), .B(n31), .Q(ML_int_3__2_) );
  NOR22 U45 ( .A(n53), .B(n27), .Q(ML_int_4__3_) );
  CLKIN0 U46 ( .A(ML_int_4__8_), .Q(n14) );
  CLKIN0 U47 ( .A(ML_int_4__3_), .Q(n19) );
  INV1 U48 ( .A(ML_int_4__5_), .Q(n17) );
  BUF2 U49 ( .A(SH[4]), .Q(n60) );
  NOR21 U50 ( .A(n54), .B(n25), .Q(ML_int_4__5_) );
  INV3 U51 ( .A(ML_int_3__5_), .Q(n25) );
  NOR21 U52 ( .A(n54), .B(n24), .Q(ML_int_4__6_) );
  INV3 U53 ( .A(ML_int_3__6_), .Q(n24) );
  NOR21 U54 ( .A(n53), .B(n29), .Q(ML_int_4__1_) );
  INV3 U55 ( .A(ML_int_3__1_), .Q(n29) );
  INV3 U56 ( .A(ML_int_3__3_), .Q(n27) );
  INV3 U57 ( .A(ML_int_3__4_), .Q(n26) );
  NOR21 U58 ( .A(n61), .B(n12), .Q(B[10]) );
  BUF2 U59 ( .A(SH[0]), .Q(n39) );
  NOR21 U60 ( .A(n61), .B(n10), .Q(B[12]) );
  NOR21 U61 ( .A(n61), .B(n16), .Q(B[6]) );
  NOR21 U62 ( .A(n61), .B(n15), .Q(B[7]) );
  NOR21 U63 ( .A(n61), .B(n14), .Q(B[8]) );
  NOR21 U64 ( .A(n61), .B(n13), .Q(B[9]) );
  INV3 U65 ( .A(ML_int_4__11_), .Q(n11) );
  NOR21 U66 ( .A(n61), .B(n9), .Q(B[13]) );
  NOR21 U67 ( .A(n61), .B(n22), .Q(B[0]) );
  BUF2 U68 ( .A(SH[0]), .Q(n36) );
  BUF2 U69 ( .A(SH[0]), .Q(n38) );
  NOR21 U70 ( .A(n61), .B(n21), .Q(B[1]) );
  NOR21 U71 ( .A(n61), .B(n20), .Q(B[2]) );
  NOR21 U72 ( .A(n61), .B(n19), .Q(B[3]) );
  NOR21 U73 ( .A(n61), .B(n18), .Q(B[4]) );
  NOR21 U74 ( .A(n61), .B(n17), .Q(B[5]) );
  BUF2 U75 ( .A(SH[0]), .Q(n37) );
  BUF2 U76 ( .A(SH[0]), .Q(n41) );
  BUF2 U77 ( .A(SH[1]), .Q(n47) );
  BUF2 U78 ( .A(SH[1]), .Q(n45) );
  BUF2 U79 ( .A(SH[1]), .Q(n46) );
  BUF2 U80 ( .A(SH[1]), .Q(n43) );
  BUF2 U81 ( .A(SH[1]), .Q(n44) );
  BUF2 U82 ( .A(SH[1]), .Q(n42) );
  BUF2 U83 ( .A(SH[4]), .Q(n61) );
  BUF2 U84 ( .A(SH[2]), .Q(n52) );
  LOGIC0 U85 ( .Q(n_Logic0_) );
  BUF2 U86 ( .A(SH[3]), .Q(n59) );
  BUF2 U87 ( .A(SH[3]), .Q(n57) );
  BUF2 U88 ( .A(SH[3]), .Q(n58) );
  BUF2 U89 ( .A(SH[3]), .Q(n54) );
  BUF2 U90 ( .A(SH[3]), .Q(n53) );
  BUF2 U91 ( .A(SH[3]), .Q(n56) );
  BUF2 U92 ( .A(SH[3]), .Q(n55) );
  BUF2 U93 ( .A(SH[2]), .Q(n48) );
  BUF2 U94 ( .A(SH[2]), .Q(n50) );
  BUF2 U95 ( .A(SH[2]), .Q(n49) );
  BUF2 U96 ( .A(SH[2]), .Q(n51) );
endmodule


module E_alu_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421;

  CLKIN3 U3 ( .A(n361), .Q(n357) );
  CLKIN8 U4 ( .A(n211), .Q(n187) );
  INV6 U5 ( .A(n50), .Q(n51) );
  INV3 U6 ( .A(n82), .Q(n1) );
  IMUX22 U7 ( .A(n311), .B(n312), .S(n313), .Q(DIFF[16]) );
  INV6 U8 ( .A(n169), .Q(n164) );
  INV6 U9 ( .A(n57), .Q(n58) );
  NAND28 U10 ( .A(n387), .B(n388), .Q(n113) );
  INV6 U11 ( .A(n355), .Q(n2) );
  CLKIN6 U12 ( .A(n341), .Q(n355) );
  AOI211 U13 ( .A(B[23]), .B(n240), .C(n241), .Q(n233) );
  INV2 U14 ( .A(n242), .Q(n241) );
  CLKIN12 U15 ( .A(n118), .Q(n403) );
  NAND23 U16 ( .A(B[2]), .B(n404), .Q(n118) );
  BUF2 U17 ( .A(n221), .Q(n30) );
  INV12 U18 ( .A(n221), .Q(n317) );
  INV10 U19 ( .A(n386), .Q(n348) );
  NAND23 U20 ( .A(n385), .B(n386), .Q(n382) );
  CLKIN1 U21 ( .A(B[14]), .Q(n351) );
  NAND26 U22 ( .A(n24), .B(B[7]), .Q(n23) );
  INV3 U23 ( .A(A[7]), .Q(n24) );
  INV6 U24 ( .A(B[15]), .Q(n325) );
  NOR22 U25 ( .A(A[27]), .B(n186), .Q(n185) );
  NOR22 U26 ( .A(n159), .B(n403), .Q(n398) );
  INV6 U27 ( .A(B[13]), .Q(n324) );
  NAND22 U28 ( .A(n155), .B(n156), .Q(n140) );
  CLKIN6 U29 ( .A(n340), .Q(n334) );
  NOR22 U30 ( .A(n126), .B(n140), .Q(n122) );
  INV6 U31 ( .A(n62), .Q(n86) );
  INV6 U32 ( .A(n89), .Q(n374) );
  NAND26 U33 ( .A(n228), .B(n229), .Q(n175) );
  NAND24 U34 ( .A(A[18]), .B(n304), .Q(n275) );
  XNR21 U35 ( .A(n115), .B(n116), .Q(DIFF[3]) );
  INV6 U36 ( .A(n373), .Q(n376) );
  INV6 U37 ( .A(B[20]), .Q(n247) );
  CLKIN3 U38 ( .A(n22), .Q(n25) );
  INV3 U39 ( .A(n325), .Q(n22) );
  NOR23 U40 ( .A(A[19]), .B(n278), .Q(n282) );
  NOR24 U41 ( .A(A[20]), .B(n247), .Q(n284) );
  NAND28 U42 ( .A(B[17]), .B(n310), .Q(n270) );
  NOR24 U43 ( .A(A[0]), .B(n289), .Q(n288) );
  INV8 U44 ( .A(B[9]), .Q(n372) );
  INV6 U45 ( .A(n318), .Q(n8) );
  NAND26 U46 ( .A(n7), .B(n137), .Q(n315) );
  NOR21 U47 ( .A(n46), .B(n26), .Q(n19) );
  NAND24 U48 ( .A(B[22]), .B(n258), .Q(n242) );
  CLKIN2 U49 ( .A(B[22]), .Q(n257) );
  CLKIN4 U50 ( .A(B[11]), .Q(n367) );
  CLKIN6 U51 ( .A(B[12]), .Q(n326) );
  NAND24 U52 ( .A(n15), .B(B[4]), .Q(n14) );
  INV6 U53 ( .A(B[4]), .Q(n110) );
  NOR21 U54 ( .A(n30), .B(n210), .Q(n214) );
  NAND22 U55 ( .A(A[14]), .B(n351), .Q(n332) );
  NAND26 U56 ( .A(n73), .B(n187), .Q(n154) );
  NAND22 U57 ( .A(n250), .B(n71), .Q(n67) );
  INV3 U58 ( .A(n306), .Q(n33) );
  INV3 U59 ( .A(n14), .Q(n407) );
  INV3 U60 ( .A(A[4]), .Q(n15) );
  INV6 U61 ( .A(B[19]), .Q(n278) );
  NOR32 U62 ( .A(n159), .B(B[0]), .C(n403), .Q(n400) );
  NOR22 U63 ( .A(n401), .B(n402), .Q(n399) );
  INV0 U64 ( .A(n332), .Q(n339) );
  INV6 U65 ( .A(n28), .Q(n281) );
  NAND24 U66 ( .A(n29), .B(B[16]), .Q(n28) );
  INV3 U67 ( .A(A[16]), .Q(n29) );
  NAND22 U68 ( .A(B[24]), .B(n222), .Q(n204) );
  INV6 U69 ( .A(B[16]), .Q(n283) );
  NOR21 U70 ( .A(n140), .B(n154), .Q(n152) );
  NAND23 U71 ( .A(n102), .B(n103), .Q(n96) );
  NAND22 U72 ( .A(A[21]), .B(n264), .Q(n237) );
  NAND22 U73 ( .A(n243), .B(n262), .Q(n263) );
  XOR20 U74 ( .A(B[27]), .B(A[27]), .Q(n192) );
  NAND22 U75 ( .A(n184), .B(n182), .Q(n201) );
  INV6 U76 ( .A(n34), .Q(n248) );
  NAND26 U77 ( .A(n63), .B(n65), .Q(n34) );
  NAND28 U78 ( .A(n166), .B(n148), .Q(n165) );
  INV8 U79 ( .A(B[17]), .Q(n309) );
  INV6 U80 ( .A(n55), .Q(n377) );
  NAND20 U81 ( .A(n201), .B(n193), .Q(n5) );
  NAND22 U82 ( .A(n3), .B(n4), .Q(n6) );
  NAND22 U83 ( .A(n5), .B(n6), .Q(DIFF[25]) );
  INV3 U84 ( .A(n201), .Q(n3) );
  INV2 U85 ( .A(n193), .Q(n4) );
  NAND26 U86 ( .A(n203), .B(n202), .Q(n193) );
  NAND24 U87 ( .A(n358), .B(n13), .Q(n356) );
  NAND26 U88 ( .A(A[11]), .B(n80), .Q(n370) );
  OAI212 U89 ( .A(n7), .B(n217), .C(n218), .Q(n216) );
  NAND23 U90 ( .A(n187), .B(n204), .Q(n217) );
  NAND28 U91 ( .A(A[17]), .B(n309), .Q(n277) );
  NAND21 U92 ( .A(n298), .B(n277), .Q(n297) );
  NAND34 U93 ( .A(n8), .B(n19), .C(n319), .Q(n7) );
  NAND24 U94 ( .A(B[14]), .B(n352), .Q(n320) );
  INV6 U95 ( .A(n269), .Q(n231) );
  NAND33 U96 ( .A(n242), .B(n153), .C(n249), .Q(n63) );
  NAND23 U97 ( .A(n76), .B(n357), .Q(n360) );
  XOR20 U98 ( .A(B[29]), .B(A[29]), .Q(n9) );
  XOR20 U99 ( .A(B[30]), .B(A[30]), .Q(n10) );
  XNR20 U100 ( .A(n1), .B(A[23]), .Q(n11) );
  XNR20 U101 ( .A(B[28]), .B(A[28]), .Q(n12) );
  CLKIN6 U102 ( .A(n113), .Q(n107) );
  INV3 U103 ( .A(n290), .Q(n421) );
  NAND24 U104 ( .A(n317), .B(n113), .Q(n386) );
  NAND22 U105 ( .A(B[26]), .B(n200), .Q(n177) );
  CLKIN3 U106 ( .A(n177), .Q(n195) );
  CLKIN15 U107 ( .A(B[23]), .Q(n232) );
  NOR22 U108 ( .A(A[3]), .B(n392), .Q(n401) );
  CLKIN4 U109 ( .A(n137), .Q(n219) );
  NOR24 U110 ( .A(A[11]), .B(n80), .Q(n318) );
  CLKIN12 U111 ( .A(n79), .Q(n80) );
  NOR23 U112 ( .A(n350), .B(n348), .Q(n62) );
  CLKIN12 U113 ( .A(n321), .Q(n26) );
  NAND28 U114 ( .A(n77), .B(n35), .Q(n134) );
  NOR24 U115 ( .A(n46), .B(n26), .Q(n35) );
  INV12 U116 ( .A(B[3]), .Q(n392) );
  NAND28 U117 ( .A(n48), .B(n317), .Q(n57) );
  NAND24 U118 ( .A(n67), .B(n68), .Q(n65) );
  INV4 U119 ( .A(B[1]), .Q(n393) );
  NAND24 U120 ( .A(A[1]), .B(n393), .Q(n161) );
  INV1 U121 ( .A(n335), .Q(n13) );
  CLKIN6 U122 ( .A(n359), .Q(n335) );
  CLKIN12 U123 ( .A(n416), .Q(n87) );
  BUF2 U124 ( .A(n76), .Q(n16) );
  CLKIN2 U125 ( .A(n97), .Q(n100) );
  CLKIN1 U126 ( .A(n101), .Q(n98) );
  NAND28 U127 ( .A(n270), .B(n271), .Q(n17) );
  NAND28 U128 ( .A(n280), .B(n18), .Q(n279) );
  INV12 U129 ( .A(n17), .Q(n18) );
  NOR23 U130 ( .A(n281), .B(n282), .Q(n280) );
  INV12 U131 ( .A(n279), .Q(n243) );
  INV4 U132 ( .A(B[7]), .Q(n27) );
  NAND24 U133 ( .A(n356), .B(n357), .Q(n341) );
  NAND22 U134 ( .A(A[12]), .B(n326), .Q(n359) );
  OAI211 U135 ( .A(n134), .B(n136), .C(n137), .Q(n132) );
  NAND22 U136 ( .A(A[15]), .B(n25), .Q(n333) );
  NOR23 U137 ( .A(n334), .B(n335), .Q(n330) );
  NOR42 U138 ( .A(n378), .B(n376), .C(n377), .D(n375), .Q(n76) );
  NAND23 U139 ( .A(n372), .B(A[9]), .Q(n89) );
  NAND26 U140 ( .A(B[10]), .B(n419), .Q(n373) );
  CLKIN3 U141 ( .A(B[10]), .Q(n418) );
  INV3 U142 ( .A(n49), .Q(n20) );
  INV0 U143 ( .A(n326), .Q(n21) );
  NOR20 U144 ( .A(A[12]), .B(n326), .Q(n361) );
  XNR22 U145 ( .A(n94), .B(n95), .Q(DIFF[7]) );
  INV12 U146 ( .A(n42), .Q(n43) );
  AOI211 U147 ( .A(n117), .B(n118), .C(n119), .Q(n116) );
  NAND24 U148 ( .A(n410), .B(n411), .Q(n135) );
  NOR24 U149 ( .A(A[13]), .B(n324), .Q(n323) );
  NAND23 U150 ( .A(n341), .B(n340), .Q(n36) );
  INV6 U151 ( .A(n367), .Q(n79) );
  CLKIN12 U152 ( .A(n23), .Q(n408) );
  NAND23 U153 ( .A(n104), .B(n105), .Q(n102) );
  NAND28 U154 ( .A(B[5]), .B(n409), .Q(n105) );
  INV10 U155 ( .A(n45), .Q(n46) );
  NAND26 U156 ( .A(n175), .B(n73), .Q(n174) );
  NAND28 U157 ( .A(A[8]), .B(n93), .Q(n416) );
  INV3 U158 ( .A(B[24]), .Q(n190) );
  CLKIN4 U159 ( .A(B[5]), .Q(n414) );
  XOR22 U160 ( .A(n344), .B(n345), .Q(DIFF[14]) );
  NOR23 U161 ( .A(n288), .B(n391), .Q(n397) );
  INV0 U162 ( .A(n358), .Q(n366) );
  AOI212 U163 ( .A(n153), .B(n249), .C(n253), .Q(n252) );
  NAND28 U164 ( .A(n136), .B(n135), .Q(n350) );
  NAND21 U165 ( .A(n35), .B(n76), .Q(n220) );
  XOR22 U166 ( .A(n9), .B(n163), .Q(DIFF[29]) );
  NOR24 U167 ( .A(n189), .B(n185), .Q(n188) );
  NAND26 U168 ( .A(n394), .B(n395), .Q(n389) );
  NOR24 U169 ( .A(n389), .B(n390), .Q(n388) );
  XNR21 U170 ( .A(n104), .B(n106), .Q(DIFF[5]) );
  NAND28 U171 ( .A(n173), .B(n174), .Q(n123) );
  NAND24 U172 ( .A(n122), .B(n139), .Q(n129) );
  NOR24 U173 ( .A(n129), .B(n130), .Q(n124) );
  CLKIN12 U174 ( .A(B[8]), .Q(n93) );
  NAND24 U175 ( .A(n56), .B(B[8]), .Q(n55) );
  AOI211 U176 ( .A(n96), .B(n97), .C(n98), .Q(n95) );
  NAND24 U177 ( .A(n261), .B(n236), .Q(n254) );
  NAND23 U178 ( .A(A[10]), .B(n418), .Q(n371) );
  AOI311 U179 ( .A(n85), .B(n88), .C(n382), .D(n374), .Q(n381) );
  XOR22 U180 ( .A(n64), .B(n380), .Q(DIFF[11]) );
  NOR24 U181 ( .A(n210), .B(n211), .Q(n213) );
  NAND24 U182 ( .A(B[1]), .B(n405), .Q(n291) );
  NOR21 U183 ( .A(A[15]), .B(n25), .Q(n329) );
  CLKIN2 U184 ( .A(n131), .Q(n31) );
  INV3 U185 ( .A(n31), .Q(n32) );
  CLKIN6 U186 ( .A(n291), .Q(n159) );
  NOR33 U187 ( .A(n161), .B(n391), .C(n403), .Q(n390) );
  NOR24 U188 ( .A(A[3]), .B(n392), .Q(n391) );
  XOR22 U189 ( .A(n10), .B(n142), .Q(DIFF[30]) );
  INV6 U190 ( .A(n151), .Q(n143) );
  INV6 U191 ( .A(n360), .Q(n349) );
  NAND23 U192 ( .A(A[6]), .B(n413), .Q(n101) );
  NAND23 U193 ( .A(n145), .B(n127), .Q(n144) );
  XNR22 U194 ( .A(n33), .B(n307), .Q(DIFF[17]) );
  AOI312 U195 ( .A(n271), .B(n294), .C(n153), .D(n295), .Q(n292) );
  NAND21 U196 ( .A(n296), .B(n275), .Q(n295) );
  NAND22 U197 ( .A(n212), .B(n213), .Q(n207) );
  OAI210 U198 ( .A(A[13]), .B(n324), .C(n320), .Q(n331) );
  NOR23 U199 ( .A(A[24]), .B(n190), .Q(n189) );
  NOR24 U200 ( .A(n407), .B(n408), .Q(n406) );
  NAND26 U201 ( .A(n327), .B(n328), .Q(n137) );
  NAND21 U202 ( .A(A[24]), .B(n190), .Q(n181) );
  OAI212 U203 ( .A(A[9]), .B(n372), .C(n373), .Q(n369) );
  NAND28 U204 ( .A(B[6]), .B(n415), .Q(n97) );
  OAI2112 U205 ( .A(n369), .B(n368), .C(n370), .D(n371), .Q(n319) );
  CLKIN1 U206 ( .A(n416), .Q(n78) );
  NAND28 U207 ( .A(n105), .B(n97), .Q(n42) );
  NOR22 U208 ( .A(n134), .B(n136), .Q(n209) );
  NAND22 U209 ( .A(A[7]), .B(n27), .Q(n136) );
  NOR23 U210 ( .A(n44), .B(n100), .Q(n410) );
  NOR23 U211 ( .A(n27), .B(A[7]), .Q(n44) );
  XOR22 U212 ( .A(n251), .B(n252), .Q(DIFF[22]) );
  NOR24 U213 ( .A(n164), .B(n165), .Q(n163) );
  AOI212 U214 ( .A(n294), .B(n153), .C(n297), .Q(n300) );
  NAND22 U215 ( .A(n123), .B(n156), .Q(n166) );
  NAND24 U216 ( .A(n342), .B(n37), .Q(n50) );
  INV4 U217 ( .A(n36), .Q(n37) );
  NAND22 U218 ( .A(n209), .B(n213), .Q(n208) );
  NAND24 U219 ( .A(A[4]), .B(n110), .Q(n109) );
  INV12 U220 ( .A(n314), .Q(n153) );
  XOR22 U221 ( .A(n353), .B(n354), .Q(DIFF[13]) );
  INV6 U222 ( .A(B[0]), .Q(n289) );
  CLKIN3 U223 ( .A(B[6]), .Q(n413) );
  NOR21 U224 ( .A(n211), .B(n220), .Q(n215) );
  NAND28 U225 ( .A(n230), .B(n243), .Q(n211) );
  CLKIN2 U226 ( .A(B[21]), .Q(n264) );
  NAND21 U227 ( .A(n191), .B(n39), .Q(n40) );
  NAND24 U228 ( .A(n38), .B(n192), .Q(n41) );
  NAND24 U229 ( .A(n40), .B(n41), .Q(DIFF[27]) );
  CLKIN4 U230 ( .A(n191), .Q(n38) );
  INV0 U231 ( .A(n192), .Q(n39) );
  NAND28 U232 ( .A(n406), .B(n43), .Q(n221) );
  AOI212 U233 ( .A(n16), .B(n86), .C(n366), .Q(n365) );
  NAND24 U234 ( .A(n343), .B(n51), .Q(n338) );
  AOI312 U235 ( .A(n342), .B(n2), .C(n343), .D(n347), .Q(n346) );
  NOR32 U236 ( .A(n32), .B(n132), .C(n133), .Q(n130) );
  AOI222 U237 ( .A(n82), .B(A[23]), .C(n233), .D(n234), .Q(n228) );
  INV0 U238 ( .A(n109), .Q(n114) );
  AOI212 U239 ( .A(n349), .B(n86), .C(n355), .Q(n354) );
  NOR21 U240 ( .A(n154), .B(n171), .Q(n170) );
  AOI2112 U241 ( .A(n204), .B(n175), .C(n206), .D(n205), .Q(n203) );
  NAND24 U242 ( .A(n61), .B(n8), .Q(n358) );
  OAI2112 U243 ( .A(n369), .B(n368), .C(n370), .D(n371), .Q(n61) );
  AOI211 U244 ( .A(n187), .B(n153), .C(n175), .Q(n227) );
  AOI211 U245 ( .A(n243), .B(n153), .C(n231), .Q(n268) );
  NOR23 U246 ( .A(n78), .B(n350), .Q(n385) );
  NAND24 U247 ( .A(n349), .B(n350), .Q(n342) );
  AOI312 U248 ( .A(n176), .B(n177), .C(n178), .D(n179), .Q(n173) );
  INV6 U249 ( .A(n138), .Q(n131) );
  NAND23 U250 ( .A(B[25]), .B(n224), .Q(n184) );
  INV1 U251 ( .A(B[25]), .Q(n223) );
  NAND28 U252 ( .A(B[18]), .B(n305), .Q(n271) );
  NOR24 U253 ( .A(n143), .B(n144), .Q(n142) );
  AOI311 U254 ( .A(n88), .B(n85), .C(n382), .D(n374), .Q(n384) );
  NAND21 U255 ( .A(n301), .B(n270), .Q(n298) );
  CLKIN6 U256 ( .A(n320), .Q(n49) );
  NOR23 U257 ( .A(n334), .B(n346), .Q(n345) );
  NOR24 U258 ( .A(n379), .B(n49), .Q(n45) );
  NOR24 U259 ( .A(n46), .B(n26), .Q(n48) );
  AOI312 U260 ( .A(n337), .B(n338), .C(n20), .D(n339), .Q(n336) );
  INV0 U261 ( .A(n357), .Q(n47) );
  NOR24 U262 ( .A(A[12]), .B(n326), .Q(n379) );
  XNR22 U263 ( .A(n72), .B(n336), .Q(DIFF[15]) );
  IMUX22 U264 ( .A(n363), .B(n364), .S(n365), .Q(DIFF[12]) );
  NAND24 U265 ( .A(n348), .B(n349), .Q(n343) );
  NAND24 U266 ( .A(n230), .B(n231), .Q(n229) );
  XOR22 U267 ( .A(n196), .B(n197), .Q(DIFF[26]) );
  NOR24 U268 ( .A(n52), .B(n53), .Q(n54) );
  NOR24 U269 ( .A(n54), .B(n78), .Q(n84) );
  INV1 U270 ( .A(n85), .Q(n52) );
  CLKIN3 U271 ( .A(n86), .Q(n53) );
  XOR22 U272 ( .A(n83), .B(n84), .Q(DIFF[9]) );
  INV4 U273 ( .A(n59), .Q(n60) );
  NOR24 U274 ( .A(n60), .B(n377), .Q(n77) );
  INV3 U275 ( .A(A[8]), .Q(n56) );
  NAND34 U276 ( .A(n113), .B(n76), .C(n58), .Q(n138) );
  NOR32 U277 ( .A(n378), .B(n376), .C(n375), .Q(n59) );
  NAND22 U278 ( .A(A[16]), .B(n283), .Q(n276) );
  OAI222 U279 ( .A(B[19]), .B(n274), .C(n282), .D(n275), .Q(n273) );
  INV2 U280 ( .A(n284), .Q(n262) );
  AOI222 U281 ( .A(n397), .B(n398), .C(n399), .D(n400), .Q(n387) );
  INV2 U282 ( .A(n70), .Q(n71) );
  INV2 U283 ( .A(n66), .Q(n68) );
  NAND21 U284 ( .A(n250), .B(n237), .Q(n253) );
  XNR20 U285 ( .A(n158), .B(n117), .Q(DIFF[2]) );
  INV3 U286 ( .A(n184), .Q(n74) );
  NAND22 U287 ( .A(n170), .B(n153), .Q(n169) );
  NOR20 U288 ( .A(n98), .B(n100), .Q(n99) );
  NAND22 U289 ( .A(n256), .B(n239), .Q(n255) );
  INV3 U290 ( .A(n255), .Q(n249) );
  NAND20 U291 ( .A(n297), .B(n271), .Q(n296) );
  OAI2112 U292 ( .A(n74), .B(n181), .C(n182), .D(n183), .Q(n178) );
  NAND20 U293 ( .A(n177), .B(n183), .Q(n196) );
  NAND20 U294 ( .A(B[30]), .B(n128), .Q(n141) );
  NOR22 U295 ( .A(A[5]), .B(n414), .Q(n412) );
  NOR20 U296 ( .A(n92), .B(n78), .Q(n91) );
  IMUX20 U297 ( .A(n266), .B(n267), .S(n268), .Q(DIFF[20]) );
  IMUX20 U298 ( .A(n225), .B(n226), .S(n227), .Q(DIFF[24]) );
  NOR20 U299 ( .A(n308), .B(n301), .Q(n311) );
  XNR22 U300 ( .A(n12), .B(n172), .Q(DIFF[28]) );
  XNR21 U301 ( .A(n81), .B(A[11]), .Q(n64) );
  INV2 U302 ( .A(n329), .Q(n328) );
  CLKIN6 U303 ( .A(n188), .Q(n75) );
  OAI220 U304 ( .A(n147), .B(n148), .C(B[29]), .D(n149), .Q(n146) );
  INV2 U305 ( .A(n185), .Q(n176) );
  NAND22 U306 ( .A(A[22]), .B(n257), .Q(n238) );
  NOR20 U307 ( .A(n69), .B(n242), .Q(n66) );
  INV0 U308 ( .A(n238), .Q(n69) );
  NAND20 U309 ( .A(n237), .B(n238), .Q(n70) );
  XOR21 U310 ( .A(n96), .B(n99), .Q(DIFF[6]) );
  XOR20 U311 ( .A(n286), .B(n160), .Q(DIFF[1]) );
  INV3 U312 ( .A(n147), .Q(n155) );
  NAND21 U313 ( .A(B[28]), .B(n168), .Q(n156) );
  NAND22 U314 ( .A(n213), .B(n219), .Q(n218) );
  NAND20 U315 ( .A(n20), .B(n332), .Q(n344) );
  XNR22 U316 ( .A(n248), .B(n11), .Q(DIFF[23]) );
  NAND20 U317 ( .A(n337), .B(n340), .Q(n353) );
  NAND20 U318 ( .A(n239), .B(n237), .Q(n259) );
  NAND20 U319 ( .A(n242), .B(n238), .Q(n251) );
  NAND22 U320 ( .A(n254), .B(n239), .Q(n250) );
  NAND20 U321 ( .A(n271), .B(n275), .Q(n299) );
  XOR21 U322 ( .A(n299), .B(n300), .Q(DIFF[18]) );
  NAND22 U323 ( .A(n207), .B(n208), .Q(n205) );
  NAND22 U324 ( .A(n150), .B(n123), .Q(n145) );
  INV3 U325 ( .A(n167), .Q(n148) );
  NOR20 U326 ( .A(B[28]), .B(n168), .Q(n167) );
  NAND20 U327 ( .A(n303), .B(n270), .Q(n302) );
  INV3 U328 ( .A(A[13]), .Q(n362) );
  INV3 U329 ( .A(A[9]), .Q(n417) );
  INV3 U330 ( .A(A[2]), .Q(n404) );
  INV3 U331 ( .A(A[25]), .Q(n224) );
  INV3 U332 ( .A(A[21]), .Q(n265) );
  INV3 U333 ( .A(A[22]), .Q(n258) );
  INV3 U334 ( .A(A[5]), .Q(n409) );
  NAND22 U335 ( .A(A[20]), .B(n247), .Q(n236) );
  INV3 U336 ( .A(A[18]), .Q(n305) );
  INV3 U337 ( .A(A[26]), .Q(n200) );
  NOR20 U338 ( .A(A[4]), .B(n110), .Q(n108) );
  NOR21 U339 ( .A(A[29]), .B(n157), .Q(n147) );
  INV3 U340 ( .A(B[29]), .Q(n157) );
  INV3 U341 ( .A(A[14]), .Q(n352) );
  NAND22 U342 ( .A(A[25]), .B(n223), .Q(n182) );
  XOR20 U343 ( .A(B[24]), .B(A[24]), .Q(n226) );
  AOI210 U344 ( .A(B[24]), .B(n222), .C(n206), .Q(n225) );
  NAND22 U345 ( .A(A[26]), .B(n199), .Q(n183) );
  CLKIN0 U346 ( .A(B[26]), .Q(n199) );
  INV3 U347 ( .A(A[6]), .Q(n415) );
  INV3 U348 ( .A(A[17]), .Q(n310) );
  INV3 U349 ( .A(A[10]), .Q(n419) );
  NOR20 U350 ( .A(n47), .B(n335), .Q(n363) );
  IMUX20 U351 ( .A(n111), .B(n112), .S(n107), .Q(DIFF[4]) );
  NOR21 U352 ( .A(n108), .B(n114), .Q(n111) );
  IMUX20 U353 ( .A(n90), .B(n91), .S(n86), .Q(DIFF[8]) );
  NOR20 U354 ( .A(A[8]), .B(n93), .Q(n92) );
  INV3 U355 ( .A(A[29]), .Q(n149) );
  INV3 U356 ( .A(A[23]), .Q(n240) );
  NAND22 U357 ( .A(n421), .B(n288), .Q(n287) );
  INV3 U358 ( .A(A[1]), .Q(n405) );
  NOR21 U359 ( .A(n284), .B(n285), .Q(n266) );
  XOR21 U360 ( .A(n292), .B(n293), .Q(DIFF[19]) );
  XNR20 U361 ( .A(n22), .B(A[15]), .Q(n72) );
  NOR33 U362 ( .A(n195), .B(n74), .C(n75), .Q(n73) );
  INV3 U363 ( .A(n308), .Q(n303) );
  NOR20 U364 ( .A(A[16]), .B(n283), .Q(n308) );
  NAND22 U365 ( .A(n420), .B(n421), .Q(DIFF[0]) );
  NAND20 U366 ( .A(n402), .B(B[0]), .Q(n420) );
  INV6 U367 ( .A(n244), .Q(n230) );
  XOR20 U368 ( .A(B[16]), .B(A[16]), .Q(n312) );
  INV3 U369 ( .A(A[24]), .Q(n222) );
  INV3 U370 ( .A(A[28]), .Q(n168) );
  INV3 U371 ( .A(A[0]), .Q(n402) );
  INV3 U372 ( .A(A[30]), .Q(n128) );
  INV3 U373 ( .A(A[27]), .Q(n180) );
  INV3 U374 ( .A(A[19]), .Q(n274) );
  OAI211 U375 ( .A(n159), .B(n160), .C(n161), .Q(n117) );
  NOR20 U376 ( .A(B[27]), .B(n180), .Q(n179) );
  INV3 U377 ( .A(B[27]), .Q(n186) );
  INV6 U378 ( .A(n162), .Q(n119) );
  NAND24 U379 ( .A(A[5]), .B(n414), .Q(n103) );
  NAND20 U380 ( .A(n103), .B(n105), .Q(n106) );
  NAND20 U381 ( .A(B[13]), .B(n362), .Q(n337) );
  NAND20 U382 ( .A(B[8]), .B(n56), .Q(n85) );
  XOR21 U383 ( .A(n383), .B(n384), .Q(DIFF[10]) );
  NAND22 U384 ( .A(n231), .B(n262), .Q(n261) );
  INV4 U385 ( .A(B[2]), .Q(n396) );
  NAND20 U386 ( .A(n118), .B(n162), .Q(n158) );
  NAND20 U387 ( .A(n88), .B(n89), .Q(n83) );
  XNR20 U388 ( .A(B[3]), .B(A[3]), .Q(n115) );
  NAND20 U389 ( .A(B[9]), .B(n417), .Q(n88) );
  INV0 U390 ( .A(n80), .Q(n81) );
  NAND20 U391 ( .A(n291), .B(n161), .Q(n286) );
  XOR20 U392 ( .A(B[31]), .B(A[31]), .Q(n121) );
  NAND20 U393 ( .A(n373), .B(n371), .Q(n383) );
  BUF2 U394 ( .A(n232), .Q(n82) );
  NAND20 U395 ( .A(n270), .B(n277), .Q(n306) );
  INV6 U396 ( .A(n154), .Q(n139) );
  XOR20 U397 ( .A(B[19]), .B(A[19]), .Q(n293) );
  AOI312 U398 ( .A(n214), .B(n215), .C(n113), .D(n216), .Q(n202) );
  NAND34 U399 ( .A(n245), .B(n239), .C(n242), .Q(n244) );
  XNR20 U400 ( .A(B[7]), .B(A[7]), .Q(n94) );
  INV2 U401 ( .A(n153), .Q(n313) );
  XOR20 U402 ( .A(B[4]), .B(A[4]), .Q(n112) );
  NAND22 U403 ( .A(n152), .B(n153), .Q(n151) );
  XOR20 U404 ( .A(B[20]), .B(A[20]), .Q(n267) );
  NOR21 U405 ( .A(B[0]), .B(n402), .Q(n290) );
  XOR20 U406 ( .A(B[8]), .B(A[8]), .Q(n90) );
  OAI211 U407 ( .A(n134), .B(n135), .C(n7), .Q(n133) );
  NOR21 U408 ( .A(n134), .B(n135), .Q(n212) );
  XOR20 U409 ( .A(n21), .B(A[12]), .Q(n364) );
  OAI212 U410 ( .A(n107), .B(n108), .C(n109), .Q(n104) );
  XOR22 U411 ( .A(n120), .B(n121), .Q(DIFF[31]) );
  AOI2112 U412 ( .A(n122), .B(n123), .C(n124), .D(n125), .Q(n120) );
  OAI222 U413 ( .A(n126), .B(n127), .C(B[30]), .D(n128), .Q(n125) );
  CLKIN3 U414 ( .A(n141), .Q(n126) );
  CLKIN3 U415 ( .A(n146), .Q(n127) );
  CLKIN3 U416 ( .A(n140), .Q(n150) );
  CLKIN3 U417 ( .A(n156), .Q(n171) );
  AOI212 U418 ( .A(n139), .B(n153), .C(n123), .Q(n172) );
  AOI312 U419 ( .A(n177), .B(n184), .C(n193), .D(n194), .Q(n191) );
  OAI212 U420 ( .A(n195), .B(n182), .C(n183), .Q(n194) );
  AOI212 U421 ( .A(n193), .B(n184), .C(n198), .Q(n197) );
  CLKIN3 U422 ( .A(n182), .Q(n198) );
  CLKIN3 U423 ( .A(n204), .Q(n210) );
  OAI2112 U424 ( .A(n235), .B(n236), .C(n237), .D(n238), .Q(n234) );
  CLKIN3 U425 ( .A(n239), .Q(n235) );
  NOR24 U426 ( .A(n284), .B(n246), .Q(n245) );
  NOR24 U427 ( .A(A[23]), .B(n232), .Q(n246) );
  CLKIN3 U428 ( .A(n181), .Q(n206) );
  XOR22 U429 ( .A(n259), .B(n260), .Q(DIFF[21]) );
  AOI212 U430 ( .A(n256), .B(n153), .C(n254), .Q(n260) );
  CLKIN3 U431 ( .A(n263), .Q(n256) );
  NAND24 U432 ( .A(B[21]), .B(n265), .Q(n239) );
  AOI312 U433 ( .A(n270), .B(n271), .C(n272), .D(n273), .Q(n269) );
  AOI212 U434 ( .A(n276), .B(n277), .C(n282), .Q(n272) );
  CLKIN3 U435 ( .A(n236), .Q(n285) );
  CLKIN3 U436 ( .A(n287), .Q(n160) );
  CLKIN3 U437 ( .A(n302), .Q(n294) );
  CLKIN6 U438 ( .A(B[18]), .Q(n304) );
  AOI212 U439 ( .A(n303), .B(n153), .C(n301), .Q(n307) );
  NOR33 U440 ( .A(n315), .B(n131), .C(n316), .Q(n314) );
  OAI222 U441 ( .A(n134), .B(n135), .C(n134), .D(n136), .Q(n316) );
  NOR24 U442 ( .A(n322), .B(n323), .Q(n321) );
  NOR24 U443 ( .A(A[15]), .B(n325), .Q(n322) );
  OAI2112 U444 ( .A(n330), .B(n331), .C(n332), .D(n333), .Q(n327) );
  CLKIN3 U445 ( .A(n276), .Q(n301) );
  CLKIN3 U446 ( .A(n337), .Q(n347) );
  NAND24 U447 ( .A(n324), .B(A[13]), .Q(n340) );
  NOR24 U448 ( .A(n374), .B(n87), .Q(n368) );
  NOR24 U449 ( .A(A[9]), .B(n372), .Q(n378) );
  NOR24 U450 ( .A(A[11]), .B(n367), .Q(n375) );
  OAI212 U451 ( .A(n376), .B(n381), .C(n371), .Q(n380) );
  NAND24 U452 ( .A(A[3]), .B(n392), .Q(n395) );
  OAI212 U453 ( .A(A[3]), .B(n392), .C(n119), .Q(n394) );
  NAND24 U454 ( .A(A[2]), .B(n396), .Q(n162) );
  OAI2112 U455 ( .A(n412), .B(n109), .C(n103), .D(n101), .Q(n411) );
endmodule


module E_alu ( o_data_AluRes, i_data_A, i_data_B, i_con_AluCtrl, i_data_shamt
 );
  output [31:0] o_data_AluRes;
  input [31:0] i_data_A;
  input [31:0] i_data_B;
  input [3:0] i_con_AluCtrl;
  input [4:0] i_data_shamt;
  wire   N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159,
         N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N244, N245, N246,
         N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257,
         N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268,
         N269, N270, N271, N272, N273, N274, N275, N276, n13, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468;

  E_alu_DW01_add_1 add_53 ( .A(i_data_A), .B({n58, i_data_B[30:28], n33, 
        i_data_B[26], n53, n80, n86, n125, n90, i_data_B[20], n82, n122, 
        i_data_B[17], n113, i_data_B[15:12], n102, i_data_B[10:8], n87, 
        i_data_B[6], n51, i_data_B[4:3], n73, i_data_B[1:0]}), .CI(n13), .SUM(
        {N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, 
        N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, 
        N124, N123, N122, N121, N120, N119, N118, N117, N116}) );
  E_alu_DW01_cmp2_1 r65 ( .A(i_data_A), .B({n58, i_data_B[30:28], n33, 
        i_data_B[26], n54, n80, n86, n125, n90, i_data_B[20], n82, n123, 
        i_data_B[17], n113, i_data_B[15:12], n103, i_data_B[10], n95, 
        i_data_B[8], n88, n11, n50, i_data_B[4], n35, n73, i_data_B[1:0]}), 
        .LEQ(n13), .TC(n13), .LT_LE(N276) );
  E_alu_DW_rash_1 r63 ( .A({n58, i_data_B[30:28], n33, i_data_B[26], n54, n80, 
        n86, n125, n90, i_data_B[20], n82, n123, i_data_B[17], n113, n32, n27, 
        n30, n28, n103, n15, n95, i_data_B[8], n88, n29, n50, i_data_B[4], n35, 
        n73, i_data_B[1:0]}), .DATA_TC(n13), .SH(i_data_shamt), .SH_TC(n13), 
        .B({N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, 
        N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, 
        N188, N187, N186, N185, N184, N183, N182, N181, N180}) );
  E_alu_DW01_ash_1 sll_56 ( .A({n58, i_data_B[30:28], n33, i_data_B[26], n54, 
        n80, n86, n125, n90, i_data_B[20], n81, n123, i_data_B[17], n113, n26, 
        i_data_B[14:12], n103, n15, n95, i_data_B[8], n87, i_data_B[6], n50, 
        i_data_B[4:3], n73, i_data_B[1:0]}), .DATA_TC(n13), .SH(i_data_shamt), 
        .SH_TC(n13), .B({N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, 
        N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148}) );
  E_alu_DW01_sub_2 sub_62 ( .A(i_data_A), .B({n58, i_data_B[30:28], n33, 
        i_data_B[26], n54, n80, n86, n125, n90, i_data_B[20], n81, n122, 
        i_data_B[17], n113, i_data_B[15:8], n87, i_data_B[6], n51, 
        i_data_B[4:3], n79, i_data_B[1:0]}), .CI(n13), .DIFF({N275, N274, N273, 
        N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, 
        N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, 
        N248, N247, N246, N245, N244}) );
  BUF8 U2 ( .A(i_data_B[19]), .Q(n81) );
  BUF12 U3 ( .A(i_data_B[19]), .Q(n82) );
  CLKBU15 U4 ( .A(i_data_B[16]), .Q(n113) );
  BUF2 U5 ( .A(i_data_B[13]), .Q(n30) );
  BUF2 U6 ( .A(n125), .Q(n1) );
  INV12 U7 ( .A(n121), .Q(n122) );
  INV15 U8 ( .A(n121), .Q(n123) );
  NAND24 U9 ( .A(n288), .B(n62), .Q(o_data_AluRes[15]) );
  CLKIN6 U10 ( .A(n77), .Q(n2) );
  CLKIN15 U11 ( .A(n76), .Q(n77) );
  OAI211 U12 ( .A(i_data_A[1]), .B(n130), .C(n120), .Q(n164) );
  BUF2 U13 ( .A(i_data_B[26]), .Q(n3) );
  NAND22 U14 ( .A(N178), .B(n7), .Q(n444) );
  CLKBU4 U15 ( .A(i_data_B[14]), .Q(n27) );
  NAND31 U16 ( .A(n75), .B(n144), .C(n290), .Q(n145) );
  NAND33 U17 ( .A(n158), .B(n160), .C(n159), .Q(n38) );
  INV6 U18 ( .A(n14), .Q(n15) );
  NAND22 U19 ( .A(N198), .B(n456), .Q(n311) );
  NAND22 U20 ( .A(n305), .B(n303), .Q(n47) );
  NAND22 U21 ( .A(n161), .B(n39), .Q(o_data_AluRes[0]) );
  NAND31 U22 ( .A(n242), .B(n241), .C(n240), .Q(o_data_AluRes[10]) );
  INV3 U23 ( .A(n67), .Q(n68) );
  NAND42 U24 ( .A(n405), .B(n404), .C(n403), .D(n402), .Q(o_data_AluRes[26])
         );
  CLKIN12 U25 ( .A(n74), .Q(n4) );
  INV10 U26 ( .A(n4), .Q(n5) );
  INV8 U27 ( .A(n4), .Q(n6) );
  INV12 U28 ( .A(n4), .Q(n7) );
  NOR23 U29 ( .A(n146), .B(n75), .Q(n74) );
  NAND24 U30 ( .A(N273), .B(n9), .Q(n438) );
  BUF2 U31 ( .A(i_data_B[12]), .Q(n28) );
  XNR20 U32 ( .A(n1), .B(i_data_A[22]), .Q(n355) );
  IMUX22 U33 ( .A(n442), .B(n441), .S(i_data_B[30]), .Q(n446) );
  NAND22 U34 ( .A(n332), .B(n331), .Q(o_data_AluRes[19]) );
  BUF6 U35 ( .A(n464), .Q(n8) );
  CLKBU12 U36 ( .A(n464), .Q(n9) );
  INV3 U37 ( .A(n145), .Q(n464) );
  CLKIN12 U38 ( .A(n101), .Q(n102) );
  CLKIN12 U39 ( .A(n134), .Q(n133) );
  AOI220 U40 ( .A(N246), .B(n8), .C(N118), .D(n57), .Q(n175) );
  IMUX21 U41 ( .A(n302), .B(n301), .S(n20), .Q(n303) );
  NAND33 U42 ( .A(n217), .B(n216), .C(n214), .Q(n65) );
  INV8 U43 ( .A(n454), .Q(n443) );
  NAND22 U44 ( .A(N202), .B(n456), .Q(n356) );
  NAND23 U45 ( .A(N166), .B(n7), .Q(n310) );
  AOI221 U46 ( .A(N244), .B(n8), .C(N148), .D(n7), .Q(n159) );
  NAND22 U47 ( .A(n100), .B(n434), .Q(n435) );
  NAND42 U48 ( .A(n447), .B(n446), .C(n445), .D(n444), .Q(n448) );
  NAND23 U49 ( .A(n250), .B(n251), .Q(n67) );
  NAND23 U50 ( .A(n342), .B(n341), .Q(n45) );
  NAND22 U51 ( .A(n372), .B(n371), .Q(n373) );
  AOI211 U52 ( .A(N171), .B(n5), .C(n369), .Q(n372) );
  NAND22 U53 ( .A(n276), .B(n277), .Q(n91) );
  AOI211 U54 ( .A(n387), .B(n119), .C(n388), .Q(n392) );
  AOI221 U55 ( .A(i_data_A[3]), .B(n179), .C(N183), .D(n456), .Q(n185) );
  AOI221 U56 ( .A(i_data_A[2]), .B(n171), .C(N182), .D(n456), .Q(n177) );
  AOI221 U57 ( .A(N190), .B(n456), .C(N158), .D(n5), .Q(n241) );
  AOI221 U58 ( .A(i_data_A[17]), .B(n300), .C(i_data_B[1]), .D(n443), .Q(n306)
         );
  NAND22 U59 ( .A(n215), .B(n66), .Q(o_data_AluRes[7]) );
  NAND22 U60 ( .A(n443), .B(n35), .Q(n10) );
  NAND24 U61 ( .A(n10), .B(n323), .Q(n325) );
  INV4 U62 ( .A(i_data_B[3]), .Q(n324) );
  CLKIN4 U63 ( .A(i_data_B[15]), .Q(n31) );
  INV12 U64 ( .A(i_data_B[11]), .Q(n101) );
  INV3 U65 ( .A(n352), .Q(n11) );
  CLKIN4 U66 ( .A(i_data_B[6]), .Q(n352) );
  OAI211 U67 ( .A(n77), .B(n396), .C(i_data_A[26]), .Q(n405) );
  NAND23 U68 ( .A(N138), .B(n56), .Q(n353) );
  NOR32 U69 ( .A(n317), .B(n314), .C(n315), .Q(n63) );
  INV6 U70 ( .A(n101), .Q(n103) );
  NAND22 U71 ( .A(n381), .B(n380), .Q(n382) );
  NAND23 U72 ( .A(N274), .B(n9), .Q(n449) );
  INV6 U73 ( .A(n71), .Q(n72) );
  NAND34 U74 ( .A(n384), .B(n386), .C(n385), .Q(n59) );
  NAND23 U75 ( .A(n376), .B(n375), .Q(o_data_AluRes[23]) );
  NAND23 U76 ( .A(n437), .B(n438), .Q(o_data_AluRes[29]) );
  CLKBU15 U77 ( .A(n76), .Q(n120) );
  BUF6 U78 ( .A(n143), .Q(n55) );
  INV4 U79 ( .A(n55), .Q(n57) );
  INV12 U80 ( .A(n94), .Q(n95) );
  XOR20 U81 ( .A(n123), .B(i_data_A[18]), .Q(n12) );
  NAND23 U82 ( .A(n152), .B(n290), .Q(n458) );
  INV6 U83 ( .A(n458), .Q(n134) );
  CLKIN3 U84 ( .A(n458), .Q(n135) );
  NAND23 U85 ( .A(n363), .B(n362), .Q(o_data_AluRes[22]) );
  BUF15 U86 ( .A(i_data_B[21]), .Q(n90) );
  IMUX21 U87 ( .A(n126), .B(n117), .S(n34), .Q(n261) );
  AOI212 U88 ( .A(i_data_A[14]), .B(n274), .C(n273), .Q(n275) );
  NAND21 U89 ( .A(n269), .B(n119), .Q(n274) );
  IMUX21 U90 ( .A(n272), .B(n271), .S(n27), .Q(n273) );
  NAND22 U91 ( .A(n194), .B(n119), .Q(n195) );
  NAND22 U92 ( .A(n162), .B(n119), .Q(n163) );
  NAND33 U93 ( .A(n393), .B(n394), .C(n395), .Q(o_data_AluRes[25]) );
  NAND22 U94 ( .A(N208), .B(n456), .Q(n425) );
  NOR21 U95 ( .A(i_data_A[17]), .B(n132), .Q(n302) );
  AOI222 U96 ( .A(N257), .B(n9), .C(N129), .D(n56), .Q(n266) );
  NAND23 U97 ( .A(n328), .B(n327), .Q(n329) );
  IMUX21 U98 ( .A(n418), .B(n417), .S(i_data_B[28]), .Q(n419) );
  BUF15 U99 ( .A(i_data_B[27]), .Q(n33) );
  INV6 U100 ( .A(n59), .Q(n60) );
  NAND23 U101 ( .A(N259), .B(n9), .Q(n285) );
  NAND34 U102 ( .A(n298), .B(n297), .C(n295), .Q(n69) );
  NAND42 U103 ( .A(n412), .B(n411), .C(n409), .D(n410), .Q(n413) );
  IMUX22 U104 ( .A(n334), .B(n333), .S(i_data_B[20]), .Q(n342) );
  NAND32 U105 ( .A(n423), .B(n424), .C(n37), .Q(o_data_AluRes[28]) );
  CLKBU15 U106 ( .A(i_data_B[23]), .Q(n86) );
  IMUX20 U107 ( .A(n127), .B(n116), .S(i_data_B[1]), .Q(n162) );
  CLKIN2 U108 ( .A(n31), .Q(n32) );
  OAI220 U109 ( .A(n138), .B(n139), .C(n147), .D(n146), .Q(n141) );
  BUF15 U110 ( .A(i_data_B[7]), .Q(n87) );
  CLKBU4 U111 ( .A(i_data_B[7]), .Q(n88) );
  NAND22 U112 ( .A(N134), .B(n57), .Q(n309) );
  INV6 U113 ( .A(i_data_B[25]), .Q(n52) );
  CLKIN6 U114 ( .A(i_data_B[10]), .Q(n14) );
  CLKIN6 U115 ( .A(i_data_B[2]), .Q(n78) );
  NOR21 U116 ( .A(i_data_A[16]), .B(n132), .Q(n294) );
  OAI212 U117 ( .A(n454), .B(n308), .C(n307), .Q(n317) );
  CLKIN6 U118 ( .A(n65), .Q(n66) );
  NOR33 U119 ( .A(n106), .B(n359), .C(n360), .Q(n363) );
  INV6 U120 ( .A(n105), .Q(n106) );
  INV6 U121 ( .A(n49), .Q(n50) );
  INV10 U122 ( .A(i_data_B[5]), .Q(n49) );
  NAND24 U123 ( .A(n41), .B(n40), .Q(n42) );
  NAND23 U124 ( .A(n212), .B(n88), .Q(n41) );
  INV6 U125 ( .A(n47), .Q(n48) );
  NAND23 U126 ( .A(N147), .B(n57), .Q(n466) );
  BUF2 U127 ( .A(i_data_B[8]), .Q(n16) );
  OAI212 U128 ( .A(i_data_A[16]), .B(n130), .C(n120), .Q(n293) );
  OAI211 U129 ( .A(n77), .B(n335), .C(i_data_A[20]), .Q(n341) );
  AOI210 U130 ( .A(n127), .B(n364), .C(n77), .Q(n365) );
  NAND23 U131 ( .A(n148), .B(n147), .Q(n136) );
  IMUX21 U132 ( .A(n127), .B(n116), .S(n29), .Q(n202) );
  NAND41 U133 ( .A(n193), .B(n192), .C(n191), .D(n190), .Q(o_data_AluRes[4])
         );
  INV4 U134 ( .A(n149), .Q(n152) );
  BUF2 U135 ( .A(i_data_B[4]), .Q(n17) );
  NAND24 U136 ( .A(n23), .B(n120), .Q(n407) );
  IMUX20 U137 ( .A(n127), .B(n116), .S(n17), .Q(n186) );
  INV12 U138 ( .A(n52), .Q(n54) );
  CLKIN8 U139 ( .A(n52), .Q(n53) );
  CLKIN6 U140 ( .A(n61), .Q(n62) );
  NAND31 U141 ( .A(n18), .B(n420), .C(i_data_A[22]), .Q(n19) );
  NAND24 U142 ( .A(n19), .B(n356), .Q(n358) );
  INV3 U143 ( .A(n357), .Q(n18) );
  NOR24 U144 ( .A(n361), .B(n358), .Q(n105) );
  BUF2 U145 ( .A(i_data_B[17]), .Q(n20) );
  NAND22 U146 ( .A(n21), .B(n22), .Q(n23) );
  INV3 U147 ( .A(i_data_A[27]), .Q(n21) );
  INV2 U148 ( .A(n129), .Q(n22) );
  BUF12 U149 ( .A(n451), .Q(n129) );
  INV6 U150 ( .A(n78), .Q(n79) );
  BUF15 U151 ( .A(n451), .Q(n128) );
  BUF15 U152 ( .A(n420), .Q(n117) );
  NAND24 U153 ( .A(n465), .B(n112), .Q(o_data_AluRes[31]) );
  CLKIN0 U154 ( .A(n1), .Q(n357) );
  NAND21 U155 ( .A(n421), .B(n2), .Q(n422) );
  OAI210 U156 ( .A(i_data_A[12]), .B(n130), .C(n119), .Q(n255) );
  OAI210 U157 ( .A(i_data_A[9]), .B(n130), .C(n120), .Q(n228) );
  OAI210 U158 ( .A(i_data_A[13]), .B(n130), .C(n2), .Q(n263) );
  NAND21 U159 ( .A(n343), .B(n119), .Q(n344) );
  OAI210 U160 ( .A(i_data_A[26]), .B(n129), .C(n120), .Q(n397) );
  OAI210 U161 ( .A(i_data_A[6]), .B(n131), .C(n119), .Q(n204) );
  NAND23 U162 ( .A(n25), .B(n310), .Q(n315) );
  NAND24 U163 ( .A(n109), .B(n353), .Q(n360) );
  NAND22 U164 ( .A(n12), .B(n24), .Q(n25) );
  INV2 U165 ( .A(n130), .Q(n24) );
  INV6 U166 ( .A(n69), .Q(n70) );
  NAND23 U167 ( .A(N199), .B(n456), .Q(n323) );
  AOI222 U168 ( .A(N265), .B(n9), .C(N137), .D(n56), .Q(n348) );
  OAI211 U169 ( .A(n77), .B(n326), .C(i_data_A[19]), .Q(n327) );
  OAI211 U170 ( .A(n77), .B(n370), .C(i_data_A[23]), .Q(n371) );
  OAI211 U171 ( .A(n77), .B(n379), .C(i_data_A[24]), .Q(n385) );
  OAI211 U172 ( .A(n77), .B(n439), .C(i_data_A[30]), .Q(n447) );
  OAI211 U173 ( .A(n77), .B(n406), .C(i_data_A[27]), .Q(n412) );
  AOI210 U174 ( .A(n127), .B(n320), .C(n77), .Q(n321) );
  OAI211 U175 ( .A(n1), .B(i_data_A[22]), .C(n77), .Q(n351) );
  INV4 U176 ( .A(n31), .Q(n26) );
  AOI212 U177 ( .A(n430), .B(n115), .C(n429), .Q(n436) );
  AOI221 U178 ( .A(N201), .B(n456), .C(N169), .D(n5), .Q(n349) );
  NAND24 U179 ( .A(n152), .B(n85), .Q(n451) );
  AOI221 U180 ( .A(n27), .B(n443), .C(N210), .D(n456), .Q(n445) );
  CLKIN6 U181 ( .A(n352), .Q(n29) );
  CLKIN6 U182 ( .A(i_data_B[9]), .Q(n94) );
  INV15 U183 ( .A(n85), .Q(n290) );
  NAND23 U184 ( .A(n337), .B(n336), .Q(n338) );
  INV1 U185 ( .A(n132), .Q(n108) );
  NAND23 U186 ( .A(N255), .B(n9), .Q(n249) );
  INV4 U187 ( .A(n63), .Q(n64) );
  NAND33 U188 ( .A(n348), .B(n350), .C(n44), .Q(o_data_AluRes[21]) );
  OAI211 U189 ( .A(i_data_A[8]), .B(n131), .C(n119), .Q(n220) );
  OAI211 U190 ( .A(i_data_A[5]), .B(n131), .C(n120), .Q(n196) );
  OAI211 U191 ( .A(i_data_A[4]), .B(n131), .C(n120), .Q(n188) );
  OAI211 U192 ( .A(i_data_A[2]), .B(n131), .C(n120), .Q(n172) );
  INV15 U193 ( .A(n128), .Q(n126) );
  INV15 U194 ( .A(n118), .Q(n76) );
  IMUX24 U195 ( .A(n282), .B(n281), .S(n114), .Q(n283) );
  AOI221 U196 ( .A(N249), .B(n8), .C(N121), .D(n56), .Q(n199) );
  AOI222 U197 ( .A(i_data_A[5]), .B(n195), .C(N185), .D(n456), .Q(n201) );
  CLKBU12 U198 ( .A(n461), .Q(n115) );
  NAND24 U199 ( .A(n291), .B(n150), .Q(n461) );
  NAND21 U200 ( .A(n299), .B(n119), .Q(n300) );
  NAND33 U201 ( .A(n306), .B(n304), .C(n48), .Q(o_data_AluRes[17]) );
  AOI221 U202 ( .A(i_data_A[21]), .B(n344), .C(n50), .D(n443), .Q(n350) );
  NAND22 U203 ( .A(n339), .B(n72), .Q(o_data_AluRes[20]) );
  INV6 U204 ( .A(i_con_AluCtrl[2]), .Q(n147) );
  INV6 U205 ( .A(n137), .Q(n144) );
  AOI222 U206 ( .A(N200), .B(n456), .C(n17), .D(n443), .Q(n337) );
  AOI211 U207 ( .A(n127), .B(n388), .C(n77), .Q(n389) );
  AOI211 U208 ( .A(n127), .B(n235), .C(n77), .Q(n236) );
  IMUX22 U209 ( .A(n246), .B(n245), .S(n103), .Q(n247) );
  NAND21 U210 ( .A(N155), .B(n6), .Q(n216) );
  INV6 U211 ( .A(n42), .Q(n214) );
  OAI212 U212 ( .A(n454), .B(n432), .C(n431), .Q(n433) );
  CLKIN15 U213 ( .A(n49), .Q(n51) );
  IMUX22 U214 ( .A(n294), .B(n293), .S(n113), .Q(n295) );
  INV6 U215 ( .A(i_con_AluCtrl[1]), .Q(n148) );
  IMUX22 U216 ( .A(n155), .B(n154), .S(n104), .Q(n156) );
  AOI212 U217 ( .A(n126), .B(n153), .C(n77), .Q(n154) );
  AOI212 U218 ( .A(n127), .B(n244), .C(n77), .Q(n245) );
  NAND22 U219 ( .A(n400), .B(n399), .Q(n401) );
  INV1 U220 ( .A(n132), .Q(n99) );
  IMUX21 U221 ( .A(n366), .B(n365), .S(n86), .Q(n374) );
  AOI222 U222 ( .A(N130), .B(n56), .C(N194), .D(n456), .Q(n278) );
  CLKIN4 U223 ( .A(n147), .Q(n75) );
  BUF12 U224 ( .A(n440), .Q(n118) );
  AOI212 U225 ( .A(i_data_A[11]), .B(n248), .C(n247), .Q(n250) );
  CLKIN15 U226 ( .A(n124), .Q(n125) );
  CLKIN12 U227 ( .A(n83), .Q(n84) );
  AOI212 U228 ( .A(i_data_A[15]), .B(n284), .C(n283), .Q(n286) );
  AOI222 U229 ( .A(i_data_A[16]), .B(n292), .C(n104), .D(n443), .Q(n298) );
  BUF15 U230 ( .A(n76), .Q(n119) );
  NAND22 U231 ( .A(n210), .B(n119), .Q(n211) );
  NAND22 U232 ( .A(n226), .B(n119), .Q(n227) );
  NAND22 U233 ( .A(n186), .B(n119), .Q(n187) );
  NAND22 U234 ( .A(n261), .B(n119), .Q(n262) );
  IMUX22 U235 ( .A(n119), .B(n133), .S(n457), .Q(n463) );
  BUF15 U236 ( .A(i_data_B[2]), .Q(n73) );
  IMUX20 U237 ( .A(n127), .B(n116), .S(n50), .Q(n194) );
  NAND23 U238 ( .A(N266), .B(n9), .Q(n362) );
  BUF12 U239 ( .A(i_data_B[31]), .Q(n58) );
  XNR21 U240 ( .A(n58), .B(i_data_A[31]), .Q(n452) );
  BUF15 U241 ( .A(i_data_B[24]), .Q(n80) );
  INV15 U242 ( .A(n128), .Q(n127) );
  NOR21 U243 ( .A(i_data_A[20]), .B(n132), .Q(n334) );
  IMUX21 U244 ( .A(n129), .B(n115), .S(i_data_B[30]), .Q(n439) );
  BUF4 U245 ( .A(n451), .Q(n131) );
  CLKIN4 U246 ( .A(n43), .Q(n44) );
  BUF2 U247 ( .A(n30), .Q(n34) );
  OAI211 U248 ( .A(i_data_A[17]), .B(n130), .C(n120), .Q(n301) );
  NOR22 U249 ( .A(i_data_A[7]), .B(n133), .Q(n213) );
  NAND23 U250 ( .A(N270), .B(n9), .Q(n402) );
  CLKIN12 U251 ( .A(n324), .Q(n35) );
  NAND21 U252 ( .A(N159), .B(n7), .Q(n251) );
  AOI221 U253 ( .A(N197), .B(n456), .C(N165), .D(n6), .Q(n305) );
  NAND34 U254 ( .A(n285), .B(n286), .C(n287), .Q(n61) );
  OAI211 U255 ( .A(n123), .B(i_data_A[18]), .C(n77), .Q(n307) );
  NAND23 U256 ( .A(N271), .B(n9), .Q(n415) );
  NAND22 U257 ( .A(n426), .B(n425), .Q(n36) );
  INV3 U258 ( .A(n36), .Q(n37) );
  INV6 U259 ( .A(n38), .Q(n39) );
  AOI222 U260 ( .A(N180), .B(n456), .C(N116), .D(n57), .Q(n160) );
  AOI212 U261 ( .A(i_data_A[0]), .B(n157), .C(n156), .Q(n158) );
  NAND22 U262 ( .A(n213), .B(n368), .Q(n40) );
  NAND22 U263 ( .A(n349), .B(n347), .Q(n43) );
  NAND24 U264 ( .A(n340), .B(n46), .Q(n71) );
  CLKIN6 U265 ( .A(n45), .Q(n46) );
  NAND23 U266 ( .A(N262), .B(n9), .Q(n318) );
  NAND43 U267 ( .A(n233), .B(n232), .C(n230), .D(n231), .Q(o_data_AluRes[9])
         );
  AOI222 U268 ( .A(N253), .B(n9), .C(N125), .D(n57), .Q(n231) );
  NOR24 U269 ( .A(n64), .B(n316), .Q(n319) );
  OAI312 U270 ( .A(i_data_A[18]), .B(n123), .C(n132), .D(n309), .Q(n316) );
  AOI222 U271 ( .A(i_data_A[7]), .B(n211), .C(N187), .D(n456), .Q(n217) );
  AOI222 U272 ( .A(N175), .B(n6), .C(n103), .D(n443), .Q(n410) );
  CLKIN15 U273 ( .A(n142), .Q(n456) );
  NAND32 U274 ( .A(n75), .B(n148), .C(n150), .Q(n142) );
  IMUX21 U275 ( .A(n378), .B(n377), .S(n80), .Q(n386) );
  OAI211 U276 ( .A(i_data_A[24]), .B(n129), .C(n120), .Q(n377) );
  IMUX21 U277 ( .A(n127), .B(n116), .S(n88), .Q(n210) );
  IMUX20 U278 ( .A(n205), .B(n204), .S(n29), .Q(n206) );
  IMUX20 U279 ( .A(n126), .B(n117), .S(n20), .Q(n299) );
  INV12 U280 ( .A(i_data_B[18]), .Q(n121) );
  AOI222 U281 ( .A(N196), .B(n456), .C(N164), .D(n6), .Q(n297) );
  INV0 U282 ( .A(n88), .Q(n368) );
  AOI221 U283 ( .A(N176), .B(n5), .C(n110), .D(n443), .Q(n426) );
  INV6 U284 ( .A(n55), .Q(n56) );
  NAND33 U285 ( .A(n278), .B(n275), .C(n92), .Q(o_data_AluRes[14]) );
  NOR41 U286 ( .A(n84), .B(i_con_AluCtrl[2]), .C(n93), .D(n290), .Q(n440) );
  NAND22 U287 ( .A(n383), .B(n60), .Q(o_data_AluRes[24]) );
  AOI212 U288 ( .A(N140), .B(n56), .C(n382), .Q(n384) );
  AOI222 U289 ( .A(N256), .B(n9), .C(N128), .D(n56), .Q(n258) );
  NAND23 U290 ( .A(n319), .B(n318), .Q(o_data_AluRes[18]) );
  AOI221 U291 ( .A(N251), .B(n9), .C(N123), .D(n57), .Q(n215) );
  NAND32 U292 ( .A(n252), .B(n249), .C(n68), .Q(o_data_AluRes[11]) );
  AOI221 U293 ( .A(N127), .B(n56), .C(N191), .D(n456), .Q(n252) );
  NAND22 U294 ( .A(N268), .B(n9), .Q(n383) );
  AOI212 U295 ( .A(N136), .B(n56), .C(n338), .Q(n340) );
  NAND22 U296 ( .A(N264), .B(n9), .Q(n339) );
  NAND23 U297 ( .A(n296), .B(n70), .Q(o_data_AluRes[16]) );
  NAND23 U298 ( .A(N267), .B(n9), .Q(n375) );
  AOI2111 U299 ( .A(N126), .B(n56), .C(n239), .D(n238), .Q(n242) );
  AOI221 U300 ( .A(N174), .B(n6), .C(n89), .D(n443), .Q(n400) );
  NAND41 U301 ( .A(n185), .B(n184), .C(n183), .D(n182), .Q(o_data_AluRes[3])
         );
  NAND22 U302 ( .A(N170), .B(n5), .Q(n354) );
  OAI312 U303 ( .A(n313), .B(n461), .C(n312), .D(n311), .Q(n314) );
  NAND22 U304 ( .A(N206), .B(n456), .Q(n399) );
  AOI222 U305 ( .A(N131), .B(n56), .C(N195), .D(n456), .Q(n288) );
  NAND23 U306 ( .A(N275), .B(n9), .Q(n465) );
  NAND21 U307 ( .A(n170), .B(n119), .Q(n171) );
  NAND21 U308 ( .A(N162), .B(n6), .Q(n277) );
  NAND22 U309 ( .A(N258), .B(n9), .Q(n276) );
  AOI212 U310 ( .A(N144), .B(n57), .C(n419), .Q(n424) );
  NAND42 U311 ( .A(n225), .B(n224), .C(n223), .D(n222), .Q(o_data_AluRes[8])
         );
  NAND42 U312 ( .A(n260), .B(n259), .C(n258), .D(n257), .Q(o_data_AluRes[12])
         );
  NAND20 U313 ( .A(n135), .B(n235), .Q(n237) );
  NAND42 U314 ( .A(n209), .B(n208), .C(n207), .D(n206), .Q(o_data_AluRes[6])
         );
  NAND42 U315 ( .A(n268), .B(n267), .C(n266), .D(n265), .Q(o_data_AluRes[13])
         );
  NOR20 U316 ( .A(i_data_A[5]), .B(n133), .Q(n197) );
  NOR21 U317 ( .A(i_data_A[30]), .B(n132), .Q(n442) );
  IMUX21 U318 ( .A(n126), .B(n117), .S(n114), .Q(n279) );
  IMUX20 U319 ( .A(n129), .B(n115), .S(n80), .Q(n379) );
  NAND22 U320 ( .A(n289), .B(n2), .Q(n292) );
  IMUX21 U321 ( .A(n126), .B(n117), .S(n113), .Q(n289) );
  BUF6 U322 ( .A(n451), .Q(n130) );
  AOI221 U323 ( .A(N245), .B(n8), .C(N117), .D(n56), .Q(n167) );
  AOI221 U324 ( .A(N247), .B(n8), .C(N119), .D(n56), .Q(n183) );
  AOI221 U325 ( .A(N252), .B(n9), .C(N124), .D(n57), .Q(n223) );
  AOI221 U326 ( .A(N248), .B(n8), .C(N120), .D(n56), .Q(n191) );
  NAND41 U327 ( .A(n177), .B(n176), .C(n175), .D(n174), .Q(o_data_AluRes[2])
         );
  NOR31 U328 ( .A(n452), .B(n460), .C(n139), .Q(n140) );
  NOR31 U329 ( .A(n115), .B(n460), .C(n459), .Q(n462) );
  NAND22 U330 ( .A(N209), .B(n456), .Q(n431) );
  IMUX20 U331 ( .A(n126), .B(n117), .S(n27), .Q(n269) );
  IMUX20 U332 ( .A(n128), .B(n115), .S(n3), .Q(n396) );
  IMUX21 U333 ( .A(n128), .B(n115), .S(n33), .Q(n406) );
  NOR20 U334 ( .A(i_data_A[24]), .B(n132), .Q(n378) );
  NOR20 U335 ( .A(i_data_A[3]), .B(n133), .Q(n181) );
  NOR20 U336 ( .A(i_data_A[8]), .B(n133), .Q(n221) );
  NOR20 U337 ( .A(i_data_A[12]), .B(n133), .Q(n256) );
  IMUX21 U338 ( .A(n398), .B(n397), .S(n3), .Q(n404) );
  NOR20 U339 ( .A(i_data_A[4]), .B(n133), .Q(n189) );
  NOR20 U340 ( .A(i_data_A[9]), .B(n133), .Q(n229) );
  NOR20 U341 ( .A(i_data_A[26]), .B(n132), .Q(n398) );
  NOR20 U342 ( .A(i_data_A[13]), .B(n132), .Q(n264) );
  NOR20 U343 ( .A(i_data_A[21]), .B(n132), .Q(n346) );
  NOR20 U344 ( .A(i_data_A[6]), .B(n133), .Q(n205) );
  IMUX20 U345 ( .A(n126), .B(n117), .S(i_data_B[28]), .Q(n421) );
  NOR20 U346 ( .A(i_data_A[1]), .B(n132), .Q(n165) );
  NOR21 U347 ( .A(i_data_A[27]), .B(n132), .Q(n408) );
  NOR20 U348 ( .A(i_data_A[2]), .B(n133), .Q(n173) );
  CLKIN3 U349 ( .A(n91), .Q(n92) );
  AOI211 U350 ( .A(n127), .B(n416), .C(n77), .Q(n417) );
  IMUX20 U351 ( .A(n129), .B(n461), .S(n86), .Q(n370) );
  LOGIC0 U352 ( .Q(n13) );
  IMUX22 U353 ( .A(n408), .B(n407), .S(n33), .Q(n411) );
  INV6 U354 ( .A(n148), .Q(n93) );
  AOI2112 U355 ( .A(N179), .B(n7), .C(n463), .D(n462), .Q(n467) );
  CLKIN6 U356 ( .A(i_con_AluCtrl[3]), .Q(n83) );
  BUF15 U357 ( .A(i_con_AluCtrl[0]), .Q(n85) );
  NAND30 U358 ( .A(n291), .B(n85), .C(n84), .Q(n139) );
  IMUX20 U359 ( .A(n197), .B(n196), .S(n50), .Q(n198) );
  NAND41 U360 ( .A(n201), .B(n200), .C(n199), .D(n198), .Q(o_data_AluRes[5])
         );
  BUF2 U361 ( .A(n15), .Q(n89) );
  IMUX20 U362 ( .A(n264), .B(n263), .S(n34), .Q(n265) );
  CLKIN0 U363 ( .A(n34), .Q(n432) );
  IMUX21 U364 ( .A(n126), .B(n117), .S(n103), .Q(n243) );
  IMUX20 U365 ( .A(n173), .B(n172), .S(n73), .Q(n174) );
  CLKIN0 U366 ( .A(n73), .Q(n308) );
  IMUX21 U367 ( .A(n127), .B(n116), .S(n35), .Q(n178) );
  IMUX21 U368 ( .A(n181), .B(n180), .S(n35), .Q(n182) );
  IMUX20 U369 ( .A(n221), .B(n220), .S(n16), .Q(n222) );
  IMUX20 U370 ( .A(n165), .B(n164), .S(i_data_B[1]), .Q(n166) );
  NAND41 U371 ( .A(n169), .B(n168), .C(n167), .D(n166), .Q(o_data_AluRes[1])
         );
  CLKIN0 U372 ( .A(n58), .Q(n459) );
  NOR20 U373 ( .A(n58), .B(i_data_A[31]), .Q(n457) );
  IMUX21 U374 ( .A(n237), .B(n236), .S(n89), .Q(n238) );
  IMUX21 U375 ( .A(n126), .B(n116), .S(n89), .Q(n234) );
  AOI211 U376 ( .A(n234), .B(n119), .C(n235), .Q(n239) );
  BUF2 U377 ( .A(n95), .Q(n96) );
  AOI212 U378 ( .A(N276), .B(n141), .C(n140), .Q(n161) );
  INV6 U379 ( .A(n111), .Q(n112) );
  INV6 U380 ( .A(i_data_B[22]), .Q(n124) );
  NAND34 U381 ( .A(n466), .B(n467), .C(n468), .Q(n111) );
  AOI211 U382 ( .A(N211), .B(n456), .C(n455), .Q(n468) );
  IMUX21 U383 ( .A(n322), .B(n321), .S(n82), .Q(n330) );
  IMUX21 U384 ( .A(n130), .B(n461), .S(n82), .Q(n326) );
  NAND31 U385 ( .A(n97), .B(n98), .C(n99), .Q(n100) );
  INV3 U386 ( .A(i_data_A[29]), .Q(n97) );
  INV0 U387 ( .A(i_data_B[29]), .Q(n98) );
  CLKIN15 U388 ( .A(n134), .Q(n132) );
  INV6 U389 ( .A(n84), .Q(n150) );
  AOI211 U390 ( .A(n127), .B(n270), .C(n77), .Q(n271) );
  IMUX21 U391 ( .A(n127), .B(n116), .S(n73), .Q(n170) );
  IMUX21 U392 ( .A(n346), .B(n345), .S(n90), .Q(n347) );
  IMUX21 U393 ( .A(n126), .B(n117), .S(n90), .Q(n343) );
  AOI221 U394 ( .A(N204), .B(n456), .C(n16), .D(n443), .Q(n381) );
  NAND31 U395 ( .A(n84), .B(i_con_AluCtrl[2]), .C(n148), .Q(n149) );
  IMUX20 U396 ( .A(n189), .B(n188), .S(n17), .Q(n190) );
  INV6 U397 ( .A(n136), .Q(n291) );
  BUF2 U398 ( .A(i_data_B[0]), .Q(n104) );
  NAND31 U399 ( .A(n107), .B(n357), .C(n108), .Q(n109) );
  INV3 U400 ( .A(i_data_A[22]), .Q(n107) );
  BUF2 U401 ( .A(n28), .Q(n110) );
  NAND31 U402 ( .A(n144), .B(n147), .C(n290), .Q(n143) );
  IMUX21 U403 ( .A(n390), .B(n389), .S(n54), .Q(n391) );
  IMUX21 U404 ( .A(n126), .B(n117), .S(n54), .Q(n387) );
  AOI220 U405 ( .A(n96), .B(n443), .C(N205), .D(n456), .Q(n394) );
  IMUX21 U406 ( .A(n229), .B(n228), .S(n96), .Q(n230) );
  IMUX21 U407 ( .A(n126), .B(n116), .S(n96), .Q(n226) );
  IMUX21 U408 ( .A(n129), .B(n115), .S(i_data_B[20]), .Q(n335) );
  BUF2 U409 ( .A(n32), .Q(n114) );
  IMUX21 U410 ( .A(n126), .B(n116), .S(n104), .Q(n151) );
  IMUX21 U411 ( .A(n127), .B(n116), .S(n16), .Q(n218) );
  IMUX21 U412 ( .A(n256), .B(n255), .S(n110), .Q(n257) );
  IMUX21 U413 ( .A(n126), .B(n117), .S(n110), .Q(n253) );
  CLKBU15 U414 ( .A(n420), .Q(n116) );
  INV6 U415 ( .A(n461), .Q(n420) );
  CLKIN3 U416 ( .A(n452), .Q(n138) );
  NAND22 U417 ( .A(n93), .B(n150), .Q(n137) );
  NAND22 U418 ( .A(n85), .B(n144), .Q(n146) );
  CLKIN3 U419 ( .A(i_data_A[31]), .Q(n460) );
  NAND22 U420 ( .A(n151), .B(n119), .Q(n157) );
  CLKIN3 U421 ( .A(i_data_A[0]), .Q(n153) );
  NAND22 U422 ( .A(n135), .B(n153), .Q(n155) );
  AOI222 U423 ( .A(i_data_A[1]), .B(n163), .C(N181), .D(n456), .Q(n169) );
  NAND22 U424 ( .A(N149), .B(n7), .Q(n168) );
  NAND22 U425 ( .A(N150), .B(n5), .Q(n176) );
  NAND22 U426 ( .A(n178), .B(n119), .Q(n179) );
  NAND22 U427 ( .A(N151), .B(n5), .Q(n184) );
  OAI212 U428 ( .A(i_data_A[3]), .B(n131), .C(n119), .Q(n180) );
  AOI222 U429 ( .A(i_data_A[4]), .B(n187), .C(N184), .D(n456), .Q(n193) );
  NAND22 U430 ( .A(N152), .B(n6), .Q(n192) );
  NAND22 U431 ( .A(N153), .B(n7), .Q(n200) );
  NAND22 U432 ( .A(n202), .B(n119), .Q(n203) );
  AOI222 U433 ( .A(i_data_A[6]), .B(n203), .C(N186), .D(n456), .Q(n209) );
  NAND22 U434 ( .A(N154), .B(n7), .Q(n208) );
  AOI222 U435 ( .A(N250), .B(n9), .C(N122), .D(n56), .Q(n207) );
  OAI212 U436 ( .A(i_data_A[7]), .B(n131), .C(n120), .Q(n212) );
  NAND22 U437 ( .A(n218), .B(n119), .Q(n219) );
  AOI222 U438 ( .A(i_data_A[8]), .B(n219), .C(N188), .D(n456), .Q(n225) );
  NAND22 U439 ( .A(N156), .B(n6), .Q(n224) );
  AOI222 U440 ( .A(i_data_A[9]), .B(n227), .C(N189), .D(n456), .Q(n233) );
  NAND22 U441 ( .A(N157), .B(n6), .Q(n232) );
  CLKIN3 U442 ( .A(i_data_A[10]), .Q(n235) );
  NAND22 U443 ( .A(N254), .B(n9), .Q(n240) );
  NAND22 U444 ( .A(n243), .B(n119), .Q(n248) );
  CLKIN3 U445 ( .A(i_data_A[11]), .Q(n244) );
  NAND22 U446 ( .A(n135), .B(n244), .Q(n246) );
  NAND22 U447 ( .A(n253), .B(n119), .Q(n254) );
  AOI222 U448 ( .A(i_data_A[12]), .B(n254), .C(N192), .D(n456), .Q(n260) );
  NAND22 U449 ( .A(N160), .B(n5), .Q(n259) );
  AOI222 U450 ( .A(i_data_A[13]), .B(n262), .C(N193), .D(n456), .Q(n268) );
  NAND22 U451 ( .A(N161), .B(n6), .Q(n267) );
  CLKIN3 U452 ( .A(i_data_A[14]), .Q(n270) );
  NAND22 U453 ( .A(n134), .B(n270), .Q(n272) );
  NAND22 U454 ( .A(N163), .B(n7), .Q(n287) );
  NAND22 U455 ( .A(n279), .B(n119), .Q(n284) );
  CLKIN3 U456 ( .A(i_data_A[15]), .Q(n280) );
  NAND22 U457 ( .A(n134), .B(n280), .Q(n282) );
  AOI212 U458 ( .A(n127), .B(n280), .C(n77), .Q(n281) );
  NAND33 U459 ( .A(n291), .B(n84), .C(n290), .Q(n454) );
  AOI222 U460 ( .A(N260), .B(n9), .C(N132), .D(n56), .Q(n296) );
  AOI222 U461 ( .A(N261), .B(n9), .C(N133), .D(n56), .Q(n304) );
  CLKIN3 U462 ( .A(n123), .Q(n313) );
  CLKIN3 U463 ( .A(i_data_A[18]), .Q(n312) );
  CLKIN3 U464 ( .A(i_data_A[19]), .Q(n320) );
  NAND22 U465 ( .A(n134), .B(n320), .Q(n322) );
  AOI212 U466 ( .A(N167), .B(n5), .C(n325), .Q(n328) );
  AOI2112 U467 ( .A(N135), .B(n57), .C(n330), .D(n329), .Q(n332) );
  NAND22 U468 ( .A(N263), .B(n9), .Q(n331) );
  OAI212 U469 ( .A(i_data_A[20]), .B(n129), .C(n120), .Q(n333) );
  NAND22 U470 ( .A(N168), .B(n5), .Q(n336) );
  OAI212 U471 ( .A(i_data_A[21]), .B(n129), .C(n120), .Q(n345) );
  OAI212 U472 ( .A(n454), .B(n352), .C(n351), .Q(n361) );
  OAI212 U473 ( .A(n355), .B(n129), .C(n354), .Q(n359) );
  CLKIN3 U474 ( .A(i_data_A[23]), .Q(n364) );
  NAND22 U475 ( .A(n135), .B(n364), .Q(n366) );
  NAND22 U476 ( .A(N203), .B(n456), .Q(n367) );
  OAI212 U477 ( .A(n454), .B(n368), .C(n367), .Q(n369) );
  AOI2112 U478 ( .A(N139), .B(n56), .C(n374), .D(n373), .Q(n376) );
  NAND22 U479 ( .A(N172), .B(n5), .Q(n380) );
  CLKIN3 U480 ( .A(i_data_A[25]), .Q(n388) );
  NAND22 U481 ( .A(n135), .B(n388), .Q(n390) );
  AOI2112 U482 ( .A(N173), .B(n7), .C(n392), .D(n391), .Q(n395) );
  AOI222 U483 ( .A(N141), .B(n57), .C(N269), .D(n9), .Q(n393) );
  AOI212 U484 ( .A(N142), .B(n57), .C(n401), .Q(n403) );
  NAND22 U485 ( .A(N207), .B(n456), .Q(n409) );
  AOI212 U486 ( .A(N143), .B(n56), .C(n413), .Q(n414) );
  NAND22 U487 ( .A(n415), .B(n414), .Q(o_data_AluRes[27]) );
  CLKIN3 U488 ( .A(i_data_A[28]), .Q(n416) );
  NAND22 U489 ( .A(n135), .B(n416), .Q(n418) );
  AOI222 U490 ( .A(n9), .B(N272), .C(i_data_A[28]), .D(n422), .Q(n423) );
  NAND22 U491 ( .A(i_data_A[29]), .B(i_data_B[29]), .Q(n427) );
  CLKIN3 U492 ( .A(n427), .Q(n430) );
  NAND22 U493 ( .A(n2), .B(n130), .Q(n428) );
  OAI222 U494 ( .A(i_data_A[29]), .B(i_data_B[29]), .C(n430), .D(n428), .Q(
        n429) );
  AOI212 U495 ( .A(N177), .B(n6), .C(n433), .Q(n434) );
  AOI2112 U496 ( .A(N145), .B(n56), .C(n435), .D(n436), .Q(n437) );
  OAI212 U497 ( .A(i_data_A[30]), .B(n129), .C(n120), .Q(n441) );
  AOI212 U498 ( .A(N146), .B(n57), .C(n448), .Q(n450) );
  NAND22 U499 ( .A(n450), .B(n449), .Q(o_data_AluRes[30]) );
  CLKIN3 U500 ( .A(n114), .Q(n453) );
  OAI222 U501 ( .A(n454), .B(n453), .C(n452), .D(n130), .Q(n455) );
endmodule


module E_alu_control ( o_con_AluCtrl, i_con_AluOp, i_con_FuncCode );
  output [3:0] o_con_AluCtrl;
  input [5:0] i_con_AluOp;
  input [5:0] i_con_FuncCode;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59;

  INV3 U3 ( .A(n12), .Q(n8) );
  NAND22 U4 ( .A(n31), .B(n3), .Q(n4) );
  NOR41 U5 ( .A(n55), .B(i_con_FuncCode[4]), .C(n53), .D(n54), .Q(n59) );
  XNR21 U6 ( .A(i_con_FuncCode[0]), .B(i_con_FuncCode[1]), .Q(n13) );
  CLKIN6 U7 ( .A(n31), .Q(n42) );
  NAND22 U8 ( .A(i_con_FuncCode[3]), .B(n12), .Q(n52) );
  INV4 U9 ( .A(n5), .Q(n43) );
  INV3 U10 ( .A(n7), .Q(n15) );
  NOR22 U11 ( .A(n28), .B(n46), .Q(n1) );
  CLKIN6 U12 ( .A(i_con_FuncCode[3]), .Q(n29) );
  CLKIN0 U13 ( .A(n24), .Q(n6) );
  INV3 U14 ( .A(n33), .Q(n35) );
  INV3 U15 ( .A(n22), .Q(n36) );
  NAND23 U16 ( .A(n8), .B(n24), .Q(n27) );
  NAND32 U17 ( .A(i_con_FuncCode[5]), .B(n30), .C(n29), .Q(n31) );
  CLKIN4 U18 ( .A(i_con_FuncCode[0]), .Q(n12) );
  NOR31 U19 ( .A(n2), .B(n5), .C(n36), .Q(n40) );
  INV3 U20 ( .A(n1), .Q(n2) );
  CLKIN6 U21 ( .A(n11), .Q(n28) );
  NAND22 U22 ( .A(n4), .B(n6), .Q(n44) );
  CLKIN6 U23 ( .A(i_con_FuncCode[5]), .Q(n41) );
  CLKIN6 U24 ( .A(i_con_FuncCode[2]), .Q(n30) );
  INV1 U25 ( .A(n41), .Q(n3) );
  AOI211 U26 ( .A(n41), .B(n8), .C(n46), .Q(n7) );
  AOI312 U27 ( .A(n29), .B(n30), .C(n27), .D(n26), .Q(n5) );
  INV4 U28 ( .A(n23), .Q(n46) );
  NOR31 U29 ( .A(n37), .B(n36), .C(n35), .Q(n38) );
  NOR42 U30 ( .A(i_con_FuncCode[4]), .B(n28), .C(n15), .D(n14), .Q(n21) );
  NAND22 U31 ( .A(i_con_FuncCode[0]), .B(i_con_FuncCode[3]), .Q(n23) );
  CLKIN4 U32 ( .A(i_con_FuncCode[1]), .Q(n24) );
  CLKIN6 U33 ( .A(i_con_AluOp[4]), .Q(n16) );
  NAND21 U34 ( .A(n48), .B(i_con_AluOp[4]), .Q(n49) );
  INV3 U35 ( .A(n56), .Q(n50) );
  AOI311 U36 ( .A(i_con_AluOp[3]), .B(i_con_AluOp[2]), .C(i_con_AluOp[0]), .D(
        n56), .Q(n57) );
  NAND22 U37 ( .A(i_con_FuncCode[1]), .B(i_con_FuncCode[5]), .Q(n25) );
  NOR31 U38 ( .A(i_con_FuncCode[4]), .B(n53), .C(n46), .Q(n9) );
  NOR24 U39 ( .A(n10), .B(n47), .Q(n51) );
  INV6 U40 ( .A(n9), .Q(n10) );
  INV3 U41 ( .A(n45), .Q(n53) );
  NAND21 U42 ( .A(i_con_FuncCode[1]), .B(i_con_FuncCode[2]), .Q(n45) );
  NAND24 U43 ( .A(n44), .B(n43), .Q(n47) );
  NAND22 U44 ( .A(n41), .B(n24), .Q(n11) );
  OAI212 U45 ( .A(n13), .B(n30), .C(n52), .Q(n14) );
  CLKIN3 U46 ( .A(i_con_AluOp[0]), .Q(n37) );
  NAND22 U47 ( .A(i_con_AluOp[1]), .B(n37), .Q(n58) );
  NAND22 U48 ( .A(i_con_AluOp[3]), .B(n16), .Q(n32) );
  CLKIN3 U49 ( .A(i_con_AluOp[2]), .Q(n18) );
  OAI212 U50 ( .A(i_con_AluOp[3]), .B(n16), .C(i_con_AluOp[1]), .Q(n17) );
  OAI212 U51 ( .A(i_con_AluOp[5]), .B(n17), .C(i_con_AluOp[0]), .Q(n22) );
  OAI312 U52 ( .A(n32), .B(n37), .C(n18), .D(n22), .Q(n56) );
  NAND22 U53 ( .A(i_con_AluOp[0]), .B(n18), .Q(n19) );
  CLKIN3 U54 ( .A(n19), .Q(n48) );
  NAND22 U55 ( .A(n48), .B(i_con_AluOp[3]), .Q(n20) );
  OAI2112 U56 ( .A(n21), .B(n58), .C(n50), .D(n20), .Q(o_con_AluCtrl[0]) );
  OAI222 U57 ( .A(n25), .B(i_con_FuncCode[2]), .C(i_con_FuncCode[3]), .D(n41), 
        .Q(n26) );
  AOI312 U58 ( .A(n29), .B(n30), .C(n27), .D(n26), .Q(n54) );
  CLKIN3 U59 ( .A(i_con_AluOp[1]), .Q(n34) );
  NAND22 U60 ( .A(n48), .B(n32), .Q(n33) );
  NOR41 U61 ( .A(i_con_FuncCode[4]), .B(n34), .C(n42), .D(n35), .Q(n39) );
  AOI212 U62 ( .A(n40), .B(n39), .C(n38), .Q(o_con_AluCtrl[1]) );
  OAI2112 U63 ( .A(n51), .B(n58), .C(n50), .D(n49), .Q(o_con_AluCtrl[2]) );
  CLKIN3 U64 ( .A(n52), .Q(n55) );
  OAI212 U65 ( .A(n59), .B(n58), .C(n57), .Q(o_con_AluCtrl[3]) );
endmodule


module E_famux5 ( i_data_rs, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fa, o_data_alusra );
  input [31:0] i_data_rs;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fa;
  output [31:0] o_data_alusra;
  wire   N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, n1, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16;

  DLPQ3 o_data_alusra_reg_31_ ( .SN(n1), .D(N53), .GN(n11), .Q(
        o_data_alusra[31]) );
  DLPQ3 o_data_alusra_reg_30_ ( .SN(n1), .D(N52), .GN(n11), .Q(
        o_data_alusra[30]) );
  DLPQ3 o_data_alusra_reg_29_ ( .SN(n1), .D(N51), .GN(n11), .Q(
        o_data_alusra[29]) );
  DLPQ3 o_data_alusra_reg_28_ ( .SN(n1), .D(N50), .GN(n11), .Q(
        o_data_alusra[28]) );
  DLPQ3 o_data_alusra_reg_27_ ( .SN(n1), .D(N49), .GN(n10), .Q(
        o_data_alusra[27]) );
  DLPQ3 o_data_alusra_reg_26_ ( .SN(n1), .D(N48), .GN(n10), .Q(
        o_data_alusra[26]) );
  DLPQ3 o_data_alusra_reg_25_ ( .SN(n1), .D(N47), .GN(n10), .Q(
        o_data_alusra[25]) );
  DLPQ3 o_data_alusra_reg_24_ ( .SN(n1), .D(N46), .GN(n10), .Q(
        o_data_alusra[24]) );
  DLPQ3 o_data_alusra_reg_23_ ( .SN(n1), .D(N45), .GN(n10), .Q(
        o_data_alusra[23]) );
  DLPQ3 o_data_alusra_reg_22_ ( .SN(n1), .D(N44), .GN(n10), .Q(
        o_data_alusra[22]) );
  DLPQ3 o_data_alusra_reg_21_ ( .SN(n1), .D(N43), .GN(n10), .Q(
        o_data_alusra[21]) );
  DLPQ3 o_data_alusra_reg_20_ ( .SN(n1), .D(N42), .GN(n9), .Q(
        o_data_alusra[20]) );
  DLPQ3 o_data_alusra_reg_19_ ( .SN(n1), .D(N41), .GN(n9), .Q(
        o_data_alusra[19]) );
  DLPQ3 o_data_alusra_reg_18_ ( .SN(n1), .D(N40), .GN(n9), .Q(
        o_data_alusra[18]) );
  DLPQ3 o_data_alusra_reg_17_ ( .SN(n1), .D(N39), .GN(n9), .Q(
        o_data_alusra[17]) );
  DLPQ3 o_data_alusra_reg_16_ ( .SN(n1), .D(N38), .GN(n9), .Q(
        o_data_alusra[16]) );
  DLPQ3 o_data_alusra_reg_15_ ( .SN(n1), .D(N37), .GN(n9), .Q(
        o_data_alusra[15]) );
  DLPQ3 o_data_alusra_reg_14_ ( .SN(n1), .D(N36), .GN(n9), .Q(
        o_data_alusra[14]) );
  DLPQ3 o_data_alusra_reg_13_ ( .SN(n1), .D(N35), .GN(n8), .Q(
        o_data_alusra[13]) );
  DLPQ3 o_data_alusra_reg_12_ ( .SN(n1), .D(N34), .GN(n8), .Q(
        o_data_alusra[12]) );
  DLPQ3 o_data_alusra_reg_11_ ( .SN(n1), .D(N33), .GN(n8), .Q(
        o_data_alusra[11]) );
  DLPQ3 o_data_alusra_reg_10_ ( .SN(n1), .D(N32), .GN(n8), .Q(
        o_data_alusra[10]) );
  DLPQ3 o_data_alusra_reg_9_ ( .SN(n1), .D(N31), .GN(n8), .Q(o_data_alusra[9])
         );
  DLPQ3 o_data_alusra_reg_8_ ( .SN(n1), .D(N30), .GN(n8), .Q(o_data_alusra[8])
         );
  DLPQ3 o_data_alusra_reg_7_ ( .SN(n1), .D(N29), .GN(n8), .Q(o_data_alusra[7])
         );
  DLPQ3 o_data_alusra_reg_6_ ( .SN(n1), .D(N28), .GN(n138), .Q(
        o_data_alusra[6]) );
  DLPQ3 o_data_alusra_reg_5_ ( .SN(n1), .D(N27), .GN(n11), .Q(o_data_alusra[5]) );
  DLPQ3 o_data_alusra_reg_4_ ( .SN(n1), .D(N26), .GN(n138), .Q(
        o_data_alusra[4]) );
  DLPQ3 o_data_alusra_reg_3_ ( .SN(n1), .D(N25), .GN(n138), .Q(
        o_data_alusra[3]) );
  DLPQ3 o_data_alusra_reg_2_ ( .SN(n1), .D(N24), .GN(n138), .Q(
        o_data_alusra[2]) );
  DLPQ3 o_data_alusra_reg_1_ ( .SN(n1), .D(N23), .GN(n11), .Q(o_data_alusra[1]) );
  DLPQ3 o_data_alusra_reg_0_ ( .SN(n1), .D(N22), .GN(n11), .Q(o_data_alusra[0]) );
  AOI220 U2 ( .A(i_data_alures[15]), .B(n7), .C(i_data_writeres[15]), .D(n6), 
        .Q(n92) );
  AOI220 U3 ( .A(i_data_alures[16]), .B(n7), .C(i_data_writeres[16]), .D(n41), 
        .Q(n89) );
  AOI220 U4 ( .A(i_data_alures[17]), .B(n7), .C(i_data_writeres[17]), .D(n6), 
        .Q(n86) );
  AOI220 U5 ( .A(i_data_alures[19]), .B(n7), .C(i_data_writeres[19]), .D(n41), 
        .Q(n80) );
  AOI220 U6 ( .A(i_data_alures[20]), .B(n7), .C(i_data_writeres[20]), .D(n6), 
        .Q(n77) );
  AOI220 U7 ( .A(i_data_alures[21]), .B(n7), .C(i_data_writeres[21]), .D(n41), 
        .Q(n74) );
  AOI220 U8 ( .A(i_data_alures[22]), .B(n7), .C(i_data_writeres[22]), .D(n41), 
        .Q(n71) );
  AOI220 U9 ( .A(i_data_alures[23]), .B(n7), .C(i_data_writeres[23]), .D(n6), 
        .Q(n68) );
  AOI220 U10 ( .A(i_data_alures[24]), .B(n7), .C(i_data_writeres[24]), .D(n6), 
        .Q(n65) );
  AOI220 U11 ( .A(i_data_alures[25]), .B(n7), .C(i_data_writeres[25]), .D(n41), 
        .Q(n62) );
  AOI220 U12 ( .A(i_data_alures[26]), .B(n7), .C(i_data_writeres[26]), .D(n6), 
        .Q(n59) );
  AOI220 U13 ( .A(i_data_alures[27]), .B(n7), .C(i_data_writeres[27]), .D(n41), 
        .Q(n56) );
  AOI220 U14 ( .A(i_data_alures[28]), .B(n7), .C(i_data_writeres[28]), .D(n41), 
        .Q(n53) );
  AOI220 U15 ( .A(i_data_alures[29]), .B(n7), .C(i_data_writeres[29]), .D(n6), 
        .Q(n50) );
  AOI220 U16 ( .A(i_data_alures[30]), .B(n7), .C(i_data_writeres[30]), .D(n6), 
        .Q(n47) );
  AOI220 U17 ( .A(i_data_alures[31]), .B(n7), .C(i_data_writeres[31]), .D(n41), 
        .Q(n39) );
  AOI220 U18 ( .A(i_data_alures[0]), .B(n40), .C(i_data_writeres[0]), .D(n41), 
        .Q(n137) );
  AOI220 U19 ( .A(i_data_alures[1]), .B(n40), .C(i_data_writeres[1]), .D(n41), 
        .Q(n134) );
  AOI220 U20 ( .A(i_data_alures[2]), .B(n40), .C(i_data_writeres[2]), .D(n6), 
        .Q(n131) );
  AOI220 U21 ( .A(i_data_alures[3]), .B(n40), .C(i_data_writeres[3]), .D(n6), 
        .Q(n128) );
  AOI220 U22 ( .A(i_data_alures[4]), .B(n40), .C(i_data_writeres[4]), .D(n41), 
        .Q(n125) );
  AOI220 U23 ( .A(i_data_alures[5]), .B(n40), .C(i_data_writeres[5]), .D(n6), 
        .Q(n122) );
  AOI220 U24 ( .A(i_data_alures[6]), .B(n40), .C(i_data_writeres[6]), .D(n41), 
        .Q(n119) );
  NAND20 U25 ( .A(i_data_lwM[7]), .B(n12), .Q(n115) );
  AOI220 U26 ( .A(i_data_alures[7]), .B(n40), .C(i_data_writeres[7]), .D(n41), 
        .Q(n116) );
  AOI220 U27 ( .A(i_data_alures[8]), .B(n40), .C(i_data_writeres[8]), .D(n6), 
        .Q(n113) );
  AOI220 U28 ( .A(i_data_alures[9]), .B(n40), .C(i_data_writeres[9]), .D(n6), 
        .Q(n110) );
  AOI220 U29 ( .A(i_data_alures[10]), .B(n40), .C(i_data_writeres[10]), .D(n41), .Q(n107) );
  AOI220 U30 ( .A(i_data_alures[11]), .B(n40), .C(i_data_writeres[11]), .D(n6), 
        .Q(n104) );
  AOI220 U31 ( .A(i_data_alures[12]), .B(n40), .C(i_data_writeres[12]), .D(n41), .Q(n101) );
  AOI220 U32 ( .A(i_data_alures[13]), .B(n40), .C(i_data_writeres[13]), .D(n6), 
        .Q(n98) );
  AOI220 U33 ( .A(i_data_alures[14]), .B(n40), .C(i_data_writeres[14]), .D(n6), 
        .Q(n95) );
  BUF2 U34 ( .A(n138), .Q(n8) );
  BUF2 U35 ( .A(n138), .Q(n9) );
  BUF2 U36 ( .A(n138), .Q(n10) );
  BUF2 U37 ( .A(n138), .Q(n11) );
  NOR40 U38 ( .A(n2), .B(n12), .C(n14), .D(n40), .Q(n138) );
  INV3 U39 ( .A(n139), .Q(n14) );
  NOR21 U40 ( .A(n4), .B(n6), .Q(n139) );
  BUF2 U41 ( .A(n44), .Q(n2) );
  BUF2 U42 ( .A(n40), .Q(n7) );
  INV3 U43 ( .A(n5), .Q(n6) );
  INV3 U44 ( .A(n3), .Q(n4) );
  BUF2 U45 ( .A(n42), .Q(n12) );
  NOR31 U46 ( .A(i_con_fa[0]), .B(i_con_fa[1]), .C(n13), .Q(n42) );
  NOR31 U47 ( .A(n16), .B(i_con_fa[1]), .C(n13), .Q(n44) );
  NOR31 U48 ( .A(i_con_fa[0]), .B(i_con_fa[2]), .C(n15), .Q(n40) );
  INV3 U49 ( .A(i_con_fa[1]), .Q(n15) );
  NAND31 U50 ( .A(n81), .B(n82), .C(n83), .Q(N40) );
  NAND22 U51 ( .A(i_data_lwM[18]), .B(n42), .Q(n82) );
  AOI221 U52 ( .A(i_data_rs[18]), .B(n4), .C(i_data_lwW[18]), .D(n44), .Q(n81)
         );
  NAND31 U53 ( .A(n93), .B(n94), .C(n95), .Q(N36) );
  NAND22 U54 ( .A(i_data_lwM[14]), .B(n12), .Q(n94) );
  AOI221 U55 ( .A(i_data_rs[14]), .B(n43), .C(i_data_lwW[14]), .D(n2), .Q(n93)
         );
  NAND31 U56 ( .A(n87), .B(n88), .C(n89), .Q(N38) );
  NAND22 U57 ( .A(i_data_lwM[16]), .B(n42), .Q(n88) );
  AOI221 U58 ( .A(i_data_rs[16]), .B(n43), .C(i_data_lwW[16]), .D(n44), .Q(n87) );
  NAND31 U59 ( .A(n66), .B(n67), .C(n68), .Q(N45) );
  NAND22 U60 ( .A(i_data_lwM[23]), .B(n12), .Q(n67) );
  AOI221 U61 ( .A(i_data_rs[23]), .B(n43), .C(i_data_lwW[23]), .D(n44), .Q(n66) );
  NAND31 U62 ( .A(n60), .B(n61), .C(n62), .Q(N47) );
  NAND22 U63 ( .A(i_data_lwM[25]), .B(n12), .Q(n61) );
  AOI221 U64 ( .A(i_data_rs[25]), .B(n4), .C(i_data_lwW[25]), .D(n44), .Q(n60)
         );
  NAND31 U65 ( .A(n54), .B(n55), .C(n56), .Q(N49) );
  NAND22 U66 ( .A(i_data_lwM[27]), .B(n12), .Q(n55) );
  AOI221 U67 ( .A(i_data_rs[27]), .B(n4), .C(i_data_lwW[27]), .D(n44), .Q(n54)
         );
  NAND31 U68 ( .A(n51), .B(n52), .C(n53), .Q(N50) );
  NAND22 U69 ( .A(i_data_lwM[28]), .B(n12), .Q(n52) );
  AOI221 U70 ( .A(i_data_rs[28]), .B(n43), .C(i_data_lwW[28]), .D(n44), .Q(n51) );
  NAND31 U71 ( .A(n135), .B(n136), .C(n137), .Q(N22) );
  NAND22 U72 ( .A(i_data_lwM[0]), .B(n42), .Q(n136) );
  AOI221 U73 ( .A(i_data_rs[0]), .B(n4), .C(i_data_lwW[0]), .D(n2), .Q(n135)
         );
  NAND31 U74 ( .A(n132), .B(n133), .C(n134), .Q(N23) );
  NAND22 U75 ( .A(i_data_lwM[1]), .B(n42), .Q(n133) );
  AOI221 U76 ( .A(i_data_rs[1]), .B(n4), .C(i_data_lwW[1]), .D(n2), .Q(n132)
         );
  NAND31 U77 ( .A(n129), .B(n130), .C(n131), .Q(N24) );
  NAND22 U78 ( .A(i_data_lwM[2]), .B(n42), .Q(n130) );
  AOI221 U79 ( .A(i_data_rs[2]), .B(n43), .C(i_data_lwW[2]), .D(n2), .Q(n129)
         );
  NAND31 U80 ( .A(n126), .B(n127), .C(n128), .Q(N25) );
  NAND22 U81 ( .A(i_data_lwM[3]), .B(n42), .Q(n127) );
  AOI221 U82 ( .A(i_data_rs[3]), .B(n4), .C(i_data_lwW[3]), .D(n2), .Q(n126)
         );
  NAND31 U83 ( .A(n123), .B(n124), .C(n125), .Q(N26) );
  NAND22 U84 ( .A(i_data_lwM[4]), .B(n42), .Q(n124) );
  AOI221 U85 ( .A(i_data_rs[4]), .B(n43), .C(i_data_lwW[4]), .D(n2), .Q(n123)
         );
  NAND31 U86 ( .A(n120), .B(n121), .C(n122), .Q(N27) );
  NAND22 U87 ( .A(i_data_lwM[5]), .B(n42), .Q(n121) );
  AOI221 U88 ( .A(i_data_rs[5]), .B(n43), .C(i_data_lwW[5]), .D(n2), .Q(n120)
         );
  NAND31 U89 ( .A(n117), .B(n118), .C(n119), .Q(N28) );
  NAND22 U90 ( .A(i_data_lwM[6]), .B(n42), .Q(n118) );
  AOI221 U91 ( .A(i_data_rs[6]), .B(n4), .C(i_data_lwW[6]), .D(n2), .Q(n117)
         );
  NAND31 U92 ( .A(n114), .B(n115), .C(n116), .Q(N29) );
  AOI221 U93 ( .A(i_data_rs[7]), .B(n4), .C(i_data_lwW[7]), .D(n2), .Q(n114)
         );
  NAND31 U94 ( .A(n111), .B(n112), .C(n113), .Q(N30) );
  NAND22 U95 ( .A(i_data_lwM[8]), .B(n12), .Q(n112) );
  AOI221 U96 ( .A(i_data_rs[8]), .B(n43), .C(i_data_lwW[8]), .D(n2), .Q(n111)
         );
  NAND31 U97 ( .A(n108), .B(n109), .C(n110), .Q(N31) );
  NAND22 U98 ( .A(i_data_lwM[9]), .B(n42), .Q(n109) );
  AOI221 U99 ( .A(i_data_rs[9]), .B(n4), .C(i_data_lwW[9]), .D(n2), .Q(n108)
         );
  NAND31 U100 ( .A(n105), .B(n106), .C(n107), .Q(N32) );
  NAND22 U101 ( .A(i_data_lwM[10]), .B(n12), .Q(n106) );
  AOI221 U102 ( .A(i_data_rs[10]), .B(n43), .C(i_data_lwW[10]), .D(n2), .Q(
        n105) );
  NAND31 U103 ( .A(n102), .B(n103), .C(n104), .Q(N33) );
  NAND22 U104 ( .A(i_data_lwM[11]), .B(n42), .Q(n103) );
  AOI221 U105 ( .A(i_data_rs[11]), .B(n43), .C(i_data_lwW[11]), .D(n2), .Q(
        n102) );
  NAND31 U106 ( .A(n99), .B(n100), .C(n101), .Q(N34) );
  NAND22 U107 ( .A(i_data_lwM[12]), .B(n42), .Q(n100) );
  AOI221 U108 ( .A(i_data_rs[12]), .B(n4), .C(i_data_lwW[12]), .D(n2), .Q(n99)
         );
  NAND31 U109 ( .A(n96), .B(n97), .C(n98), .Q(N35) );
  NAND22 U110 ( .A(i_data_lwM[13]), .B(n12), .Q(n97) );
  AOI221 U111 ( .A(i_data_rs[13]), .B(n4), .C(i_data_lwW[13]), .D(n2), .Q(n96)
         );
  NAND31 U112 ( .A(n90), .B(n91), .C(n92), .Q(N37) );
  NAND22 U113 ( .A(i_data_lwM[15]), .B(n12), .Q(n91) );
  AOI221 U114 ( .A(i_data_rs[15]), .B(n4), .C(i_data_lwW[15]), .D(n44), .Q(n90) );
  NAND31 U115 ( .A(n84), .B(n85), .C(n86), .Q(N39) );
  NAND22 U116 ( .A(i_data_lwM[17]), .B(n12), .Q(n85) );
  AOI221 U117 ( .A(i_data_rs[17]), .B(n43), .C(i_data_lwW[17]), .D(n44), .Q(
        n84) );
  NAND31 U118 ( .A(n78), .B(n79), .C(n80), .Q(N41) );
  NAND22 U119 ( .A(i_data_lwM[19]), .B(n12), .Q(n79) );
  AOI221 U120 ( .A(i_data_rs[19]), .B(n4), .C(i_data_lwW[19]), .D(n44), .Q(n78) );
  NAND31 U121 ( .A(n75), .B(n76), .C(n77), .Q(N42) );
  NAND22 U122 ( .A(i_data_lwM[20]), .B(n12), .Q(n76) );
  AOI221 U123 ( .A(i_data_rs[20]), .B(n43), .C(i_data_lwW[20]), .D(n44), .Q(
        n75) );
  NAND31 U124 ( .A(n72), .B(n73), .C(n74), .Q(N43) );
  NAND22 U125 ( .A(i_data_lwM[21]), .B(n12), .Q(n73) );
  AOI221 U126 ( .A(i_data_rs[21]), .B(n4), .C(i_data_lwW[21]), .D(n44), .Q(n72) );
  NAND31 U127 ( .A(n69), .B(n70), .C(n71), .Q(N44) );
  NAND22 U128 ( .A(i_data_lwM[22]), .B(n12), .Q(n70) );
  AOI221 U129 ( .A(i_data_rs[22]), .B(n4), .C(i_data_lwW[22]), .D(n44), .Q(n69) );
  NAND31 U130 ( .A(n63), .B(n64), .C(n65), .Q(N46) );
  NAND22 U131 ( .A(i_data_lwM[24]), .B(n12), .Q(n64) );
  AOI221 U132 ( .A(i_data_rs[24]), .B(n4), .C(i_data_lwW[24]), .D(n44), .Q(n63) );
  NAND31 U133 ( .A(n57), .B(n58), .C(n59), .Q(N48) );
  NAND22 U134 ( .A(i_data_lwM[26]), .B(n12), .Q(n58) );
  AOI221 U135 ( .A(i_data_rs[26]), .B(n43), .C(i_data_lwW[26]), .D(n44), .Q(
        n57) );
  NAND31 U136 ( .A(n48), .B(n49), .C(n50), .Q(N51) );
  NAND22 U137 ( .A(i_data_lwM[29]), .B(n12), .Q(n49) );
  AOI221 U138 ( .A(i_data_rs[29]), .B(n43), .C(i_data_lwW[29]), .D(n44), .Q(
        n48) );
  NAND31 U139 ( .A(n45), .B(n46), .C(n47), .Q(N52) );
  NAND22 U140 ( .A(i_data_lwM[30]), .B(n12), .Q(n46) );
  AOI221 U141 ( .A(i_data_rs[30]), .B(n4), .C(i_data_lwW[30]), .D(n2), .Q(n45)
         );
  NAND31 U142 ( .A(n37), .B(n38), .C(n39), .Q(N53) );
  NAND22 U143 ( .A(i_data_lwM[31]), .B(n12), .Q(n38) );
  AOI221 U144 ( .A(i_data_rs[31]), .B(n4), .C(i_data_lwW[31]), .D(n2), .Q(n37)
         );
  INV3 U145 ( .A(n41), .Q(n5) );
  NOR31 U146 ( .A(i_con_fa[1]), .B(i_con_fa[2]), .C(n16), .Q(n41) );
  INV3 U147 ( .A(n43), .Q(n3) );
  NOR31 U148 ( .A(i_con_fa[1]), .B(i_con_fa[2]), .C(i_con_fa[0]), .Q(n43) );
  INV3 U149 ( .A(i_con_fa[0]), .Q(n16) );
  INV3 U150 ( .A(i_con_fa[2]), .Q(n13) );
  AOI221 U151 ( .A(i_data_alures[18]), .B(n7), .C(i_data_writeres[18]), .D(n41), .Q(n83) );
  LOGIC1 U152 ( .Q(n1) );
endmodule


module E_fbmux5 ( i_data_rt, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fb, o_data_alusrb );
  input [31:0] i_data_rt;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fb;
  output [31:0] o_data_alusrb;
  wire   N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, n1, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13;

  DLPQ3 o_data_alusrb_reg_31_ ( .SN(n1), .D(N53), .GN(n8), .Q(
        o_data_alusrb[31]) );
  DLPQ3 o_data_alusrb_reg_30_ ( .SN(n1), .D(N52), .GN(n8), .Q(
        o_data_alusrb[30]) );
  DLPQ3 o_data_alusrb_reg_29_ ( .SN(n1), .D(N51), .GN(n8), .Q(
        o_data_alusrb[29]) );
  DLPQ3 o_data_alusrb_reg_28_ ( .SN(n1), .D(N50), .GN(n8), .Q(
        o_data_alusrb[28]) );
  DLPQ3 o_data_alusrb_reg_27_ ( .SN(n1), .D(N49), .GN(n8), .Q(
        o_data_alusrb[27]) );
  DLPQ3 o_data_alusrb_reg_26_ ( .SN(n1), .D(N48), .GN(n138), .Q(
        o_data_alusrb[26]) );
  DLPQ3 o_data_alusrb_reg_25_ ( .SN(n1), .D(N47), .GN(n8), .Q(
        o_data_alusrb[25]) );
  DLPQ3 o_data_alusrb_reg_24_ ( .SN(n1), .D(N46), .GN(n8), .Q(
        o_data_alusrb[24]) );
  DLPQ3 o_data_alusrb_reg_23_ ( .SN(n1), .D(N45), .GN(n8), .Q(
        o_data_alusrb[23]) );
  DLPQ3 o_data_alusrb_reg_22_ ( .SN(n1), .D(N44), .GN(n8), .Q(
        o_data_alusrb[22]) );
  DLPQ3 o_data_alusrb_reg_21_ ( .SN(n1), .D(N43), .GN(n8), .Q(
        o_data_alusrb[21]) );
  DLPQ3 o_data_alusrb_reg_20_ ( .SN(n1), .D(N42), .GN(n8), .Q(
        o_data_alusrb[20]) );
  DLPQ3 o_data_alusrb_reg_19_ ( .SN(n1), .D(N41), .GN(n8), .Q(
        o_data_alusrb[19]) );
  DLPQ3 o_data_alusrb_reg_18_ ( .SN(n1), .D(N40), .GN(n8), .Q(
        o_data_alusrb[18]) );
  DLPQ3 o_data_alusrb_reg_17_ ( .SN(n1), .D(N39), .GN(n8), .Q(
        o_data_alusrb[17]) );
  DLPQ3 o_data_alusrb_reg_16_ ( .SN(n1), .D(N38), .GN(n8), .Q(
        o_data_alusrb[16]) );
  DLPQ3 o_data_alusrb_reg_15_ ( .SN(n1), .D(N37), .GN(n138), .Q(
        o_data_alusrb[15]) );
  DLPQ3 o_data_alusrb_reg_14_ ( .SN(n1), .D(N36), .GN(n8), .Q(
        o_data_alusrb[14]) );
  DLPQ3 o_data_alusrb_reg_13_ ( .SN(n1), .D(N35), .GN(n8), .Q(
        o_data_alusrb[13]) );
  DLPQ3 o_data_alusrb_reg_12_ ( .SN(n1), .D(N34), .GN(n138), .Q(
        o_data_alusrb[12]) );
  DLPQ3 o_data_alusrb_reg_11_ ( .SN(n1), .D(N33), .GN(n8), .Q(
        o_data_alusrb[11]) );
  DLPQ3 o_data_alusrb_reg_10_ ( .SN(n1), .D(N32), .GN(n8), .Q(
        o_data_alusrb[10]) );
  DLPQ3 o_data_alusrb_reg_9_ ( .SN(n1), .D(N31), .GN(n8), .Q(o_data_alusrb[9])
         );
  DLPQ3 o_data_alusrb_reg_8_ ( .SN(n1), .D(N30), .GN(n8), .Q(o_data_alusrb[8])
         );
  DLPQ3 o_data_alusrb_reg_7_ ( .SN(n1), .D(N29), .GN(n138), .Q(
        o_data_alusrb[7]) );
  DLPQ3 o_data_alusrb_reg_6_ ( .SN(n1), .D(N28), .GN(n138), .Q(
        o_data_alusrb[6]) );
  DLPQ3 o_data_alusrb_reg_5_ ( .SN(n1), .D(N27), .GN(n8), .Q(o_data_alusrb[5])
         );
  DLPQ3 o_data_alusrb_reg_4_ ( .SN(n1), .D(N26), .GN(n138), .Q(
        o_data_alusrb[4]) );
  DLPQ3 o_data_alusrb_reg_3_ ( .SN(n1), .D(N25), .GN(n8), .Q(o_data_alusrb[3])
         );
  DLPQ3 o_data_alusrb_reg_2_ ( .SN(n1), .D(N24), .GN(n138), .Q(
        o_data_alusrb[2]) );
  DLPQ3 o_data_alusrb_reg_1_ ( .SN(n1), .D(N23), .GN(n138), .Q(
        o_data_alusrb[1]) );
  DLPQ3 o_data_alusrb_reg_0_ ( .SN(n1), .D(N22), .GN(n8), .Q(o_data_alusrb[0])
         );
  AOI220 U2 ( .A(i_data_alures[15]), .B(n7), .C(i_data_writeres[15]), .D(n6), 
        .Q(n92) );
  AOI220 U3 ( .A(i_data_alures[16]), .B(n7), .C(i_data_writeres[16]), .D(n41), 
        .Q(n89) );
  AOI220 U4 ( .A(i_data_alures[17]), .B(n7), .C(i_data_writeres[17]), .D(n6), 
        .Q(n86) );
  AOI220 U5 ( .A(i_data_alures[19]), .B(n7), .C(i_data_writeres[19]), .D(n41), 
        .Q(n80) );
  AOI220 U6 ( .A(i_data_alures[20]), .B(n7), .C(i_data_writeres[20]), .D(n6), 
        .Q(n77) );
  AOI220 U7 ( .A(i_data_alures[21]), .B(n7), .C(i_data_writeres[21]), .D(n41), 
        .Q(n74) );
  AOI220 U8 ( .A(i_data_alures[22]), .B(n7), .C(i_data_writeres[22]), .D(n41), 
        .Q(n71) );
  AOI220 U9 ( .A(i_data_alures[23]), .B(n7), .C(i_data_writeres[23]), .D(n6), 
        .Q(n68) );
  AOI220 U10 ( .A(i_data_alures[24]), .B(n7), .C(i_data_writeres[24]), .D(n6), 
        .Q(n65) );
  AOI220 U11 ( .A(i_data_alures[25]), .B(n7), .C(i_data_writeres[25]), .D(n41), 
        .Q(n62) );
  AOI220 U12 ( .A(i_data_alures[26]), .B(n7), .C(i_data_writeres[26]), .D(n6), 
        .Q(n59) );
  AOI220 U13 ( .A(i_data_alures[27]), .B(n7), .C(i_data_writeres[27]), .D(n41), 
        .Q(n56) );
  AOI220 U14 ( .A(i_data_alures[28]), .B(n7), .C(i_data_writeres[28]), .D(n41), 
        .Q(n53) );
  AOI220 U15 ( .A(i_data_alures[29]), .B(n7), .C(i_data_writeres[29]), .D(n6), 
        .Q(n50) );
  AOI220 U16 ( .A(i_data_alures[30]), .B(n7), .C(i_data_writeres[30]), .D(n6), 
        .Q(n47) );
  AOI220 U17 ( .A(i_data_alures[31]), .B(n7), .C(i_data_writeres[31]), .D(n41), 
        .Q(n39) );
  AOI220 U18 ( .A(i_data_alures[0]), .B(n40), .C(i_data_writeres[0]), .D(n41), 
        .Q(n137) );
  AOI220 U19 ( .A(i_data_alures[1]), .B(n40), .C(i_data_writeres[1]), .D(n41), 
        .Q(n134) );
  AOI220 U20 ( .A(i_data_alures[2]), .B(n40), .C(i_data_writeres[2]), .D(n6), 
        .Q(n131) );
  AOI220 U21 ( .A(i_data_alures[3]), .B(n40), .C(i_data_writeres[3]), .D(n6), 
        .Q(n128) );
  AOI220 U22 ( .A(i_data_alures[4]), .B(n40), .C(i_data_writeres[4]), .D(n41), 
        .Q(n125) );
  AOI220 U23 ( .A(i_data_alures[5]), .B(n40), .C(i_data_writeres[5]), .D(n6), 
        .Q(n122) );
  AOI220 U24 ( .A(i_data_alures[6]), .B(n40), .C(i_data_writeres[6]), .D(n41), 
        .Q(n119) );
  NAND20 U25 ( .A(i_data_lwM[7]), .B(n9), .Q(n115) );
  AOI220 U26 ( .A(i_data_alures[7]), .B(n40), .C(i_data_writeres[7]), .D(n41), 
        .Q(n116) );
  AOI220 U27 ( .A(i_data_alures[8]), .B(n40), .C(i_data_writeres[8]), .D(n6), 
        .Q(n113) );
  AOI220 U28 ( .A(i_data_alures[9]), .B(n40), .C(i_data_writeres[9]), .D(n6), 
        .Q(n110) );
  AOI220 U29 ( .A(i_data_alures[10]), .B(n40), .C(i_data_writeres[10]), .D(n41), .Q(n107) );
  AOI220 U30 ( .A(i_data_alures[11]), .B(n40), .C(i_data_writeres[11]), .D(n6), 
        .Q(n104) );
  AOI220 U31 ( .A(i_data_alures[12]), .B(n40), .C(i_data_writeres[12]), .D(n41), .Q(n101) );
  AOI220 U32 ( .A(i_data_alures[13]), .B(n40), .C(i_data_writeres[13]), .D(n6), 
        .Q(n98) );
  AOI220 U33 ( .A(i_data_alures[14]), .B(n40), .C(i_data_writeres[14]), .D(n6), 
        .Q(n95) );
  BUF2 U34 ( .A(n138), .Q(n8) );
  NOR40 U35 ( .A(n2), .B(n9), .C(n11), .D(n40), .Q(n138) );
  INV3 U36 ( .A(n139), .Q(n11) );
  NOR21 U37 ( .A(n4), .B(n6), .Q(n139) );
  BUF2 U38 ( .A(n44), .Q(n2) );
  BUF2 U39 ( .A(n40), .Q(n7) );
  INV3 U40 ( .A(n5), .Q(n6) );
  INV3 U41 ( .A(n3), .Q(n4) );
  BUF2 U42 ( .A(n42), .Q(n9) );
  NOR31 U43 ( .A(i_con_fb[0]), .B(i_con_fb[1]), .C(n10), .Q(n42) );
  NOR31 U44 ( .A(n13), .B(i_con_fb[1]), .C(n10), .Q(n44) );
  NOR31 U45 ( .A(i_con_fb[0]), .B(i_con_fb[2]), .C(n12), .Q(n40) );
  INV3 U46 ( .A(i_con_fb[1]), .Q(n12) );
  NAND31 U47 ( .A(n81), .B(n82), .C(n83), .Q(N40) );
  NAND22 U48 ( .A(i_data_lwM[18]), .B(n42), .Q(n82) );
  AOI221 U49 ( .A(i_data_rt[18]), .B(n4), .C(i_data_lwW[18]), .D(n44), .Q(n81)
         );
  NAND31 U50 ( .A(n93), .B(n94), .C(n95), .Q(N36) );
  NAND22 U51 ( .A(i_data_lwM[14]), .B(n9), .Q(n94) );
  AOI221 U52 ( .A(i_data_rt[14]), .B(n43), .C(i_data_lwW[14]), .D(n2), .Q(n93)
         );
  NAND31 U53 ( .A(n87), .B(n88), .C(n89), .Q(N38) );
  NAND22 U54 ( .A(i_data_lwM[16]), .B(n42), .Q(n88) );
  AOI221 U55 ( .A(i_data_rt[16]), .B(n43), .C(i_data_lwW[16]), .D(n44), .Q(n87) );
  NAND31 U56 ( .A(n66), .B(n67), .C(n68), .Q(N45) );
  NAND22 U57 ( .A(i_data_lwM[23]), .B(n9), .Q(n67) );
  AOI221 U58 ( .A(i_data_rt[23]), .B(n43), .C(i_data_lwW[23]), .D(n44), .Q(n66) );
  NAND31 U59 ( .A(n60), .B(n61), .C(n62), .Q(N47) );
  NAND22 U60 ( .A(i_data_lwM[25]), .B(n9), .Q(n61) );
  AOI221 U61 ( .A(i_data_rt[25]), .B(n4), .C(i_data_lwW[25]), .D(n44), .Q(n60)
         );
  NAND31 U62 ( .A(n54), .B(n55), .C(n56), .Q(N49) );
  NAND22 U63 ( .A(i_data_lwM[27]), .B(n9), .Q(n55) );
  AOI221 U64 ( .A(i_data_rt[27]), .B(n4), .C(i_data_lwW[27]), .D(n44), .Q(n54)
         );
  NAND31 U65 ( .A(n51), .B(n52), .C(n53), .Q(N50) );
  NAND22 U66 ( .A(i_data_lwM[28]), .B(n9), .Q(n52) );
  AOI221 U67 ( .A(i_data_rt[28]), .B(n43), .C(i_data_lwW[28]), .D(n44), .Q(n51) );
  NAND31 U68 ( .A(n135), .B(n136), .C(n137), .Q(N22) );
  NAND22 U69 ( .A(i_data_lwM[0]), .B(n42), .Q(n136) );
  AOI221 U70 ( .A(i_data_rt[0]), .B(n4), .C(i_data_lwW[0]), .D(n2), .Q(n135)
         );
  NAND31 U71 ( .A(n132), .B(n133), .C(n134), .Q(N23) );
  NAND22 U72 ( .A(i_data_lwM[1]), .B(n42), .Q(n133) );
  AOI221 U73 ( .A(i_data_rt[1]), .B(n4), .C(i_data_lwW[1]), .D(n2), .Q(n132)
         );
  NAND31 U74 ( .A(n129), .B(n130), .C(n131), .Q(N24) );
  NAND22 U75 ( .A(i_data_lwM[2]), .B(n42), .Q(n130) );
  AOI221 U76 ( .A(i_data_rt[2]), .B(n43), .C(i_data_lwW[2]), .D(n2), .Q(n129)
         );
  NAND31 U77 ( .A(n126), .B(n127), .C(n128), .Q(N25) );
  NAND22 U78 ( .A(i_data_lwM[3]), .B(n42), .Q(n127) );
  AOI221 U79 ( .A(i_data_rt[3]), .B(n4), .C(i_data_lwW[3]), .D(n2), .Q(n126)
         );
  NAND31 U80 ( .A(n123), .B(n124), .C(n125), .Q(N26) );
  NAND22 U81 ( .A(i_data_lwM[4]), .B(n42), .Q(n124) );
  AOI221 U82 ( .A(i_data_rt[4]), .B(n43), .C(i_data_lwW[4]), .D(n2), .Q(n123)
         );
  NAND31 U83 ( .A(n120), .B(n121), .C(n122), .Q(N27) );
  NAND22 U84 ( .A(i_data_lwM[5]), .B(n42), .Q(n121) );
  AOI221 U85 ( .A(i_data_rt[5]), .B(n43), .C(i_data_lwW[5]), .D(n2), .Q(n120)
         );
  NAND31 U86 ( .A(n117), .B(n118), .C(n119), .Q(N28) );
  NAND22 U87 ( .A(i_data_lwM[6]), .B(n42), .Q(n118) );
  AOI221 U88 ( .A(i_data_rt[6]), .B(n4), .C(i_data_lwW[6]), .D(n2), .Q(n117)
         );
  NAND31 U89 ( .A(n114), .B(n115), .C(n116), .Q(N29) );
  AOI221 U90 ( .A(i_data_rt[7]), .B(n4), .C(i_data_lwW[7]), .D(n2), .Q(n114)
         );
  NAND31 U91 ( .A(n111), .B(n112), .C(n113), .Q(N30) );
  NAND22 U92 ( .A(i_data_lwM[8]), .B(n9), .Q(n112) );
  AOI221 U93 ( .A(i_data_rt[8]), .B(n43), .C(i_data_lwW[8]), .D(n2), .Q(n111)
         );
  NAND31 U94 ( .A(n108), .B(n109), .C(n110), .Q(N31) );
  NAND22 U95 ( .A(i_data_lwM[9]), .B(n42), .Q(n109) );
  AOI221 U96 ( .A(i_data_rt[9]), .B(n4), .C(i_data_lwW[9]), .D(n2), .Q(n108)
         );
  NAND31 U97 ( .A(n105), .B(n106), .C(n107), .Q(N32) );
  NAND22 U98 ( .A(i_data_lwM[10]), .B(n9), .Q(n106) );
  AOI221 U99 ( .A(i_data_rt[10]), .B(n43), .C(i_data_lwW[10]), .D(n2), .Q(n105) );
  NAND31 U100 ( .A(n102), .B(n103), .C(n104), .Q(N33) );
  NAND22 U101 ( .A(i_data_lwM[11]), .B(n42), .Q(n103) );
  AOI221 U102 ( .A(i_data_rt[11]), .B(n43), .C(i_data_lwW[11]), .D(n2), .Q(
        n102) );
  NAND31 U103 ( .A(n99), .B(n100), .C(n101), .Q(N34) );
  NAND22 U104 ( .A(i_data_lwM[12]), .B(n42), .Q(n100) );
  AOI221 U105 ( .A(i_data_rt[12]), .B(n4), .C(i_data_lwW[12]), .D(n2), .Q(n99)
         );
  NAND31 U106 ( .A(n96), .B(n97), .C(n98), .Q(N35) );
  NAND22 U107 ( .A(i_data_lwM[13]), .B(n9), .Q(n97) );
  AOI221 U108 ( .A(i_data_rt[13]), .B(n4), .C(i_data_lwW[13]), .D(n2), .Q(n96)
         );
  NAND31 U109 ( .A(n90), .B(n91), .C(n92), .Q(N37) );
  NAND22 U110 ( .A(i_data_lwM[15]), .B(n9), .Q(n91) );
  AOI221 U111 ( .A(i_data_rt[15]), .B(n4), .C(i_data_lwW[15]), .D(n44), .Q(n90) );
  NAND31 U112 ( .A(n84), .B(n85), .C(n86), .Q(N39) );
  NAND22 U113 ( .A(i_data_lwM[17]), .B(n9), .Q(n85) );
  AOI221 U114 ( .A(i_data_rt[17]), .B(n43), .C(i_data_lwW[17]), .D(n44), .Q(
        n84) );
  NAND31 U115 ( .A(n78), .B(n79), .C(n80), .Q(N41) );
  NAND22 U116 ( .A(i_data_lwM[19]), .B(n9), .Q(n79) );
  AOI221 U117 ( .A(i_data_rt[19]), .B(n4), .C(i_data_lwW[19]), .D(n44), .Q(n78) );
  NAND31 U118 ( .A(n75), .B(n76), .C(n77), .Q(N42) );
  NAND22 U119 ( .A(i_data_lwM[20]), .B(n9), .Q(n76) );
  AOI221 U120 ( .A(i_data_rt[20]), .B(n43), .C(i_data_lwW[20]), .D(n44), .Q(
        n75) );
  NAND31 U121 ( .A(n72), .B(n73), .C(n74), .Q(N43) );
  NAND22 U122 ( .A(i_data_lwM[21]), .B(n9), .Q(n73) );
  AOI221 U123 ( .A(i_data_rt[21]), .B(n4), .C(i_data_lwW[21]), .D(n44), .Q(n72) );
  NAND31 U124 ( .A(n69), .B(n70), .C(n71), .Q(N44) );
  NAND22 U125 ( .A(i_data_lwM[22]), .B(n9), .Q(n70) );
  AOI221 U126 ( .A(i_data_rt[22]), .B(n4), .C(i_data_lwW[22]), .D(n44), .Q(n69) );
  NAND31 U127 ( .A(n63), .B(n64), .C(n65), .Q(N46) );
  NAND22 U128 ( .A(i_data_lwM[24]), .B(n9), .Q(n64) );
  AOI221 U129 ( .A(i_data_rt[24]), .B(n4), .C(i_data_lwW[24]), .D(n44), .Q(n63) );
  NAND31 U130 ( .A(n57), .B(n58), .C(n59), .Q(N48) );
  NAND22 U131 ( .A(i_data_lwM[26]), .B(n9), .Q(n58) );
  AOI221 U132 ( .A(i_data_rt[26]), .B(n43), .C(i_data_lwW[26]), .D(n44), .Q(
        n57) );
  NAND31 U133 ( .A(n48), .B(n49), .C(n50), .Q(N51) );
  NAND22 U134 ( .A(i_data_lwM[29]), .B(n9), .Q(n49) );
  AOI221 U135 ( .A(i_data_rt[29]), .B(n43), .C(i_data_lwW[29]), .D(n44), .Q(
        n48) );
  NAND31 U136 ( .A(n45), .B(n46), .C(n47), .Q(N52) );
  NAND22 U137 ( .A(i_data_lwM[30]), .B(n9), .Q(n46) );
  AOI221 U138 ( .A(i_data_rt[30]), .B(n4), .C(i_data_lwW[30]), .D(n2), .Q(n45)
         );
  NAND31 U139 ( .A(n37), .B(n38), .C(n39), .Q(N53) );
  NAND22 U140 ( .A(i_data_lwM[31]), .B(n9), .Q(n38) );
  AOI221 U141 ( .A(i_data_rt[31]), .B(n4), .C(i_data_lwW[31]), .D(n2), .Q(n37)
         );
  INV3 U142 ( .A(n41), .Q(n5) );
  NOR31 U143 ( .A(i_con_fb[1]), .B(i_con_fb[2]), .C(n13), .Q(n41) );
  INV3 U144 ( .A(n43), .Q(n3) );
  NOR31 U145 ( .A(i_con_fb[1]), .B(i_con_fb[2]), .C(i_con_fb[0]), .Q(n43) );
  INV3 U146 ( .A(i_con_fb[0]), .Q(n13) );
  INV3 U147 ( .A(i_con_fb[2]), .Q(n10) );
  AOI221 U148 ( .A(i_data_alures[18]), .B(n7), .C(i_data_writeres[18]), .D(n41), .Q(n83) );
  LOGIC1 U149 ( .Q(n1) );
endmodule


module E_alubmux ( i_data_fb, i_data_imm, i_con_imm, o_data_alub );
  input [31:0] i_data_fb;
  input [31:0] i_data_imm;
  output [31:0] o_data_alub;
  input i_con_imm;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52;

  CLKIN6 U1 ( .A(n48), .Q(o_data_alub[9]) );
  CLKIN15 U2 ( .A(i_con_imm), .Q(n42) );
  INV3 U3 ( .A(i_data_fb[16]), .Q(n9) );
  INV3 U4 ( .A(i_data_imm[16]), .Q(n10) );
  NAND28 U5 ( .A(n17), .B(n18), .Q(n30) );
  CLKIN12 U6 ( .A(n11), .Q(o_data_alub[20]) );
  INV3 U7 ( .A(i_data_fb[13]), .Q(n13) );
  INV3 U8 ( .A(i_data_imm[13]), .Q(n14) );
  INV3 U9 ( .A(i_data_fb[0]), .Q(n24) );
  INV3 U10 ( .A(i_data_fb[23]), .Q(n4) );
  INV3 U11 ( .A(i_data_imm[23]), .Q(n5) );
  CLKIN3 U12 ( .A(i_data_imm[0]), .Q(n25) );
  INV3 U13 ( .A(i_data_fb[8]), .Q(n29) );
  INV3 U14 ( .A(i_data_imm[8]), .Q(n27) );
  INV2 U15 ( .A(n15), .Q(n1) );
  CLKIN12 U16 ( .A(n49), .Q(o_data_alub[10]) );
  CLKIN15 U17 ( .A(n39), .Q(n15) );
  CLKIN12 U18 ( .A(n52), .Q(o_data_alub[14]) );
  CLKIN8 U19 ( .A(n50), .Q(o_data_alub[11]) );
  CLKIN6 U20 ( .A(n47), .Q(o_data_alub[6]) );
  INV10 U21 ( .A(n44), .Q(o_data_alub[1]) );
  MUX26 U22 ( .A(n2), .B(n3), .S(n40), .Q(n33) );
  INV15 U23 ( .A(i_data_fb[4]), .Q(n2) );
  INV15 U24 ( .A(i_data_imm[4]), .Q(n3) );
  CLKIN4 U25 ( .A(i_data_imm[5]), .Q(n7) );
  IMUX23 U26 ( .A(n7), .B(n6), .S(n15), .Q(o_data_alub[5]) );
  IMUX21 U27 ( .A(n4), .B(n5), .S(n40), .Q(o_data_alub[23]) );
  INV15 U28 ( .A(i_data_fb[5]), .Q(n6) );
  INV2 U29 ( .A(n40), .Q(n38) );
  NAND24 U30 ( .A(n22), .B(n20), .Q(n18) );
  INV8 U31 ( .A(n28), .Q(n20) );
  BUF12 U32 ( .A(n35), .Q(o_data_alub[15]) );
  NAND24 U33 ( .A(n21), .B(n16), .Q(n17) );
  IMUX21 U34 ( .A(n9), .B(n10), .S(n39), .Q(o_data_alub[16]) );
  CLKIN15 U35 ( .A(n33), .Q(o_data_alub[4]) );
  MUX26 U36 ( .A(i_data_fb[30]), .B(i_data_imm[30]), .S(n20), .Q(
        o_data_alub[30]) );
  INV6 U37 ( .A(n45), .Q(o_data_alub[2]) );
  INV15 U38 ( .A(n43), .Q(o_data_alub[0]) );
  MUX24 U39 ( .A(i_data_fb[29]), .B(i_data_imm[29]), .S(n20), .Q(
        o_data_alub[29]) );
  IMUX22 U40 ( .A(i_data_fb[20]), .B(i_data_imm[20]), .S(n39), .Q(n11) );
  OAI222 U41 ( .A(n13), .B(n41), .C(n14), .D(n28), .Q(o_data_alub[13]) );
  CLKIN15 U42 ( .A(n40), .Q(n28) );
  INV2 U43 ( .A(n20), .Q(n16) );
  MUX22 U44 ( .A(i_data_fb[27]), .B(i_data_imm[27]), .S(n40), .Q(
        o_data_alub[27]) );
  INV8 U45 ( .A(n46), .Q(o_data_alub[3]) );
  INV15 U46 ( .A(n30), .Q(o_data_alub[17]) );
  MUX22 U47 ( .A(i_data_fb[26]), .B(i_data_imm[26]), .S(n40), .Q(
        o_data_alub[26]) );
  MUX24 U48 ( .A(i_data_fb[7]), .B(i_data_imm[7]), .S(n40), .Q(o_data_alub[7])
         );
  INV3 U49 ( .A(i_data_fb[17]), .Q(n21) );
  INV3 U50 ( .A(i_data_imm[17]), .Q(n22) );
  BUF12 U51 ( .A(n51), .Q(n19) );
  INV15 U52 ( .A(n34), .Q(n41) );
  AOI222 U53 ( .A(n39), .B(i_data_imm[2]), .C(n34), .D(i_data_fb[2]), .Q(n45)
         );
  AOI221 U54 ( .A(i_data_fb[6]), .B(n15), .C(n40), .D(i_data_imm[6]), .Q(n47)
         );
  MUX22 U55 ( .A(i_data_fb[25]), .B(i_data_imm[25]), .S(n40), .Q(
        o_data_alub[25]) );
  MUX22 U56 ( .A(i_data_fb[22]), .B(i_data_imm[22]), .S(n40), .Q(
        o_data_alub[22]) );
  INV15 U57 ( .A(n19), .Q(o_data_alub[12]) );
  MUX24 U58 ( .A(i_data_fb[28]), .B(i_data_imm[28]), .S(n41), .Q(
        o_data_alub[28]) );
  CLKIN6 U59 ( .A(n23), .Q(n43) );
  MUX24 U60 ( .A(i_data_fb[21]), .B(i_data_imm[21]), .S(n41), .Q(
        o_data_alub[21]) );
  MUX21 U61 ( .A(i_data_fb[31]), .B(i_data_imm[31]), .S(n41), .Q(
        o_data_alub[31]) );
  AOI222 U62 ( .A(i_data_fb[11]), .B(n28), .C(n40), .D(i_data_imm[11]), .Q(n50) );
  OAI221 U63 ( .A(n40), .B(n36), .C(n37), .D(n15), .Q(n35) );
  AOI222 U64 ( .A(n15), .B(i_data_fb[3]), .C(n41), .D(i_data_imm[3]), .Q(n46)
         );
  CLKIN15 U65 ( .A(n39), .Q(n34) );
  AOI221 U66 ( .A(n42), .B(i_data_fb[12]), .C(i_data_imm[12]), .D(n40), .Q(n51) );
  OAI222 U67 ( .A(n40), .B(n24), .C(n25), .D(n38), .Q(n23) );
  INV15 U68 ( .A(n42), .Q(n40) );
  OAI222 U69 ( .A(n27), .B(n28), .C(n29), .D(n40), .Q(o_data_alub[8]) );
  INV15 U70 ( .A(n42), .Q(n39) );
  INV3 U71 ( .A(i_data_fb[15]), .Q(n36) );
  INV3 U72 ( .A(i_data_imm[15]), .Q(n37) );
  MUX22 U73 ( .A(i_data_fb[24]), .B(i_data_imm[24]), .S(n40), .Q(
        o_data_alub[24]) );
  MUX24 U74 ( .A(i_data_fb[19]), .B(i_data_imm[19]), .S(n39), .Q(
        o_data_alub[19]) );
  MUX24 U75 ( .A(i_data_fb[18]), .B(i_data_imm[18]), .S(n41), .Q(
        o_data_alub[18]) );
  AOI222 U76 ( .A(n28), .B(i_data_fb[14]), .C(n1), .D(i_data_imm[14]), .Q(n52)
         );
  AOI222 U77 ( .A(i_data_fb[1]), .B(n15), .C(n40), .D(i_data_imm[1]), .Q(n44)
         );
  AOI222 U78 ( .A(i_data_fb[9]), .B(n15), .C(n40), .D(i_data_imm[9]), .Q(n48)
         );
  AOI222 U79 ( .A(n40), .B(i_data_imm[10]), .C(n28), .D(i_data_fb[10]), .Q(n49) );
endmodule


module E_rdmux ( i_data_rtE, i_data_rdE, i_con_regdst, i_con_aluPC4, 
        o_data_writeE );
  input [4:0] i_data_rtE;
  input [4:0] i_data_rdE;
  output [4:0] o_data_writeE;
  input i_con_regdst, i_con_aluPC4;
  wire   n7, n8, n9, n10, n11, n1, n2, n3, n4, n5, n6, n12;

  BUF6 U2 ( .A(i_con_regdst), .Q(n1) );
  OAI2111 U3 ( .A(n1), .B(n6), .C(n12), .D(n11), .Q(o_data_writeE[0]) );
  INV3 U4 ( .A(i_data_rtE[0]), .Q(n6) );
  NAND22 U5 ( .A(i_data_rdE[0]), .B(n1), .Q(n11) );
  OAI2111 U6 ( .A(n1), .B(n5), .C(n12), .D(n10), .Q(o_data_writeE[1]) );
  INV3 U7 ( .A(i_data_rtE[1]), .Q(n5) );
  NAND22 U8 ( .A(i_data_rdE[1]), .B(n1), .Q(n10) );
  OAI2111 U9 ( .A(n1), .B(n2), .C(n12), .D(n7), .Q(o_data_writeE[4]) );
  INV3 U10 ( .A(i_data_rtE[4]), .Q(n2) );
  NAND22 U11 ( .A(i_data_rdE[4]), .B(n1), .Q(n7) );
  OAI2111 U12 ( .A(n1), .B(n3), .C(n12), .D(n8), .Q(o_data_writeE[3]) );
  INV3 U13 ( .A(i_data_rtE[3]), .Q(n3) );
  NAND22 U14 ( .A(i_data_rdE[3]), .B(n1), .Q(n8) );
  OAI2111 U15 ( .A(n1), .B(n4), .C(n12), .D(n9), .Q(o_data_writeE[2]) );
  INV3 U16 ( .A(i_data_rtE[2]), .Q(n4) );
  NAND22 U17 ( .A(i_data_rdE[2]), .B(n1), .Q(n9) );
  INV3 U18 ( .A(i_con_aluPC4), .Q(n12) );
endmodule


module D_compare_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  INV3 U1 ( .A(NE), .Q(EQ) );
  INV3 U2 ( .A(n27), .Q(n2) );
  INV3 U3 ( .A(A[1]), .Q(n4) );
  INV3 U4 ( .A(B[0]), .Q(n3) );
  NAND20 U5 ( .A(n5), .B(n6), .Q(NE) );
  NOR40 U6 ( .A(n7), .B(n8), .C(n9), .D(n10), .Q(n6) );
  NAND40 U7 ( .A(n11), .B(n12), .C(n13), .D(n14), .Q(n10) );
  XNR20 U8 ( .A(B[11]), .B(A[11]), .Q(n14) );
  XNR20 U9 ( .A(B[12]), .B(A[12]), .Q(n13) );
  XNR20 U10 ( .A(B[13]), .B(A[13]), .Q(n12) );
  XNR20 U11 ( .A(B[14]), .B(A[14]), .Q(n11) );
  NAND40 U12 ( .A(n15), .B(n16), .C(n17), .D(n18), .Q(n9) );
  XNR20 U13 ( .A(B[7]), .B(A[7]), .Q(n18) );
  XNR20 U14 ( .A(B[8]), .B(A[8]), .Q(n17) );
  XNR20 U15 ( .A(B[9]), .B(A[9]), .Q(n16) );
  XNR20 U16 ( .A(B[10]), .B(A[10]), .Q(n15) );
  NAND40 U17 ( .A(n19), .B(n20), .C(n21), .D(n22), .Q(n8) );
  XNR20 U18 ( .A(B[3]), .B(A[3]), .Q(n22) );
  XNR20 U19 ( .A(B[4]), .B(A[4]), .Q(n21) );
  XNR20 U20 ( .A(B[5]), .B(A[5]), .Q(n20) );
  XNR20 U21 ( .A(B[6]), .B(A[6]), .Q(n19) );
  NAND40 U22 ( .A(n23), .B(n24), .C(n2), .D(n25), .Q(n7) );
  OAI220 U23 ( .A(n26), .B(n4), .C(B[1]), .D(n26), .Q(n25) );
  NOR20 U24 ( .A(n3), .B(A[0]), .Q(n26) );
  AOI220 U25 ( .A(n4), .B(n28), .C(n28), .D(B[1]), .Q(n27) );
  NAND20 U26 ( .A(A[0]), .B(n3), .Q(n28) );
  XNR20 U27 ( .A(B[31]), .B(A[31]), .Q(n24) );
  XNR20 U28 ( .A(B[2]), .B(A[2]), .Q(n23) );
  NOR40 U29 ( .A(n29), .B(n30), .C(n31), .D(n32), .Q(n5) );
  NAND40 U30 ( .A(n33), .B(n34), .C(n35), .D(n36), .Q(n32) );
  XNR20 U31 ( .A(B[27]), .B(A[27]), .Q(n36) );
  XNR20 U32 ( .A(B[28]), .B(A[28]), .Q(n35) );
  XNR20 U33 ( .A(B[29]), .B(A[29]), .Q(n34) );
  XNR20 U34 ( .A(B[30]), .B(A[30]), .Q(n33) );
  NAND40 U35 ( .A(n37), .B(n38), .C(n39), .D(n40), .Q(n31) );
  XNR20 U36 ( .A(B[23]), .B(A[23]), .Q(n40) );
  XNR20 U37 ( .A(B[24]), .B(A[24]), .Q(n39) );
  XNR20 U38 ( .A(B[25]), .B(A[25]), .Q(n38) );
  XNR20 U39 ( .A(B[26]), .B(A[26]), .Q(n37) );
  NAND40 U40 ( .A(n41), .B(n42), .C(n43), .D(n44), .Q(n30) );
  XNR20 U41 ( .A(B[19]), .B(A[19]), .Q(n44) );
  XNR20 U42 ( .A(B[20]), .B(A[20]), .Q(n43) );
  XNR20 U43 ( .A(B[21]), .B(A[21]), .Q(n42) );
  XNR20 U44 ( .A(B[22]), .B(A[22]), .Q(n41) );
  NAND40 U45 ( .A(n45), .B(n46), .C(n47), .D(n48), .Q(n29) );
  XNR20 U46 ( .A(B[15]), .B(A[15]), .Q(n48) );
  XNR20 U47 ( .A(B[16]), .B(A[16]), .Q(n47) );
  XNR20 U48 ( .A(B[17]), .B(A[17]), .Q(n46) );
  XNR20 U49 ( .A(B[18]), .B(A[18]), .Q(n45) );
endmodule


module D_compare ( o_con_ifbranch, i_data_rs, i_data_rt, i_con_bop );
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [2:0] i_con_bop;
  output o_con_ifbranch;
  wire   N32, N33, n4, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n1, n2, n3, n5, n6;

  D_compare_DW01_cmp6_0 r49 ( .A(i_data_rs), .B(i_data_rt), .TC(n4), .EQ(N32), 
        .NE(N33) );
  CLKIN3 U2 ( .A(i_con_bop[2]), .Q(n3) );
  AOI211 U3 ( .A(n15), .B(n5), .C(n3), .Q(n12) );
  INV3 U4 ( .A(n15), .Q(n2) );
  OAI311 U5 ( .A(n5), .B(i_con_bop[2]), .C(n10), .D(n11), .Q(o_con_ifbranch)
         );
  AOI211 U6 ( .A(N33), .B(n6), .C(n16), .Q(n10) );
  AOI311 U7 ( .A(n6), .B(n1), .C(n12), .D(n13), .Q(n11) );
  AOI211 U8 ( .A(n1), .B(n2), .C(n6), .Q(n16) );
  INV3 U9 ( .A(i_con_bop[0]), .Q(n6) );
  NOR31 U10 ( .A(n6), .B(i_con_bop[1]), .C(n14), .Q(n13) );
  AOI221 U11 ( .A(N32), .B(n3), .C(i_data_rs[31]), .D(i_con_bop[2]), .Q(n14)
         );
  INV3 U12 ( .A(i_con_bop[1]), .Q(n5) );
  NOR40 U13 ( .A(i_data_rs[9]), .B(i_data_rs[8]), .C(i_data_rs[7]), .D(
        i_data_rs[6]), .Q(n26) );
  NOR40 U14 ( .A(i_data_rs[26]), .B(i_data_rs[25]), .C(i_data_rs[24]), .D(
        i_data_rs[23]), .Q(n23) );
  NOR40 U15 ( .A(i_data_rs[5]), .B(i_data_rs[4]), .C(i_data_rs[3]), .D(
        i_data_rs[30]), .Q(n25) );
  NOR40 U16 ( .A(i_data_rs[15]), .B(i_data_rs[14]), .C(i_data_rs[13]), .D(
        i_data_rs[12]), .Q(n20) );
  NOR40 U17 ( .A(i_data_rs[22]), .B(i_data_rs[21]), .C(i_data_rs[20]), .D(
        i_data_rs[1]), .Q(n22) );
  NOR40 U18 ( .A(i_data_rs[19]), .B(i_data_rs[18]), .C(i_data_rs[17]), .D(
        i_data_rs[16]), .Q(n21) );
  NOR40 U19 ( .A(i_data_rs[2]), .B(i_data_rs[29]), .C(i_data_rs[28]), .D(
        i_data_rs[27]), .Q(n24) );
  NOR21 U20 ( .A(n17), .B(n18), .Q(n15) );
  NAND41 U21 ( .A(n19), .B(n20), .C(n21), .D(n22), .Q(n18) );
  NAND41 U22 ( .A(n23), .B(n24), .C(n25), .D(n26), .Q(n17) );
  NOR31 U23 ( .A(i_data_rs[0]), .B(i_data_rs[11]), .C(i_data_rs[10]), .Q(n19)
         );
  INV3 U24 ( .A(i_data_rs[31]), .Q(n1) );
  LOGIC0 U25 ( .Q(n4) );
endmodule


module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Ealuop, i_con_Ealusrc, 
        i_con_Eregdst, i_con_Mmemread, i_con_Mmemwrite, i_con_Wloadmux, 
        i_con_Walupc8, i_con_Wmemtoreg, i_con_Wregwrite, i_con_Efamux, 
        i_con_Efbmux, i_con_bop, o_data_pc4, o_data_alures, o_data_rt, 
        o_addr_regdst, o_con_Mmemread, o_con_Mmemwrite, o_con_Wloadmux, 
        o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_addr_Erd, 
        o_addr_Mrt, o_FaluresE, o_con_ifbranch );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [5:0] i_con_Ealuop;
  input [1:0] i_con_Wloadmux;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [2:0] i_con_bop;
  output [31:0] o_data_pc4;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [1:0] o_con_Wloadmux;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  output [31:0] o_FaluresE;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Walupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Walupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;

  DFC3 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[0]) );
  DFC3 pipe_alures_reg_13_ ( .D(o_FaluresE[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[13]) );
  DFC3 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC3 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC3 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC3 pipe_rt_reg_28_ ( .D(compare_i_data_rt[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[28]) );
  DFC3 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  DFC3 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC3 pipe_rt_reg_25_ ( .D(compare_i_data_rt[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[25]) );
  DFC3 pipe_rt_reg_24_ ( .D(compare_i_data_rt[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[24]) );
  DFC3 pipe_rt_reg_23_ ( .D(compare_i_data_rt[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[23]) );
  DFC3 pipe_rt_reg_22_ ( .D(compare_i_data_rt[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[22]) );
  DFC3 pipe_rt_reg_21_ ( .D(compare_i_data_rt[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[21]) );
  DFC3 pipe_rt_reg_20_ ( .D(compare_i_data_rt[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[20]) );
  DFC3 pipe_rt_reg_19_ ( .D(compare_i_data_rt[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[19]) );
  DFC3 pipe_rt_reg_18_ ( .D(compare_i_data_rt[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[18]) );
  DFC3 pipe_rt_reg_17_ ( .D(compare_i_data_rt[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[17]) );
  DFC3 pipe_rt_reg_16_ ( .D(compare_i_data_rt[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[16]) );
  DFC3 pipe_rt_reg_15_ ( .D(compare_i_data_rt[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[15]) );
  DFC3 pipe_rt_reg_14_ ( .D(compare_i_data_rt[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[14]) );
  DFC3 pipe_rt_reg_13_ ( .D(compare_i_data_rt[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[13]) );
  DFC3 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC3 pipe_rt_reg_11_ ( .D(compare_i_data_rt[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[11]) );
  DFC3 pipe_rt_reg_10_ ( .D(compare_i_data_rt[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[10]) );
  DFC3 pipe_rt_reg_9_ ( .D(compare_i_data_rt[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[9]) );
  DFC3 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC3 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC3 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC3 pipe_rt_reg_5_ ( .D(compare_i_data_rt[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[5]) );
  DFC3 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(compare_i_data_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[2]) );
  DFC3 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC3 pipe_rt_reg_0_ ( .D(compare_i_data_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[0]) );
  DFC3 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wloadmux_reg_1_ ( .D(i_con_Wloadmux[1]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[1]) );
  DFC3 pipe_con_Wloadmux_reg_0_ ( .D(i_con_Wloadmux[0]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[0]) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  E_alu u_alu ( .o_data_AluRes(o_FaluresE), .i_data_A(compare_i_data_rs), 
        .i_data_B({alu_i_data_B[31:30], n6, alu_i_data_B[28:27], n9, 
        alu_i_data_B[25:14], n3, alu_i_data_B[12:9], n10, alu_i_data_B[7:0]}), 
        .i_con_AluCtrl(alu_i_con_AluCtrl), .i_data_shamt({i_data_immext[10:7], 
        n5}) );
  E_alu_control u_alu_control ( .o_con_AluCtrl(alu_i_con_AluCtrl), 
        .i_con_AluOp(i_con_Ealuop), .i_con_FuncCode(i_data_immext[5:0]) );
  E_famux5 u_famux5 ( .i_data_rs(i_data_rs), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fa(i_con_Efamux), .o_data_alusra(
        compare_i_data_rs) );
  E_fbmux5 u_fbmux ( .i_data_rt(i_data_rt), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fb(i_con_Efbmux), .o_data_alusrb(
        compare_i_data_rt) );
  E_alubmux u_alubmux ( .i_data_fb(compare_i_data_rt), .i_data_imm({
        i_data_immext[31:7], n5, n1, i_data_immext[4], n2, i_data_immext[2], 
        n8, n7}), .i_con_imm(i_con_Ealusrc), .o_data_alub(alu_i_data_B) );
  E_rdmux u_rdmux ( .i_data_rtE(i_addr_rt), .i_data_rdE(i_addr_rd), 
        .i_con_regdst(i_con_Eregdst), .i_con_aluPC4(i_con_Walupc8), 
        .o_data_writeE(o_addr_Erd) );
  D_compare u_compare ( .o_con_ifbranch(o_con_ifbranch), .i_data_rs(
        compare_i_data_rs), .i_data_rt(compare_i_data_rt), .i_con_bop(
        i_con_bop) );
  DFC1 pipe_alures_reg_16_ ( .D(o_FaluresE[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[16]) );
  DFC1 pipe_alures_reg_25_ ( .D(o_FaluresE[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[25]) );
  DFC1 pipe_alures_reg_28_ ( .D(o_FaluresE[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[28]) );
  DFC1 pipe_alures_reg_14_ ( .D(o_FaluresE[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[14]) );
  DFC1 pipe_alures_reg_27_ ( .D(o_FaluresE[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[27]) );
  DFC1 pipe_alures_reg_23_ ( .D(o_FaluresE[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[23]) );
  DFC1 pipe_alures_reg_18_ ( .D(o_FaluresE[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[18]) );
  DFC1 pipe_alures_reg_26_ ( .D(o_FaluresE[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[26]) );
  DFC1 pipe_alures_reg_24_ ( .D(o_FaluresE[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[24]) );
  DFC1 pipe_alures_reg_21_ ( .D(o_FaluresE[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[21]) );
  DFC1 pipe_alures_reg_20_ ( .D(o_FaluresE[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[20]) );
  DFC1 pipe_alures_reg_15_ ( .D(o_FaluresE[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[15]) );
  DFC1 pipe_alures_reg_11_ ( .D(o_FaluresE[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[11]) );
  DFC1 pipe_alures_reg_7_ ( .D(o_FaluresE[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[7]) );
  DFC1 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC1 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC1 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC1 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC1 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC1 pipe_alures_reg_30_ ( .D(o_FaluresE[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[30]) );
  DFC1 pipe_alures_reg_29_ ( .D(o_FaluresE[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[29]) );
  DFC1 pipe_alures_reg_22_ ( .D(o_FaluresE[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[22]) );
  DFC1 pipe_alures_reg_19_ ( .D(o_FaluresE[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[19]) );
  DFC1 pipe_alures_reg_17_ ( .D(o_FaluresE[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[17]) );
  DFC1 pipe_alures_reg_10_ ( .D(o_FaluresE[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[10]) );
  DFC1 pipe_alures_reg_5_ ( .D(o_FaluresE[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[5]) );
  DFC1 pipe_alures_reg_2_ ( .D(o_FaluresE[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[2]) );
  DFC1 pipe_alures_reg_1_ ( .D(o_FaluresE[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[1]) );
  DFC1 pipe_alures_reg_0_ ( .D(o_FaluresE[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[0]) );
  DFC1 pipe_con_Walupc8_reg ( .D(i_con_Walupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Walupc8) );
  DFC1 pipe_alures_reg_9_ ( .D(o_FaluresE[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[9]) );
  DFC1 pipe_alures_reg_3_ ( .D(o_FaluresE[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[3]) );
  DFC1 pipe_alures_reg_6_ ( .D(o_FaluresE[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[6]) );
  DFC1 pipe_alures_reg_8_ ( .D(o_FaluresE[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[8]) );
  DFC1 pipe_alures_reg_4_ ( .D(o_FaluresE[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[4]) );
  DFC1 pipe_alures_reg_12_ ( .D(o_FaluresE[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[12]) );
  DFC1 pipe_alures_reg_31_ ( .D(o_FaluresE[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[31]) );
  INV12 U3 ( .A(n4), .Q(n5) );
  BUF6 U4 ( .A(i_data_immext[3]), .Q(n2) );
  BUF4 U5 ( .A(i_data_immext[0]), .Q(n7) );
  BUF2 U6 ( .A(i_data_immext[1]), .Q(n8) );
  BUF2 U7 ( .A(i_data_immext[5]), .Q(n1) );
  BUF15 U8 ( .A(alu_i_data_B[29]), .Q(n6) );
  BUF15 U9 ( .A(alu_i_data_B[13]), .Q(n3) );
  CLKIN6 U10 ( .A(i_data_immext[6]), .Q(n4) );
  BUF15 U11 ( .A(alu_i_data_B[8]), .Q(n10) );
  BUF15 U12 ( .A(alu_i_data_B[26]), .Q(n9) );
endmodule


module mem_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  NAND22 U2 ( .A(A[8]), .B(n2), .Q(n1) );
  NAND22 U3 ( .A(n71), .B(n2), .Q(n87) );
  NAND22 U4 ( .A(n81), .B(A[13]), .Q(n82) );
  NOR21 U5 ( .A(n41), .B(n68), .Q(n69) );
  NOR21 U6 ( .A(n41), .B(n54), .Q(n55) );
  NAND22 U7 ( .A(n19), .B(n21), .Q(n20) );
  INV3 U8 ( .A(n29), .Q(n53) );
  INV3 U9 ( .A(n85), .Q(n2) );
  NAND41 U10 ( .A(n96), .B(n70), .C(n71), .D(n72), .Q(n29) );
  NOR31 U11 ( .A(n73), .B(n74), .C(n75), .Q(n72) );
  NOR31 U12 ( .A(SUM[2]), .B(n14), .C(n76), .Q(n70) );
  XNR21 U13 ( .A(n69), .B(n61), .Q(SUM[17]) );
  XOR21 U14 ( .A(n66), .B(A[18]), .Q(SUM[18]) );
  NOR21 U15 ( .A(n41), .B(n67), .Q(n66) );
  INV3 U16 ( .A(n65), .Q(n67) );
  XNR21 U17 ( .A(n55), .B(n45), .Q(SUM[21]) );
  INV3 U18 ( .A(n25), .Q(n21) );
  NAND31 U19 ( .A(n26), .B(n53), .C(n27), .Q(n25) );
  NOR21 U20 ( .A(n30), .B(n31), .Q(n26) );
  INV3 U21 ( .A(n28), .Q(n27) );
  NOR21 U22 ( .A(n61), .B(n68), .Q(n65) );
  XNR21 U23 ( .A(n92), .B(n89), .Q(SUM[10]) );
  XNR21 U24 ( .A(n81), .B(n73), .Q(SUM[13]) );
  XOR21 U25 ( .A(n51), .B(A[22]), .Q(SUM[22]) );
  NOR21 U26 ( .A(n45), .B(n52), .Q(n51) );
  NAND22 U27 ( .A(n49), .B(n53), .Q(n52) );
  XNR21 U28 ( .A(n9), .B(n10), .Q(SUM[5]) );
  XNR21 U29 ( .A(n6), .B(n7), .Q(SUM[6]) );
  XOR21 U30 ( .A(n36), .B(n33), .Q(SUM[25]) );
  XOR21 U31 ( .A(A[26]), .B(n37), .Q(SUM[26]) );
  NOR21 U32 ( .A(n85), .B(n93), .Q(n92) );
  INV3 U33 ( .A(n94), .Q(n93) );
  NOR21 U34 ( .A(n4), .B(n3), .Q(n94) );
  XNR21 U35 ( .A(A[9]), .B(n1), .Q(SUM[9]) );
  XNR21 U36 ( .A(A[14]), .B(n82), .Q(SUM[14]) );
  INV3 U37 ( .A(n83), .Q(n81) );
  NAND22 U38 ( .A(n84), .B(n2), .Q(n83) );
  NOR21 U39 ( .A(n74), .B(n86), .Q(n84) );
  NAND22 U40 ( .A(n95), .B(n96), .Q(n85) );
  NOR21 U41 ( .A(n14), .B(SUM[2]), .Q(n95) );
  NOR21 U42 ( .A(n36), .B(n33), .Q(n37) );
  INV3 U43 ( .A(n11), .Q(n9) );
  NAND22 U44 ( .A(n12), .B(A[2]), .Q(n11) );
  NOR21 U45 ( .A(n13), .B(n14), .Q(n12) );
  INV3 U46 ( .A(n8), .Q(n6) );
  NAND22 U47 ( .A(n9), .B(A[5]), .Q(n8) );
  INV3 U48 ( .A(n71), .Q(n86) );
  INV3 U49 ( .A(n32), .Q(n31) );
  NOR21 U50 ( .A(n33), .B(n34), .Q(n32) );
  NOR21 U51 ( .A(n73), .B(n75), .Q(n80) );
  NOR31 U52 ( .A(n89), .B(n88), .C(n4), .Q(n71) );
  NAND22 U53 ( .A(A[11]), .B(A[8]), .Q(n88) );
  NAND22 U54 ( .A(n42), .B(n43), .Q(n28) );
  NOR31 U55 ( .A(n46), .B(n44), .C(n45), .Q(n42) );
  NAND22 U56 ( .A(A[23]), .B(A[20]), .Q(n44) );
  INV3 U57 ( .A(A[3]), .Q(n14) );
  INV3 U58 ( .A(A[2]), .Q(SUM[2]) );
  INV3 U59 ( .A(A[13]), .Q(n73) );
  NAND22 U60 ( .A(n58), .B(n59), .Q(n56) );
  NOR21 U61 ( .A(n61), .B(n62), .Q(n58) );
  INV3 U62 ( .A(n60), .Q(n59) );
  NAND22 U63 ( .A(A[19]), .B(A[16]), .Q(n60) );
  NAND22 U64 ( .A(n97), .B(n98), .Q(n77) );
  NOR21 U65 ( .A(n99), .B(n13), .Q(n97) );
  NOR21 U66 ( .A(n10), .B(n7), .Q(n98) );
  INV3 U67 ( .A(A[7]), .Q(n99) );
  INV3 U68 ( .A(A[10]), .Q(n89) );
  INV3 U69 ( .A(A[17]), .Q(n61) );
  INV3 U70 ( .A(A[18]), .Q(n62) );
  INV3 U71 ( .A(A[9]), .Q(n4) );
  INV3 U72 ( .A(A[14]), .Q(n75) );
  XOR21 U73 ( .A(n57), .B(A[20]), .Q(SUM[20]) );
  NOR21 U74 ( .A(n41), .B(n56), .Q(n57) );
  XOR21 U75 ( .A(n40), .B(A[24]), .Q(SUM[24]) );
  NOR21 U76 ( .A(n41), .B(n28), .Q(n40) );
  XOR21 U77 ( .A(n24), .B(A[29]), .Q(SUM[29]) );
  NOR21 U78 ( .A(n25), .B(n22), .Q(n24) );
  XOR21 U79 ( .A(n17), .B(A[31]), .Q(SUM[31]) );
  NOR21 U80 ( .A(n25), .B(n18), .Q(n17) );
  NAND22 U81 ( .A(A[30]), .B(n19), .Q(n18) );
  XOR21 U82 ( .A(n47), .B(n48), .Q(SUM[23]) );
  INV3 U83 ( .A(A[23]), .Q(n47) );
  NAND31 U84 ( .A(n50), .B(n53), .C(n49), .Q(n48) );
  NOR21 U85 ( .A(n45), .B(n46), .Q(n50) );
  INV3 U86 ( .A(A[5]), .Q(n10) );
  INV3 U87 ( .A(A[6]), .Q(n7) );
  INV3 U88 ( .A(A[12]), .Q(n74) );
  INV3 U89 ( .A(A[4]), .Q(n13) );
  INV3 U90 ( .A(A[15]), .Q(n76) );
  INV3 U91 ( .A(A[21]), .Q(n45) );
  INV3 U92 ( .A(A[25]), .Q(n33) );
  NAND22 U93 ( .A(A[20]), .B(n43), .Q(n54) );
  INV3 U94 ( .A(A[22]), .Q(n46) );
  INV3 U95 ( .A(A[26]), .Q(n34) );
  XOR21 U96 ( .A(n53), .B(A[16]), .Q(SUM[16]) );
  XOR21 U97 ( .A(n2), .B(A[8]), .Q(SUM[8]) );
  XOR21 U98 ( .A(n21), .B(A[28]), .Q(SUM[28]) );
  XOR21 U99 ( .A(n63), .B(A[19]), .Q(SUM[19]) );
  NOR21 U100 ( .A(n62), .B(n64), .Q(n63) );
  NAND22 U101 ( .A(n65), .B(n53), .Q(n64) );
  XOR21 U102 ( .A(n78), .B(A[15]), .Q(SUM[15]) );
  NOR21 U103 ( .A(n83), .B(n79), .Q(n78) );
  INV3 U104 ( .A(n80), .Q(n79) );
  XOR21 U105 ( .A(A[27]), .B(n35), .Q(SUM[27]) );
  NOR31 U106 ( .A(n34), .B(n36), .C(n33), .Q(n35) );
  XNR21 U107 ( .A(A[30]), .B(n20), .Q(SUM[30]) );
  NAND22 U108 ( .A(A[27]), .B(A[24]), .Q(n30) );
  XNR21 U109 ( .A(A[12]), .B(n87), .Q(SUM[12]) );
  INV3 U110 ( .A(A[16]), .Q(n68) );
  XOR21 U111 ( .A(n90), .B(n91), .Q(SUM[11]) );
  INV3 U112 ( .A(A[11]), .Q(n90) );
  NAND22 U113 ( .A(n92), .B(A[10]), .Q(n91) );
  XOR21 U114 ( .A(n99), .B(n5), .Q(SUM[7]) );
  NAND22 U115 ( .A(n6), .B(A[6]), .Q(n5) );
  INV3 U116 ( .A(A[8]), .Q(n3) );
  NAND22 U117 ( .A(n38), .B(n53), .Q(n36) );
  NOR21 U118 ( .A(n39), .B(n28), .Q(n38) );
  INV3 U119 ( .A(A[24]), .Q(n39) );
  NOR21 U120 ( .A(n22), .B(n23), .Q(n19) );
  INV3 U121 ( .A(A[29]), .Q(n23) );
  XOR21 U122 ( .A(A[4]), .B(n15), .Q(SUM[4]) );
  NOR21 U123 ( .A(SUM[2]), .B(n14), .Q(n15) );
  INV3 U124 ( .A(A[28]), .Q(n22) );
  XOR21 U125 ( .A(A[3]), .B(A[2]), .Q(SUM[3]) );
  CLKIN3 U126 ( .A(n54), .Q(n49) );
  CLKIN3 U127 ( .A(n56), .Q(n43) );
  CLKIN3 U128 ( .A(n53), .Q(n41) );
  CLKIN3 U129 ( .A(n77), .Q(n96) );
endmodule


module mem ( i_clk, i_nrst, i_data_pc4, i_data_alures, i_data_memout, 
        i_addr_regdst, i_con_Wloadmux, i_con_Walupc8, i_con_Wmemtoreg, 
        i_con_Wregwrite, i_con_FWmemread, i_addr_Mrt, o_data_pc8, 
        o_data_alures, o_data_memout, o_addr_regdst, o_con_Wloadmux, 
        o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread, 
        o_addr_Wrt );
  input [31:0] i_data_pc4;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [4:0] i_addr_regdst;
  input [1:0] i_con_Wloadmux;
  input [4:0] i_addr_Mrt;
  output [31:0] o_data_pc8;
  output [31:0] o_data_alures;
  output [31:0] o_data_memout;
  output [4:0] o_addr_regdst;
  output [1:0] o_con_Wloadmux;
  output [4:0] o_addr_Wrt;
  input i_clk, i_nrst, i_con_Walupc8, i_con_Wmemtoreg, i_con_Wregwrite,
         i_con_FWmemread;
  output o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread;
  wire   n_Logic1_, n_Logic0_;
  wire   [31:0] pc8;

  DFC3 pipe_rt_reg_4_ ( .D(i_addr_Mrt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(i_addr_Mrt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(i_addr_Mrt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[2]) );
  DFC3 pipe_rt_reg_1_ ( .D(i_addr_Mrt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[1]) );
  DFC3 pipe_rt_reg_0_ ( .D(i_addr_Mrt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[0]) );
  DFC3 pipe_data_pc8_reg_31_ ( .D(pc8[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[31]) );
  DFC3 pipe_data_pc8_reg_30_ ( .D(pc8[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[30]) );
  DFC3 pipe_data_pc8_reg_29_ ( .D(pc8[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[29]) );
  DFC3 pipe_data_pc8_reg_28_ ( .D(pc8[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[28]) );
  DFC3 pipe_data_pc8_reg_27_ ( .D(pc8[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[27]) );
  DFC3 pipe_data_pc8_reg_26_ ( .D(pc8[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[26]) );
  DFC3 pipe_data_pc8_reg_25_ ( .D(pc8[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[25]) );
  DFC3 pipe_data_pc8_reg_24_ ( .D(pc8[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[24]) );
  DFC3 pipe_data_pc8_reg_23_ ( .D(pc8[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[23]) );
  DFC3 pipe_data_pc8_reg_22_ ( .D(pc8[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[22]) );
  DFC3 pipe_data_pc8_reg_21_ ( .D(pc8[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[21]) );
  DFC3 pipe_data_pc8_reg_20_ ( .D(pc8[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[20]) );
  DFC3 pipe_data_pc8_reg_19_ ( .D(pc8[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[19]) );
  DFC3 pipe_data_pc8_reg_18_ ( .D(pc8[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[18]) );
  DFC3 pipe_data_pc8_reg_17_ ( .D(pc8[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[17]) );
  DFC3 pipe_data_pc8_reg_16_ ( .D(pc8[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[16]) );
  DFC3 pipe_data_pc8_reg_15_ ( .D(pc8[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[15]) );
  DFC3 pipe_data_pc8_reg_14_ ( .D(pc8[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[14]) );
  DFC3 pipe_data_pc8_reg_13_ ( .D(pc8[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[13]) );
  DFC3 pipe_data_pc8_reg_12_ ( .D(pc8[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[12]) );
  DFC3 pipe_data_pc8_reg_11_ ( .D(pc8[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[11]) );
  DFC3 pipe_data_pc8_reg_10_ ( .D(pc8[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[10]) );
  DFC3 pipe_data_pc8_reg_9_ ( .D(pc8[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[9]) );
  DFC3 pipe_data_pc8_reg_8_ ( .D(pc8[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[8]) );
  DFC3 pipe_data_pc8_reg_7_ ( .D(pc8[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[7]) );
  DFC3 pipe_data_pc8_reg_6_ ( .D(pc8[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[6]) );
  DFC3 pipe_data_pc8_reg_5_ ( .D(pc8[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[5]) );
  DFC3 pipe_data_pc8_reg_4_ ( .D(pc8[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[4]) );
  DFC3 pipe_data_pc8_reg_3_ ( .D(pc8[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[3]) );
  DFC3 pipe_data_pc8_reg_2_ ( .D(pc8[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[2]) );
  DFC3 pipe_data_pc8_reg_1_ ( .D(pc8[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[1]) );
  DFC3 pipe_data_pc8_reg_0_ ( .D(pc8[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[0]) );
  DFC3 pipe_data_alures_reg_31_ ( .D(i_data_alures[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[31]) );
  DFC3 pipe_data_alures_reg_30_ ( .D(i_data_alures[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[30]) );
  DFC3 pipe_data_alures_reg_29_ ( .D(i_data_alures[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[29]) );
  DFC3 pipe_data_alures_reg_28_ ( .D(i_data_alures[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[28]) );
  DFC3 pipe_data_alures_reg_27_ ( .D(i_data_alures[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[27]) );
  DFC3 pipe_data_alures_reg_26_ ( .D(i_data_alures[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[26]) );
  DFC3 pipe_data_alures_reg_25_ ( .D(i_data_alures[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[25]) );
  DFC3 pipe_data_alures_reg_24_ ( .D(i_data_alures[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[24]) );
  DFC3 pipe_data_alures_reg_23_ ( .D(i_data_alures[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[23]) );
  DFC3 pipe_data_alures_reg_22_ ( .D(i_data_alures[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[22]) );
  DFC3 pipe_data_alures_reg_21_ ( .D(i_data_alures[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[21]) );
  DFC3 pipe_data_alures_reg_20_ ( .D(i_data_alures[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[20]) );
  DFC3 pipe_data_alures_reg_19_ ( .D(i_data_alures[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[19]) );
  DFC3 pipe_data_alures_reg_18_ ( .D(i_data_alures[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[18]) );
  DFC3 pipe_data_alures_reg_17_ ( .D(i_data_alures[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[17]) );
  DFC3 pipe_data_alures_reg_16_ ( .D(i_data_alures[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[16]) );
  DFC3 pipe_data_alures_reg_15_ ( .D(i_data_alures[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[15]) );
  DFC3 pipe_data_alures_reg_14_ ( .D(i_data_alures[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[14]) );
  DFC3 pipe_data_alures_reg_13_ ( .D(i_data_alures[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[13]) );
  DFC3 pipe_data_alures_reg_12_ ( .D(i_data_alures[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[12]) );
  DFC3 pipe_data_alures_reg_11_ ( .D(i_data_alures[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[11]) );
  DFC3 pipe_data_alures_reg_10_ ( .D(i_data_alures[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[10]) );
  DFC3 pipe_data_alures_reg_9_ ( .D(i_data_alures[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC3 pipe_data_alures_reg_8_ ( .D(i_data_alures[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC3 pipe_data_alures_reg_7_ ( .D(i_data_alures[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC3 pipe_data_alures_reg_6_ ( .D(i_data_alures[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC3 pipe_data_alures_reg_5_ ( .D(i_data_alures[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC3 pipe_data_alures_reg_4_ ( .D(i_data_alures[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC3 pipe_data_alures_reg_3_ ( .D(i_data_alures[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC3 pipe_data_alures_reg_2_ ( .D(i_data_alures[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC3 pipe_data_alures_reg_1_ ( .D(i_data_alures[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC3 pipe_data_alures_reg_0_ ( .D(i_data_alures[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC3 pipe_data_memout_reg_31_ ( .D(i_data_memout[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[31]) );
  DFC3 pipe_data_memout_reg_30_ ( .D(i_data_memout[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[30]) );
  DFC3 pipe_data_memout_reg_29_ ( .D(i_data_memout[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[29]) );
  DFC3 pipe_data_memout_reg_28_ ( .D(i_data_memout[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[28]) );
  DFC3 pipe_data_memout_reg_27_ ( .D(i_data_memout[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[27]) );
  DFC3 pipe_data_memout_reg_26_ ( .D(i_data_memout[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[26]) );
  DFC3 pipe_data_memout_reg_25_ ( .D(i_data_memout[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[25]) );
  DFC3 pipe_data_memout_reg_24_ ( .D(i_data_memout[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[24]) );
  DFC3 pipe_data_memout_reg_23_ ( .D(i_data_memout[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[23]) );
  DFC3 pipe_data_memout_reg_22_ ( .D(i_data_memout[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[22]) );
  DFC3 pipe_data_memout_reg_21_ ( .D(i_data_memout[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[21]) );
  DFC3 pipe_data_memout_reg_20_ ( .D(i_data_memout[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[20]) );
  DFC3 pipe_data_memout_reg_19_ ( .D(i_data_memout[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[19]) );
  DFC3 pipe_data_memout_reg_18_ ( .D(i_data_memout[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[18]) );
  DFC3 pipe_data_memout_reg_17_ ( .D(i_data_memout[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[17]) );
  DFC3 pipe_data_memout_reg_16_ ( .D(i_data_memout[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[16]) );
  DFC3 pipe_data_memout_reg_15_ ( .D(i_data_memout[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[15]) );
  DFC3 pipe_data_memout_reg_14_ ( .D(i_data_memout[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[14]) );
  DFC3 pipe_data_memout_reg_13_ ( .D(i_data_memout[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[13]) );
  DFC3 pipe_data_memout_reg_12_ ( .D(i_data_memout[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[12]) );
  DFC3 pipe_data_memout_reg_11_ ( .D(i_data_memout[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[11]) );
  DFC3 pipe_data_memout_reg_10_ ( .D(i_data_memout[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[10]) );
  DFC3 pipe_data_memout_reg_9_ ( .D(i_data_memout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[9]) );
  DFC3 pipe_data_memout_reg_8_ ( .D(i_data_memout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[8]) );
  DFC3 pipe_data_memout_reg_7_ ( .D(i_data_memout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[7]) );
  DFC3 pipe_data_memout_reg_6_ ( .D(i_data_memout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[6]) );
  DFC3 pipe_data_memout_reg_5_ ( .D(i_data_memout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[5]) );
  DFC3 pipe_data_memout_reg_4_ ( .D(i_data_memout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[4]) );
  DFC3 pipe_data_memout_reg_3_ ( .D(i_data_memout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[3]) );
  DFC3 pipe_data_memout_reg_2_ ( .D(i_data_memout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[2]) );
  DFC3 pipe_data_memout_reg_1_ ( .D(i_data_memout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[1]) );
  DFC3 pipe_data_memout_reg_0_ ( .D(i_data_memout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[0]) );
  DFC3 pipe_addr_regdst_reg_4_ ( .D(i_addr_regdst[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[4]) );
  DFC3 pipe_addr_regdst_reg_3_ ( .D(i_addr_regdst[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[3]) );
  DFC3 pipe_addr_regdst_reg_2_ ( .D(i_addr_regdst[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[2]) );
  DFC3 pipe_addr_regdst_reg_1_ ( .D(i_addr_regdst[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[1]) );
  DFC3 pipe_addr_regdst_reg_0_ ( .D(i_addr_regdst[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[0]) );
  DFC3 pipe_con_Wloadmux_reg_1_ ( .D(i_con_Wloadmux[1]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[1]) );
  DFC3 pipe_con_Wloadmux_reg_0_ ( .D(i_con_Wloadmux[0]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[0]) );
  DFC3 pipe_con_Walupc8_reg ( .D(i_con_Walupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Walupc8) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_con_FWmemread_reg ( .D(i_con_FWmemread), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_FWmemread) );
  mem_DW01_add_1 add_31 ( .A(i_data_pc4), .B({n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic1_, n_Logic0_, n_Logic0_}), .CI(n_Logic0_), .SUM(pc8) );
  LOGIC0 U3 ( .Q(n_Logic0_) );
  LOGIC1 U4 ( .Q(n_Logic1_) );
endmodule


module W_resmux ( i_data_alures, i_data_pc8, i_con_pc8, o_data_alu );
  input [31:0] i_data_alures;
  input [31:0] i_data_pc8;
  output [31:0] o_data_alu;
  input i_con_pc8;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n1, n2, n3, n4, n5, n6, n7;

  CLKIN3 U1 ( .A(n35), .Q(o_data_alu[8]) );
  CLKIN3 U2 ( .A(n34), .Q(o_data_alu[9]) );
  CLKIN3 U3 ( .A(n36), .Q(o_data_alu[7]) );
  INV3 U4 ( .A(n7), .Q(n1) );
  INV3 U5 ( .A(n7), .Q(n2) );
  INV3 U6 ( .A(n65), .Q(o_data_alu[0]) );
  INV3 U7 ( .A(n54), .Q(o_data_alu[1]) );
  INV3 U8 ( .A(n43), .Q(o_data_alu[2]) );
  INV3 U9 ( .A(n40), .Q(o_data_alu[3]) );
  INV3 U10 ( .A(n58), .Q(o_data_alu[16]) );
  INV3 U11 ( .A(n57), .Q(o_data_alu[17]) );
  INV3 U12 ( .A(n55), .Q(o_data_alu[19]) );
  INV3 U13 ( .A(n53), .Q(o_data_alu[20]) );
  INV3 U14 ( .A(n52), .Q(o_data_alu[21]) );
  INV3 U15 ( .A(n51), .Q(o_data_alu[22]) );
  INV3 U16 ( .A(n50), .Q(o_data_alu[23]) );
  INV3 U17 ( .A(n49), .Q(o_data_alu[24]) );
  INV3 U18 ( .A(n48), .Q(o_data_alu[25]) );
  INV3 U19 ( .A(n47), .Q(o_data_alu[26]) );
  INV3 U20 ( .A(n46), .Q(o_data_alu[27]) );
  INV3 U21 ( .A(n45), .Q(o_data_alu[28]) );
  INV3 U22 ( .A(n44), .Q(o_data_alu[29]) );
  INV3 U23 ( .A(n42), .Q(o_data_alu[30]) );
  INV3 U24 ( .A(n41), .Q(o_data_alu[31]) );
  INV3 U25 ( .A(n56), .Q(o_data_alu[18]) );
  INV3 U26 ( .A(n39), .Q(o_data_alu[4]) );
  INV3 U27 ( .A(n38), .Q(o_data_alu[5]) );
  INV3 U28 ( .A(n37), .Q(o_data_alu[6]) );
  BUF2 U29 ( .A(n7), .Q(n3) );
  BUF2 U30 ( .A(n7), .Q(n4) );
  BUF2 U31 ( .A(n7), .Q(n5) );
  BUF2 U32 ( .A(n7), .Q(n6) );
  AOI221 U33 ( .A(i_data_alures[0]), .B(n3), .C(i_data_pc8[0]), .D(n1), .Q(n65) );
  AOI221 U34 ( .A(i_data_alures[1]), .B(n4), .C(i_data_pc8[1]), .D(n1), .Q(n54) );
  AOI221 U35 ( .A(i_data_alures[2]), .B(n5), .C(i_data_pc8[2]), .D(n2), .Q(n43) );
  AOI221 U36 ( .A(i_data_alures[3]), .B(n6), .C(i_data_pc8[3]), .D(n2), .Q(n40) );
  AOI221 U37 ( .A(i_data_alures[16]), .B(n3), .C(i_data_pc8[16]), .D(n1), .Q(
        n58) );
  AOI221 U38 ( .A(i_data_alures[17]), .B(n4), .C(i_data_pc8[17]), .D(n1), .Q(
        n57) );
  AOI221 U39 ( .A(i_data_alures[18]), .B(n4), .C(i_data_pc8[18]), .D(n1), .Q(
        n56) );
  AOI221 U40 ( .A(i_data_alures[19]), .B(n4), .C(i_data_pc8[19]), .D(n1), .Q(
        n55) );
  AOI221 U41 ( .A(i_data_alures[20]), .B(n4), .C(i_data_pc8[20]), .D(n1), .Q(
        n53) );
  AOI221 U42 ( .A(i_data_alures[21]), .B(n4), .C(i_data_pc8[21]), .D(n2), .Q(
        n52) );
  AOI221 U43 ( .A(i_data_alures[22]), .B(n4), .C(i_data_pc8[22]), .D(n2), .Q(
        n51) );
  AOI221 U44 ( .A(i_data_alures[23]), .B(n4), .C(i_data_pc8[23]), .D(n2), .Q(
        n50) );
  AOI221 U45 ( .A(i_data_alures[24]), .B(n5), .C(i_data_pc8[24]), .D(n2), .Q(
        n49) );
  AOI221 U46 ( .A(i_data_alures[25]), .B(n5), .C(i_data_pc8[25]), .D(n2), .Q(
        n48) );
  AOI221 U47 ( .A(i_data_alures[26]), .B(n5), .C(i_data_pc8[26]), .D(n2), .Q(
        n47) );
  AOI221 U48 ( .A(i_data_alures[27]), .B(n5), .C(i_data_pc8[27]), .D(n2), .Q(
        n46) );
  AOI221 U49 ( .A(i_data_alures[28]), .B(n5), .C(i_data_pc8[28]), .D(n2), .Q(
        n45) );
  AOI221 U50 ( .A(i_data_alures[29]), .B(n5), .C(i_data_pc8[29]), .D(n2), .Q(
        n44) );
  AOI221 U51 ( .A(i_data_alures[30]), .B(n5), .C(i_data_pc8[30]), .D(n2), .Q(
        n42) );
  AOI221 U52 ( .A(i_data_alures[31]), .B(n6), .C(i_data_pc8[31]), .D(n2), .Q(
        n41) );
  INV3 U53 ( .A(i_con_pc8), .Q(n7) );
  INV3 U54 ( .A(n64), .Q(o_data_alu[10]) );
  AOI221 U55 ( .A(i_data_alures[10]), .B(n3), .C(i_data_pc8[10]), .D(n1), .Q(
        n64) );
  INV3 U56 ( .A(n63), .Q(o_data_alu[11]) );
  AOI221 U57 ( .A(i_data_alures[11]), .B(n3), .C(i_data_pc8[11]), .D(n1), .Q(
        n63) );
  INV3 U58 ( .A(n62), .Q(o_data_alu[12]) );
  AOI221 U59 ( .A(i_data_alures[12]), .B(n3), .C(i_data_pc8[12]), .D(n1), .Q(
        n62) );
  INV3 U60 ( .A(n61), .Q(o_data_alu[13]) );
  AOI221 U61 ( .A(i_data_alures[13]), .B(n3), .C(i_data_pc8[13]), .D(n1), .Q(
        n61) );
  INV3 U62 ( .A(n60), .Q(o_data_alu[14]) );
  AOI221 U63 ( .A(i_data_alures[14]), .B(n3), .C(i_data_pc8[14]), .D(n1), .Q(
        n60) );
  INV3 U64 ( .A(n59), .Q(o_data_alu[15]) );
  AOI221 U65 ( .A(i_data_alures[15]), .B(n3), .C(i_data_pc8[15]), .D(n1), .Q(
        n59) );
  AOI221 U66 ( .A(i_data_alures[4]), .B(n6), .C(i_data_pc8[4]), .D(n1), .Q(n39) );
  AOI221 U67 ( .A(i_data_alures[5]), .B(n6), .C(i_data_pc8[5]), .D(n2), .Q(n38) );
  AOI221 U68 ( .A(i_data_alures[6]), .B(n6), .C(i_data_pc8[6]), .D(n1), .Q(n37) );
  AOI221 U69 ( .A(i_data_alures[7]), .B(n6), .C(i_data_pc8[7]), .D(n2), .Q(n36) );
  AOI221 U70 ( .A(i_data_alures[8]), .B(n6), .C(i_data_pc8[8]), .D(n1), .Q(n35) );
  AOI221 U71 ( .A(i_data_alures[9]), .B(n6), .C(i_data_pc8[9]), .D(n2), .Q(n34) );
endmodule


module W_loadmux3 ( i_data_Rdata, i_con_loadsig, o_data_Wdata );
  input [31:0] i_data_Rdata;
  input [1:0] i_con_loadsig;
  output [31:0] o_data_Wdata;
  wire   n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n1, n2, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n51, n52;

  INV3 U2 ( .A(i_con_loadsig[0]), .Q(n52) );
  NOR21 U3 ( .A(n41), .B(n25), .Q(n49) );
  BUF6 U4 ( .A(n23), .Q(n2) );
  NOR22 U5 ( .A(i_con_loadsig[0]), .B(i_con_loadsig[1]), .Q(n25) );
  NOR22 U6 ( .A(n11), .B(n48), .Q(n21) );
  NAND22 U7 ( .A(i_con_loadsig[1]), .B(n52), .Q(n48) );
  AOI211 U8 ( .A(n41), .B(i_data_Rdata[15]), .C(n21), .Q(n23) );
  NOR21 U9 ( .A(n52), .B(i_con_loadsig[1]), .Q(n41) );
  NOR20 U10 ( .A(n51), .B(n11), .Q(o_data_Wdata[7]) );
  AOI210 U11 ( .A(n19), .B(i_data_Rdata[10]), .C(n21), .Q(n47) );
  AOI210 U12 ( .A(n19), .B(i_data_Rdata[11]), .C(n21), .Q(n46) );
  AOI210 U13 ( .A(n19), .B(i_data_Rdata[12]), .C(n21), .Q(n45) );
  AOI210 U14 ( .A(n19), .B(i_data_Rdata[13]), .C(n21), .Q(n44) );
  AOI210 U15 ( .A(n19), .B(i_data_Rdata[14]), .C(n21), .Q(n43) );
  AOI210 U16 ( .A(n19), .B(i_data_Rdata[15]), .C(n21), .Q(n42) );
  NAND20 U17 ( .A(i_data_Rdata[16]), .B(n25), .Q(n40) );
  NAND20 U18 ( .A(i_data_Rdata[17]), .B(n25), .Q(n39) );
  NAND20 U19 ( .A(i_data_Rdata[18]), .B(n25), .Q(n38) );
  NAND20 U20 ( .A(i_data_Rdata[19]), .B(n25), .Q(n37) );
  NAND20 U21 ( .A(i_data_Rdata[20]), .B(n25), .Q(n36) );
  NAND20 U22 ( .A(i_data_Rdata[21]), .B(n25), .Q(n35) );
  NAND20 U23 ( .A(i_data_Rdata[22]), .B(n25), .Q(n34) );
  CLKIN3 U24 ( .A(n22), .Q(o_data_Wdata[8]) );
  AOI210 U25 ( .A(n19), .B(i_data_Rdata[8]), .C(n21), .Q(n22) );
  CLKIN3 U26 ( .A(n20), .Q(o_data_Wdata[9]) );
  AOI210 U27 ( .A(n19), .B(i_data_Rdata[9]), .C(n21), .Q(n20) );
  INV3 U28 ( .A(n49), .Q(n19) );
  INV3 U29 ( .A(n50), .Q(n51) );
  NAND22 U30 ( .A(n49), .B(n48), .Q(n50) );
  INV3 U31 ( .A(n47), .Q(o_data_Wdata[10]) );
  INV3 U32 ( .A(n46), .Q(o_data_Wdata[11]) );
  INV3 U33 ( .A(n45), .Q(o_data_Wdata[12]) );
  INV3 U34 ( .A(n44), .Q(o_data_Wdata[13]) );
  INV3 U35 ( .A(n43), .Q(o_data_Wdata[14]) );
  INV3 U36 ( .A(n42), .Q(o_data_Wdata[15]) );
  BUF2 U37 ( .A(n25), .Q(n1) );
  INV3 U38 ( .A(i_data_Rdata[7]), .Q(n11) );
  NOR21 U39 ( .A(n51), .B(n18), .Q(o_data_Wdata[0]) );
  INV3 U40 ( .A(i_data_Rdata[0]), .Q(n18) );
  NOR21 U41 ( .A(n51), .B(n17), .Q(o_data_Wdata[1]) );
  INV3 U42 ( .A(i_data_Rdata[1]), .Q(n17) );
  NOR21 U43 ( .A(n51), .B(n16), .Q(o_data_Wdata[2]) );
  INV3 U44 ( .A(i_data_Rdata[2]), .Q(n16) );
  NOR21 U45 ( .A(n51), .B(n15), .Q(o_data_Wdata[3]) );
  INV3 U46 ( .A(i_data_Rdata[3]), .Q(n15) );
  NOR21 U47 ( .A(n51), .B(n14), .Q(o_data_Wdata[4]) );
  INV3 U48 ( .A(i_data_Rdata[4]), .Q(n14) );
  NOR21 U49 ( .A(n51), .B(n13), .Q(o_data_Wdata[5]) );
  INV3 U50 ( .A(i_data_Rdata[5]), .Q(n13) );
  NOR21 U51 ( .A(n51), .B(n12), .Q(o_data_Wdata[6]) );
  INV3 U52 ( .A(i_data_Rdata[6]), .Q(n12) );
  NAND22 U53 ( .A(n2), .B(n40), .Q(o_data_Wdata[16]) );
  NAND22 U54 ( .A(n2), .B(n39), .Q(o_data_Wdata[17]) );
  NAND22 U55 ( .A(n2), .B(n38), .Q(o_data_Wdata[18]) );
  NAND22 U56 ( .A(n2), .B(n37), .Q(o_data_Wdata[19]) );
  NAND22 U57 ( .A(n2), .B(n36), .Q(o_data_Wdata[20]) );
  NAND22 U58 ( .A(n2), .B(n35), .Q(o_data_Wdata[21]) );
  NAND22 U59 ( .A(n2), .B(n34), .Q(o_data_Wdata[22]) );
  NAND22 U60 ( .A(n2), .B(n33), .Q(o_data_Wdata[23]) );
  NAND22 U61 ( .A(i_data_Rdata[23]), .B(n1), .Q(n33) );
  NAND22 U62 ( .A(n2), .B(n32), .Q(o_data_Wdata[24]) );
  NAND22 U63 ( .A(i_data_Rdata[24]), .B(n1), .Q(n32) );
  NAND22 U64 ( .A(n2), .B(n31), .Q(o_data_Wdata[25]) );
  NAND22 U65 ( .A(i_data_Rdata[25]), .B(n1), .Q(n31) );
  NAND22 U66 ( .A(n2), .B(n30), .Q(o_data_Wdata[26]) );
  NAND22 U67 ( .A(i_data_Rdata[26]), .B(n1), .Q(n30) );
  NAND22 U68 ( .A(n2), .B(n29), .Q(o_data_Wdata[27]) );
  NAND22 U69 ( .A(i_data_Rdata[27]), .B(n1), .Q(n29) );
  NAND22 U70 ( .A(n2), .B(n28), .Q(o_data_Wdata[28]) );
  NAND22 U71 ( .A(i_data_Rdata[28]), .B(n1), .Q(n28) );
  NAND22 U72 ( .A(n2), .B(n27), .Q(o_data_Wdata[29]) );
  NAND22 U73 ( .A(i_data_Rdata[29]), .B(n1), .Q(n27) );
  NAND22 U74 ( .A(n2), .B(n26), .Q(o_data_Wdata[30]) );
  NAND22 U75 ( .A(i_data_Rdata[30]), .B(n1), .Q(n26) );
  NAND22 U76 ( .A(n2), .B(n24), .Q(o_data_Wdata[31]) );
  NAND22 U77 ( .A(i_data_Rdata[31]), .B(n1), .Q(n24) );
endmodule


module W_datamux ( i_data_alu, i_data_load, i_con_memtoreg, o_data_toreg );
  input [31:0] i_data_alu;
  input [31:0] i_data_load;
  output [31:0] o_data_toreg;
  input i_con_memtoreg;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n1, n2, n3, n4, n5, n6;

  INV3 U1 ( .A(n35), .Q(o_data_toreg[8]) );
  INV3 U2 ( .A(n38), .Q(o_data_toreg[5]) );
  INV3 U3 ( .A(n37), .Q(o_data_toreg[6]) );
  INV3 U4 ( .A(n52), .Q(o_data_toreg[21]) );
  INV3 U5 ( .A(n65), .Q(o_data_toreg[0]) );
  INV3 U6 ( .A(n34), .Q(o_data_toreg[9]) );
  INV3 U7 ( .A(n40), .Q(o_data_toreg[3]) );
  INV3 U8 ( .A(n51), .Q(o_data_toreg[22]) );
  INV3 U9 ( .A(n39), .Q(o_data_toreg[4]) );
  INV3 U10 ( .A(n43), .Q(o_data_toreg[2]) );
  CLKIN3 U11 ( .A(n54), .Q(o_data_toreg[1]) );
  CLKIN3 U12 ( .A(n58), .Q(o_data_toreg[16]) );
  CLKIN3 U13 ( .A(n57), .Q(o_data_toreg[17]) );
  CLKIN3 U14 ( .A(n56), .Q(o_data_toreg[18]) );
  CLKIN3 U15 ( .A(n55), .Q(o_data_toreg[19]) );
  CLKIN3 U16 ( .A(n53), .Q(o_data_toreg[20]) );
  CLKIN3 U17 ( .A(n50), .Q(o_data_toreg[23]) );
  CLKIN3 U18 ( .A(n49), .Q(o_data_toreg[24]) );
  CLKIN3 U19 ( .A(n48), .Q(o_data_toreg[25]) );
  CLKIN3 U20 ( .A(n47), .Q(o_data_toreg[26]) );
  CLKIN3 U21 ( .A(n46), .Q(o_data_toreg[27]) );
  CLKIN3 U22 ( .A(n45), .Q(o_data_toreg[28]) );
  CLKIN3 U23 ( .A(n44), .Q(o_data_toreg[29]) );
  CLKIN3 U24 ( .A(n42), .Q(o_data_toreg[30]) );
  CLKIN3 U25 ( .A(n41), .Q(o_data_toreg[31]) );
  CLKIN3 U26 ( .A(n64), .Q(o_data_toreg[10]) );
  CLKIN3 U27 ( .A(n63), .Q(o_data_toreg[11]) );
  CLKIN3 U28 ( .A(n62), .Q(o_data_toreg[12]) );
  CLKIN3 U29 ( .A(n61), .Q(o_data_toreg[13]) );
  CLKIN3 U30 ( .A(n60), .Q(o_data_toreg[14]) );
  CLKIN3 U31 ( .A(n59), .Q(o_data_toreg[15]) );
  CLKIN3 U32 ( .A(n36), .Q(o_data_toreg[7]) );
  AOI221 U33 ( .A(i_data_alu[0]), .B(n2), .C(i_data_load[0]), .D(n1), .Q(n65)
         );
  AOI221 U34 ( .A(i_data_alu[1]), .B(n3), .C(i_data_load[1]), .D(
        i_con_memtoreg), .Q(n54) );
  AOI221 U35 ( .A(i_data_alu[2]), .B(n4), .C(i_data_load[2]), .D(n1), .Q(n43)
         );
  AOI221 U36 ( .A(i_data_alu[3]), .B(n5), .C(i_data_load[3]), .D(n1), .Q(n40)
         );
  AOI221 U37 ( .A(i_data_alu[10]), .B(n2), .C(i_data_load[10]), .D(
        i_con_memtoreg), .Q(n64) );
  AOI221 U38 ( .A(i_data_alu[11]), .B(n2), .C(i_data_load[11]), .D(
        i_con_memtoreg), .Q(n63) );
  AOI221 U39 ( .A(i_data_alu[12]), .B(n2), .C(i_data_load[12]), .D(
        i_con_memtoreg), .Q(n62) );
  AOI221 U40 ( .A(i_data_alu[13]), .B(n2), .C(i_data_load[13]), .D(
        i_con_memtoreg), .Q(n61) );
  AOI221 U41 ( .A(i_data_alu[14]), .B(n2), .C(i_data_load[14]), .D(
        i_con_memtoreg), .Q(n60) );
  AOI221 U42 ( .A(i_data_alu[15]), .B(n2), .C(i_data_load[15]), .D(
        i_con_memtoreg), .Q(n59) );
  AOI221 U43 ( .A(i_data_alu[16]), .B(n2), .C(i_data_load[16]), .D(
        i_con_memtoreg), .Q(n58) );
  AOI221 U44 ( .A(i_data_alu[17]), .B(n3), .C(i_data_load[17]), .D(
        i_con_memtoreg), .Q(n57) );
  AOI221 U45 ( .A(i_data_alu[19]), .B(n3), .C(i_data_load[19]), .D(
        i_con_memtoreg), .Q(n55) );
  AOI221 U46 ( .A(i_data_alu[20]), .B(n3), .C(i_data_load[20]), .D(
        i_con_memtoreg), .Q(n53) );
  AOI221 U47 ( .A(i_data_alu[21]), .B(n3), .C(i_data_load[21]), .D(n1), .Q(n52) );
  AOI221 U48 ( .A(i_data_alu[22]), .B(n3), .C(i_data_load[22]), .D(n1), .Q(n51) );
  AOI221 U49 ( .A(i_data_alu[23]), .B(n3), .C(i_data_load[23]), .D(n1), .Q(n50) );
  AOI221 U50 ( .A(i_data_alu[24]), .B(n4), .C(i_data_load[24]), .D(n1), .Q(n49) );
  AOI221 U51 ( .A(i_data_alu[25]), .B(n4), .C(i_data_load[25]), .D(n1), .Q(n48) );
  AOI221 U52 ( .A(i_data_alu[26]), .B(n4), .C(i_data_load[26]), .D(n1), .Q(n47) );
  AOI221 U53 ( .A(i_data_alu[27]), .B(n4), .C(i_data_load[27]), .D(n1), .Q(n46) );
  AOI221 U54 ( .A(i_data_alu[28]), .B(n4), .C(i_data_load[28]), .D(n1), .Q(n45) );
  AOI221 U55 ( .A(i_data_alu[29]), .B(n4), .C(i_data_load[29]), .D(n1), .Q(n44) );
  AOI221 U56 ( .A(i_data_alu[30]), .B(n4), .C(i_data_load[30]), .D(n1), .Q(n42) );
  AOI221 U57 ( .A(i_data_alu[31]), .B(n5), .C(i_data_load[31]), .D(n1), .Q(n41) );
  AOI221 U58 ( .A(i_data_alu[18]), .B(n3), .C(i_data_load[18]), .D(n1), .Q(n56) );
  AOI221 U59 ( .A(i_data_alu[4]), .B(n5), .C(i_data_load[4]), .D(n1), .Q(n39)
         );
  AOI221 U60 ( .A(i_data_alu[5]), .B(n5), .C(i_data_load[5]), .D(n1), .Q(n38)
         );
  AOI221 U61 ( .A(i_data_alu[6]), .B(n5), .C(i_data_load[6]), .D(n1), .Q(n37)
         );
  AOI221 U62 ( .A(i_data_alu[7]), .B(n5), .C(i_data_load[7]), .D(n1), .Q(n36)
         );
  INV3 U63 ( .A(n6), .Q(n1) );
  BUF2 U64 ( .A(n6), .Q(n2) );
  BUF2 U65 ( .A(n6), .Q(n3) );
  BUF2 U66 ( .A(n6), .Q(n4) );
  BUF2 U67 ( .A(n6), .Q(n5) );
  AOI221 U68 ( .A(i_data_alu[8]), .B(n5), .C(i_data_load[8]), .D(n1), .Q(n35)
         );
  AOI221 U69 ( .A(i_data_alu[9]), .B(n5), .C(i_data_load[9]), .D(n1), .Q(n34)
         );
  INV3 U70 ( .A(i_con_memtoreg), .Q(n6) );
endmodule


module writeback ( i_data_pc8, i_data_alures, i_data_memout, i_con_Wloadmux, 
        i_con_Walupc8, i_con_Wmemtoreg, o_data_regwrite );
  input [31:0] i_data_pc8;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [1:0] i_con_Wloadmux;
  output [31:0] o_data_regwrite;
  input i_con_Walupc8, i_con_Wmemtoreg;

  wire   [31:0] datamux_i_data_alu;
  wire   [31:0] datamux_i_data_load;

  W_resmux u_resmux ( .i_data_alures(i_data_alures), .i_data_pc8(i_data_pc8), 
        .i_con_pc8(i_con_Walupc8), .o_data_alu(datamux_i_data_alu) );
  W_loadmux3 u_loadmux ( .i_data_Rdata(i_data_memout), .i_con_loadsig(
        i_con_Wloadmux), .o_data_Wdata(datamux_i_data_load) );
  W_datamux u_datamux ( .i_data_alu(datamux_i_data_alu), .i_data_load(
        datamux_i_data_load), .i_con_memtoreg(i_con_Wmemtoreg), .o_data_toreg(
        o_data_regwrite) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Mmemread, ex_con_Mmemwrite, ex_con_Walupc8, ex_con_Wmemtoreg,
         mem_con_Walupc8, mem_con_Wmemtoreg, wb_con_Walupc8, wb_con_Wmemtoreg,
         n1, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26,
         SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28,
         SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30,
         SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32,
         SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34;
  wire   [31:0] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [31:0] id_addr_pc4;
  wire   [31:0] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [1:0] ex_con_Wloadmux;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] wb_data_memout;
  wire   [31:0] mem_data_pc4;
  wire   [1:0] mem_con_Wloadmux;
  wire   [31:0] wb_data_pc8;
  wire   [31:0] mem_data_alures;
  wire   [1:0] wb_con_Wloadmux;

  fetch u_fetch ( .i_clk(clk), .i_nrst(rst_n), .i_addr_b(if_addr_b), 
        .i_addr_j({if_addr_j, n1, n1}), .i_addr_jr(id_data_jr), .i_con_b(
        if_con_b), .i_con_j(if_con_j), .i_data_instr(read_instruction), 
        .i_con_ifstall(if_con_ifstall), .o_addr_pc(instruction_address), 
        .o_addr_pc4(id_addr_pc4), .o_data_instr(id_data_instr) );
  decode u_decode ( .i_clk(clk), .i_nrst(rst_n), .i_addr_pc4(id_addr_pc4), 
        .i_data_instr(id_data_instr), .i_con_Wregwrite(id_con_Wregwrite), 
        .i_data_Wregwrite(id_data_Wregwrite), .i_addr_Wregwrite(
        id_addr_Wregwrite), .i_addr_Erd(for_o_addr_Erd), .i_addr_Mrd(
        mem_addr_regdst), .i_con_Eregwrite(ex_con_Wregwrite), 
        .i_con_Mregwrite(mem_con_Wregwrite), .i_addr_rtM(for_addr_rtM), 
        .i_addr_rtW(for_addr_rtW), .i_con_memreadM(mem_read), .i_con_memreadW(
        for_FWmemread), .o_data_rs(id_data_rs), .o_data_rt(ex_data_rt), 
        .o_addr_rd(ex_addr_rd), .o_addr_rt(ex_addr_rt), .o_data_jr(id_data_jr), 
        .o_con_jump(if_con_j), .o_addr_pc4(ex_data_pc4), .o_addr_branch(
        if_addr_b), .o_addr_jump({if_addr_j, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .o_con_Ealuop(ex_con_Ealuop), 
        .o_con_Ealusrc(ex_con_Ealusrc), .o_con_Eregdst(ex_con_Eregdst), 
        .o_con_Mmemread(ex_con_Mmemread), .o_con_Mmemwrite(ex_con_Mmemwrite), 
        .o_con_Wloadmux(ex_con_Wloadmux), .o_con_Walupc8(ex_con_Walupc8), 
        .o_con_Wmemtoreg(ex_con_Wmemtoreg), .o_con_Wregwrite(ex_con_Wregwrite), 
        .o_con_ifstall(if_con_ifstall), .o_con_Ebop(ex_con_bop), 
        .o_data_signext(ex_data_immext), .o_con_Efamux(for_o_con_Efamux), 
        .o_con_Efbmux(for_o_con_Efbmux), .o_data_Fmemout(for_memout) );
  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext(
        ex_data_immext), .i_addr_rt(ex_addr_rt), .i_addr_rd(ex_addr_rd), 
        .i_data_FEalures(data_address), .i_data_FMalures(id_data_Wregwrite), 
        .i_data_FMmemout(wb_data_memout), .i_data_FWmemout(for_memout), 
        .i_con_Ealuop(ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), 
        .i_con_Mmemwrite(ex_con_Mmemwrite), .i_con_Wloadmux(ex_con_Wloadmux), 
        .i_con_Walupc8(ex_con_Walupc8), .i_con_Wmemtoreg(ex_con_Wmemtoreg), 
        .i_con_Wregwrite(ex_con_Wregwrite), .i_con_Efamux(for_o_con_Efamux), 
        .i_con_Efbmux(for_o_con_Efbmux), .i_con_bop(ex_con_bop), .o_data_pc4(
        mem_data_pc4), .o_data_alures(data_address), .o_data_rt(write_data), 
        .o_addr_regdst(mem_addr_regdst), .o_con_Mmemread(mem_read), 
        .o_con_Mmemwrite(mem_write), .o_con_Wloadmux(mem_con_Wloadmux), 
        .o_con_Walupc8(mem_con_Walupc8), .o_con_Wmemtoreg(mem_con_Wmemtoreg), 
        .o_con_Wregwrite(mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), 
        .o_addr_Mrt(for_addr_rtM), .o_FaluresE({SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, 
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, 
        SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, 
        SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, 
        SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, 
        SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, 
        SYNOPSYS_UNCONNECTED_34}), .o_con_ifbranch(if_con_b) );
  mem u_mem ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(mem_data_pc4), 
        .i_data_alures(data_address), .i_data_memout(read_data), 
        .i_addr_regdst(mem_addr_regdst), .i_con_Wloadmux(mem_con_Wloadmux), 
        .i_con_Walupc8(mem_con_Walupc8), .i_con_Wmemtoreg(mem_con_Wmemtoreg), 
        .i_con_Wregwrite(mem_con_Wregwrite), .i_con_FWmemread(ex_con_Mmemread), 
        .i_addr_Mrt(for_addr_rtM), .o_data_pc8(wb_data_pc8), .o_data_alures(
        mem_data_alures), .o_data_memout(wb_data_memout), .o_addr_regdst(
        id_addr_Wregwrite), .o_con_Wloadmux(wb_con_Wloadmux), .o_con_Walupc8(
        wb_con_Walupc8), .o_con_Wmemtoreg(wb_con_Wmemtoreg), .o_con_Wregwrite(
        id_con_Wregwrite), .o_con_FWmemread(for_FWmemread), .o_addr_Wrt(
        for_addr_rtW) );
  writeback u_writeback ( .i_data_pc8(wb_data_pc8), .i_data_alures(
        mem_data_alures), .i_data_memout(wb_data_memout), .i_con_Wloadmux(
        wb_con_Wloadmux), .i_con_Walupc8(wb_con_Walupc8), .i_con_Wmemtoreg(
        wb_con_Wmemtoreg), .o_data_regwrite(id_data_Wregwrite) );
  LOGIC0 U1 ( .Q(n1) );
endmodule

