// Verilog simulation library for c35_IOLIB_ANA_3B_3M
// Owner: austriamicrosystems AG  HIT-Kit: Digital
module APRIO1K5P_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO200P_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO50P_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO500P_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module AVSUBP_3B (A);
  input A ;
endmodule
module APRIOWP_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module AGNDALLP_3B (A);
  input A ;
endmodule
module AVDDALLP_3B (A);
  input A ;
endmodule
module APRIOP_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
