module FILLANT25 (ANT1);
  input ANT1 ;
endmodule
module FILLANT10 (ANT1);
  input ANT1 ;
endmodule
module FILLANT1 (ANT1);
  input ANT1 ;
endmodule
module FILLANT2 (ANT1);
  input ANT1 ;
endmodule
module FILLANT5 (ANT1);
  input ANT1 ;
endmodule
module FILLANT25_3B (ANT1);
  input ANT1 ;
endmodule
module FILLANT10_3B (ANT1);
  input ANT1 ;
endmodule
module FILLANT1_3B (ANT1);
  input ANT1 ;
endmodule
module FILLANT2_3B (ANT1);
  input ANT1 ;
endmodule
module FILLANT5_3B (ANT1);
  input ANT1 ;
endmodule
