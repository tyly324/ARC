
module F_jumpmux ( i_addr_j, i_addr_jr, i_addr_pc4, i_con_jump, o_addr_jumpmux
 );
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [31:0] i_addr_pc4;
  input [1:0] i_con_jump;
  output [31:0] o_addr_jumpmux;
  wire   n3, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n23,
         n24, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n1, n2, n5, n6, n19, n20,
         n21, n22, n25, n26, n27, n28, n29, n30, n31, n32, n69, n70, n71, n72;

  BUF2 U1 ( .A(n71), .Q(n1) );
  AOI221 U2 ( .A(i_addr_pc4[3]), .B(n1), .C(i_addr_jr[3]), .D(n70), .Q(n17) );
  AOI221 U3 ( .A(i_addr_pc4[4]), .B(n1), .C(i_addr_jr[4]), .D(n70), .Q(n15) );
  AOI221 U4 ( .A(i_addr_pc4[5]), .B(n71), .C(i_addr_jr[5]), .D(n70), .Q(n13)
         );
  AOI221 U5 ( .A(i_addr_pc4[6]), .B(n71), .C(i_addr_jr[6]), .D(n70), .Q(n11)
         );
  AOI221 U6 ( .A(i_addr_pc4[7]), .B(n1), .C(i_addr_jr[7]), .D(n70), .Q(n9) );
  AOI221 U7 ( .A(i_addr_pc4[8]), .B(n1), .C(i_addr_jr[8]), .D(n70), .Q(n7) );
  AOI221 U8 ( .A(i_addr_pc4[9]), .B(n1), .C(i_addr_jr[9]), .D(n70), .Q(n3) );
  AOI221 U9 ( .A(i_addr_pc4[2]), .B(n71), .C(i_addr_jr[2]), .D(n70), .Q(n23)
         );
  AOI221 U10 ( .A(i_addr_pc4[15]), .B(n1), .C(i_addr_jr[15]), .D(n70), .Q(n55)
         );
  AOI221 U11 ( .A(i_addr_pc4[16]), .B(n71), .C(i_addr_jr[16]), .D(n70), .Q(n53) );
  AOI221 U12 ( .A(i_addr_pc4[17]), .B(n71), .C(i_addr_jr[17]), .D(n70), .Q(n51) );
  AOI221 U13 ( .A(i_addr_pc4[18]), .B(n71), .C(i_addr_jr[18]), .D(n70), .Q(n49) );
  AOI221 U14 ( .A(i_addr_pc4[19]), .B(n71), .C(i_addr_jr[19]), .D(n70), .Q(n47) );
  AOI221 U15 ( .A(i_addr_pc4[20]), .B(n71), .C(i_addr_jr[20]), .D(n70), .Q(n43) );
  AOI221 U16 ( .A(i_addr_pc4[21]), .B(n1), .C(i_addr_jr[21]), .D(n70), .Q(n41)
         );
  AOI221 U17 ( .A(i_addr_pc4[22]), .B(n1), .C(i_addr_jr[22]), .D(n70), .Q(n39)
         );
  AOI221 U18 ( .A(i_addr_pc4[23]), .B(n1), .C(i_addr_jr[23]), .D(n70), .Q(n37)
         );
  AOI221 U19 ( .A(i_addr_pc4[24]), .B(n1), .C(i_addr_jr[24]), .D(n70), .Q(n35)
         );
  AOI221 U20 ( .A(i_addr_pc4[25]), .B(n1), .C(i_addr_jr[25]), .D(n70), .Q(n33)
         );
  AOI221 U21 ( .A(i_addr_pc4[10]), .B(n1), .C(i_addr_jr[10]), .D(n70), .Q(n65)
         );
  AOI221 U22 ( .A(i_addr_pc4[11]), .B(n1), .C(i_addr_jr[11]), .D(n70), .Q(n63)
         );
  AOI221 U23 ( .A(i_addr_pc4[12]), .B(n1), .C(i_addr_jr[12]), .D(n70), .Q(n61)
         );
  AOI221 U24 ( .A(i_addr_pc4[13]), .B(n1), .C(i_addr_jr[13]), .D(n70), .Q(n59)
         );
  AOI221 U25 ( .A(i_addr_pc4[14]), .B(n1), .C(i_addr_jr[14]), .D(n70), .Q(n57)
         );
  INV3 U26 ( .A(n19), .Q(n70) );
  NAND22 U27 ( .A(n67), .B(n68), .Q(o_addr_jumpmux[0]) );
  NAND22 U28 ( .A(i_addr_j[0]), .B(n72), .Q(n68) );
  NAND22 U29 ( .A(n65), .B(n66), .Q(o_addr_jumpmux[10]) );
  NAND22 U30 ( .A(i_addr_j[10]), .B(n72), .Q(n66) );
  NAND22 U31 ( .A(n63), .B(n64), .Q(o_addr_jumpmux[11]) );
  NAND22 U32 ( .A(i_addr_j[11]), .B(n72), .Q(n64) );
  NAND22 U33 ( .A(n61), .B(n62), .Q(o_addr_jumpmux[12]) );
  NAND22 U34 ( .A(i_addr_j[12]), .B(n72), .Q(n62) );
  NAND22 U35 ( .A(n59), .B(n60), .Q(o_addr_jumpmux[13]) );
  NAND22 U36 ( .A(i_addr_j[13]), .B(n72), .Q(n60) );
  NAND22 U37 ( .A(n57), .B(n58), .Q(o_addr_jumpmux[14]) );
  NAND22 U38 ( .A(i_addr_j[14]), .B(n72), .Q(n58) );
  NAND22 U39 ( .A(n55), .B(n56), .Q(o_addr_jumpmux[15]) );
  NAND22 U40 ( .A(i_addr_j[15]), .B(n72), .Q(n56) );
  NAND22 U41 ( .A(n53), .B(n54), .Q(o_addr_jumpmux[16]) );
  NAND22 U42 ( .A(i_addr_j[16]), .B(n72), .Q(n54) );
  NAND22 U43 ( .A(n51), .B(n52), .Q(o_addr_jumpmux[17]) );
  NAND22 U44 ( .A(i_addr_j[17]), .B(n72), .Q(n52) );
  NAND22 U45 ( .A(n49), .B(n50), .Q(o_addr_jumpmux[18]) );
  NAND22 U46 ( .A(i_addr_j[18]), .B(n72), .Q(n50) );
  NAND22 U47 ( .A(n47), .B(n48), .Q(o_addr_jumpmux[19]) );
  NAND22 U48 ( .A(i_addr_j[19]), .B(n72), .Q(n48) );
  NAND22 U49 ( .A(n3), .B(n4), .Q(o_addr_jumpmux[9]) );
  NAND22 U50 ( .A(i_addr_j[9]), .B(n72), .Q(n4) );
  NAND22 U51 ( .A(n45), .B(n46), .Q(o_addr_jumpmux[1]) );
  NAND22 U52 ( .A(i_addr_j[1]), .B(n72), .Q(n46) );
  NAND22 U53 ( .A(n23), .B(n24), .Q(o_addr_jumpmux[2]) );
  NAND22 U54 ( .A(i_addr_j[2]), .B(n72), .Q(n24) );
  NAND22 U55 ( .A(n17), .B(n18), .Q(o_addr_jumpmux[3]) );
  NAND22 U56 ( .A(i_addr_j[3]), .B(n72), .Q(n18) );
  NAND22 U57 ( .A(n15), .B(n16), .Q(o_addr_jumpmux[4]) );
  NAND22 U58 ( .A(i_addr_j[4]), .B(n72), .Q(n16) );
  NAND22 U59 ( .A(n13), .B(n14), .Q(o_addr_jumpmux[5]) );
  NAND22 U60 ( .A(i_addr_j[5]), .B(n72), .Q(n14) );
  NAND22 U61 ( .A(n11), .B(n12), .Q(o_addr_jumpmux[6]) );
  NAND22 U62 ( .A(i_addr_j[6]), .B(n72), .Q(n12) );
  NAND22 U63 ( .A(n9), .B(n10), .Q(o_addr_jumpmux[7]) );
  NAND22 U64 ( .A(i_addr_j[7]), .B(n72), .Q(n10) );
  NAND22 U65 ( .A(n7), .B(n8), .Q(o_addr_jumpmux[8]) );
  NAND22 U66 ( .A(i_addr_j[8]), .B(n72), .Q(n8) );
  NAND22 U67 ( .A(n43), .B(n44), .Q(o_addr_jumpmux[20]) );
  NAND22 U68 ( .A(i_addr_j[20]), .B(n72), .Q(n44) );
  NAND22 U69 ( .A(n41), .B(n42), .Q(o_addr_jumpmux[21]) );
  NAND22 U70 ( .A(i_addr_j[21]), .B(n72), .Q(n42) );
  NAND22 U71 ( .A(n39), .B(n40), .Q(o_addr_jumpmux[22]) );
  NAND22 U72 ( .A(i_addr_j[22]), .B(n72), .Q(n40) );
  NAND22 U73 ( .A(n37), .B(n38), .Q(o_addr_jumpmux[23]) );
  NAND22 U74 ( .A(i_addr_j[23]), .B(n72), .Q(n38) );
  NAND22 U75 ( .A(n35), .B(n36), .Q(o_addr_jumpmux[24]) );
  NAND22 U76 ( .A(i_addr_j[24]), .B(n72), .Q(n36) );
  NAND22 U77 ( .A(n33), .B(n34), .Q(o_addr_jumpmux[25]) );
  NAND22 U78 ( .A(i_addr_j[25]), .B(n72), .Q(n34) );
  AOI221 U79 ( .A(i_addr_j[26]), .B(n72), .C(i_addr_pc4[26]), .D(n71), .Q(n21)
         );
  AOI221 U80 ( .A(i_addr_j[27]), .B(n72), .C(i_addr_pc4[27]), .D(n71), .Q(n25)
         );
  AOI221 U81 ( .A(i_addr_j[28]), .B(n72), .C(i_addr_pc4[28]), .D(n71), .Q(n27)
         );
  AOI221 U82 ( .A(i_addr_j[29]), .B(n72), .C(i_addr_pc4[29]), .D(n71), .Q(n29)
         );
  AOI221 U83 ( .A(i_addr_j[30]), .B(n72), .C(i_addr_pc4[30]), .D(n71), .Q(n31)
         );
  AOI221 U84 ( .A(i_addr_j[31]), .B(n72), .C(i_addr_pc4[31]), .D(n71), .Q(n69)
         );
  AOI221 U85 ( .A(i_addr_pc4[1]), .B(n1), .C(i_addr_jr[1]), .D(n70), .Q(n45)
         );
  AOI221 U86 ( .A(i_addr_pc4[0]), .B(n1), .C(i_addr_jr[0]), .D(n70), .Q(n67)
         );
  CLKIN3 U87 ( .A(i_con_jump[1]), .Q(n2) );
  NAND22 U88 ( .A(i_con_jump[0]), .B(n2), .Q(n5) );
  CLKIN3 U89 ( .A(n5), .Q(n72) );
  XNR21 U90 ( .A(i_con_jump[0]), .B(i_con_jump[1]), .Q(n71) );
  CLKIN3 U91 ( .A(i_con_jump[0]), .Q(n6) );
  NAND22 U92 ( .A(i_con_jump[1]), .B(n6), .Q(n19) );
  NAND22 U93 ( .A(i_addr_jr[26]), .B(n70), .Q(n20) );
  NAND22 U94 ( .A(n21), .B(n20), .Q(o_addr_jumpmux[26]) );
  NAND22 U95 ( .A(i_addr_jr[27]), .B(n70), .Q(n22) );
  NAND22 U96 ( .A(n25), .B(n22), .Q(o_addr_jumpmux[27]) );
  NAND22 U97 ( .A(i_addr_jr[28]), .B(n70), .Q(n26) );
  NAND22 U98 ( .A(n27), .B(n26), .Q(o_addr_jumpmux[28]) );
  NAND22 U99 ( .A(i_addr_jr[29]), .B(n70), .Q(n28) );
  NAND22 U100 ( .A(n29), .B(n28), .Q(o_addr_jumpmux[29]) );
  NAND22 U101 ( .A(i_addr_jr[30]), .B(n70), .Q(n30) );
  NAND22 U102 ( .A(n31), .B(n30), .Q(o_addr_jumpmux[30]) );
  NAND22 U103 ( .A(i_addr_jr[31]), .B(n70), .Q(n32) );
  NAND22 U104 ( .A(n69), .B(n32), .Q(o_addr_jumpmux[31]) );
endmodule


module F_branchmux ( i_addr_jumpmux, i_addr_b, i_con_ifbranch, o_addr_nextpc
 );
  input [31:0] i_addr_jumpmux;
  input [31:0] i_addr_b;
  output [31:0] o_addr_nextpc;
  input i_con_ifbranch;
  wire   n34, n35, n36, n37, n38, n39, n40, n43, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n1, n2,
         n3, n4, n5;

  INV3 U1 ( .A(i_con_ifbranch), .Q(n5) );
  INV3 U2 ( .A(n3), .Q(n2) );
  INV2 U3 ( .A(n5), .Q(n1) );
  INV2 U4 ( .A(n65), .Q(o_addr_nextpc[0]) );
  INV2 U5 ( .A(n64), .Q(o_addr_nextpc[10]) );
  INV2 U6 ( .A(n63), .Q(o_addr_nextpc[11]) );
  INV2 U7 ( .A(n62), .Q(o_addr_nextpc[12]) );
  INV2 U8 ( .A(n61), .Q(o_addr_nextpc[13]) );
  INV2 U9 ( .A(n60), .Q(o_addr_nextpc[14]) );
  INV2 U10 ( .A(n59), .Q(o_addr_nextpc[15]) );
  INV2 U11 ( .A(n58), .Q(o_addr_nextpc[16]) );
  INV2 U12 ( .A(n57), .Q(o_addr_nextpc[17]) );
  INV2 U13 ( .A(n56), .Q(o_addr_nextpc[18]) );
  INV2 U14 ( .A(n55), .Q(o_addr_nextpc[19]) );
  INV2 U15 ( .A(n34), .Q(o_addr_nextpc[9]) );
  AOI220 U16 ( .A(n2), .B(i_addr_b[9]), .C(i_addr_jumpmux[9]), .D(n3), .Q(n34)
         );
  INV2 U17 ( .A(n54), .Q(o_addr_nextpc[1]) );
  INV2 U18 ( .A(n43), .Q(o_addr_nextpc[2]) );
  INV2 U19 ( .A(n40), .Q(o_addr_nextpc[3]) );
  INV2 U20 ( .A(n39), .Q(o_addr_nextpc[4]) );
  INV2 U21 ( .A(n38), .Q(o_addr_nextpc[5]) );
  INV2 U22 ( .A(n37), .Q(o_addr_nextpc[6]) );
  INV2 U23 ( .A(n36), .Q(o_addr_nextpc[7]) );
  AOI220 U24 ( .A(i_addr_b[7]), .B(n2), .C(i_addr_jumpmux[7]), .D(n3), .Q(n36)
         );
  INV2 U25 ( .A(n35), .Q(o_addr_nextpc[8]) );
  AOI220 U26 ( .A(i_addr_b[8]), .B(n2), .C(i_addr_jumpmux[8]), .D(n3), .Q(n35)
         );
  INV2 U27 ( .A(n53), .Q(o_addr_nextpc[20]) );
  INV2 U28 ( .A(n52), .Q(o_addr_nextpc[21]) );
  INV2 U29 ( .A(n51), .Q(o_addr_nextpc[22]) );
  INV2 U30 ( .A(n50), .Q(o_addr_nextpc[23]) );
  INV2 U31 ( .A(n49), .Q(o_addr_nextpc[24]) );
  INV2 U32 ( .A(n48), .Q(o_addr_nextpc[25]) );
  BUF2 U33 ( .A(n5), .Q(n3) );
  BUF2 U34 ( .A(n5), .Q(n4) );
  AOI221 U35 ( .A(i_addr_b[0]), .B(n1), .C(i_addr_jumpmux[0]), .D(n4), .Q(n65)
         );
  AOI221 U36 ( .A(i_addr_b[10]), .B(n1), .C(i_addr_jumpmux[10]), .D(n4), .Q(
        n64) );
  AOI221 U37 ( .A(i_addr_b[11]), .B(n1), .C(i_addr_jumpmux[11]), .D(n4), .Q(
        n63) );
  AOI221 U38 ( .A(i_addr_b[12]), .B(n1), .C(i_addr_jumpmux[12]), .D(n4), .Q(
        n62) );
  AOI221 U39 ( .A(i_addr_b[13]), .B(n1), .C(i_addr_jumpmux[13]), .D(n4), .Q(
        n61) );
  AOI221 U40 ( .A(i_addr_b[14]), .B(n1), .C(i_addr_jumpmux[14]), .D(n4), .Q(
        n60) );
  AOI221 U41 ( .A(i_addr_b[15]), .B(n1), .C(i_addr_jumpmux[15]), .D(n3), .Q(
        n59) );
  AOI221 U42 ( .A(i_addr_b[16]), .B(n1), .C(i_addr_jumpmux[16]), .D(n4), .Q(
        n58) );
  AOI221 U43 ( .A(i_addr_b[17]), .B(n1), .C(i_addr_jumpmux[17]), .D(n4), .Q(
        n57) );
  AOI221 U44 ( .A(i_addr_b[18]), .B(n1), .C(i_addr_jumpmux[18]), .D(n4), .Q(
        n56) );
  AOI221 U45 ( .A(i_addr_b[19]), .B(n1), .C(i_addr_jumpmux[19]), .D(n4), .Q(
        n55) );
  AOI221 U46 ( .A(i_addr_b[1]), .B(n2), .C(i_addr_jumpmux[1]), .D(n4), .Q(n54)
         );
  AOI221 U47 ( .A(i_addr_b[2]), .B(n2), .C(i_addr_jumpmux[2]), .D(n4), .Q(n43)
         );
  AOI221 U48 ( .A(i_addr_b[3]), .B(n2), .C(i_addr_jumpmux[3]), .D(n3), .Q(n40)
         );
  AOI221 U49 ( .A(i_addr_b[4]), .B(n2), .C(i_addr_jumpmux[4]), .D(n4), .Q(n39)
         );
  AOI221 U50 ( .A(i_addr_b[5]), .B(n2), .C(i_addr_jumpmux[5]), .D(n4), .Q(n38)
         );
  AOI221 U51 ( .A(i_addr_b[6]), .B(n2), .C(i_addr_jumpmux[6]), .D(n4), .Q(n37)
         );
  AOI221 U52 ( .A(i_addr_b[20]), .B(n2), .C(i_addr_jumpmux[20]), .D(n4), .Q(
        n53) );
  AOI221 U53 ( .A(i_addr_b[21]), .B(n2), .C(i_addr_jumpmux[21]), .D(n4), .Q(
        n52) );
  AOI221 U54 ( .A(i_addr_b[22]), .B(n2), .C(i_addr_jumpmux[22]), .D(n4), .Q(
        n51) );
  AOI221 U55 ( .A(i_addr_b[23]), .B(n2), .C(i_addr_jumpmux[23]), .D(n3), .Q(
        n50) );
  AOI221 U56 ( .A(i_addr_b[24]), .B(n2), .C(i_addr_jumpmux[24]), .D(n4), .Q(
        n49) );
  AOI221 U57 ( .A(i_addr_b[25]), .B(n2), .C(i_addr_jumpmux[25]), .D(n4), .Q(
        n48) );
  MUX22 U58 ( .A(i_addr_jumpmux[26]), .B(i_addr_b[26]), .S(n1), .Q(
        o_addr_nextpc[26]) );
  MUX22 U59 ( .A(i_addr_jumpmux[27]), .B(i_addr_b[27]), .S(n1), .Q(
        o_addr_nextpc[27]) );
  MUX22 U60 ( .A(i_addr_jumpmux[28]), .B(i_addr_b[28]), .S(n1), .Q(
        o_addr_nextpc[28]) );
  MUX22 U61 ( .A(i_addr_jumpmux[29]), .B(i_addr_b[29]), .S(n1), .Q(
        o_addr_nextpc[29]) );
  MUX22 U62 ( .A(i_addr_jumpmux[30]), .B(i_addr_b[30]), .S(n1), .Q(
        o_addr_nextpc[30]) );
  MUX22 U63 ( .A(i_addr_jumpmux[31]), .B(i_addr_b[31]), .S(n1), .Q(
        o_addr_nextpc[31]) );
endmodule


module F_pc ( i_clk, i_rst_n, i_con_stall, i_addr_next_pc, o_addr_pc );
  input [31:0] i_addr_next_pc;
  output [31:0] o_addr_pc;
  input i_clk, i_rst_n, i_con_stall;


  DFEC1 program_counter_reg_31_ ( .D(i_addr_next_pc[31]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[31]) );
  DFEC1 program_counter_reg_1_ ( .D(i_addr_next_pc[1]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[1]) );
  DFEC1 program_counter_reg_0_ ( .D(i_addr_next_pc[0]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[0]) );
  DFEC1 program_counter_reg_30_ ( .D(i_addr_next_pc[30]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[30]) );
  DFEC1 program_counter_reg_29_ ( .D(i_addr_next_pc[29]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[29]) );
  DFEC1 program_counter_reg_26_ ( .D(i_addr_next_pc[26]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[26]) );
  DFEC1 program_counter_reg_25_ ( .D(i_addr_next_pc[25]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[25]) );
  DFEC1 program_counter_reg_27_ ( .D(i_addr_next_pc[27]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[27]) );
  DFEC1 program_counter_reg_28_ ( .D(i_addr_next_pc[28]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[28]) );
  DFEC1 program_counter_reg_22_ ( .D(i_addr_next_pc[22]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[22]) );
  DFEC1 program_counter_reg_21_ ( .D(i_addr_next_pc[21]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[21]) );
  DFEC1 program_counter_reg_18_ ( .D(i_addr_next_pc[18]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[18]) );
  DFEC1 program_counter_reg_17_ ( .D(i_addr_next_pc[17]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[17]) );
  DFEC1 program_counter_reg_14_ ( .D(i_addr_next_pc[14]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[14]) );
  DFEC1 program_counter_reg_13_ ( .D(i_addr_next_pc[13]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[13]) );
  DFEC1 program_counter_reg_10_ ( .D(i_addr_next_pc[10]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[10]) );
  DFEC1 program_counter_reg_9_ ( .D(i_addr_next_pc[9]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[9]) );
  DFEC1 program_counter_reg_23_ ( .D(i_addr_next_pc[23]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[23]) );
  DFEC1 program_counter_reg_19_ ( .D(i_addr_next_pc[19]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[19]) );
  DFEC1 program_counter_reg_15_ ( .D(i_addr_next_pc[15]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[15]) );
  DFEC1 program_counter_reg_11_ ( .D(i_addr_next_pc[11]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[11]) );
  DFEC1 program_counter_reg_24_ ( .D(i_addr_next_pc[24]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[24]) );
  DFEC1 program_counter_reg_20_ ( .D(i_addr_next_pc[20]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[20]) );
  DFEC1 program_counter_reg_16_ ( .D(i_addr_next_pc[16]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[16]) );
  DFEC1 program_counter_reg_12_ ( .D(i_addr_next_pc[12]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[12]) );
  DFEC1 program_counter_reg_6_ ( .D(i_addr_next_pc[6]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[6]) );
  DFEC1 program_counter_reg_5_ ( .D(i_addr_next_pc[5]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[5]) );
  DFEC1 program_counter_reg_2_ ( .D(i_addr_next_pc[2]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[2]) );
  DFEC1 program_counter_reg_7_ ( .D(i_addr_next_pc[7]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[7]) );
  DFEC1 program_counter_reg_3_ ( .D(i_addr_next_pc[3]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[3]) );
  DFEC1 program_counter_reg_8_ ( .D(i_addr_next_pc[8]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[8]) );
  DFEC1 program_counter_reg_4_ ( .D(i_addr_next_pc[4]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[4]) );
endmodule


module F_add4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  NOR21 U2 ( .A(n81), .B(n82), .Q(n80) );
  INV3 U3 ( .A(n83), .Q(n81) );
  NOR31 U4 ( .A(n10), .B(n84), .C(n7), .Q(n83) );
  NAND22 U5 ( .A(n34), .B(n35), .Q(n33) );
  NOR31 U6 ( .A(n38), .B(n36), .C(n37), .Q(n35) );
  NOR21 U7 ( .A(n22), .B(n33), .Q(n21) );
  INV3 U8 ( .A(n23), .Q(n22) );
  NOR31 U9 ( .A(n26), .B(n24), .C(n25), .Q(n23) );
  XNR21 U10 ( .A(n29), .B(n25), .Q(SUM[26]) );
  NOR21 U11 ( .A(n26), .B(n30), .Q(n29) );
  INV3 U12 ( .A(n57), .Q(n46) );
  NAND31 U13 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  NOR21 U14 ( .A(n62), .B(n63), .Q(n58) );
  INV3 U15 ( .A(n61), .Q(n59) );
  XNR21 U16 ( .A(n31), .B(n26), .Q(SUM[25]) );
  XNR21 U17 ( .A(n68), .B(n63), .Q(SUM[13]) );
  XNR21 U18 ( .A(n55), .B(n50), .Q(SUM[17]) );
  XNR21 U19 ( .A(n43), .B(n38), .Q(SUM[21]) );
  XNR21 U20 ( .A(n66), .B(n62), .Q(SUM[14]) );
  XNR21 U21 ( .A(n53), .B(n49), .Q(SUM[18]) );
  XNR21 U22 ( .A(n41), .B(n37), .Q(SUM[22]) );
  XNR21 U23 ( .A(n77), .B(n74), .Q(SUM[10]) );
  NOR21 U24 ( .A(n78), .B(n2), .Q(n77) );
  NOR21 U25 ( .A(n50), .B(n54), .Q(n53) );
  NOR21 U26 ( .A(n63), .B(n67), .Q(n66) );
  NOR21 U27 ( .A(n38), .B(n42), .Q(n41) );
  XNR21 U28 ( .A(n1), .B(n2), .Q(SUM[9]) );
  XNR21 U29 ( .A(n9), .B(n10), .Q(SUM[5]) );
  XNR21 U30 ( .A(n6), .B(n7), .Q(SUM[6]) );
  INV3 U31 ( .A(n8), .Q(n6) );
  NAND22 U32 ( .A(n9), .B(A[5]), .Q(n8) );
  NAND22 U33 ( .A(A[3]), .B(A[2]), .Q(n82) );
  XNR21 U34 ( .A(A[29]), .B(n15), .Q(SUM[29]) );
  XOR21 U35 ( .A(A[30]), .B(n14), .Q(SUM[30]) );
  XOR21 U36 ( .A(n27), .B(n28), .Q(SUM[27]) );
  INV3 U37 ( .A(A[27]), .Q(n27) );
  NAND22 U38 ( .A(n29), .B(A[26]), .Q(n28) );
  XOR21 U39 ( .A(n12), .B(n13), .Q(SUM[31]) );
  INV3 U40 ( .A(A[31]), .Q(n12) );
  NAND22 U41 ( .A(A[30]), .B(n14), .Q(n13) );
  NOR21 U42 ( .A(n19), .B(n20), .Q(n18) );
  INV3 U43 ( .A(A[28]), .Q(n20) );
  NOR21 U44 ( .A(n71), .B(n3), .Q(n60) );
  INV3 U45 ( .A(n72), .Q(n71) );
  NOR31 U46 ( .A(n2), .B(n73), .C(n74), .Q(n72) );
  NAND22 U47 ( .A(A[11]), .B(A[8]), .Q(n73) );
  NOR21 U48 ( .A(n33), .B(n32), .Q(n31) );
  INV3 U49 ( .A(A[24]), .Q(n32) );
  INV3 U50 ( .A(A[5]), .Q(n10) );
  NOR21 U51 ( .A(n15), .B(n16), .Q(n14) );
  INV3 U52 ( .A(A[29]), .Q(n16) );
  INV3 U53 ( .A(A[6]), .Q(n7) );
  NAND22 U54 ( .A(A[7]), .B(A[4]), .Q(n84) );
  INV3 U55 ( .A(A[2]), .Q(SUM[2]) );
  INV3 U56 ( .A(n45), .Q(n34) );
  NAND22 U57 ( .A(n46), .B(n47), .Q(n45) );
  NOR31 U58 ( .A(n50), .B(n48), .C(n49), .Q(n47) );
  NAND22 U59 ( .A(A[19]), .B(A[16]), .Q(n48) );
  XNR21 U60 ( .A(A[28]), .B(n19), .Q(SUM[28]) );
  XNR21 U61 ( .A(A[12]), .B(n69), .Q(SUM[12]) );
  XNR21 U62 ( .A(A[16]), .B(n57), .Q(SUM[16]) );
  XNR21 U63 ( .A(A[20]), .B(n45), .Q(SUM[20]) );
  XNR21 U64 ( .A(A[24]), .B(n33), .Q(SUM[24]) );
  XOR21 U65 ( .A(n75), .B(n76), .Q(SUM[11]) );
  INV3 U66 ( .A(A[11]), .Q(n75) );
  NAND22 U67 ( .A(n77), .B(A[10]), .Q(n76) );
  XOR21 U68 ( .A(n64), .B(n65), .Q(SUM[15]) );
  INV3 U69 ( .A(A[15]), .Q(n64) );
  NAND22 U70 ( .A(n66), .B(A[14]), .Q(n65) );
  XOR21 U71 ( .A(n51), .B(n52), .Q(SUM[19]) );
  INV3 U72 ( .A(A[19]), .Q(n51) );
  NAND22 U73 ( .A(n53), .B(A[18]), .Q(n52) );
  XOR21 U74 ( .A(n39), .B(n40), .Q(SUM[23]) );
  INV3 U75 ( .A(A[23]), .Q(n39) );
  NAND22 U76 ( .A(n41), .B(A[22]), .Q(n40) );
  INV3 U77 ( .A(A[17]), .Q(n50) );
  INV3 U78 ( .A(A[21]), .Q(n38) );
  NOR21 U79 ( .A(n3), .B(n79), .Q(n1) );
  INV3 U80 ( .A(A[8]), .Q(n79) );
  INV3 U81 ( .A(A[9]), .Q(n2) );
  INV3 U82 ( .A(A[13]), .Q(n63) );
  INV3 U83 ( .A(A[14]), .Q(n62) );
  NOR21 U84 ( .A(n69), .B(n70), .Q(n68) );
  INV3 U85 ( .A(A[12]), .Q(n70) );
  INV3 U86 ( .A(A[10]), .Q(n74) );
  INV3 U87 ( .A(A[18]), .Q(n49) );
  INV3 U88 ( .A(A[22]), .Q(n37) );
  NOR21 U89 ( .A(n57), .B(n56), .Q(n55) );
  INV3 U90 ( .A(A[16]), .Q(n56) );
  NOR21 U91 ( .A(n45), .B(n44), .Q(n43) );
  INV3 U92 ( .A(A[20]), .Q(n44) );
  NAND22 U93 ( .A(A[23]), .B(A[20]), .Q(n36) );
  NAND22 U94 ( .A(A[27]), .B(A[24]), .Q(n24) );
  NAND22 U95 ( .A(A[15]), .B(A[12]), .Q(n61) );
  XNR21 U96 ( .A(A[4]), .B(n82), .Q(SUM[4]) );
  XNR21 U97 ( .A(A[8]), .B(n3), .Q(SUM[8]) );
  XOR21 U98 ( .A(n4), .B(n5), .Q(SUM[7]) );
  INV3 U99 ( .A(A[7]), .Q(n4) );
  NAND22 U100 ( .A(n6), .B(A[6]), .Q(n5) );
  NOR21 U101 ( .A(n82), .B(n11), .Q(n9) );
  INV3 U102 ( .A(A[4]), .Q(n11) );
  INV3 U103 ( .A(A[25]), .Q(n26) );
  INV3 U104 ( .A(A[26]), .Q(n25) );
  XOR21 U105 ( .A(A[3]), .B(A[2]), .Q(SUM[3]) );
  CLKIN3 U106 ( .A(n18), .Q(n15) );
  CLKIN3 U107 ( .A(n21), .Q(n19) );
  CLKIN3 U108 ( .A(n31), .Q(n30) );
  CLKIN3 U109 ( .A(n43), .Q(n42) );
  CLKIN3 U110 ( .A(n55), .Q(n54) );
  CLKIN3 U111 ( .A(n68), .Q(n67) );
  CLKIN3 U112 ( .A(n60), .Q(n69) );
  CLKIN3 U113 ( .A(n1), .Q(n78) );
  CLKIN3 U114 ( .A(n80), .Q(n3) );
endmodule


module F_add4 ( i_addr_pc, o_addr_pcadd4 );
  input [31:0] i_addr_pc;
  output [31:0] o_addr_pcadd4;
  wire   n2, n1;

  F_add4_DW01_add_1 add_5 ( .A(i_addr_pc), .B({n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n2, n1, n1}), .CI(n1), .SUM(o_addr_pcadd4) );
  LOGIC0 U3 ( .Q(n1) );
  LOGIC1 U4 ( .Q(n2) );
endmodule


module fetch ( i_clk, i_nrst, i_addr_b, i_addr_j, i_addr_jr, i_con_b, i_con_j, 
        i_data_instr, i_con_ifstall, o_addr_pc, o_addr_pc4, o_data_instr );
  input [31:0] i_addr_b;
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [1:0] i_con_j;
  input [31:0] i_data_instr;
  output [31:0] o_addr_pc;
  output [31:0] o_addr_pc4;
  output [31:0] o_data_instr;
  input i_clk, i_nrst, i_con_b, i_con_ifstall;

  wire   [31:0] jmux_i_addr_pc4;
  wire   [31:0] bmux_i_addr_jumpmux;
  wire   [31:0] pc_i_addr_next_pc;

  DFC3 pipe_instr_reg_31_ ( .D(i_data_instr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[31]) );
  DFC3 pipe_instr_reg_30_ ( .D(i_data_instr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[30]) );
  DFC3 pipe_instr_reg_29_ ( .D(i_data_instr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[29]) );
  DFC3 pipe_instr_reg_28_ ( .D(i_data_instr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[28]) );
  DFC3 pipe_instr_reg_27_ ( .D(i_data_instr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[27]) );
  DFC3 pipe_instr_reg_26_ ( .D(i_data_instr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[26]) );
  DFC3 pipe_instr_reg_25_ ( .D(i_data_instr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[25]) );
  DFC3 pipe_instr_reg_24_ ( .D(i_data_instr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[24]) );
  DFC3 pipe_instr_reg_23_ ( .D(i_data_instr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[23]) );
  DFC3 pipe_instr_reg_22_ ( .D(i_data_instr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[22]) );
  DFC3 pipe_instr_reg_21_ ( .D(i_data_instr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[21]) );
  DFC3 pipe_instr_reg_20_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[20]) );
  DFC3 pipe_instr_reg_19_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[19]) );
  DFC3 pipe_instr_reg_18_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[18]) );
  DFC3 pipe_instr_reg_17_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[17]) );
  DFC3 pipe_instr_reg_16_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[16]) );
  DFC3 pipe_instr_reg_15_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[15]) );
  DFC3 pipe_instr_reg_14_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[14]) );
  DFC3 pipe_instr_reg_13_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[13]) );
  DFC3 pipe_instr_reg_12_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[12]) );
  DFC3 pipe_instr_reg_11_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[11]) );
  DFC3 pipe_instr_reg_10_ ( .D(i_data_instr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[10]) );
  DFC3 pipe_instr_reg_9_ ( .D(i_data_instr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[9]) );
  DFC3 pipe_instr_reg_8_ ( .D(i_data_instr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[8]) );
  DFC3 pipe_instr_reg_7_ ( .D(i_data_instr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[7]) );
  DFC3 pipe_instr_reg_6_ ( .D(i_data_instr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[6]) );
  DFC3 pipe_instr_reg_5_ ( .D(i_data_instr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[5]) );
  DFC3 pipe_instr_reg_4_ ( .D(i_data_instr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[4]) );
  DFC3 pipe_instr_reg_3_ ( .D(i_data_instr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[3]) );
  DFC3 pipe_instr_reg_2_ ( .D(i_data_instr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[2]) );
  DFC3 pipe_instr_reg_1_ ( .D(i_data_instr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[1]) );
  DFC3 pipe_instr_reg_0_ ( .D(i_data_instr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(jmux_i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(jmux_i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(jmux_i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(jmux_i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(jmux_i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(jmux_i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(jmux_i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(jmux_i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(jmux_i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(jmux_i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(jmux_i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(jmux_i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(jmux_i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(jmux_i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(jmux_i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(jmux_i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(jmux_i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(jmux_i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(jmux_i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(jmux_i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(jmux_i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(jmux_i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(jmux_i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(jmux_i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(jmux_i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(jmux_i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(jmux_i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(jmux_i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(jmux_i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(jmux_i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(jmux_i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(jmux_i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  F_jumpmux u_jumpmux ( .i_addr_j(i_addr_j), .i_addr_jr(i_addr_jr), 
        .i_addr_pc4(jmux_i_addr_pc4), .i_con_jump(i_con_j), .o_addr_jumpmux(
        bmux_i_addr_jumpmux) );
  F_branchmux u_branchmux ( .i_addr_jumpmux(bmux_i_addr_jumpmux), .i_addr_b(
        i_addr_b), .i_con_ifbranch(i_con_b), .o_addr_nextpc(pc_i_addr_next_pc)
         );
  F_pc u_pc ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_con_stall(i_con_ifstall), 
        .i_addr_next_pc(pc_i_addr_next_pc), .o_addr_pc(o_addr_pc) );
  F_add4 u_add4 ( .i_addr_pc(o_addr_pc), .o_addr_pcadd4(jmux_i_addr_pc4) );
endmodule


module D_control ( o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite, 
        o_con_alusrc, o_con_regwrite, o_con_ifsign, o_con_loadsig, o_con_aluop, 
        i_con_instru );
  output [1:0] o_con_loadsig;
  output [5:0] o_con_aluop;
  input [5:0] i_con_instru;
  output o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite,
         o_con_alusrc, o_con_regwrite, o_con_ifsign;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n1, n2, n4, n5, n6, n7, n8, n9, n11, n12, n13, n15,
         n16, n17, n18, n19, n20;

  OAI212 U8 ( .A(i_con_instru[4]), .B(n26), .C(n25), .Q(o_con_memread) );
  OAI212 U24 ( .A(i_con_instru[4]), .B(n9), .C(n16), .Q(o_con_aluop[2]) );
  OAI2111 U2 ( .A(i_con_instru[4]), .B(n7), .C(n43), .D(n16), .Q(
        o_con_aluop[1]) );
  INV3 U3 ( .A(n46), .Q(n13) );
  NOR21 U4 ( .A(n27), .B(i_con_instru[4]), .Q(o_con_loadsig[1]) );
  INV3 U5 ( .A(o_con_aluop[5]), .Q(n16) );
  NAND22 U6 ( .A(n25), .B(n2), .Q(o_con_memtoreg) );
  INV3 U7 ( .A(o_con_memwrite), .Q(n2) );
  INV3 U9 ( .A(n43), .Q(o_con_aluop[4]) );
  INV3 U10 ( .A(n42), .Q(o_con_aluop[3]) );
  AOI211 U11 ( .A(n1), .B(n32), .C(o_con_aluop[4]), .Q(n42) );
  NAND31 U12 ( .A(n38), .B(n20), .C(n39), .Q(n27) );
  NAND31 U13 ( .A(n23), .B(n19), .C(n50), .Q(n34) );
  AOI2111 U14 ( .A(n1), .B(n6), .C(o_con_loadsig[0]), .D(o_con_loadsig[1]), 
        .Q(n25) );
  NAND22 U15 ( .A(n13), .B(n39), .Q(n40) );
  AOI311 U16 ( .A(n12), .B(n41), .C(n9), .D(i_con_instru[4]), .Q(
        o_con_aluop[0]) );
  NAND22 U17 ( .A(n50), .B(n20), .Q(n46) );
  NAND22 U18 ( .A(n44), .B(n45), .Q(n32) );
  NAND22 U19 ( .A(n13), .B(n18), .Q(n35) );
  NAND22 U20 ( .A(n36), .B(n1), .Q(n43) );
  NOR21 U21 ( .A(n41), .B(i_con_instru[4]), .Q(o_con_aluop[5]) );
  NOR21 U22 ( .A(n28), .B(i_con_instru[4]), .Q(o_con_loadsig[0]) );
  INV3 U23 ( .A(n41), .Q(n15) );
  INV3 U25 ( .A(n51), .Q(n12) );
  NAND31 U26 ( .A(n35), .B(n44), .C(n34), .Q(n51) );
  NOR21 U27 ( .A(i_con_instru[4]), .B(n31), .Q(o_con_alusrc) );
  NOR40 U28 ( .A(n15), .B(n11), .C(n32), .D(n30), .Q(n31) );
  INV3 U29 ( .A(n40), .Q(n11) );
  INV3 U30 ( .A(n47), .Q(n7) );
  NAND41 U31 ( .A(n12), .B(n48), .C(n45), .D(n40), .Q(n47) );
  NAND41 U32 ( .A(n20), .B(n19), .C(n18), .D(n8), .Q(n48) );
  INV3 U33 ( .A(n49), .Q(n9) );
  NAND31 U34 ( .A(n40), .B(n26), .C(n45), .Q(n49) );
  NOR40 U35 ( .A(n36), .B(n4), .C(n5), .D(n6), .Q(n21) );
  INV3 U36 ( .A(n27), .Q(n5) );
  INV3 U37 ( .A(n28), .Q(n4) );
  NOR31 U38 ( .A(n17), .B(i_con_instru[4]), .C(n8), .Q(o_con_memwrite) );
  NAND41 U39 ( .A(i_con_instru[2]), .B(i_con_instru[1]), .C(n50), .D(
        i_con_instru[0]), .Q(n26) );
  NAND41 U40 ( .A(n21), .B(n33), .C(n34), .D(n35), .Q(n30) );
  NAND22 U41 ( .A(i_con_instru[5]), .B(i_con_instru[3]), .Q(n33) );
  NAND31 U42 ( .A(n50), .B(n23), .C(i_con_instru[1]), .Q(n41) );
  OAI311 U43 ( .A(n46), .B(i_con_instru[2]), .C(n19), .D(n26), .Q(n36) );
  NAND31 U44 ( .A(i_con_instru[2]), .B(i_con_instru[1]), .C(n13), .Q(n45) );
  NOR21 U45 ( .A(n18), .B(i_con_instru[1]), .Q(n39) );
  NAND31 U46 ( .A(n38), .B(i_con_instru[0]), .C(n39), .Q(n28) );
  NOR21 U47 ( .A(n17), .B(i_con_instru[5]), .Q(n50) );
  INV3 U48 ( .A(i_con_instru[2]), .Q(n18) );
  NOR21 U49 ( .A(n20), .B(i_con_instru[2]), .Q(n23) );
  NAND31 U50 ( .A(n50), .B(i_con_instru[0]), .C(n39), .Q(n44) );
  INV3 U51 ( .A(i_con_instru[0]), .Q(n20) );
  INV3 U52 ( .A(i_con_instru[1]), .Q(n19) );
  AOI311 U53 ( .A(n21), .B(n7), .C(n22), .D(i_con_instru[4]), .Q(
        o_con_regwrite) );
  AOI311 U54 ( .A(n23), .B(n17), .C(i_con_instru[1]), .D(n15), .Q(n22) );
  NOR21 U55 ( .A(n8), .B(i_con_instru[3]), .Q(n38) );
  INV3 U56 ( .A(i_con_instru[3]), .Q(n17) );
  INV3 U57 ( .A(i_con_instru[5]), .Q(n8) );
  INV3 U58 ( .A(n29), .Q(o_con_ifsign) );
  NAND22 U59 ( .A(n1), .B(n30), .Q(n29) );
  INV3 U60 ( .A(n37), .Q(n6) );
  NAND31 U61 ( .A(i_con_instru[1]), .B(n23), .C(n38), .Q(n37) );
  NOR40 U62 ( .A(n24), .B(i_con_instru[3]), .C(i_con_instru[5]), .D(
        i_con_instru[4]), .Q(o_con_regdst) );
  NAND31 U63 ( .A(n19), .B(n18), .C(n20), .Q(n24) );
  INV3 U64 ( .A(i_con_instru[4]), .Q(n1) );
endmodule


module D_jb_control ( o_con_jump, o_con_bop, o_con_aluPC4, o_con_ifstall, 
        i_con_instru, i_con_func, i_con_rt );
  output [1:0] o_con_jump;
  output [2:0] o_con_bop;
  input [5:0] i_con_instru;
  input [5:0] i_con_func;
  input i_con_rt;
  output o_con_aluPC4, o_con_ifstall;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n2, n3, n4,
         n5, n6;

  OAI222 U13 ( .A(n5), .B(n16), .C(n14), .D(n17), .Q(o_con_bop[1]) );
  NAND31 U3 ( .A(n5), .B(n3), .C(n6), .Q(n8) );
  NAND22 U4 ( .A(n7), .B(n8), .Q(o_con_jump[1]) );
  INV3 U5 ( .A(n7), .Q(n2) );
  INV3 U6 ( .A(n13), .Q(o_con_ifstall) );
  AOI211 U7 ( .A(n3), .B(n14), .C(n2), .Q(n13) );
  NAND22 U8 ( .A(n7), .B(n4), .Q(n17) );
  OAI311 U9 ( .A(n4), .B(n2), .C(n14), .D(n16), .Q(o_con_bop[0]) );
  OAI2111 U10 ( .A(n9), .B(n8), .C(n10), .D(n7), .Q(o_con_jump[0]) );
  NOR40 U11 ( .A(n11), .B(i_con_func[2]), .C(i_con_func[5]), .D(i_con_func[4]), 
        .Q(n9) );
  NAND22 U12 ( .A(i_con_instru[1]), .B(n3), .Q(n10) );
  NAND22 U14 ( .A(n12), .B(i_con_func[3]), .Q(n11) );
  NOR31 U15 ( .A(i_con_instru[3]), .B(i_con_instru[5]), .C(i_con_instru[4]), 
        .Q(n7) );
  INV3 U16 ( .A(i_con_instru[1]), .Q(n5) );
  INV3 U17 ( .A(i_con_instru[2]), .Q(n3) );
  INV3 U18 ( .A(i_con_instru[0]), .Q(n6) );
  NOR21 U19 ( .A(i_con_func[1]), .B(i_con_func[0]), .Q(n12) );
  NAND22 U20 ( .A(i_con_instru[0]), .B(n5), .Q(n14) );
  NOR40 U21 ( .A(i_con_instru[2]), .B(n2), .C(n5), .D(n6), .Q(o_con_aluPC4) );
  NAND31 U22 ( .A(n7), .B(n6), .C(i_con_instru[2]), .Q(n16) );
  NOR31 U23 ( .A(n15), .B(n2), .C(n6), .Q(o_con_bop[2]) );
  XNR21 U24 ( .A(n5), .B(i_con_instru[2]), .Q(n15) );
  INV3 U25 ( .A(n18), .Q(n4) );
  NOR21 U26 ( .A(i_con_instru[2]), .B(i_con_rt), .Q(n18) );
endmodule


module D_pcadd_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258;

  NAND22 U2 ( .A(n30), .B(n27), .Q(n31) );
  NAND22 U3 ( .A(n204), .B(n214), .Q(n221) );
  NAND22 U4 ( .A(n169), .B(n179), .Q(n188) );
  NAND22 U5 ( .A(n133), .B(n143), .Q(n154) );
  NAND22 U6 ( .A(n100), .B(n108), .Q(n119) );
  NAND22 U7 ( .A(n79), .B(n82), .Q(n89) );
  INV3 U8 ( .A(B[23]), .Q(n6) );
  XOR21 U9 ( .A(n22), .B(n24), .Q(SUM[6]) );
  NOR21 U10 ( .A(n248), .B(n25), .Q(n24) );
  INV3 U11 ( .A(B[30]), .Q(n9) );
  NAND31 U12 ( .A(n230), .B(n231), .C(n232), .Q(n228) );
  NOR21 U13 ( .A(n244), .B(n245), .Q(n231) );
  NOR21 U14 ( .A(n25), .B(n246), .Q(n230) );
  NAND31 U15 ( .A(n71), .B(n72), .C(n73), .Q(n70) );
  NOR21 U16 ( .A(n75), .B(n76), .Q(n72) );
  NOR21 U17 ( .A(n77), .B(n78), .Q(n71) );
  INV3 U18 ( .A(n74), .Q(n73) );
  AOI211 U19 ( .A(n237), .B(n42), .C(n43), .Q(n233) );
  XNR21 U20 ( .A(n89), .B(n88), .Q(SUM[26]) );
  INV3 U21 ( .A(n211), .Q(n210) );
  AOI211 U22 ( .A(n212), .B(n204), .C(n213), .Q(n211) );
  INV3 U23 ( .A(n214), .Q(n213) );
  INV3 U24 ( .A(n176), .Q(n175) );
  AOI211 U25 ( .A(n177), .B(n169), .C(n178), .Q(n176) );
  INV3 U26 ( .A(n179), .Q(n178) );
  INV3 U27 ( .A(n140), .Q(n139) );
  AOI211 U28 ( .A(n141), .B(n133), .C(n142), .Q(n140) );
  INV3 U29 ( .A(n143), .Q(n142) );
  INV3 U30 ( .A(n26), .Q(n248) );
  AOI211 U31 ( .A(n80), .B(n79), .C(n81), .Q(n68) );
  INV3 U32 ( .A(n82), .Q(n81) );
  AOI211 U33 ( .A(n106), .B(n100), .C(n107), .Q(n103) );
  INV3 U34 ( .A(n108), .Q(n107) );
  XNR21 U35 ( .A(n188), .B(n187), .Q(SUM[14]) );
  XNR21 U36 ( .A(n221), .B(n220), .Q(SUM[10]) );
  XOR21 U37 ( .A(n193), .B(n189), .Q(SUM[13]) );
  NAND22 U38 ( .A(n190), .B(n181), .Q(n193) );
  XOR21 U39 ( .A(n158), .B(n155), .Q(SUM[17]) );
  NAND22 U40 ( .A(n156), .B(n145), .Q(n158) );
  XOR21 U41 ( .A(n123), .B(n120), .Q(SUM[21]) );
  NAND22 U42 ( .A(n121), .B(n111), .Q(n123) );
  XOR21 U43 ( .A(n93), .B(n90), .Q(SUM[25]) );
  NAND22 U44 ( .A(n91), .B(n84), .Q(n93) );
  NAND22 U45 ( .A(n144), .B(n160), .Q(n159) );
  NAND22 U46 ( .A(n161), .B(n134), .Q(n160) );
  INV3 U47 ( .A(n162), .Q(n161) );
  XNR21 U48 ( .A(n154), .B(n153), .Q(SUM[18]) );
  XNR21 U49 ( .A(n119), .B(n118), .Q(SUM[22]) );
  INV3 U50 ( .A(n79), .Q(n78) );
  XNR21 U51 ( .A(n31), .B(n29), .Q(SUM[5]) );
  XOR21 U52 ( .A(n10), .B(n11), .Q(SUM[9]) );
  NAND22 U53 ( .A(n12), .B(n13), .Q(n10) );
  NAND22 U54 ( .A(n27), .B(n28), .Q(n22) );
  NAND22 U55 ( .A(n29), .B(n30), .Q(n28) );
  XOR21 U56 ( .A(n41), .B(n54), .Q(SUM[2]) );
  NOR21 U57 ( .A(n43), .B(n55), .Q(n54) );
  XNR21 U58 ( .A(n58), .B(n149), .Q(SUM[1]) );
  NAND22 U59 ( .A(n59), .B(n56), .Q(n149) );
  INV3 U60 ( .A(n144), .Q(n184) );
  NAND22 U61 ( .A(n56), .B(n57), .Q(n41) );
  NAND22 U62 ( .A(n58), .B(n59), .Q(n57) );
  INV3 U63 ( .A(n150), .Q(n58) );
  AOI311 U64 ( .A(n99), .B(n100), .C(n101), .D(n102), .Q(n74) );
  NOR31 U65 ( .A(n109), .B(n112), .C(n113), .Q(n99) );
  NOR21 U66 ( .A(B[20]), .B(A[20]), .Q(n112) );
  OAI2111 U67 ( .A(n226), .B(n227), .C(n228), .D(n229), .Q(n205) );
  NOR21 U68 ( .A(A[7]), .B(B[7]), .Q(n227) );
  NAND22 U69 ( .A(B[7]), .B(A[7]), .Q(n229) );
  AOI211 U70 ( .A(n247), .B(n23), .C(n248), .Q(n226) );
  NAND22 U71 ( .A(B[29]), .B(A[29]), .Q(n53) );
  NOR21 U72 ( .A(A[29]), .B(B[29]), .Q(n52) );
  NAND22 U73 ( .A(n253), .B(n254), .Q(n204) );
  INV3 U74 ( .A(A[10]), .Q(n254) );
  INV3 U75 ( .A(B[10]), .Q(n253) );
  NOR21 U76 ( .A(n66), .B(n67), .Q(n62) );
  INV3 U77 ( .A(n85), .Q(n66) );
  NAND22 U78 ( .A(B[27]), .B(A[27]), .Q(n85) );
  NAND22 U79 ( .A(B[2]), .B(A[2]), .Q(n238) );
  NAND22 U80 ( .A(B[10]), .B(A[10]), .Q(n214) );
  XOR21 U81 ( .A(n44), .B(n45), .Q(SUM[31]) );
  XNR21 U82 ( .A(B[31]), .B(A[31]), .Q(n44) );
  AOI211 U83 ( .A(n46), .B(n47), .C(n48), .Q(n45) );
  NOR21 U84 ( .A(n49), .B(n9), .Q(n48) );
  XOR21 U85 ( .A(n86), .B(n87), .Q(SUM[27]) );
  XNR21 U86 ( .A(B[27]), .B(A[27]), .Q(n86) );
  AOI211 U87 ( .A(n88), .B(n79), .C(n81), .Q(n87) );
  XOR21 U88 ( .A(n116), .B(n117), .Q(SUM[23]) );
  XNR21 U89 ( .A(B[23]), .B(A[23]), .Q(n116) );
  AOI211 U90 ( .A(n118), .B(n100), .C(n107), .Q(n117) );
  NAND22 U91 ( .A(n130), .B(n131), .Q(n101) );
  AOI221 U92 ( .A(A[19]), .B(B[19]), .C(n138), .D(n139), .Q(n130) );
  NAND31 U93 ( .A(n132), .B(n133), .C(n134), .Q(n131) );
  INV3 U94 ( .A(n146), .Q(n138) );
  NAND22 U95 ( .A(n166), .B(n167), .Q(n134) );
  AOI221 U96 ( .A(A[15]), .B(B[15]), .C(n174), .D(n175), .Q(n166) );
  NAND31 U97 ( .A(n168), .B(n169), .C(n170), .Q(n167) );
  INV3 U98 ( .A(n182), .Q(n174) );
  NAND22 U99 ( .A(B[5]), .B(A[5]), .Q(n27) );
  NAND22 U100 ( .A(B[4]), .B(A[4]), .Q(n34) );
  NAND22 U101 ( .A(B[8]), .B(A[8]), .Q(n19) );
  NAND22 U102 ( .A(B[12]), .B(A[12]), .Q(n180) );
  NOR21 U103 ( .A(A[24]), .B(B[24]), .Q(n95) );
  NOR21 U104 ( .A(B[4]), .B(A[4]), .Q(n244) );
  NAND22 U105 ( .A(B[9]), .B(A[9]), .Q(n13) );
  NAND22 U106 ( .A(B[17]), .B(A[17]), .Q(n145) );
  NAND22 U107 ( .A(n249), .B(n250), .Q(n23) );
  INV3 U108 ( .A(A[6]), .Q(n250) );
  INV3 U109 ( .A(B[6]), .Q(n249) );
  NOR21 U110 ( .A(A[20]), .B(B[20]), .Q(n126) );
  NAND22 U111 ( .A(B[28]), .B(A[28]), .Q(n64) );
  NOR21 U112 ( .A(A[28]), .B(B[28]), .Q(n63) );
  NOR21 U113 ( .A(B[7]), .B(A[7]), .Q(n245) );
  NAND22 U114 ( .A(B[6]), .B(A[6]), .Q(n26) );
  NAND22 U115 ( .A(n201), .B(n202), .Q(n170) );
  AOI221 U116 ( .A(A[11]), .B(B[11]), .C(n209), .D(n210), .Q(n201) );
  NAND31 U117 ( .A(n203), .B(n204), .C(n205), .Q(n202) );
  INV3 U118 ( .A(n215), .Q(n209) );
  INV3 U119 ( .A(n232), .Q(n32) );
  INV3 U120 ( .A(A[3]), .Q(n235) );
  INV3 U121 ( .A(B[3]), .Q(n236) );
  NOR31 U122 ( .A(n135), .B(n136), .C(n137), .Q(n132) );
  NOR21 U123 ( .A(B[16]), .B(A[16]), .Q(n136) );
  NOR21 U124 ( .A(B[19]), .B(A[19]), .Q(n137) );
  NOR31 U125 ( .A(n206), .B(n207), .C(n208), .Q(n203) );
  NOR21 U126 ( .A(B[11]), .B(A[11]), .Q(n207) );
  NOR21 U127 ( .A(B[8]), .B(A[8]), .Q(n208) );
  NAND22 U128 ( .A(n222), .B(n223), .Q(n12) );
  INV3 U129 ( .A(A[9]), .Q(n223) );
  INV3 U130 ( .A(B[9]), .Q(n222) );
  NAND22 U131 ( .A(n197), .B(n198), .Q(n190) );
  INV3 U132 ( .A(A[13]), .Q(n198) );
  INV3 U133 ( .A(B[13]), .Q(n197) );
  XOR21 U134 ( .A(n65), .B(n62), .Q(SUM[28]) );
  XNR21 U135 ( .A(B[28]), .B(A[28]), .Q(n65) );
  XOR21 U136 ( .A(n60), .B(n51), .Q(SUM[29]) );
  XNR21 U137 ( .A(B[29]), .B(A[29]), .Q(n60) );
  XOR21 U138 ( .A(n1), .B(n47), .Q(SUM[30]) );
  XOR21 U139 ( .A(B[30]), .B(A[30]), .Q(n1) );
  NOR21 U140 ( .A(A[3]), .B(B[3]), .Q(n234) );
  NAND22 U141 ( .A(n251), .B(n252), .Q(n30) );
  INV3 U142 ( .A(A[5]), .Q(n252) );
  INV3 U143 ( .A(B[5]), .Q(n251) );
  NAND22 U144 ( .A(n2), .B(n163), .Q(n156) );
  INV3 U145 ( .A(A[17]), .Q(n163) );
  INV3 U146 ( .A(B[17]), .Q(n2) );
  NAND22 U147 ( .A(n191), .B(n192), .Q(n169) );
  INV3 U148 ( .A(A[14]), .Q(n192) );
  INV3 U149 ( .A(B[14]), .Q(n191) );
  NAND22 U150 ( .A(B[16]), .B(A[16]), .Q(n144) );
  NAND22 U151 ( .A(B[14]), .B(A[14]), .Q(n179) );
  NAND22 U152 ( .A(B[18]), .B(A[18]), .Q(n143) );
  NAND22 U153 ( .A(B[22]), .B(A[22]), .Q(n108) );
  NAND22 U154 ( .A(B[26]), .B(A[26]), .Q(n82) );
  XOR21 U155 ( .A(n185), .B(n186), .Q(SUM[15]) );
  XNR21 U156 ( .A(B[15]), .B(A[15]), .Q(n185) );
  AOI211 U157 ( .A(n187), .B(n169), .C(n178), .Q(n186) );
  XOR21 U158 ( .A(n151), .B(n152), .Q(SUM[19]) );
  XNR21 U159 ( .A(B[19]), .B(A[19]), .Q(n151) );
  AOI211 U160 ( .A(n153), .B(n133), .C(n142), .Q(n152) );
  NAND22 U161 ( .A(B[20]), .B(A[20]), .Q(n110) );
  NAND22 U162 ( .A(B[24]), .B(A[24]), .Q(n83) );
  NAND22 U163 ( .A(B[13]), .B(A[13]), .Q(n181) );
  NAND22 U164 ( .A(B[21]), .B(A[21]), .Q(n111) );
  NAND22 U165 ( .A(B[25]), .B(A[25]), .Q(n84) );
  NOR21 U166 ( .A(A[8]), .B(B[8]), .Q(n225) );
  NOR21 U167 ( .A(A[12]), .B(B[12]), .Q(n196) );
  NOR31 U168 ( .A(n171), .B(n172), .C(n173), .Q(n168) );
  NOR21 U169 ( .A(B[15]), .B(A[15]), .Q(n173) );
  NOR21 U170 ( .A(B[12]), .B(A[12]), .Q(n172) );
  NAND22 U171 ( .A(n4), .B(n127), .Q(n121) );
  INV3 U172 ( .A(A[21]), .Q(n127) );
  INV3 U173 ( .A(B[21]), .Q(n4) );
  XOR21 U174 ( .A(n218), .B(n219), .Q(SUM[11]) );
  XNR21 U175 ( .A(B[11]), .B(A[11]), .Q(n218) );
  AOI211 U176 ( .A(n220), .B(n204), .C(n213), .Q(n219) );
  NOR21 U177 ( .A(B[23]), .B(A[23]), .Q(n113) );
  NOR21 U178 ( .A(A[15]), .B(B[15]), .Q(n182) );
  NOR21 U179 ( .A(A[11]), .B(B[11]), .Q(n215) );
  NOR21 U180 ( .A(A[19]), .B(B[19]), .Q(n146) );
  NOR21 U181 ( .A(A[23]), .B(B[23]), .Q(n104) );
  IMUX21 U182 ( .A(n97), .B(n98), .S(n74), .Q(SUM[24]) );
  XNR21 U183 ( .A(B[24]), .B(A[24]), .Q(n98) );
  NOR21 U184 ( .A(n114), .B(n115), .Q(n97) );
  NOR21 U185 ( .A(B[24]), .B(A[24]), .Q(n114) );
  IMUX21 U186 ( .A(n128), .B(n129), .S(n125), .Q(SUM[20]) );
  XNR21 U187 ( .A(B[20]), .B(A[20]), .Q(n129) );
  NOR21 U188 ( .A(n147), .B(n148), .Q(n128) );
  NOR21 U189 ( .A(B[20]), .B(A[20]), .Q(n147) );
  NAND22 U190 ( .A(n5), .B(n122), .Q(n100) );
  INV3 U191 ( .A(A[22]), .Q(n122) );
  INV3 U192 ( .A(B[22]), .Q(n5) );
  NAND22 U193 ( .A(n8), .B(n92), .Q(n79) );
  INV3 U194 ( .A(A[26]), .Q(n92) );
  INV3 U195 ( .A(B[26]), .Q(n8) );
  NAND22 U196 ( .A(n3), .B(n157), .Q(n133) );
  INV3 U197 ( .A(A[18]), .Q(n157) );
  INV3 U198 ( .A(B[18]), .Q(n3) );
  NAND22 U199 ( .A(n7), .B(n96), .Q(n91) );
  INV3 U200 ( .A(A[25]), .Q(n96) );
  INV3 U201 ( .A(B[25]), .Q(n7) );
  NOR21 U202 ( .A(A[4]), .B(B[4]), .Q(n33) );
  NOR21 U203 ( .A(A[16]), .B(B[16]), .Q(n162) );
  NOR21 U204 ( .A(B[24]), .B(A[24]), .Q(n75) );
  XOR21 U205 ( .A(n20), .B(n21), .Q(SUM[7]) );
  XNR21 U206 ( .A(B[7]), .B(A[7]), .Q(n20) );
  AOI211 U207 ( .A(n22), .B(n23), .C(n248), .Q(n21) );
  NOR21 U208 ( .A(B[27]), .B(A[27]), .Q(n76) );
  NOR21 U209 ( .A(A[27]), .B(B[27]), .Q(n69) );
  IMUX21 U210 ( .A(n164), .B(n165), .S(n134), .Q(SUM[16]) );
  NOR21 U211 ( .A(n183), .B(n184), .Q(n165) );
  XNR21 U212 ( .A(B[16]), .B(A[16]), .Q(n164) );
  NOR21 U213 ( .A(B[16]), .B(A[16]), .Q(n183) );
  IMUX21 U214 ( .A(n14), .B(n15), .S(n16), .Q(SUM[8]) );
  NOR21 U215 ( .A(n17), .B(n18), .Q(n14) );
  XNR21 U216 ( .A(B[8]), .B(A[8]), .Q(n15) );
  NOR21 U217 ( .A(B[8]), .B(A[8]), .Q(n17) );
  IMUX21 U218 ( .A(n199), .B(n200), .S(n195), .Q(SUM[12]) );
  NOR21 U219 ( .A(n216), .B(n217), .Q(n199) );
  XNR21 U220 ( .A(B[12]), .B(A[12]), .Q(n200) );
  NOR21 U221 ( .A(B[12]), .B(A[12]), .Q(n216) );
  INV3 U222 ( .A(A[23]), .Q(n105) );
  INV3 U223 ( .A(n50), .Q(n46) );
  NOR21 U224 ( .A(A[30]), .B(B[30]), .Q(n50) );
  NAND22 U225 ( .A(n242), .B(n243), .Q(n42) );
  INV3 U226 ( .A(A[2]), .Q(n243) );
  INV3 U227 ( .A(B[2]), .Q(n242) );
  XOR21 U228 ( .A(n39), .B(n40), .Q(SUM[3]) );
  XNR21 U229 ( .A(B[3]), .B(A[3]), .Q(n39) );
  AOI211 U230 ( .A(n41), .B(n42), .C(n43), .Q(n40) );
  IMUX21 U231 ( .A(n35), .B(n36), .S(n32), .Q(SUM[4]) );
  NOR21 U232 ( .A(n37), .B(n38), .Q(n35) );
  XNR21 U233 ( .A(B[4]), .B(A[4]), .Q(n36) );
  NOR21 U234 ( .A(B[4]), .B(A[4]), .Q(n37) );
  INV3 U235 ( .A(B[0]), .Q(n255) );
  INV3 U236 ( .A(n257), .Q(n256) );
  NOR21 U237 ( .A(B[0]), .B(n258), .Q(n257) );
  INV3 U238 ( .A(A[30]), .Q(n49) );
  INV3 U239 ( .A(A[0]), .Q(n258) );
  NAND22 U240 ( .A(n240), .B(n241), .Q(n59) );
  INV3 U241 ( .A(B[1]), .Q(n240) );
  INV3 U242 ( .A(A[1]), .Q(n241) );
  NAND22 U243 ( .A(B[1]), .B(A[1]), .Q(n56) );
  NAND22 U244 ( .A(B[0]), .B(A[0]), .Q(n150) );
  CLKIN3 U245 ( .A(n19), .Q(n18) );
  OAI212 U246 ( .A(n32), .B(n33), .C(n34), .Q(n29) );
  CLKIN3 U247 ( .A(n34), .Q(n38) );
  OAI212 U248 ( .A(n51), .B(n52), .C(n53), .Q(n47) );
  CLKIN3 U249 ( .A(n42), .Q(n55) );
  CLKIN3 U250 ( .A(n61), .Q(n51) );
  OAI212 U251 ( .A(n62), .B(n63), .C(n64), .Q(n61) );
  OAI212 U252 ( .A(n68), .B(n69), .C(n70), .Q(n67) );
  OAI212 U253 ( .A(n77), .B(n83), .C(n84), .Q(n80) );
  OAI212 U254 ( .A(n77), .B(n90), .C(n84), .Q(n88) );
  CLKIN3 U255 ( .A(n91), .Q(n77) );
  CLKIN3 U256 ( .A(n94), .Q(n90) );
  OAI212 U257 ( .A(n74), .B(n95), .C(n83), .Q(n94) );
  OAI222 U258 ( .A(n103), .B(n104), .C(n6), .D(n105), .Q(n102) );
  OAI212 U259 ( .A(n109), .B(n110), .C(n111), .Q(n106) );
  CLKIN3 U260 ( .A(n83), .Q(n115) );
  OAI212 U261 ( .A(n109), .B(n120), .C(n111), .Q(n118) );
  CLKIN3 U262 ( .A(n121), .Q(n109) );
  CLKIN3 U263 ( .A(n124), .Q(n120) );
  OAI212 U264 ( .A(n125), .B(n126), .C(n110), .Q(n124) );
  CLKIN3 U265 ( .A(n101), .Q(n125) );
  OAI212 U266 ( .A(n135), .B(n144), .C(n145), .Q(n141) );
  CLKIN3 U267 ( .A(n110), .Q(n148) );
  OAI212 U268 ( .A(n135), .B(n155), .C(n145), .Q(n153) );
  CLKIN3 U269 ( .A(n156), .Q(n135) );
  CLKIN3 U270 ( .A(n159), .Q(n155) );
  OAI212 U271 ( .A(n171), .B(n180), .C(n181), .Q(n177) );
  OAI212 U272 ( .A(n171), .B(n189), .C(n181), .Q(n187) );
  CLKIN3 U273 ( .A(n190), .Q(n171) );
  CLKIN3 U274 ( .A(n194), .Q(n189) );
  OAI212 U275 ( .A(n195), .B(n196), .C(n180), .Q(n194) );
  CLKIN3 U276 ( .A(n170), .Q(n195) );
  OAI212 U277 ( .A(n206), .B(n19), .C(n13), .Q(n212) );
  CLKIN3 U278 ( .A(n180), .Q(n217) );
  OAI212 U279 ( .A(n11), .B(n206), .C(n13), .Q(n220) );
  CLKIN3 U280 ( .A(n12), .Q(n206) );
  CLKIN3 U281 ( .A(n224), .Q(n11) );
  OAI212 U282 ( .A(n16), .B(n225), .C(n19), .Q(n224) );
  CLKIN3 U283 ( .A(n205), .Q(n16) );
  OAI222 U284 ( .A(n233), .B(n234), .C(n235), .D(n236), .Q(n232) );
  CLKIN3 U285 ( .A(n238), .Q(n43) );
  OAI212 U286 ( .A(n239), .B(n150), .C(n56), .Q(n237) );
  CLKIN3 U287 ( .A(n59), .Q(n239) );
  CLKIN3 U288 ( .A(n23), .Q(n25) );
  OAI212 U289 ( .A(n246), .B(n34), .C(n27), .Q(n247) );
  CLKIN3 U290 ( .A(n30), .Q(n246) );
  OAI212 U291 ( .A(A[0]), .B(n255), .C(n256), .Q(SUM[0]) );
endmodule


module D_pcadd ( i_addr_pcadd4E, i_data_immshiftl, o_addr_pcbranchE );
  input [31:0] i_addr_pcadd4E;
  input [31:0] i_data_immshiftl;
  output [31:0] o_addr_pcbranchE;
  wire   n1;

  D_pcadd_DW01_add_1 add_5 ( .A(i_addr_pcadd4E), .B(i_data_immshiftl), .CI(n1), 
        .SUM(o_addr_pcbranchE) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_addr_Rt, i_con_RegWr, 
        i_addr_Rd, i_data_Rd, o_data_Rs, o_data_Rt );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rt;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr;
  wire   n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883;
  wire   [1023:0] regs;

  DFEC1 regs_reg_30__31_ ( .D(i_data_Rd[31]), .E(n854), .C(i_clk), .RN(n829), 
        .Q(regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(i_data_Rd[30]), .E(n854), .C(i_clk), .RN(n829), 
        .Q(regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(n820), .E(n854), .C(i_clk), .RN(n829), .Q(
        regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(i_data_Rd[28]), .E(n854), .C(i_clk), .RN(n829), 
        .Q(regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(i_data_Rd[27]), .E(n854), .C(i_clk), .RN(n830), 
        .Q(regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(i_data_Rd[26]), .E(n854), .C(i_clk), .RN(n830), 
        .Q(regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(i_data_Rd[25]), .E(n854), .C(i_clk), .RN(n830), 
        .Q(regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(i_data_Rd[24]), .E(n854), .C(i_clk), .RN(n830), 
        .Q(regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(n806), .E(n854), .C(i_clk), .RN(n830), .Q(
        regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(i_data_Rd[22]), .E(n854), .C(i_clk), .RN(n830), 
        .Q(regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(n801), .E(n854), .C(i_clk), .RN(n830), .Q(
        regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(n797), .E(n854), .C(i_clk), .RN(n830), .Q(
        regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n854), .C(i_clk), .RN(n830), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(i_data_Rd[18]), .E(n854), .C(i_clk), .RN(n831), 
        .Q(regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(n787), .E(n854), .C(i_clk), .RN(n831), .Q(
        regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(n783), .E(n854), .C(i_clk), .RN(n831), .Q(
        regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(n779), .E(n854), .C(i_clk), .RN(n831), .Q(
        regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(n775), .E(n854), .C(i_clk), .RN(n831), .Q(
        regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(i_data_Rd[13]), .E(n854), .C(i_clk), .RN(n831), 
        .Q(regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(n772), .E(n854), .C(i_clk), .RN(n831), .Q(
        regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(n768), .E(n854), .C(i_clk), .RN(n831), .Q(
        regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(n765), .E(n854), .C(i_clk), .RN(n831), .Q(
        regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(i_data_Rd[9]), .E(n854), .C(i_clk), .RN(n832), 
        .Q(regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(i_data_Rd[8]), .E(n854), .C(i_clk), .RN(n832), 
        .Q(regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(i_data_Rd[7]), .E(n854), .C(i_clk), .RN(n832), 
        .Q(regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n854), .C(i_clk), .RN(n832), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(i_data_Rd[5]), .E(n854), .C(i_clk), .RN(n832), 
        .Q(regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(i_data_Rd[4]), .E(n854), .C(i_clk), .RN(n832), 
        .Q(regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(n744), .E(n854), .C(i_clk), .RN(n832), .Q(
        regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(i_data_Rd[2]), .E(n854), .C(i_clk), .RN(n832), 
        .Q(regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n854), .C(i_clk), .RN(n832), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(n734), .E(n854), .C(i_clk), .RN(n833), .Q(
        regs[960]) );
  DFEC1 regs_reg_26__31_ ( .D(i_data_Rd[31]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(i_data_Rd[30]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(n820), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(i_data_Rd[28]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(i_data_Rd[27]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(i_data_Rd[26]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(i_data_Rd[25]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(i_data_Rd[24]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(n806), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(i_data_Rd[22]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(n801), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(n797), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(i_data_Rd[18]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(n787), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(n783), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(n779), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(n775), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(i_data_Rd[13]), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(n772), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(n768), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(n765), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(i_data_Rd[9]), .E(n858), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(i_data_Rd[8]), .E(n858), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(i_data_Rd[7]), .E(n858), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n858), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(i_data_Rd[5]), .E(n858), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(i_data_Rd[4]), .E(n858), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(n744), .E(n858), .C(i_clk), .RN(i_rst_n), .Q(
        regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(i_data_Rd[2]), .E(n858), .C(i_clk), .RN(n833), 
        .Q(regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n858), .C(i_clk), .RN(n834), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(n734), .E(n858), .C(i_clk), .RN(n826), .Q(
        regs[832]) );
  DFEC1 regs_reg_22__31_ ( .D(i_data_Rd[31]), .E(n847), .C(i_clk), .RN(n840), 
        .Q(regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(i_data_Rd[30]), .E(n847), .C(i_clk), .RN(n826), 
        .Q(regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(n819), .E(n847), .C(i_clk), .RN(n827), .Q(
        regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(i_data_Rd[28]), .E(n847), .C(i_clk), .RN(n828), 
        .Q(regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(n815), .E(n847), .C(i_clk), .RN(n829), .Q(
        regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(i_data_Rd[26]), .E(n847), .C(i_clk), .RN(n830), 
        .Q(regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(i_data_Rd[25]), .E(n847), .C(i_clk), .RN(n831), 
        .Q(regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(n809), .E(n847), .C(i_clk), .RN(n832), .Q(
        regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(n805), .E(n847), .C(i_clk), .RN(n833), .Q(
        regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(n804), .E(n847), .C(i_clk), .RN(n837), .Q(
        regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(n800), .E(n847), .C(i_clk), .RN(n838), .Q(
        regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(n796), .E(n847), .C(i_clk), .RN(n839), .Q(
        regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(n793), .E(n847), .C(i_clk), .RN(n840), .Q(
        regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(n790), .E(n847), .C(i_clk), .RN(n826), .Q(
        regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(n786), .E(n847), .C(i_clk), .RN(n829), .Q(
        regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(n782), .E(n847), .C(i_clk), .RN(n830), .Q(
        regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(n778), .E(n847), .C(i_clk), .RN(n827), .Q(
        regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(i_data_Rd[14]), .E(n847), .C(i_clk), .RN(n828), 
        .Q(regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(i_data_Rd[13]), .E(n847), .C(i_clk), .RN(i_rst_n), .Q(regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(n771), .E(n847), .C(i_clk), .RN(n845), .Q(
        regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(i_data_Rd[11]), .E(n847), .C(i_clk), .RN(i_rst_n), .Q(regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(n764), .E(n847), .C(i_clk), .RN(n842), .Q(
        regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(n762), .E(n847), .C(i_clk), .RN(n832), .Q(
        regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(n759), .E(n847), .C(i_clk), .RN(n844), .Q(
        regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(n756), .E(n847), .C(i_clk), .RN(n843), .Q(
        regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(n753), .E(n847), .C(i_clk), .RN(n842), .Q(
        regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(n750), .E(n847), .C(i_clk), .RN(i_rst_n), .Q(
        regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(n747), .E(n847), .C(i_clk), .RN(n831), .Q(
        regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(n743), .E(n847), .C(i_clk), .RN(n832), .Q(
        regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(n740), .E(n847), .C(i_clk), .RN(n833), .Q(
        regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(n737), .E(n847), .C(i_clk), .RN(n834), .Q(
        regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(n733), .E(n847), .C(i_clk), .RN(n835), .Q(
        regs[704]) );
  DFEC1 regs_reg_18__31_ ( .D(i_data_Rd[31]), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(i_data_Rd[30]), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(n819), .E(n851), .C(i_clk), .RN(n840), .Q(
        regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(i_data_Rd[28]), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(n815), .E(n851), .C(i_clk), .RN(n829), .Q(
        regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(i_data_Rd[26]), .E(n851), .C(i_clk), .RN(n830), 
        .Q(regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(i_data_Rd[25]), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(n809), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(n805), .E(n851), .C(i_clk), .RN(n837), .Q(
        regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(n804), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(n800), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(n796), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(n793), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(n790), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(n786), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(n782), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(n778), .E(n851), .C(i_clk), .RN(n836), .Q(
        regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(i_data_Rd[14]), .E(n851), .C(i_clk), .RN(n834), 
        .Q(regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(i_data_Rd[13]), .E(n851), .C(i_clk), .RN(n842), 
        .Q(regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(n771), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(i_data_Rd[11]), .E(n851), .C(i_clk), .RN(n844), 
        .Q(regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(n764), .E(n851), .C(i_clk), .RN(n843), .Q(
        regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(n762), .E(n851), .C(i_clk), .RN(n842), .Q(
        regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(n759), .E(n851), .C(i_clk), .RN(n845), .Q(
        regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(n756), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(n753), .E(n851), .C(i_clk), .RN(n837), .Q(
        regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(n750), .E(n851), .C(i_clk), .RN(n827), .Q(
        regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(n747), .E(n851), .C(i_clk), .RN(n828), .Q(
        regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(n743), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(n740), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(n737), .E(n851), .C(i_clk), .RN(i_rst_n), .Q(
        regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(n733), .E(n851), .C(i_clk), .RN(n834), .Q(
        regs[576]) );
  DFEC1 regs_reg_14__31_ ( .D(n824), .E(n864), .C(i_clk), .RN(n837), .Q(
        regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(n822), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(n818), .E(n864), .C(i_clk), .RN(n845), .Q(
        regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(n816), .E(n864), .C(i_clk), .RN(n845), .Q(
        regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(n814), .E(n864), .C(i_clk), .RN(n833), .Q(
        regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(n812), .E(n864), .C(i_clk), .RN(n842), .Q(
        regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(i_data_Rd[25]), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(n808), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(i_data_Rd[23]), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(n803), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(n799), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(n795), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(n792), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(n789), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(n785), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(n781), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(n777), .E(n864), .C(i_clk), .RN(n825), .Q(
        regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n864), .C(i_clk), .RN(n841), 
        .Q(regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(n774), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(n770), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(n767), .E(n864), .C(i_clk), .RN(n841), .Q(
        regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(n761), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(n758), .E(n864), .C(i_clk), .RN(n843), .Q(
        regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(n755), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(n752), .E(n864), .C(i_clk), .RN(n833), .Q(
        regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(n749), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(n746), .E(n864), .C(i_clk), .RN(n843), .Q(
        regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(n742), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(n739), .E(n864), .C(i_clk), .RN(i_rst_n), .Q(
        regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(n736), .E(n864), .C(i_clk), .RN(n831), .Q(
        regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(n732), .E(n864), .C(i_clk), .RN(n829), .Q(
        regs[448]) );
  DFEC1 regs_reg_10__31_ ( .D(n824), .E(n868), .C(i_clk), .RN(n835), .Q(
        regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(n822), .E(n868), .C(i_clk), .RN(n845), .Q(
        regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(n818), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(n816), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(n814), .E(n868), .C(i_clk), .RN(n834), .Q(
        regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(n812), .E(n868), .C(i_clk), .RN(n825), .Q(
        regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(i_data_Rd[25]), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(n808), .E(n868), .C(i_clk), .RN(n845), .Q(
        regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(i_data_Rd[23]), .E(n868), .C(i_clk), .RN(n844), 
        .Q(regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(n803), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(n799), .E(n868), .C(i_clk), .RN(n832), .Q(
        regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(n795), .E(n868), .C(i_clk), .RN(n844), .Q(
        regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(n792), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(n789), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(n785), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(n781), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(n777), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n868), .C(i_clk), .RN(n845), 
        .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(n774), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(n770), .E(n868), .C(i_clk), .RN(n825), .Q(
        regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(n767), .E(n868), .C(i_clk), .RN(n836), .Q(
        regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n868), .C(i_clk), .RN(n844), 
        .Q(regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(n761), .E(n868), .C(i_clk), .RN(n839), .Q(
        regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(n758), .E(n868), .C(i_clk), .RN(n837), .Q(
        regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(n755), .E(n868), .C(i_clk), .RN(n835), .Q(
        regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(n752), .E(n868), .C(i_clk), .RN(n825), .Q(
        regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(n749), .E(n868), .C(i_clk), .RN(n839), .Q(
        regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(n746), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(n742), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(n739), .E(n868), .C(i_clk), .RN(n830), .Q(
        regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(n736), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(n732), .E(n868), .C(i_clk), .RN(i_rst_n), .Q(
        regs[320]) );
  DFEC1 regs_reg_6__31_ ( .D(n823), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(n821), .E(n872), .C(i_clk), .RN(n845), .Q(
        regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(n817), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(i_data_Rd[28]), .E(n872), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(n813), .E(n872), .C(i_clk), .RN(n838), .Q(
        regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(n811), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(n810), .E(n872), .C(i_clk), .RN(n831), .Q(
        regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(n807), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(i_data_Rd[23]), .E(n872), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(n802), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(n798), .E(n872), .C(i_clk), .RN(n842), .Q(
        regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(n794), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(n791), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(n788), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(n784), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(n780), .E(n872), .C(i_clk), .RN(n845), .Q(
        regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(n776), .E(n872), .C(i_clk), .RN(n834), .Q(
        regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(i_data_Rd[14]), .E(n872), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(n773), .E(n872), .C(i_clk), .RN(n837), .Q(
        regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(n769), .E(n872), .C(i_clk), .RN(n843), .Q(
        regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(n766), .E(n872), .C(i_clk), .RN(n839), .Q(
        regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(n763), .E(n872), .C(i_clk), .RN(n840), .Q(
        regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(n760), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(n757), .E(n872), .C(i_clk), .RN(n844), .Q(
        regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(n754), .E(n872), .C(i_clk), .RN(n843), .Q(
        regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(n751), .E(n872), .C(i_clk), .RN(n842), .Q(
        regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(n748), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(n745), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(n741), .E(n872), .C(i_clk), .RN(n837), .Q(
        regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(n738), .E(n872), .C(i_clk), .RN(n828), .Q(
        regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(n735), .E(n872), .C(i_clk), .RN(n826), .Q(
        regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(n731), .E(n872), .C(i_clk), .RN(n827), .Q(
        regs[192]) );
  DFEC1 regs_reg_2__31_ ( .D(n823), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(n821), .E(n876), .C(i_clk), .RN(n827), .Q(
        regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(n817), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(i_data_Rd[28]), .E(n876), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(n813), .E(n876), .C(i_clk), .RN(n827), .Q(
        regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(n811), .E(n876), .C(i_clk), .RN(n840), .Q(
        regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(n810), .E(n876), .C(i_clk), .RN(n828), .Q(
        regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(n807), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(i_data_Rd[23]), .E(n876), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(n802), .E(n876), .C(i_clk), .RN(n836), .Q(
        regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(n798), .E(n876), .C(i_clk), .RN(n841), .Q(
        regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(n794), .E(n876), .C(i_clk), .RN(n839), .Q(
        regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(n791), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(n788), .E(n876), .C(i_clk), .RN(n825), .Q(
        regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(n784), .E(n876), .C(i_clk), .RN(n841), .Q(
        regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(n780), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(n776), .E(n876), .C(i_clk), .RN(n841), .Q(
        regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(i_data_Rd[14]), .E(n876), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(n773), .E(n876), .C(i_clk), .RN(n836), .Q(
        regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(n769), .E(n876), .C(i_clk), .RN(n835), .Q(
        regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(n766), .E(n876), .C(i_clk), .RN(n843), .Q(
        regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(n763), .E(n876), .C(i_clk), .RN(n825), .Q(
        regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(n760), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(n757), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(n754), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(n751), .E(n876), .C(i_clk), .RN(n842), .Q(regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(n748), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(n745), .E(n876), .C(i_clk), .RN(n825), .Q(regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(n741), .E(n876), .C(i_clk), .RN(n842), .Q(regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(n738), .E(n876), .C(i_clk), .RN(n835), .Q(regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(n735), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(n731), .E(n876), .C(i_clk), .RN(n834), .Q(regs[64]) );
  DFEC1 regs_reg_31__31_ ( .D(i_data_Rd[31]), .E(n861), .C(i_clk), .RN(n826), 
        .Q(regs[1023]) );
  DFEC1 regs_reg_31__30_ ( .D(i_data_Rd[30]), .E(n861), .C(i_clk), .RN(n826), 
        .Q(regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(n820), .E(n861), .C(i_clk), .RN(n826), .Q(
        regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(i_data_Rd[28]), .E(n861), .C(i_clk), .RN(n826), 
        .Q(regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(i_data_Rd[27]), .E(n861), .C(i_clk), .RN(n826), 
        .Q(regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(i_data_Rd[26]), .E(n861), .C(i_clk), .RN(n826), 
        .Q(regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(i_data_Rd[25]), .E(n861), .C(i_clk), .RN(n826), 
        .Q(regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(n809), .E(n861), .C(i_clk), .RN(n826), .Q(
        regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(n806), .E(n861), .C(i_clk), .RN(n826), .Q(
        regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(i_data_Rd[22]), .E(n861), .C(i_clk), .RN(n827), 
        .Q(regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(n801), .E(n861), .C(i_clk), .RN(n827), .Q(
        regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(n797), .E(n861), .C(i_clk), .RN(n827), .Q(
        regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n861), .C(i_clk), .RN(n827), 
        .Q(regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(i_data_Rd[18]), .E(n861), .C(i_clk), .RN(n827), 
        .Q(regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(n787), .E(n861), .C(i_clk), .RN(n827), .Q(
        regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(n783), .E(n861), .C(i_clk), .RN(n827), .Q(
        regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(n779), .E(n861), .C(i_clk), .RN(n827), .Q(
        regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(n775), .E(n861), .C(i_clk), .RN(n827), .Q(
        regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(i_data_Rd[13]), .E(n861), .C(i_clk), .RN(n828), 
        .Q(regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(n772), .E(n861), .C(i_clk), .RN(n828), .Q(
        regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(n768), .E(n861), .C(i_clk), .RN(n828), .Q(
        regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(n765), .E(n861), .C(i_clk), .RN(n828), .Q(
        regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(i_data_Rd[9]), .E(n861), .C(i_clk), .RN(n828), 
        .Q(regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(i_data_Rd[8]), .E(n861), .C(i_clk), .RN(n828), 
        .Q(regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(i_data_Rd[7]), .E(n861), .C(i_clk), .RN(n828), 
        .Q(regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n861), .C(i_clk), .RN(n828), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(i_data_Rd[5]), .E(n861), .C(i_clk), .RN(n828), 
        .Q(regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(i_data_Rd[4]), .E(n861), .C(i_clk), .RN(n829), 
        .Q(regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(n744), .E(n861), .C(i_clk), .RN(n829), .Q(
        regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(i_data_Rd[2]), .E(n861), .C(i_clk), .RN(n829), 
        .Q(regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n861), .C(i_clk), .RN(n829), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(n734), .E(n861), .C(i_clk), .RN(n829), .Q(
        regs[992]) );
  DFEC1 regs_reg_29__31_ ( .D(i_data_Rd[31]), .E(n855), .C(i_clk), .RN(n833), 
        .Q(regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(i_data_Rd[30]), .E(n855), .C(i_clk), .RN(n833), 
        .Q(regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(n820), .E(n855), .C(i_clk), .RN(n833), .Q(
        regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(i_data_Rd[28]), .E(n855), .C(i_clk), .RN(n833), 
        .Q(regs[956]) );
  DFEC1 regs_reg_29__27_ ( .D(i_data_Rd[27]), .E(n855), .C(i_clk), .RN(n833), 
        .Q(regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(i_data_Rd[26]), .E(n855), .C(i_clk), .RN(n833), 
        .Q(regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(i_data_Rd[25]), .E(n855), .C(i_clk), .RN(n833), 
        .Q(regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(n808), .E(n855), .C(i_clk), .RN(n833), .Q(
        regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(n806), .E(n855), .C(i_clk), .RN(n834), .Q(
        regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(i_data_Rd[22]), .E(n855), .C(i_clk), .RN(n834), 
        .Q(regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(n801), .E(n855), .C(i_clk), .RN(n834), .Q(
        regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(n797), .E(n855), .C(i_clk), .RN(n834), .Q(
        regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n855), .C(i_clk), .RN(n834), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(i_data_Rd[18]), .E(n855), .C(i_clk), .RN(n834), 
        .Q(regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(n787), .E(n855), .C(i_clk), .RN(n834), .Q(
        regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(n783), .E(n855), .C(i_clk), .RN(n834), .Q(
        regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(n779), .E(n855), .C(i_clk), .RN(n834), .Q(
        regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(n775), .E(n855), .C(i_clk), .RN(n835), .Q(
        regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(i_data_Rd[13]), .E(n855), .C(i_clk), .RN(n835), 
        .Q(regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(n772), .E(n855), .C(i_clk), .RN(n835), .Q(
        regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(n768), .E(n855), .C(i_clk), .RN(n835), .Q(
        regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(n765), .E(n855), .C(i_clk), .RN(n835), .Q(
        regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(i_data_Rd[9]), .E(n855), .C(i_clk), .RN(n835), 
        .Q(regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(i_data_Rd[8]), .E(n855), .C(i_clk), .RN(n835), 
        .Q(regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(i_data_Rd[7]), .E(n855), .C(i_clk), .RN(n835), 
        .Q(regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n855), .C(i_clk), .RN(n835), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(i_data_Rd[5]), .E(n855), .C(i_clk), .RN(n836), 
        .Q(regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(i_data_Rd[4]), .E(n855), .C(i_clk), .RN(n836), 
        .Q(regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(n744), .E(n855), .C(i_clk), .RN(n836), .Q(
        regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(i_data_Rd[2]), .E(n855), .C(i_clk), .RN(n836), 
        .Q(regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n855), .C(i_clk), .RN(n836), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(n734), .E(n855), .C(i_clk), .RN(n836), .Q(
        regs[928]) );
  DFEC1 regs_reg_28__31_ ( .D(i_data_Rd[31]), .E(n856), .C(i_clk), .RN(n836), 
        .Q(regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(i_data_Rd[30]), .E(n856), .C(i_clk), .RN(n836), 
        .Q(regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(n820), .E(n856), .C(i_clk), .RN(n836), .Q(
        regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(i_data_Rd[28]), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(i_data_Rd[27]), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(i_data_Rd[26]), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(i_data_Rd[25]), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(n807), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(
        regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(n806), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(
        regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(i_data_Rd[22]), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(n801), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(
        regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(n797), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(
        regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n856), .C(i_clk), .RN(n837), 
        .Q(regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(i_data_Rd[18]), .E(n856), .C(i_clk), .RN(n837), 
        .Q(regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(n787), .E(n856), .C(i_clk), .RN(n837), .Q(
        regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(n783), .E(n856), .C(i_clk), .RN(n837), .Q(
        regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(n779), .E(n856), .C(i_clk), .RN(n837), .Q(
        regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(n775), .E(n856), .C(i_clk), .RN(n837), .Q(
        regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(i_data_Rd[13]), .E(n856), .C(i_clk), .RN(n837), 
        .Q(regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(n772), .E(n856), .C(i_clk), .RN(n837), .Q(
        regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(n768), .E(n856), .C(i_clk), .RN(n837), .Q(
        regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(n765), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(
        regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(i_data_Rd[9]), .E(n856), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(i_data_Rd[8]), .E(n856), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(i_data_Rd[7]), .E(n856), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n856), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(i_data_Rd[5]), .E(n856), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(i_data_Rd[4]), .E(n856), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(n744), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(
        regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(i_data_Rd[2]), .E(n856), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n856), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(n734), .E(n856), .C(i_clk), .RN(i_rst_n), .Q(
        regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(i_data_Rd[31]), .E(n857), .C(i_clk), .RN(n838), 
        .Q(regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(i_data_Rd[30]), .E(n857), .C(i_clk), .RN(n837), 
        .Q(regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(n820), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(n816), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(i_data_Rd[27]), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(i_data_Rd[26]), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(i_data_Rd[25]), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(n809), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(n806), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(i_data_Rd[22]), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(n801), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(n797), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(i_data_Rd[18]), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(n787), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(n783), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(n779), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(n775), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(i_data_Rd[13]), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(n772), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(n768), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(n765), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(n762), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(i_data_Rd[8]), .E(n857), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(i_data_Rd[7]), .E(n857), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n857), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(i_data_Rd[5]), .E(n857), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(i_data_Rd[4]), .E(n857), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(n744), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(n740), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(n737), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(n734), .E(n857), .C(i_clk), .RN(i_rst_n), .Q(
        regs[864]) );
  DFEC1 regs_reg_25__31_ ( .D(i_data_Rd[31]), .E(n859), .C(i_clk), .RN(n827), 
        .Q(regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(i_data_Rd[30]), .E(n859), .C(i_clk), .RN(n828), 
        .Q(regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(n820), .E(n859), .C(i_clk), .RN(n829), .Q(
        regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(i_data_Rd[28]), .E(n859), .C(i_clk), .RN(n830), 
        .Q(regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(i_data_Rd[27]), .E(n859), .C(i_clk), .RN(n831), 
        .Q(regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(i_data_Rd[26]), .E(n859), .C(i_clk), .RN(n835), 
        .Q(regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(i_data_Rd[25]), .E(n859), .C(i_clk), .RN(i_rst_n), .Q(regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(n808), .E(n859), .C(i_clk), .RN(i_rst_n), .Q(
        regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(n806), .E(n859), .C(i_clk), .RN(i_rst_n), .Q(
        regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(i_data_Rd[22]), .E(n859), .C(i_clk), .RN(i_rst_n), .Q(regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(n801), .E(n859), .C(i_clk), .RN(i_rst_n), .Q(
        regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(n797), .E(n859), .C(i_clk), .RN(n844), .Q(
        regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(i_data_Rd[19]), .E(n859), .C(i_clk), .RN(i_rst_n), .Q(regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(i_data_Rd[18]), .E(n859), .C(i_clk), .RN(i_rst_n), .Q(regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(n787), .E(n859), .C(i_clk), .RN(n845), .Q(
        regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(n783), .E(n859), .C(i_clk), .RN(n828), .Q(
        regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(n779), .E(n859), .C(i_clk), .RN(i_rst_n), .Q(
        regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(n775), .E(n859), .C(i_clk), .RN(n842), .Q(
        regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(i_data_Rd[13]), .E(n859), .C(i_clk), .RN(n839), 
        .Q(regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(n772), .E(n859), .C(i_clk), .RN(n832), .Q(
        regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(n768), .E(n859), .C(i_clk), .RN(n833), .Q(
        regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(n765), .E(n859), .C(i_clk), .RN(n834), .Q(
        regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(n761), .E(n859), .C(i_clk), .RN(n826), .Q(
        regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(i_data_Rd[8]), .E(n859), .C(i_clk), .RN(n827), 
        .Q(regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(i_data_Rd[7]), .E(n859), .C(i_clk), .RN(n842), 
        .Q(regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(i_data_Rd[6]), .E(n859), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(i_data_Rd[5]), .E(n859), .C(i_clk), .RN(n826), 
        .Q(regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(i_data_Rd[4]), .E(n859), .C(i_clk), .RN(n827), 
        .Q(regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(n744), .E(n859), .C(i_clk), .RN(n838), .Q(
        regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(n739), .E(n859), .C(i_clk), .RN(n839), .Q(
        regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(n736), .E(n859), .C(i_clk), .RN(n840), .Q(
        regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(n734), .E(n859), .C(i_clk), .RN(n837), .Q(
        regs[800]) );
  DFEC1 regs_reg_24__31_ ( .D(i_data_Rd[31]), .E(n860), .C(i_clk), .RN(i_rst_n), .Q(regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(i_data_Rd[30]), .E(n860), .C(i_clk), .RN(i_rst_n), .Q(regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(n820), .E(n860), .C(i_clk), .RN(i_rst_n), .Q(
        regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(n816), .E(n860), .C(i_clk), .RN(n832), .Q(
        regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(i_data_Rd[27]), .E(n860), .C(i_clk), .RN(n825), 
        .Q(regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(i_data_Rd[26]), .E(n860), .C(i_clk), .RN(n833), 
        .Q(regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(n810), .E(n860), .C(i_clk), .RN(i_rst_n), .Q(
        regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(n807), .E(n860), .C(i_clk), .RN(n845), .Q(
        regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(n806), .E(n860), .C(i_clk), .RN(n844), .Q(
        regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(i_data_Rd[22]), .E(n860), .C(i_clk), .RN(n843), 
        .Q(regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(n801), .E(n860), .C(i_clk), .RN(n834), .Q(
        regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(n797), .E(n860), .C(i_clk), .RN(n826), .Q(
        regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(i_data_Rd[19]), .E(n860), .C(i_clk), .RN(n827), 
        .Q(regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(i_data_Rd[18]), .E(n860), .C(i_clk), .RN(n828), 
        .Q(regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(n787), .E(n860), .C(i_clk), .RN(n835), .Q(
        regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(n783), .E(n860), .C(i_clk), .RN(n836), .Q(
        regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(n779), .E(n860), .C(i_clk), .RN(n829), .Q(
        regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(n775), .E(n860), .C(i_clk), .RN(n830), .Q(
        regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(i_data_Rd[13]), .E(n860), .C(i_clk), .RN(n831), 
        .Q(regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(n772), .E(n860), .C(i_clk), .RN(n826), .Q(
        regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(n768), .E(n860), .C(i_clk), .RN(n827), .Q(
        regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(n765), .E(n860), .C(i_clk), .RN(n828), .Q(
        regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(n760), .E(n860), .C(i_clk), .RN(n829), .Q(
        regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(i_data_Rd[8]), .E(n860), .C(i_clk), .RN(n830), 
        .Q(regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(i_data_Rd[7]), .E(n860), .C(i_clk), .RN(n831), 
        .Q(regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(i_data_Rd[6]), .E(n860), .C(i_clk), .RN(n835), 
        .Q(regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(i_data_Rd[5]), .E(n860), .C(i_clk), .RN(n836), 
        .Q(regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(i_data_Rd[4]), .E(n860), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(n744), .E(n860), .C(i_clk), .RN(n842), .Q(
        regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(n738), .E(n860), .C(i_clk), .RN(i_rst_n), .Q(
        regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(n735), .E(n860), .C(i_clk), .RN(i_rst_n), .Q(
        regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(n734), .E(n860), .C(i_clk), .RN(i_rst_n), .Q(
        regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(i_data_Rd[31]), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(i_data_Rd[30]), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(n819), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(i_data_Rd[28]), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(n815), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(i_data_Rd[26]), .E(n846), .C(i_clk), .RN(n826), 
        .Q(regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(i_data_Rd[25]), .E(n846), .C(i_clk), .RN(n827), 
        .Q(regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(n809), .E(n846), .C(i_clk), .RN(n828), .Q(
        regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(n805), .E(n846), .C(i_clk), .RN(n829), .Q(
        regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(n804), .E(n846), .C(i_clk), .RN(n830), .Q(
        regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(n800), .E(n846), .C(i_clk), .RN(n831), .Q(
        regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(n796), .E(n846), .C(i_clk), .RN(n832), .Q(
        regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(n793), .E(n846), .C(i_clk), .RN(n833), .Q(
        regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(n790), .E(n846), .C(i_clk), .RN(n834), .Q(
        regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(n786), .E(n846), .C(i_clk), .RN(n842), .Q(
        regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(n782), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(n778), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(i_data_Rd[14]), .E(n846), .C(i_clk), .RN(n839), 
        .Q(regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(i_data_Rd[13]), .E(n846), .C(i_clk), .RN(n841), 
        .Q(regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(n771), .E(n846), .C(i_clk), .RN(n839), .Q(
        regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(i_data_Rd[11]), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(n764), .E(n846), .C(i_clk), .RN(n837), .Q(
        regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(n762), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(n759), .E(n846), .C(i_clk), .RN(n841), .Q(
        regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(n756), .E(n846), .C(i_clk), .RN(n844), .Q(
        regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(n753), .E(n846), .C(i_clk), .RN(n843), .Q(
        regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(n750), .E(n846), .C(i_clk), .RN(n842), .Q(
        regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(n747), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(n743), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(n740), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(n737), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(n733), .E(n846), .C(i_clk), .RN(i_rst_n), .Q(
        regs[736]) );
  DFEC1 regs_reg_21__31_ ( .D(i_data_Rd[31]), .E(n848), .C(i_clk), .RN(n836), 
        .Q(regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(i_data_Rd[30]), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(n819), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(i_data_Rd[28]), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(n815), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(i_data_Rd[26]), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(i_data_Rd[25]), .E(n848), .C(i_clk), .RN(n840), 
        .Q(regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(n809), .E(n848), .C(i_clk), .RN(n828), .Q(
        regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(n805), .E(n848), .C(i_clk), .RN(n840), .Q(
        regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(n804), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(n800), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(n796), .E(n848), .C(i_clk), .RN(n825), .Q(
        regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(n793), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(n790), .E(n848), .C(i_clk), .RN(n835), .Q(
        regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(n786), .E(n848), .C(i_clk), .RN(n844), .Q(
        regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(n782), .E(n848), .C(i_clk), .RN(n843), .Q(
        regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(n778), .E(n848), .C(i_clk), .RN(n845), .Q(
        regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(i_data_Rd[14]), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(i_data_Rd[13]), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(n771), .E(n848), .C(i_clk), .RN(n843), .Q(
        regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(i_data_Rd[11]), .E(n848), .C(i_clk), .RN(n834), 
        .Q(regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(n764), .E(n848), .C(i_clk), .RN(n841), .Q(
        regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(n762), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(n759), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(n756), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(n753), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(n750), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(n747), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(n743), .E(n848), .C(i_clk), .RN(n837), .Q(
        regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(n740), .E(n848), .C(i_clk), .RN(n838), .Q(
        regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(n737), .E(n848), .C(i_clk), .RN(i_rst_n), .Q(
        regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(n733), .E(n848), .C(i_clk), .RN(n837), .Q(
        regs[672]) );
  DFEC1 regs_reg_20__31_ ( .D(i_data_Rd[31]), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(i_data_Rd[30]), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(n819), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(
        regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(i_data_Rd[28]), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(n815), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(
        regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(i_data_Rd[26]), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(i_data_Rd[25]), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(n809), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(
        regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(n805), .E(n849), .C(i_clk), .RN(n838), .Q(
        regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(n804), .E(n849), .C(i_clk), .RN(n839), .Q(
        regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(n800), .E(n849), .C(i_clk), .RN(n840), .Q(
        regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(n796), .E(n849), .C(i_clk), .RN(n826), .Q(
        regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(n793), .E(n849), .C(i_clk), .RN(n827), .Q(
        regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(n790), .E(n849), .C(i_clk), .RN(n828), .Q(
        regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(n786), .E(n849), .C(i_clk), .RN(n830), .Q(
        regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(n782), .E(n849), .C(i_clk), .RN(n831), .Q(
        regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(n778), .E(n849), .C(i_clk), .RN(n829), .Q(
        regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(i_data_Rd[14]), .E(n849), .C(i_clk), .RN(n836), 
        .Q(regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(i_data_Rd[13]), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(n771), .E(n849), .C(i_clk), .RN(n837), .Q(
        regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(i_data_Rd[11]), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(n764), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(
        regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(n762), .E(n849), .C(i_clk), .RN(n825), .Q(
        regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(n759), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(
        regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(n756), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(
        regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(n753), .E(n849), .C(i_clk), .RN(n841), .Q(
        regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(n750), .E(n849), .C(i_clk), .RN(i_rst_n), .Q(
        regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(n747), .E(n849), .C(i_clk), .RN(n826), .Q(
        regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(n743), .E(n849), .C(i_clk), .RN(n827), .Q(
        regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(n740), .E(n849), .C(i_clk), .RN(n828), .Q(
        regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(n737), .E(n849), .C(i_clk), .RN(n829), .Q(
        regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(n733), .E(n849), .C(i_clk), .RN(n830), .Q(
        regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(i_data_Rd[31]), .E(n850), .C(i_clk), .RN(n831), 
        .Q(regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(i_data_Rd[30]), .E(n850), .C(i_clk), .RN(n832), 
        .Q(regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(n819), .E(n850), .C(i_clk), .RN(n833), .Q(
        regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(i_data_Rd[28]), .E(n850), .C(i_clk), .RN(n844), 
        .Q(regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(n815), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(
        regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(i_data_Rd[26]), .E(n850), .C(i_clk), .RN(n836), 
        .Q(regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(i_data_Rd[25]), .E(n850), .C(i_clk), .RN(n832), 
        .Q(regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(n809), .E(n850), .C(i_clk), .RN(n838), .Q(
        regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(n805), .E(n850), .C(i_clk), .RN(n839), .Q(
        regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(n804), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(
        regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(n800), .E(n850), .C(i_clk), .RN(n836), .Q(
        regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(n796), .E(n850), .C(i_clk), .RN(n838), .Q(
        regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(n793), .E(n850), .C(i_clk), .RN(n838), .Q(
        regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(n790), .E(n850), .C(i_clk), .RN(n837), .Q(
        regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(n786), .E(n850), .C(i_clk), .RN(n826), .Q(
        regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(n782), .E(n850), .C(i_clk), .RN(n842), .Q(
        regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(n778), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(
        regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(i_data_Rd[14]), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(i_data_Rd[13]), .E(n850), .C(i_clk), .RN(n845), 
        .Q(regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(n771), .E(n850), .C(i_clk), .RN(n825), .Q(
        regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(i_data_Rd[11]), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(n764), .E(n850), .C(i_clk), .RN(n841), .Q(
        regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(n762), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(
        regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(n759), .E(n850), .C(i_clk), .RN(n844), .Q(
        regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(n756), .E(n850), .C(i_clk), .RN(n843), .Q(
        regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(n753), .E(n850), .C(i_clk), .RN(n842), .Q(
        regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(n750), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(
        regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(n747), .E(n850), .C(i_clk), .RN(n826), .Q(
        regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(n743), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(
        regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(n740), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(
        regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(n737), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(
        regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(n733), .E(n850), .C(i_clk), .RN(i_rst_n), .Q(
        regs[608]) );
  DFEC1 regs_reg_17__31_ ( .D(n824), .E(n852), .C(i_clk), .RN(n839), .Q(
        regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(n822), .E(n852), .C(i_clk), .RN(n845), .Q(
        regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(n819), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(i_data_Rd[28]), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(n815), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(n811), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(i_data_Rd[25]), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(n809), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(n805), .E(n852), .C(i_clk), .RN(n841), .Q(
        regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(n804), .E(n852), .C(i_clk), .RN(n835), .Q(
        regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(n800), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(n796), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(n793), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(n790), .E(n852), .C(i_clk), .RN(n838), .Q(
        regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(n786), .E(n852), .C(i_clk), .RN(n831), .Q(
        regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(n782), .E(n852), .C(i_clk), .RN(n841), .Q(
        regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(n778), .E(n852), .C(i_clk), .RN(n839), .Q(
        regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(i_data_Rd[14]), .E(n852), .C(i_clk), .RN(n840), 
        .Q(regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(n774), .E(n852), .C(i_clk), .RN(n845), .Q(
        regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(n771), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(i_data_Rd[11]), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(n764), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(n762), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(n759), .E(n852), .C(i_clk), .RN(n838), .Q(
        regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(n756), .E(n852), .C(i_clk), .RN(n842), .Q(
        regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(n753), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(n750), .E(n852), .C(i_clk), .RN(n839), .Q(
        regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(n747), .E(n852), .C(i_clk), .RN(n825), .Q(
        regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(n743), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(n740), .E(n852), .C(i_clk), .RN(n841), .Q(
        regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(n737), .E(n852), .C(i_clk), .RN(i_rst_n), .Q(
        regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(n733), .E(n852), .C(i_clk), .RN(n835), .Q(
        regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(n823), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(n821), .E(n853), .C(i_clk), .RN(n844), .Q(
        regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(n819), .E(n853), .C(i_clk), .RN(n843), .Q(
        regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(n816), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(n815), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(n812), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(i_data_Rd[25]), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(n809), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(n805), .E(n853), .C(i_clk), .RN(n844), .Q(
        regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(n804), .E(n853), .C(i_clk), .RN(n843), .Q(
        regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(n800), .E(n853), .C(i_clk), .RN(n826), .Q(
        regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(n796), .E(n853), .C(i_clk), .RN(n827), .Q(
        regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(n793), .E(n853), .C(i_clk), .RN(n828), .Q(
        regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(n790), .E(n853), .C(i_clk), .RN(n829), .Q(
        regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(n786), .E(n853), .C(i_clk), .RN(n830), .Q(
        regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(n782), .E(n853), .C(i_clk), .RN(n836), .Q(
        regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(n778), .E(n853), .C(i_clk), .RN(n842), .Q(
        regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(i_data_Rd[14]), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(n773), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(n771), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(i_data_Rd[11]), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(n764), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(n762), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(n759), .E(n853), .C(i_clk), .RN(n838), .Q(
        regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(n756), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(n753), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(n750), .E(n853), .C(i_clk), .RN(n845), .Q(
        regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(n747), .E(n853), .C(i_clk), .RN(n841), .Q(
        regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(n743), .E(n853), .C(i_clk), .RN(n845), .Q(
        regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(n740), .E(n853), .C(i_clk), .RN(n833), .Q(
        regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(n737), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(n733), .E(n853), .C(i_clk), .RN(i_rst_n), .Q(
        regs[512]) );
  DFEC1 regs_reg_15__31_ ( .D(n824), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(n822), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(n818), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(n816), .E(n863), .C(i_clk), .RN(n831), .Q(
        regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(n814), .E(n863), .C(i_clk), .RN(n845), .Q(
        regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(n812), .E(n863), .C(i_clk), .RN(n833), .Q(
        regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(i_data_Rd[25]), .E(n863), .C(i_clk), .RN(n834), 
        .Q(regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(n808), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(i_data_Rd[23]), .E(n863), .C(i_clk), .RN(n843), 
        .Q(regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(n803), .E(n863), .C(i_clk), .RN(n832), .Q(
        regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(n799), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(n795), .E(n863), .C(i_clk), .RN(n837), .Q(
        regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(n792), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(n789), .E(n863), .C(i_clk), .RN(n844), .Q(
        regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(n785), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(n781), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(n777), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(n774), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(n770), .E(n863), .C(i_clk), .RN(n826), .Q(
        regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(n767), .E(n863), .C(i_clk), .RN(n827), .Q(
        regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n863), .C(i_clk), .RN(n828), 
        .Q(regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(n761), .E(n863), .C(i_clk), .RN(n829), .Q(
        regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(n758), .E(n863), .C(i_clk), .RN(n830), .Q(
        regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(n755), .E(n863), .C(i_clk), .RN(n831), .Q(
        regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(n752), .E(n863), .C(i_clk), .RN(n832), .Q(
        regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(n749), .E(n863), .C(i_clk), .RN(n833), .Q(
        regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(n746), .E(n863), .C(i_clk), .RN(n834), .Q(
        regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(n742), .E(n863), .C(i_clk), .RN(n825), .Q(
        regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(n739), .E(n863), .C(i_clk), .RN(i_rst_n), .Q(
        regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(n736), .E(n863), .C(i_clk), .RN(n832), .Q(
        regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(n732), .E(n863), .C(i_clk), .RN(n834), .Q(
        regs[480]) );
  DFEC1 regs_reg_13__31_ ( .D(n824), .E(n865), .C(i_clk), .RN(n839), .Q(
        regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(n822), .E(n865), .C(i_clk), .RN(n834), .Q(
        regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(n818), .E(n865), .C(i_clk), .RN(n844), .Q(
        regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(n816), .E(n865), .C(i_clk), .RN(n843), .Q(
        regs[444]) );
  DFEC1 regs_reg_13__27_ ( .D(n814), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(n812), .E(n865), .C(i_clk), .RN(n840), .Q(
        regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(i_data_Rd[25]), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(n808), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(i_data_Rd[23]), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(n803), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(n799), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(n795), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(n792), .E(n865), .C(i_clk), .RN(n833), .Q(
        regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(n789), .E(n865), .C(i_clk), .RN(n839), .Q(
        regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(n785), .E(n865), .C(i_clk), .RN(n840), .Q(
        regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(n781), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(n777), .E(n865), .C(i_clk), .RN(n835), .Q(
        regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n865), .C(i_clk), .RN(n840), 
        .Q(regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(n774), .E(n865), .C(i_clk), .RN(n830), .Q(
        regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(n770), .E(n865), .C(i_clk), .RN(n836), .Q(
        regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(n767), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(n761), .E(n865), .C(i_clk), .RN(n835), .Q(
        regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(n758), .E(n865), .C(i_clk), .RN(n841), .Q(
        regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(n755), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(n752), .E(n865), .C(i_clk), .RN(n836), .Q(
        regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(n749), .E(n865), .C(i_clk), .RN(n832), .Q(
        regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(n746), .E(n865), .C(i_clk), .RN(n835), .Q(
        regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(n742), .E(n865), .C(i_clk), .RN(n832), .Q(
        regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(n739), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(n736), .E(n865), .C(i_clk), .RN(n843), .Q(
        regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(n732), .E(n865), .C(i_clk), .RN(i_rst_n), .Q(
        regs[416]) );
  DFEC1 regs_reg_12__31_ ( .D(n824), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(n822), .E(n866), .C(i_clk), .RN(n836), .Q(
        regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(n818), .E(n866), .C(i_clk), .RN(n841), .Q(
        regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(n816), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(n814), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(n812), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(i_data_Rd[25]), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(n808), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(n805), .E(n866), .C(i_clk), .RN(n843), .Q(
        regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(n803), .E(n866), .C(i_clk), .RN(n830), .Q(
        regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(n799), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(n795), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(n792), .E(n866), .C(i_clk), .RN(n838), .Q(
        regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(n789), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(n785), .E(n866), .C(i_clk), .RN(n829), .Q(
        regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(n781), .E(n866), .C(i_clk), .RN(n830), .Q(
        regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(n777), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n866), .C(i_clk), .RN(n832), 
        .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(n774), .E(n866), .C(i_clk), .RN(n833), .Q(
        regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(n770), .E(n866), .C(i_clk), .RN(n826), .Q(
        regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(n767), .E(n866), .C(i_clk), .RN(n827), .Q(
        regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n866), .C(i_clk), .RN(n828), 
        .Q(regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(n761), .E(n866), .C(i_clk), .RN(n840), .Q(
        regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(n758), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(n755), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(n752), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(n749), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(n746), .E(n866), .C(i_clk), .RN(n842), .Q(
        regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(n742), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(n739), .E(n866), .C(i_clk), .RN(n840), .Q(
        regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(n736), .E(n866), .C(i_clk), .RN(n832), .Q(
        regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(n732), .E(n866), .C(i_clk), .RN(i_rst_n), .Q(
        regs[384]) );
  DFEC1 regs_reg_11__31_ ( .D(n824), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(n822), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(n818), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(n816), .E(n867), .C(i_clk), .RN(n836), .Q(
        regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(n814), .E(n867), .C(i_clk), .RN(n844), .Q(
        regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(n812), .E(n867), .C(i_clk), .RN(n829), .Q(
        regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(i_data_Rd[25]), .E(n867), .C(i_clk), .RN(n838), 
        .Q(regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(n808), .E(n867), .C(i_clk), .RN(n839), .Q(
        regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(n806), .E(n867), .C(i_clk), .RN(n831), .Q(
        regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(n803), .E(n867), .C(i_clk), .RN(n834), .Q(
        regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(n799), .E(n867), .C(i_clk), .RN(n843), .Q(
        regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(n795), .E(n867), .C(i_clk), .RN(n833), .Q(
        regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(n792), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(n789), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(n785), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(n781), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(n777), .E(n867), .C(i_clk), .RN(n830), .Q(
        regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n867), .C(i_clk), .RN(n841), 
        .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(n774), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(n770), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(n767), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(n765), .E(n867), .C(i_clk), .RN(n834), .Q(
        regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(n761), .E(n867), .C(i_clk), .RN(n825), .Q(
        regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(n758), .E(n867), .C(i_clk), .RN(n841), .Q(
        regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(n755), .E(n867), .C(i_clk), .RN(n835), .Q(
        regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(n752), .E(n867), .C(i_clk), .RN(n834), .Q(
        regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(n749), .E(n867), .C(i_clk), .RN(n831), .Q(
        regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(n746), .E(n867), .C(i_clk), .RN(n836), .Q(
        regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(n742), .E(n867), .C(i_clk), .RN(n844), .Q(
        regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(n739), .E(n867), .C(i_clk), .RN(n836), .Q(
        regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(n736), .E(n867), .C(i_clk), .RN(i_rst_n), .Q(
        regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(n732), .E(n867), .C(i_clk), .RN(n835), .Q(
        regs[352]) );
  DFEC1 regs_reg_9__31_ ( .D(n824), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(n822), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(n818), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(n816), .E(n869), .C(i_clk), .RN(n844), .Q(
        regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(n814), .E(n869), .C(i_clk), .RN(n843), .Q(
        regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(n812), .E(n869), .C(i_clk), .RN(n842), .Q(
        regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(i_data_Rd[25]), .E(n869), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(n808), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(n805), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(n803), .E(n869), .C(i_clk), .RN(n845), .Q(
        regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(n799), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(n795), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(n792), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(n789), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(n785), .E(n869), .C(i_clk), .RN(n832), .Q(
        regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(n781), .E(n869), .C(i_clk), .RN(n842), .Q(
        regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(n777), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(n775), .E(n869), .C(i_clk), .RN(n842), .Q(
        regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(n774), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(n770), .E(n869), .C(i_clk), .RN(n845), .Q(
        regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(n767), .E(n869), .C(i_clk), .RN(n831), .Q(
        regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(n764), .E(n869), .C(i_clk), .RN(n825), .Q(
        regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(n761), .E(n869), .C(i_clk), .RN(n834), .Q(
        regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(n758), .E(n869), .C(i_clk), .RN(n825), .Q(
        regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(n755), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(n752), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(n749), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(n746), .E(n869), .C(i_clk), .RN(n829), .Q(
        regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(n742), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(n739), .E(n869), .C(i_clk), .RN(i_rst_n), .Q(
        regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(n736), .E(n869), .C(i_clk), .RN(n838), .Q(
        regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(n732), .E(n869), .C(i_clk), .RN(n831), .Q(
        regs[288]) );
  DFEC1 regs_reg_8__31_ ( .D(n824), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(n822), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(n818), .E(n870), .C(i_clk), .RN(n841), .Q(
        regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(n816), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(n814), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(n812), .E(n870), .C(i_clk), .RN(n844), .Q(
        regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(n810), .E(n870), .C(i_clk), .RN(n843), .Q(
        regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(n808), .E(n870), .C(i_clk), .RN(n842), .Q(
        regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(n806), .E(n870), .C(i_clk), .RN(n825), .Q(
        regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(n803), .E(n870), .C(i_clk), .RN(n845), .Q(
        regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(n799), .E(n870), .C(i_clk), .RN(n845), .Q(
        regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(n795), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(n792), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(n789), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(n785), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(n781), .E(n870), .C(i_clk), .RN(n833), .Q(
        regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(n777), .E(n870), .C(i_clk), .RN(n844), .Q(
        regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(i_data_Rd[14]), .E(n870), .C(i_clk), .RN(n843), 
        .Q(regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(n774), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(n770), .E(n870), .C(i_clk), .RN(n841), .Q(
        regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(n767), .E(n870), .C(i_clk), .RN(n842), .Q(
        regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(n763), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(n761), .E(n870), .C(i_clk), .RN(n829), .Q(
        regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(n758), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(n755), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(n752), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(n749), .E(n870), .C(i_clk), .RN(n830), .Q(
        regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(n746), .E(n870), .C(i_clk), .RN(n845), .Q(
        regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(n742), .E(n870), .C(i_clk), .RN(n836), .Q(
        regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(n739), .E(n870), .C(i_clk), .RN(n841), .Q(
        regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(n736), .E(n870), .C(i_clk), .RN(n835), .Q(
        regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(n732), .E(n870), .C(i_clk), .RN(n833), .Q(
        regs[256]) );
  DFEC1 regs_reg_7__31_ ( .D(n823), .E(n871), .C(i_clk), .RN(n828), .Q(
        regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(n821), .E(n871), .C(i_clk), .RN(n825), .Q(
        regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(n817), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(i_data_Rd[28]), .E(n871), .C(i_clk), .RN(n825), 
        .Q(regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(n813), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(n811), .E(n871), .C(i_clk), .RN(n835), .Q(
        regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(n810), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(n807), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(i_data_Rd[23]), .E(n871), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(n802), .E(n871), .C(i_clk), .RN(n832), .Q(
        regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(n798), .E(n871), .C(i_clk), .RN(n828), .Q(
        regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(n794), .E(n871), .C(i_clk), .RN(n842), .Q(
        regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(n791), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(n788), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(n784), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(n780), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(n776), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(i_data_Rd[14]), .E(n871), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(n773), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(n769), .E(n871), .C(i_clk), .RN(n825), .Q(
        regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(n766), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(n763), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(n760), .E(n871), .C(i_clk), .RN(n829), .Q(
        regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(n757), .E(n871), .C(i_clk), .RN(n830), .Q(
        regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(n754), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(n751), .E(n871), .C(i_clk), .RN(n841), .Q(
        regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(n748), .E(n871), .C(i_clk), .RN(n831), .Q(
        regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(n745), .E(n871), .C(i_clk), .RN(n825), .Q(
        regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(n741), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(n738), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(n735), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(n731), .E(n871), .C(i_clk), .RN(i_rst_n), .Q(
        regs[224]) );
  DFEC1 regs_reg_5__31_ ( .D(n823), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(n821), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(n817), .E(n873), .C(i_clk), .RN(n831), .Q(
        regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(i_data_Rd[28]), .E(n873), .C(i_clk), .RN(n838), 
        .Q(regs[188]) );
  DFEC1 regs_reg_5__27_ ( .D(n813), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(n811), .E(n873), .C(i_clk), .RN(n841), .Q(
        regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(n810), .E(n873), .C(i_clk), .RN(n841), .Q(
        regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(n807), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(n805), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(n802), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(n798), .E(n873), .C(i_clk), .RN(n828), .Q(
        regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(n794), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(n791), .E(n873), .C(i_clk), .RN(n845), .Q(
        regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(n788), .E(n873), .C(i_clk), .RN(n835), .Q(
        regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(n784), .E(n873), .C(i_clk), .RN(n843), .Q(
        regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(n780), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(n776), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(i_data_Rd[14]), .E(n873), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(n773), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(n769), .E(n873), .C(i_clk), .RN(n840), .Q(
        regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(n766), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(n763), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(n760), .E(n873), .C(i_clk), .RN(n825), .Q(
        regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(n757), .E(n873), .C(i_clk), .RN(n829), .Q(
        regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(n754), .E(n873), .C(i_clk), .RN(n827), .Q(
        regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(n751), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(n748), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(n745), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(n741), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(n738), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(n735), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(n731), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[160]) );
  DFEC1 regs_reg_4__31_ ( .D(n823), .E(n874), .C(i_clk), .RN(n837), .Q(
        regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(n821), .E(n874), .C(i_clk), .RN(n840), .Q(
        regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(n817), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(i_data_Rd[28]), .E(n874), .C(i_clk), .RN(n826), 
        .Q(regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(n813), .E(n874), .C(i_clk), .RN(n833), .Q(
        regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(n811), .E(n874), .C(i_clk), .RN(n844), .Q(
        regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(n810), .E(n874), .C(i_clk), .RN(n843), .Q(
        regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(n807), .E(n874), .C(i_clk), .RN(n842), .Q(
        regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(n806), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(n802), .E(n874), .C(i_clk), .RN(n844), .Q(
        regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(n798), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(n794), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(n791), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(n788), .E(n874), .C(i_clk), .RN(n830), .Q(
        regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(n784), .E(n874), .C(i_clk), .RN(n838), .Q(
        regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(n780), .E(n874), .C(i_clk), .RN(n837), .Q(
        regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(n776), .E(n874), .C(i_clk), .RN(n833), .Q(
        regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(i_data_Rd[14]), .E(n874), .C(i_clk), .RN(n826), 
        .Q(regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(n773), .E(n874), .C(i_clk), .RN(n836), .Q(
        regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(n769), .E(n874), .C(i_clk), .RN(n825), .Q(
        regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(n766), .E(n874), .C(i_clk), .RN(n838), .Q(
        regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(n763), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(n760), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(n757), .E(n874), .C(i_clk), .RN(n843), .Q(
        regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(n754), .E(n874), .C(i_clk), .RN(n841), .Q(
        regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(n751), .E(n874), .C(i_clk), .RN(n838), .Q(
        regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(n748), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(n745), .E(n874), .C(i_clk), .RN(n842), .Q(
        regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(n741), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(n738), .E(n874), .C(i_clk), .RN(n843), .Q(
        regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(n735), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(n731), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[128]) );
  DFEC1 regs_reg_3__31_ ( .D(n823), .E(n875), .C(i_clk), .RN(n837), .Q(
        regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(n821), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(n817), .E(n875), .C(i_clk), .RN(n840), .Q(
        regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(i_data_Rd[28]), .E(n875), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(n813), .E(n875), .C(i_clk), .RN(n825), .Q(
        regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(n811), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(n810), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(n807), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(i_data_Rd[23]), .E(n875), .C(i_clk), .RN(n841), 
        .Q(regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(n802), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(n798), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(n794), .E(n875), .C(i_clk), .RN(n843), .Q(
        regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(n791), .E(n875), .C(i_clk), .RN(n841), .Q(
        regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(n788), .E(n875), .C(i_clk), .RN(n844), .Q(
        regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(n784), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(n780), .E(n875), .C(i_clk), .RN(n844), .Q(
        regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(n776), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(i_data_Rd[14]), .E(n875), .C(i_clk), .RN(n844), 
        .Q(regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(n773), .E(n875), .C(i_clk), .RN(n827), .Q(
        regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(n769), .E(n875), .C(i_clk), .RN(n825), .Q(
        regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(n766), .E(n875), .C(i_clk), .RN(n845), .Q(
        regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(n763), .E(n875), .C(i_clk), .RN(n825), .Q(
        regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(n760), .E(n875), .C(i_clk), .RN(n829), .Q(
        regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(n757), .E(n875), .C(i_clk), .RN(n839), .Q(
        regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(n754), .E(n875), .C(i_clk), .RN(n837), .Q(
        regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(n751), .E(n875), .C(i_clk), .RN(n845), .Q(
        regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(n748), .E(n875), .C(i_clk), .RN(n845), .Q(
        regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(n745), .E(n875), .C(i_clk), .RN(n839), .Q(
        regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(n741), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(n738), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(n735), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(n731), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[96]) );
  DFEC1 regs_reg_1__31_ ( .D(n823), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(n821), .E(n877), .C(i_clk), .RN(n832), .Q(
        regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(n817), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(i_data_Rd[28]), .E(n877), .C(i_clk), .RN(n844), 
        .Q(regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(n813), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(n811), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(n810), .E(n877), .C(i_clk), .RN(n840), .Q(
        regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(n807), .E(n877), .C(i_clk), .RN(n825), .Q(
        regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(n805), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(n802), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(n798), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(n794), .E(n877), .C(i_clk), .RN(n826), .Q(
        regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(n791), .E(n877), .C(i_clk), .RN(n838), .Q(
        regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(n788), .E(n877), .C(i_clk), .RN(n838), .Q(
        regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(n784), .E(n877), .C(i_clk), .RN(n838), .Q(
        regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(n780), .E(n877), .C(i_clk), .RN(n838), .Q(
        regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(n776), .E(n877), .C(i_clk), .RN(n838), .Q(
        regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(i_data_Rd[14]), .E(n877), .C(i_clk), .RN(n838), 
        .Q(regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(n773), .E(n877), .C(i_clk), .RN(n838), .Q(
        regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(n769), .E(n877), .C(i_clk), .RN(n838), .Q(
        regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(n766), .E(n877), .C(i_clk), .RN(n838), .Q(
        regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(n763), .E(n877), .C(i_clk), .RN(n839), .Q(
        regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(n760), .E(n877), .C(i_clk), .RN(n839), .Q(regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(n757), .E(n877), .C(i_clk), .RN(n839), .Q(regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(n754), .E(n877), .C(i_clk), .RN(n839), .Q(regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(n751), .E(n877), .C(i_clk), .RN(n839), .Q(regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(n748), .E(n877), .C(i_clk), .RN(n839), .Q(regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(n745), .E(n877), .C(i_clk), .RN(n839), .Q(regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(n741), .E(n877), .C(i_clk), .RN(n839), .Q(regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(n738), .E(n877), .C(i_clk), .RN(n839), .Q(regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(n735), .E(n877), .C(i_clk), .RN(n840), .Q(regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(n731), .E(n877), .C(i_clk), .RN(n840), .Q(regs[32]) );
  DFEC1 regs_reg_0__31_ ( .D(n823), .E(n878), .C(i_clk), .RN(n840), .Q(
        regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(n821), .E(n878), .C(i_clk), .RN(n840), .Q(
        regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(n817), .E(n878), .C(i_clk), .RN(n840), .Q(
        regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(i_data_Rd[28]), .E(n878), .C(i_clk), .RN(n840), 
        .Q(regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(n813), .E(n878), .C(i_clk), .RN(n840), .Q(
        regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(n811), .E(n878), .C(i_clk), .RN(n840), .Q(
        regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(n810), .E(n878), .C(i_clk), .RN(n840), .Q(
        regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(n807), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(n806), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(n802), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(n798), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(n794), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(n791), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(n788), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(n784), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(n780), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(n776), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(n775), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(n773), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(n769), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(n766), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(n763), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(n760), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(n757), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(n754), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(n751), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(n748), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(n745), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(n741), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(n738), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(n735), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(n731), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(
        regs[0]) );
  BUF2 U2 ( .A(n840), .Q(n837) );
  BUF2 U3 ( .A(n825), .Q(n836) );
  BUF2 U4 ( .A(n845), .Q(n835) );
  BUF2 U5 ( .A(n842), .Q(n834) );
  BUF2 U6 ( .A(n842), .Q(n833) );
  BUF2 U7 ( .A(n842), .Q(n832) );
  BUF2 U8 ( .A(n843), .Q(n831) );
  BUF2 U9 ( .A(n843), .Q(n830) );
  BUF2 U10 ( .A(n843), .Q(n829) );
  BUF2 U11 ( .A(n844), .Q(n828) );
  BUF2 U12 ( .A(n844), .Q(n827) );
  BUF2 U13 ( .A(n844), .Q(n826) );
  BUF2 U14 ( .A(n841), .Q(n840) );
  BUF2 U15 ( .A(n841), .Q(n839) );
  BUF2 U16 ( .A(n841), .Q(n838) );
  BUF2 U17 ( .A(n845), .Q(n842) );
  BUF2 U18 ( .A(n835), .Q(n843) );
  BUF2 U19 ( .A(n836), .Q(n844) );
  BUF2 U20 ( .A(n845), .Q(n841) );
  BUF2 U21 ( .A(n385), .Q(n376) );
  BUF2 U22 ( .A(i_addr_Rt[0]), .Q(n377) );
  BUF2 U23 ( .A(n385), .Q(n378) );
  BUF2 U24 ( .A(n386), .Q(n379) );
  BUF2 U25 ( .A(n386), .Q(n380) );
  BUF2 U26 ( .A(n387), .Q(n381) );
  BUF2 U27 ( .A(n387), .Q(n382) );
  BUF2 U28 ( .A(n388), .Q(n383) );
  BUF2 U29 ( .A(n388), .Q(n384) );
  BUF2 U30 ( .A(n730), .Q(n719) );
  BUF2 U31 ( .A(i_addr_Rs[0]), .Q(n720) );
  BUF2 U32 ( .A(i_addr_Rs[0]), .Q(n721) );
  BUF2 U33 ( .A(n729), .Q(n722) );
  BUF2 U34 ( .A(n729), .Q(n723) );
  BUF2 U35 ( .A(n730), .Q(n724) );
  BUF2 U36 ( .A(n730), .Q(n725) );
  INV3 U37 ( .A(n40), .Q(n861) );
  NAND22 U38 ( .A(n41), .B(n42), .Q(n40) );
  BUF2 U39 ( .A(i_addr_Rt[1]), .Q(n371) );
  BUF2 U40 ( .A(n370), .Q(n372) );
  BUF2 U41 ( .A(n718), .Q(n714) );
  BUF2 U42 ( .A(n713), .Q(n715) );
  BUF2 U43 ( .A(n713), .Q(n716) );
  BUF2 U44 ( .A(n825), .Q(n845) );
  BUF2 U45 ( .A(i_rst_n), .Q(n825) );
  BUF2 U46 ( .A(i_data_Rd[0]), .Q(n731) );
  BUF2 U47 ( .A(i_data_Rd[1]), .Q(n735) );
  BUF2 U48 ( .A(i_data_Rd[2]), .Q(n738) );
  BUF2 U49 ( .A(i_data_Rd[3]), .Q(n741) );
  BUF2 U50 ( .A(i_data_Rd[4]), .Q(n745) );
  BUF2 U51 ( .A(i_data_Rd[5]), .Q(n748) );
  BUF2 U52 ( .A(i_data_Rd[6]), .Q(n751) );
  BUF2 U53 ( .A(i_data_Rd[7]), .Q(n754) );
  BUF2 U54 ( .A(i_data_Rd[8]), .Q(n757) );
  BUF2 U55 ( .A(i_data_Rd[9]), .Q(n760) );
  BUF2 U56 ( .A(i_data_Rd[10]), .Q(n763) );
  BUF2 U57 ( .A(i_data_Rd[11]), .Q(n766) );
  BUF2 U58 ( .A(i_data_Rd[12]), .Q(n769) );
  BUF2 U59 ( .A(i_data_Rd[13]), .Q(n773) );
  BUF2 U60 ( .A(i_data_Rd[15]), .Q(n776) );
  BUF2 U61 ( .A(i_data_Rd[0]), .Q(n732) );
  BUF2 U62 ( .A(i_data_Rd[1]), .Q(n736) );
  BUF2 U63 ( .A(i_data_Rd[2]), .Q(n739) );
  BUF2 U64 ( .A(i_data_Rd[3]), .Q(n742) );
  BUF2 U65 ( .A(i_data_Rd[4]), .Q(n746) );
  BUF2 U66 ( .A(i_data_Rd[5]), .Q(n749) );
  BUF2 U67 ( .A(i_data_Rd[6]), .Q(n752) );
  BUF2 U68 ( .A(i_data_Rd[7]), .Q(n755) );
  BUF2 U69 ( .A(i_data_Rd[8]), .Q(n758) );
  BUF2 U70 ( .A(i_data_Rd[9]), .Q(n761) );
  BUF2 U71 ( .A(i_data_Rd[11]), .Q(n767) );
  BUF2 U72 ( .A(i_data_Rd[12]), .Q(n770) );
  BUF2 U73 ( .A(i_data_Rd[13]), .Q(n774) );
  BUF2 U74 ( .A(i_data_Rd[15]), .Q(n777) );
  BUF2 U75 ( .A(i_data_Rd[0]), .Q(n733) );
  BUF2 U76 ( .A(i_data_Rd[1]), .Q(n737) );
  BUF2 U77 ( .A(i_data_Rd[2]), .Q(n740) );
  BUF2 U78 ( .A(i_data_Rd[3]), .Q(n743) );
  BUF2 U79 ( .A(i_data_Rd[4]), .Q(n747) );
  BUF2 U80 ( .A(i_data_Rd[5]), .Q(n750) );
  BUF2 U81 ( .A(i_data_Rd[6]), .Q(n753) );
  BUF2 U82 ( .A(i_data_Rd[7]), .Q(n756) );
  BUF2 U83 ( .A(i_data_Rd[8]), .Q(n759) );
  BUF2 U84 ( .A(i_data_Rd[9]), .Q(n762) );
  BUF2 U85 ( .A(i_data_Rd[10]), .Q(n764) );
  BUF2 U86 ( .A(i_data_Rd[12]), .Q(n771) );
  BUF2 U87 ( .A(i_data_Rd[15]), .Q(n778) );
  BUF2 U88 ( .A(i_data_Rd[0]), .Q(n734) );
  BUF2 U89 ( .A(i_data_Rd[3]), .Q(n744) );
  BUF2 U90 ( .A(i_data_Rd[10]), .Q(n765) );
  BUF2 U91 ( .A(i_data_Rd[11]), .Q(n768) );
  BUF2 U92 ( .A(i_data_Rd[12]), .Q(n772) );
  BUF2 U93 ( .A(i_data_Rd[14]), .Q(n775) );
  BUF2 U94 ( .A(i_data_Rd[15]), .Q(n779) );
  NOR31 U95 ( .A(n862), .B(n879), .C(n883), .Q(n42) );
  NOR31 U96 ( .A(n880), .B(n881), .C(n882), .Q(n41) );
  INV3 U97 ( .A(n77), .Q(n860) );
  NAND22 U98 ( .A(n45), .B(n42), .Q(n77) );
  INV3 U99 ( .A(n78), .Q(n859) );
  NAND22 U100 ( .A(n47), .B(n42), .Q(n78) );
  INV3 U101 ( .A(n79), .Q(n858) );
  NAND22 U102 ( .A(n49), .B(n42), .Q(n79) );
  INV3 U103 ( .A(n80), .Q(n857) );
  NAND22 U104 ( .A(n51), .B(n42), .Q(n80) );
  INV3 U105 ( .A(n81), .Q(n856) );
  NAND22 U106 ( .A(n53), .B(n42), .Q(n81) );
  INV3 U107 ( .A(n82), .Q(n855) );
  NAND22 U108 ( .A(n55), .B(n42), .Q(n82) );
  INV3 U109 ( .A(n56), .Q(n872) );
  NAND22 U110 ( .A(n44), .B(n57), .Q(n56) );
  INV3 U111 ( .A(n58), .Q(n871) );
  NAND22 U112 ( .A(n44), .B(n41), .Q(n58) );
  INV3 U113 ( .A(n46), .Q(n877) );
  NAND22 U114 ( .A(n47), .B(n44), .Q(n46) );
  INV3 U115 ( .A(n61), .Q(n869) );
  NAND22 U116 ( .A(n60), .B(n47), .Q(n61) );
  INV3 U117 ( .A(n62), .Q(n868) );
  NAND22 U118 ( .A(n60), .B(n49), .Q(n62) );
  INV3 U119 ( .A(n64), .Q(n866) );
  NAND22 U120 ( .A(n60), .B(n53), .Q(n64) );
  INV3 U121 ( .A(n65), .Q(n865) );
  NAND22 U122 ( .A(n60), .B(n55), .Q(n65) );
  INV3 U123 ( .A(n67), .Q(n863) );
  NAND22 U124 ( .A(n60), .B(n41), .Q(n67) );
  INV3 U125 ( .A(n70), .Q(n852) );
  NAND22 U126 ( .A(n69), .B(n47), .Q(n70) );
  INV3 U127 ( .A(n71), .Q(n851) );
  NAND22 U128 ( .A(n69), .B(n49), .Q(n71) );
  INV3 U129 ( .A(n73), .Q(n849) );
  NAND22 U130 ( .A(n69), .B(n53), .Q(n73) );
  INV3 U131 ( .A(n74), .Q(n848) );
  NAND22 U132 ( .A(n69), .B(n55), .Q(n74) );
  INV3 U133 ( .A(n76), .Q(n846) );
  NAND22 U134 ( .A(n69), .B(n41), .Q(n76) );
  INV3 U135 ( .A(n39), .Q(n854) );
  NAND22 U136 ( .A(n42), .B(n57), .Q(n39) );
  INV3 U137 ( .A(n48), .Q(n876) );
  NAND22 U138 ( .A(n49), .B(n44), .Q(n48) );
  INV3 U139 ( .A(n50), .Q(n875) );
  NAND22 U140 ( .A(n51), .B(n44), .Q(n50) );
  INV3 U141 ( .A(n52), .Q(n874) );
  NAND22 U142 ( .A(n53), .B(n44), .Q(n52) );
  INV3 U143 ( .A(n54), .Q(n873) );
  NAND22 U144 ( .A(n55), .B(n44), .Q(n54) );
  INV3 U145 ( .A(n43), .Q(n878) );
  NAND22 U146 ( .A(n44), .B(n45), .Q(n43) );
  INV3 U147 ( .A(n59), .Q(n870) );
  NAND22 U148 ( .A(n60), .B(n45), .Q(n59) );
  INV3 U149 ( .A(n68), .Q(n853) );
  NAND22 U150 ( .A(n69), .B(n45), .Q(n68) );
  INV3 U151 ( .A(n66), .Q(n864) );
  NAND22 U152 ( .A(n60), .B(n57), .Q(n66) );
  INV3 U153 ( .A(n75), .Q(n847) );
  NAND22 U154 ( .A(n69), .B(n57), .Q(n75) );
  INV3 U155 ( .A(n72), .Q(n850) );
  NAND22 U156 ( .A(n69), .B(n51), .Q(n72) );
  INV3 U157 ( .A(n63), .Q(n867) );
  NAND22 U158 ( .A(n60), .B(n51), .Q(n63) );
  BUF2 U159 ( .A(n369), .Q(n373) );
  BUF2 U160 ( .A(n369), .Q(n374) );
  BUF2 U161 ( .A(n712), .Q(n717) );
  BUF2 U162 ( .A(i_data_Rd[16]), .Q(n780) );
  BUF2 U163 ( .A(i_data_Rd[16]), .Q(n781) );
  BUF2 U164 ( .A(i_data_Rd[16]), .Q(n782) );
  BUF2 U165 ( .A(i_data_Rd[16]), .Q(n783) );
  BUF2 U166 ( .A(i_data_Rd[17]), .Q(n784) );
  BUF2 U167 ( .A(i_data_Rd[17]), .Q(n785) );
  BUF2 U168 ( .A(i_data_Rd[17]), .Q(n786) );
  BUF2 U169 ( .A(i_data_Rd[17]), .Q(n787) );
  BUF2 U170 ( .A(i_data_Rd[18]), .Q(n788) );
  BUF2 U171 ( .A(i_data_Rd[18]), .Q(n789) );
  BUF2 U172 ( .A(i_data_Rd[18]), .Q(n790) );
  BUF2 U173 ( .A(i_data_Rd[19]), .Q(n791) );
  BUF2 U174 ( .A(i_data_Rd[20]), .Q(n794) );
  BUF2 U175 ( .A(i_data_Rd[21]), .Q(n798) );
  BUF2 U176 ( .A(i_data_Rd[22]), .Q(n802) );
  BUF2 U177 ( .A(i_data_Rd[24]), .Q(n807) );
  BUF2 U178 ( .A(i_data_Rd[25]), .Q(n810) );
  BUF2 U179 ( .A(i_data_Rd[26]), .Q(n811) );
  BUF2 U180 ( .A(i_data_Rd[27]), .Q(n813) );
  BUF2 U181 ( .A(i_data_Rd[29]), .Q(n817) );
  BUF2 U182 ( .A(i_data_Rd[30]), .Q(n821) );
  BUF2 U183 ( .A(i_data_Rd[31]), .Q(n823) );
  BUF2 U184 ( .A(i_data_Rd[19]), .Q(n792) );
  BUF2 U185 ( .A(i_data_Rd[20]), .Q(n795) );
  BUF2 U186 ( .A(i_data_Rd[21]), .Q(n799) );
  BUF2 U187 ( .A(i_data_Rd[22]), .Q(n803) );
  BUF2 U188 ( .A(i_data_Rd[24]), .Q(n808) );
  BUF2 U189 ( .A(i_data_Rd[26]), .Q(n812) );
  BUF2 U190 ( .A(i_data_Rd[27]), .Q(n814) );
  BUF2 U191 ( .A(i_data_Rd[28]), .Q(n816) );
  BUF2 U192 ( .A(i_data_Rd[29]), .Q(n818) );
  BUF2 U193 ( .A(i_data_Rd[30]), .Q(n822) );
  BUF2 U194 ( .A(i_data_Rd[31]), .Q(n824) );
  BUF2 U195 ( .A(i_data_Rd[19]), .Q(n793) );
  BUF2 U196 ( .A(i_data_Rd[20]), .Q(n796) );
  BUF2 U197 ( .A(i_data_Rd[21]), .Q(n800) );
  BUF2 U198 ( .A(i_data_Rd[22]), .Q(n804) );
  BUF2 U199 ( .A(i_data_Rd[23]), .Q(n805) );
  BUF2 U200 ( .A(i_data_Rd[24]), .Q(n809) );
  BUF2 U201 ( .A(i_data_Rd[27]), .Q(n815) );
  BUF2 U202 ( .A(i_data_Rd[29]), .Q(n819) );
  BUF2 U203 ( .A(i_data_Rd[20]), .Q(n797) );
  BUF2 U204 ( .A(i_data_Rd[21]), .Q(n801) );
  BUF2 U205 ( .A(i_data_Rd[23]), .Q(n806) );
  BUF2 U206 ( .A(i_data_Rd[29]), .Q(n820) );
  BUF2 U207 ( .A(i_addr_Rt[0]), .Q(n385) );
  BUF2 U208 ( .A(i_addr_Rt[0]), .Q(n386) );
  BUF2 U209 ( .A(i_addr_Rt[0]), .Q(n387) );
  BUF2 U210 ( .A(i_addr_Rt[0]), .Q(n388) );
  BUF2 U211 ( .A(i_addr_Rs[0]), .Q(n726) );
  BUF2 U212 ( .A(i_addr_Rs[0]), .Q(n727) );
  BUF2 U213 ( .A(i_addr_Rs[0]), .Q(n728) );
  BUF2 U214 ( .A(i_addr_Rs[0]), .Q(n729) );
  BUF2 U215 ( .A(i_addr_Rs[0]), .Q(n730) );
  BUF2 U216 ( .A(i_addr_Rt[1]), .Q(n370) );
  BUF2 U217 ( .A(i_addr_Rs[1]), .Q(n713) );
  NOR31 U218 ( .A(i_addr_Rd[3]), .B(i_addr_Rd[4]), .C(n883), .Q(n44) );
  NOR31 U219 ( .A(n862), .B(i_addr_Rd[3]), .C(n883), .Q(n69) );
  NOR31 U220 ( .A(n879), .B(i_addr_Rd[4]), .C(n883), .Q(n60) );
  MUX22 U221 ( .A(n394), .B(n389), .S(i_addr_Rs[4]), .Q(o_data_Rs[0]) );
  IMUX40 U222 ( .A(n390), .B(n391), .C(n392), .D(n393), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n389) );
  IMUX40 U223 ( .A(n395), .B(n396), .C(n397), .D(n398), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n394) );
  NOR31 U224 ( .A(n881), .B(i_addr_Rd[0]), .C(n880), .Q(n57) );
  NOR31 U225 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(i_addr_Rd[0]), .Q(n45)
         );
  NOR31 U226 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n880), .Q(n53) );
  NOR31 U227 ( .A(n880), .B(i_addr_Rd[1]), .C(n882), .Q(n55) );
  NOR31 U228 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(n882), .Q(n47) );
  NOR31 U229 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[2]), .C(n881), .Q(n49) );
  NOR31 U230 ( .A(n881), .B(i_addr_Rd[2]), .C(n882), .Q(n51) );
  IMUX40 U231 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n387), .S1(n372), .Q(n10) );
  IMUX40 U232 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n386), .S1(i_addr_Rt[1]), .Q(n8) );
  IMUX40 U233 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n388), .S1(i_addr_Rt[1]), .Q(n7) );
  IMUX40 U234 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(i_addr_Rt[0]), .S1(n375), .Q(n5) );
  IMUX40 U235 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(i_addr_Rt[0]), .S1(n371), .Q(n3) );
  IMUX40 U236 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n2) );
  IMUX40 U237 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n387), .S1(n369), .Q(n15) );
  IMUX40 U238 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n388), .S1(i_addr_Rt[1]), .Q(n13) );
  IMUX40 U239 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n383), .S1(i_addr_Rt[1]), .Q(n12) );
  IMUX40 U240 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n388), .S1(n375), .Q(n20) );
  IMUX40 U241 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n18) );
  IMUX40 U242 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(i_addr_Rt[0]), .S1(n369), .Q(n25) );
  IMUX40 U243 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n388), .S1(n374), .Q(n23) );
  IMUX40 U244 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n388), .S1(i_addr_Rt[1]), .Q(n22) );
  IMUX40 U245 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n380), .S1(n375), .Q(n30) );
  IMUX40 U246 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n386), .S1(i_addr_Rt[1]), .Q(n28) );
  IMUX40 U247 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n378), .S1(n371), .Q(n35) );
  IMUX40 U248 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n376), .S1(i_addr_Rt[1]), .Q(n33) );
  IMUX40 U249 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n386), .S1(i_addr_Rt[1]), .Q(n32) );
  IMUX40 U250 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n383), .S1(n369), .Q(n84) );
  IMUX40 U251 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n387), .S1(i_addr_Rt[1]), .Q(n38) );
  IMUX40 U252 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(i_addr_Rt[0]), .S1(n375), .Q(n89) );
  IMUX40 U253 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n386), .S1(n370), .Q(n87) );
  IMUX40 U254 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n86) );
  IMUX40 U255 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(i_addr_Rt[0]), .S1(n371), .Q(n94) );
  IMUX40 U256 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n92) );
  IMUX40 U257 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n376), .S1(n375), .Q(n99) );
  IMUX40 U258 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n97) );
  IMUX40 U259 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n387), .S1(n373), .Q(n96) );
  IMUX40 U260 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n388), .S1(n375), .Q(n104) );
  IMUX40 U261 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n386), .S1(i_addr_Rt[1]), .Q(n102) );
  IMUX40 U262 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n387), .S1(n373), .Q(n109) );
  IMUX40 U263 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n376), .S1(n372), .Q(n107) );
  IMUX40 U264 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n106) );
  IMUX40 U265 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n388), .S1(i_addr_Rt[1]), .Q(n114) );
  IMUX40 U266 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n386), .S1(i_addr_Rt[1]), .Q(n112) );
  IMUX40 U267 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n388), .S1(n375), .Q(n119) );
  IMUX40 U268 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n117) );
  IMUX40 U269 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n379), .S1(n370), .Q(n116) );
  IMUX40 U270 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n386), .S1(n375), .Q(n124) );
  IMUX40 U271 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n387), .S1(n372), .Q(n122) );
  IMUX40 U272 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n387), .S1(n375), .Q(n129) );
  IMUX40 U273 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n387), .S1(n371), .Q(n127) );
  IMUX40 U274 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n378), .S1(i_addr_Rt[1]), .Q(n126) );
  IMUX40 U275 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n388), .S1(n369), .Q(n134) );
  IMUX40 U276 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n387), .S1(n375), .Q(n132) );
  IMUX40 U277 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n384), .S1(n375), .Q(n139) );
  IMUX40 U278 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n388), .S1(n369), .Q(n137) );
  IMUX40 U279 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n136) );
  IMUX40 U280 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n377), .S1(i_addr_Rt[1]), .Q(n144) );
  IMUX40 U281 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n142) );
  IMUX40 U282 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n385), .S1(n370), .Q(n149) );
  IMUX40 U283 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n387), .S1(n374), .Q(n147) );
  IMUX40 U284 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n388), .S1(i_addr_Rt[1]), .Q(n146) );
  IMUX40 U285 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n376), .S1(n371), .Q(n154) );
  IMUX40 U286 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n378), .S1(n375), .Q(n152) );
  IMUX40 U287 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n376), .S1(n369), .Q(n159) );
  IMUX40 U288 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n376), .S1(n369), .Q(n157) );
  IMUX40 U289 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n376), .S1(i_addr_Rt[1]), .Q(n156) );
  IMUX40 U290 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n376), .S1(i_addr_Rt[1]), .Q(n164) );
  IMUX40 U291 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n376), .S1(n369), .Q(n162) );
  IMUX40 U292 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n376), .S1(n371), .Q(n169) );
  IMUX40 U293 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n376), .S1(n375), .Q(n167) );
  IMUX40 U294 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n376), .S1(n374), .Q(n166) );
  IMUX40 U295 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n377), .S1(i_addr_Rt[1]), .Q(n174) );
  IMUX40 U296 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n377), .S1(n372), .Q(n172) );
  IMUX40 U297 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n377), .S1(n375), .Q(n179) );
  IMUX40 U298 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n377), .S1(n369), .Q(n177) );
  IMUX40 U299 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n377), .S1(i_addr_Rt[1]), .Q(n176) );
  IMUX40 U300 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n377), .S1(n375), .Q(n184) );
  IMUX40 U301 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n377), .S1(i_addr_Rt[1]), .Q(n182) );
  IMUX40 U302 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n378), .S1(n371), .Q(n189) );
  IMUX40 U303 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n378), .S1(n371), .Q(n187) );
  IMUX40 U304 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n378), .S1(n371), .Q(n186) );
  IMUX40 U305 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n378), .S1(n371), .Q(n194) );
  IMUX40 U306 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n378), .S1(n371), .Q(n192) );
  IMUX40 U307 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n378), .S1(n371), .Q(n199) );
  IMUX40 U308 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n378), .S1(i_addr_Rt[1]), .Q(n197) );
  IMUX40 U309 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n378), .S1(i_addr_Rt[1]), .Q(n196) );
  IMUX40 U310 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n380), .S1(i_addr_Rt[1]), .Q(n204) );
  IMUX40 U311 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n382), .S1(i_addr_Rt[1]), .Q(n202) );
  IMUX40 U312 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n385), .S1(n371), .Q(n209) );
  IMUX40 U313 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n384), .S1(i_addr_Rt[1]), .Q(n207) );
  IMUX40 U314 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n384), .S1(n372), .Q(n206) );
  IMUX40 U315 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n379), .S1(n373), .Q(n214) );
  IMUX40 U316 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n380), .S1(n369), .Q(n212) );
  IMUX40 U317 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n383), .S1(n372), .Q(n219) );
  IMUX40 U318 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(i_addr_Rt[0]), .S1(n372), .Q(n217) );
  IMUX40 U319 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n385), .S1(n370), .Q(n216) );
  IMUX40 U320 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n382), .S1(n370), .Q(n224) );
  IMUX40 U321 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n378), .S1(n370), .Q(n222) );
  IMUX40 U322 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n229) );
  IMUX40 U323 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n227) );
  IMUX40 U324 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n386), .S1(n370), .Q(n226) );
  IMUX40 U325 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n379), .S1(n370), .Q(n234) );
  IMUX40 U326 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n379), .S1(n370), .Q(n232) );
  IMUX40 U327 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n379), .S1(n370), .Q(n239) );
  IMUX40 U328 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n379), .S1(n370), .Q(n237) );
  IMUX40 U329 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n379), .S1(n370), .Q(n236) );
  IMUX40 U330 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n379), .S1(n370), .Q(n244) );
  IMUX40 U331 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n379), .S1(n372), .Q(n242) );
  IMUX40 U332 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n380), .S1(n369), .Q(n249) );
  IMUX40 U333 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n380), .S1(n375), .Q(n247) );
  IMUX40 U334 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n380), .S1(n375), .Q(n246) );
  IMUX40 U335 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n380), .S1(n375), .Q(n254) );
  IMUX40 U336 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n380), .S1(n370), .Q(n252) );
  IMUX40 U337 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n380), .S1(n369), .Q(n259) );
  IMUX40 U338 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n380), .S1(n370), .Q(n257) );
  IMUX40 U339 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n380), .S1(n372), .Q(n256) );
  IMUX40 U340 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n385), .S1(n370), .Q(n264) );
  IMUX40 U341 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n386), .S1(n370), .Q(n262) );
  IMUX40 U342 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n380), .S1(n371), .Q(n269) );
  IMUX40 U343 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n386), .S1(n371), .Q(n267) );
  IMUX40 U344 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n376), .S1(n371), .Q(n266) );
  IMUX40 U345 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(i_addr_Rt[0]), .S1(n371), .Q(n274) );
  IMUX40 U346 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n387), .S1(n371), .Q(n272) );
  IMUX40 U347 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n381), .S1(n369), .Q(n279) );
  IMUX40 U348 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n381), .S1(n369), .Q(n277) );
  IMUX40 U349 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n381), .S1(n369), .Q(n276) );
  IMUX40 U350 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n381), .S1(n373), .Q(n284) );
  IMUX40 U351 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n381), .S1(n373), .Q(n282) );
  IMUX40 U352 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n381), .S1(n372), .Q(n289) );
  IMUX40 U353 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n381), .S1(n369), .Q(n287) );
  IMUX40 U354 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n381), .S1(n373), .Q(n286) );
  IMUX40 U355 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n382), .S1(n372), .Q(n294) );
  IMUX40 U356 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n382), .S1(n372), .Q(n292) );
  IMUX40 U357 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n382), .S1(n373), .Q(n299) );
  IMUX40 U358 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n382), .S1(n372), .Q(n297) );
  IMUX40 U359 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n382), .S1(n374), .Q(n296) );
  IMUX40 U360 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n382), .S1(n374), .Q(n304) );
  IMUX40 U361 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n382), .S1(n372), .Q(n302) );
  IMUX40 U362 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n387), .S1(n371), .Q(n309) );
  IMUX40 U363 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n386), .S1(n372), .Q(n307) );
  IMUX40 U364 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n378), .S1(n372), .Q(n306) );
  IMUX40 U365 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n376), .S1(n372), .Q(n314) );
  IMUX40 U366 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n377), .S1(n372), .Q(n312) );
  IMUX40 U367 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n377), .S1(n372), .Q(n319) );
  IMUX40 U368 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n385), .S1(n372), .Q(n317) );
  IMUX40 U369 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n381), .S1(n372), .Q(n316) );
  IMUX40 U370 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n383), .S1(n374), .Q(n324) );
  IMUX40 U371 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n383), .S1(n373), .Q(n322) );
  IMUX40 U372 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n383), .S1(n370), .Q(n329) );
  IMUX40 U373 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n383), .S1(n369), .Q(n327) );
  IMUX40 U374 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n383), .S1(n374), .Q(n326) );
  IMUX40 U375 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n383), .S1(n373), .Q(n334) );
  IMUX40 U376 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n383), .S1(n374), .Q(n332) );
  IMUX40 U377 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n384), .S1(n372), .Q(n339) );
  IMUX40 U378 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n384), .S1(n372), .Q(n337) );
  IMUX40 U379 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n384), .S1(n369), .Q(n336) );
  IMUX40 U380 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n384), .S1(n374), .Q(n344) );
  IMUX40 U381 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n384), .S1(n369), .Q(n342) );
  IMUX40 U382 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n384), .S1(n373), .Q(n349) );
  IMUX40 U383 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n384), .S1(n373), .Q(n347) );
  IMUX40 U384 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n384), .S1(n373), .Q(n346) );
  IMUX40 U385 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(i_addr_Rt[0]), .S1(n373), .Q(n354) );
  IMUX40 U386 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(i_addr_Rt[0]), .S1(n373), .Q(n352) );
  IMUX40 U387 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n384), .S1(n374), .Q(n359) );
  IMUX40 U388 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n388), .S1(n374), .Q(n357) );
  IMUX40 U389 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n356) );
  IMUX40 U390 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n364) );
  IMUX40 U391 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n362) );
  IMUX40 U392 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n726), .S1(n718), .Q(n398) );
  IMUX40 U393 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n726), .S1(n714), .Q(n396) );
  IMUX40 U394 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n726), .S1(n713), .Q(n395) );
  IMUX40 U395 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(n724), .S1(i_addr_Rs[1]), .Q(n393) );
  IMUX40 U396 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(n725), .S1(n714), .Q(n391) );
  IMUX40 U397 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(n727), .S1(i_addr_Rs[1]), .Q(n390) );
  IMUX40 U398 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n726), .S1(i_addr_Rs[1]), .Q(n403) );
  IMUX40 U399 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n726), .S1(n714), .Q(n401) );
  IMUX40 U400 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n726), .S1(i_addr_Rs[1]), .Q(n400) );
  IMUX40 U401 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n726), .S1(n714), .Q(n408) );
  IMUX40 U402 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n726), .S1(i_addr_Rs[1]), .Q(n406) );
  IMUX40 U403 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n730), .S1(n712), .Q(n413) );
  IMUX40 U404 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n729), .S1(n718), .Q(n411) );
  IMUX40 U405 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n730), .S1(n714), .Q(n410) );
  IMUX40 U406 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n720), .S1(n713), .Q(n418) );
  IMUX40 U407 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n721), .S1(n718), .Q(n416) );
  IMUX40 U408 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n730), .S1(n718), .Q(n423) );
  IMUX40 U409 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n722), .S1(n716), .Q(n421) );
  IMUX40 U410 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n729), .S1(i_addr_Rs[1]), .Q(n420) );
  IMUX40 U411 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n428) );
  IMUX40 U412 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n426) );
  IMUX40 U413 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n726), .S1(n714), .Q(n433) );
  IMUX40 U414 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n729), .S1(n712), .Q(n431) );
  IMUX40 U415 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(i_addr_Rs[0]), .S1(n714), .Q(n430) );
  IMUX40 U416 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n438) );
  IMUX40 U417 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(i_addr_Rs[0]), .S1(n712), .Q(n436) );
  IMUX40 U418 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n727), .S1(n718), .Q(n443) );
  IMUX40 U419 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n727), .S1(n718), .Q(n441) );
  IMUX40 U420 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n727), .S1(n718), .Q(n440) );
  IMUX40 U421 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n727), .S1(n718), .Q(n448) );
  IMUX40 U422 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n727), .S1(n716), .Q(n446) );
  IMUX40 U423 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n727), .S1(n718), .Q(n453) );
  IMUX40 U424 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n727), .S1(n713), .Q(n451) );
  IMUX40 U425 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n727), .S1(n712), .Q(n450) );
  IMUX40 U426 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n720), .S1(n713), .Q(n458) );
  IMUX40 U427 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n730), .S1(n713), .Q(n456) );
  IMUX40 U428 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n729), .S1(n713), .Q(n463) );
  IMUX40 U429 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(i_addr_Rs[0]), .S1(n713), .Q(n461) );
  IMUX40 U430 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n460) );
  IMUX40 U431 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n468) );
  IMUX40 U432 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(i_addr_Rs[0]), .S1(n712), .Q(n466) );
  IMUX40 U433 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n727), .S1(n718), .Q(n473) );
  IMUX40 U434 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n721), .S1(i_addr_Rs[1]), .Q(n471) );
  IMUX40 U435 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(i_addr_Rs[0]), .S1(n713), .Q(n470) );
  IMUX40 U436 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(i_addr_Rs[0]), .S1(n713), .Q(n478) );
  IMUX40 U437 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(i_addr_Rs[0]), .S1(n715), .Q(n476) );
  IMUX40 U438 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n728), .S1(i_addr_Rs[1]), .Q(n483) );
  IMUX40 U439 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n727), .S1(i_addr_Rs[1]), .Q(n481) );
  IMUX40 U440 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n726), .S1(n713), .Q(n480) );
  IMUX40 U441 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n728), .S1(n714), .Q(n488) );
  IMUX40 U442 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n730), .S1(n712), .Q(n486) );
  IMUX40 U443 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n724), .S1(n715), .Q(n493) );
  IMUX40 U444 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n729), .S1(n713), .Q(n491) );
  IMUX40 U445 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n726), .S1(i_addr_Rs[1]), .Q(n490) );
  IMUX40 U446 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(i_addr_Rs[0]), .S1(n718), .Q(n498) );
  IMUX40 U447 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n727), .S1(n715), .Q(n496) );
  IMUX40 U448 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n719), .S1(n713), .Q(n503) );
  IMUX40 U449 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n501) );
  IMUX40 U450 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n719), .S1(n718), .Q(n500) );
  IMUX40 U451 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n719), .S1(n715), .Q(n508) );
  IMUX40 U452 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n506) );
  IMUX40 U453 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n719), .S1(n716), .Q(n513) );
  IMUX40 U454 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n719), .S1(n713), .Q(n511) );
  IMUX40 U455 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n719), .S1(n714), .Q(n510) );
  IMUX40 U456 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n730), .S1(n714), .Q(n518) );
  IMUX40 U457 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n728), .S1(n712), .Q(n516) );
  IMUX40 U458 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n723), .S1(n712), .Q(n523) );
  IMUX40 U459 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n722), .S1(n718), .Q(n521) );
  IMUX40 U460 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n719), .S1(n713), .Q(n520) );
  IMUX40 U461 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n728), .S1(n713), .Q(n528) );
  IMUX40 U462 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n723), .S1(n713), .Q(n526) );
  IMUX40 U463 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n720), .S1(n716), .Q(n533) );
  IMUX40 U464 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n720), .S1(n716), .Q(n531) );
  IMUX40 U465 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n720), .S1(n712), .Q(n530) );
  IMUX40 U466 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n720), .S1(n716), .Q(n538) );
  IMUX40 U467 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n720), .S1(n718), .Q(n536) );
  IMUX40 U468 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n720), .S1(n715), .Q(n543) );
  IMUX40 U469 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n720), .S1(n712), .Q(n541) );
  IMUX40 U470 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n720), .S1(n714), .Q(n540) );
  IMUX40 U471 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n721), .S1(n712), .Q(n548) );
  IMUX40 U472 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n721), .S1(n713), .Q(n546) );
  IMUX40 U473 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n721), .S1(n712), .Q(n553) );
  IMUX40 U474 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n721), .S1(n713), .Q(n551) );
  IMUX40 U475 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n721), .S1(i_addr_Rs[1]), .Q(n550) );
  IMUX40 U476 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n721), .S1(i_addr_Rs[1]), .Q(n558) );
  IMUX40 U477 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n721), .S1(i_addr_Rs[1]), .Q(n556) );
  IMUX40 U478 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n725), .S1(i_addr_Rs[1]), .Q(n563) );
  IMUX40 U479 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n561) );
  IMUX40 U480 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n730), .S1(n714), .Q(n560) );
  IMUX40 U481 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n729), .S1(n713), .Q(n568) );
  IMUX40 U482 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n724), .S1(n712), .Q(n566) );
  IMUX40 U483 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n730), .S1(n712), .Q(n573) );
  IMUX40 U484 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n729), .S1(n714), .Q(n571) );
  IMUX40 U485 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n729), .S1(i_addr_Rs[1]), .Q(n570) );
  IMUX40 U486 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n728), .S1(n712), .Q(n578) );
  IMUX40 U487 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n728), .S1(i_addr_Rs[1]), .Q(n576) );
  IMUX40 U488 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n730), .S1(n718), .Q(n583) );
  IMUX40 U489 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n730), .S1(i_addr_Rs[1]), .Q(n581) );
  IMUX40 U490 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n727), .S1(i_addr_Rs[1]), .Q(n580) );
  IMUX40 U491 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n728), .S1(n718), .Q(n588) );
  IMUX40 U492 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n730), .S1(n713), .Q(n586) );
  IMUX40 U493 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n728), .S1(n712), .Q(n593) );
  IMUX40 U494 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n728), .S1(n712), .Q(n591) );
  IMUX40 U495 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n723), .S1(i_addr_Rs[1]), .Q(n590) );
  IMUX40 U496 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n728), .S1(i_addr_Rs[1]), .Q(n598) );
  IMUX40 U497 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n728), .S1(i_addr_Rs[1]), .Q(n596) );
  IMUX40 U498 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n719), .S1(n712), .Q(n603) );
  IMUX40 U499 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n724), .S1(n718), .Q(n601) );
  IMUX40 U500 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n723), .S1(n712), .Q(n600) );
  IMUX40 U501 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n724), .S1(n716), .Q(n608) );
  IMUX40 U502 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n730), .S1(n718), .Q(n606) );
  IMUX40 U503 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n719), .S1(n714), .Q(n613) );
  IMUX40 U504 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n722), .S1(n714), .Q(n611) );
  IMUX40 U505 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n729), .S1(n714), .Q(n610) );
  IMUX40 U506 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n728), .S1(n714), .Q(n618) );
  IMUX40 U507 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n729), .S1(n714), .Q(n616) );
  IMUX40 U508 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n722), .S1(n715), .Q(n623) );
  IMUX40 U509 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n722), .S1(n715), .Q(n621) );
  IMUX40 U510 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n722), .S1(n715), .Q(n620) );
  IMUX40 U511 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n722), .S1(n715), .Q(n628) );
  IMUX40 U512 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n722), .S1(n715), .Q(n626) );
  IMUX40 U513 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n722), .S1(n715), .Q(n633) );
  IMUX40 U514 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n722), .S1(n716), .Q(n631) );
  IMUX40 U515 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n722), .S1(n716), .Q(n630) );
  IMUX40 U516 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n725), .S1(n716), .Q(n638) );
  IMUX40 U517 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n720), .S1(n716), .Q(n636) );
  IMUX40 U518 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n726), .S1(n716), .Q(n643) );
  IMUX40 U519 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n726), .S1(n716), .Q(n641) );
  IMUX40 U520 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n727), .S1(n716), .Q(n640) );
  IMUX40 U521 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n719), .S1(n714), .Q(n648) );
  IMUX40 U522 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n726), .S1(n715), .Q(n646) );
  IMUX40 U523 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n723), .S1(n716), .Q(n653) );
  IMUX40 U524 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n723), .S1(n715), .Q(n651) );
  IMUX40 U525 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n723), .S1(n715), .Q(n650) );
  IMUX40 U526 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n723), .S1(n716), .Q(n658) );
  IMUX40 U527 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n723), .S1(n715), .Q(n656) );
  IMUX40 U528 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n723), .S1(n714), .Q(n663) );
  IMUX40 U529 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n723), .S1(n716), .Q(n661) );
  IMUX40 U530 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n723), .S1(n715), .Q(n660) );
  IMUX40 U531 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n724), .S1(n716), .Q(n668) );
  IMUX40 U532 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n724), .S1(n716), .Q(n666) );
  IMUX40 U533 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n724), .S1(n715), .Q(n673) );
  IMUX40 U534 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n724), .S1(n714), .Q(n671) );
  IMUX40 U535 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n724), .S1(n718), .Q(n670) );
  IMUX40 U536 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n724), .S1(n714), .Q(n678) );
  IMUX40 U537 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n724), .S1(n715), .Q(n676) );
  IMUX40 U538 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n725), .S1(n715), .Q(n683) );
  IMUX40 U539 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n725), .S1(n712), .Q(n681) );
  IMUX40 U540 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n725), .S1(n712), .Q(n680) );
  IMUX40 U541 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n725), .S1(n715), .Q(n688) );
  IMUX40 U542 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n725), .S1(n718), .Q(n686) );
  IMUX40 U543 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n725), .S1(n717), .Q(n685) );
  IMUX40 U544 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n725), .S1(n717), .Q(n693) );
  IMUX40 U545 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n725), .S1(n717), .Q(n691) );
  IMUX40 U546 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n725), .S1(n717), .Q(n690) );
  IMUX40 U547 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n730), .S1(n717), .Q(n698) );
  IMUX40 U548 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n723), .S1(n717), .Q(n695) );
  IMUX40 U549 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(i_addr_Rs[0]), .S1(n717), .Q(n696) );
  IMUX40 U550 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(i_addr_Rs[0]), .S1(n715), .Q(n703) );
  IMUX40 U551 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n725), .S1(n717), .Q(n701) );
  IMUX40 U552 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n719), .S1(n717), .Q(n700) );
  IMUX40 U553 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n729), .S1(n714), .Q(n708) );
  IMUX40 U554 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n727), .S1(n717), .Q(n705) );
  IMUX40 U555 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n730), .S1(n717), .Q(n706) );
  IMUX40 U556 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n387), .S1(n371), .Q(n9) );
  IMUX40 U557 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(i_addr_Rt[0]), .S1(n375), .Q(n4) );
  IMUX40 U558 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n387), .S1(n375), .Q(n14) );
  IMUX40 U559 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n388), .S1(n370), .Q(n19) );
  IMUX40 U560 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n387), .S1(n371), .Q(n24) );
  IMUX40 U561 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n387), .S1(n375), .Q(n29) );
  IMUX40 U562 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n386), .S1(n375), .Q(n34) );
  IMUX40 U563 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n387), .S1(n375), .Q(n83) );
  IMUX40 U564 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n376), .S1(n375), .Q(n88) );
  IMUX40 U565 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n388), .S1(n369), .Q(n93) );
  IMUX40 U566 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n377), .S1(n369), .Q(n98) );
  IMUX40 U567 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n386), .S1(n369), .Q(n103) );
  IMUX40 U568 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n377), .S1(n369), .Q(n108) );
  IMUX40 U569 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n385), .S1(n369), .Q(n113) );
  IMUX40 U570 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n387), .S1(n375), .Q(n118) );
  IMUX40 U571 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n379), .S1(n373), .Q(n123) );
  IMUX40 U572 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n388), .S1(n375), .Q(n128) );
  IMUX40 U573 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n386), .S1(n370), .Q(n133) );
  IMUX40 U574 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n386), .S1(n375), .Q(n138) );
  IMUX40 U575 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n388), .S1(n372), .Q(n143) );
  IMUX40 U576 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n377), .S1(n372), .Q(n148) );
  IMUX40 U577 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n386), .S1(n369), .Q(n153) );
  IMUX40 U578 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n376), .S1(n372), .Q(n158) );
  IMUX40 U579 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n376), .S1(i_addr_Rt[1]), .Q(n163) );
  IMUX40 U580 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n376), .S1(n371), .Q(n168) );
  IMUX40 U581 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n377), .S1(n371), .Q(n173) );
  IMUX40 U582 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n377), .S1(n375), .Q(n178) );
  IMUX40 U583 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n377), .S1(n369), .Q(n183) );
  IMUX40 U584 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n378), .S1(n371), .Q(n188) );
  IMUX40 U585 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n378), .S1(n371), .Q(n193) );
  IMUX40 U586 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n378), .S1(n369), .Q(n198) );
  IMUX40 U587 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n381), .S1(i_addr_Rt[1]), .Q(n203) );
  IMUX40 U588 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n383), .S1(n370), .Q(n208) );
  IMUX40 U589 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n385), .S1(n374), .Q(n213) );
  IMUX40 U590 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n377), .S1(n375), .Q(n218) );
  IMUX40 U591 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n223) );
  IMUX40 U592 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n387), .S1(n370), .Q(n228) );
  IMUX40 U593 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n379), .S1(n370), .Q(n233) );
  IMUX40 U594 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n379), .S1(n370), .Q(n238) );
  IMUX40 U595 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n379), .S1(n371), .Q(n243) );
  IMUX40 U596 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n380), .S1(n375), .Q(n248) );
  IMUX40 U597 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n380), .S1(n372), .Q(n253) );
  IMUX40 U598 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n380), .S1(n370), .Q(n258) );
  IMUX40 U599 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n386), .S1(n372), .Q(n263) );
  IMUX40 U600 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n379), .S1(n371), .Q(n268) );
  IMUX40 U601 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n385), .S1(n371), .Q(n273) );
  IMUX40 U602 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n381), .S1(n369), .Q(n278) );
  IMUX40 U603 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n381), .S1(n372), .Q(n283) );
  IMUX40 U604 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n381), .S1(n372), .Q(n288) );
  IMUX40 U605 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n382), .S1(n373), .Q(n293) );
  IMUX40 U606 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n382), .S1(n371), .Q(n298) );
  IMUX40 U607 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n382), .S1(n374), .Q(n303) );
  IMUX40 U608 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n381), .S1(n371), .Q(n308) );
  IMUX40 U609 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n378), .S1(n372), .Q(n313) );
  IMUX40 U610 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n382), .S1(n372), .Q(n318) );
  IMUX40 U611 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n383), .S1(n373), .Q(n323) );
  IMUX40 U612 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n383), .S1(n369), .Q(n328) );
  IMUX40 U613 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n383), .S1(n374), .Q(n333) );
  IMUX40 U614 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n384), .S1(n369), .Q(n338) );
  IMUX40 U615 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n384), .S1(n373), .Q(n343) );
  IMUX40 U616 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n384), .S1(n373), .Q(n348) );
  IMUX40 U617 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(i_addr_Rt[0]), .S1(n373), .Q(n353) );
  IMUX40 U618 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n383), .S1(n374), .Q(n358) );
  IMUX40 U619 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n363) );
  IMUX40 U620 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n726), .S1(n716), .Q(n397) );
  IMUX40 U621 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(n723), .S1(n716), .Q(n392) );
  IMUX40 U622 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n726), .S1(i_addr_Rs[1]), .Q(n402) );
  IMUX40 U623 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n726), .S1(i_addr_Rs[1]), .Q(n407) );
  IMUX40 U624 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n721), .S1(n712), .Q(n412) );
  IMUX40 U625 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n728), .S1(n714), .Q(n417) );
  IMUX40 U626 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n422) );
  IMUX40 U627 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n427) );
  IMUX40 U628 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n727), .S1(n716), .Q(n432) );
  IMUX40 U629 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(i_addr_Rs[0]), .S1(n715), .Q(n437) );
  IMUX40 U630 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n727), .S1(n712), .Q(n442) );
  IMUX40 U631 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n727), .S1(n715), .Q(n447) );
  IMUX40 U632 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n727), .S1(n712), .Q(n452) );
  IMUX40 U633 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n728), .S1(n718), .Q(n457) );
  IMUX40 U634 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n729), .S1(n712), .Q(n462) );
  IMUX40 U635 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(i_addr_Rs[0]), .S1(n713), .Q(n467) );
  IMUX40 U636 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n726), .S1(n715), .Q(n472) );
  IMUX40 U637 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n728), .S1(n713), .Q(n477) );
  IMUX40 U638 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n729), .S1(i_addr_Rs[1]), .Q(n482) );
  IMUX40 U639 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n729), .S1(n713), .Q(n487) );
  IMUX40 U640 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n723), .S1(n714), .Q(n492) );
  IMUX40 U641 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n725), .S1(i_addr_Rs[1]), .Q(n497) );
  IMUX40 U642 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n719), .S1(n712), .Q(n502) );
  IMUX40 U643 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n719), .S1(n713), .Q(n507) );
  IMUX40 U644 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n719), .S1(n713), .Q(n512) );
  IMUX40 U645 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n725), .S1(n714), .Q(n517) );
  IMUX40 U646 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n721), .S1(n712), .Q(n522) );
  IMUX40 U647 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n724), .S1(n712), .Q(n527) );
  IMUX40 U648 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n720), .S1(n715), .Q(n532) );
  IMUX40 U649 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n720), .S1(n715), .Q(n537) );
  IMUX40 U650 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n720), .S1(n713), .Q(n542) );
  IMUX40 U651 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n721), .S1(n713), .Q(n547) );
  IMUX40 U652 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n721), .S1(n712), .Q(n552) );
  IMUX40 U653 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n721), .S1(i_addr_Rs[1]), .Q(n557) );
  IMUX40 U654 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n719), .S1(n713), .Q(n562) );
  IMUX40 U655 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n730), .S1(n713), .Q(n567) );
  IMUX40 U656 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n729), .S1(n713), .Q(n572) );
  IMUX40 U657 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n720), .S1(n718), .Q(n577) );
  IMUX40 U658 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n725), .S1(n714), .Q(n582) );
  IMUX40 U659 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n729), .S1(n714), .Q(n587) );
  IMUX40 U660 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n728), .S1(n713), .Q(n592) );
  IMUX40 U661 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n728), .S1(n718), .Q(n597) );
  IMUX40 U662 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n720), .S1(n714), .Q(n602) );
  IMUX40 U663 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n730), .S1(n715), .Q(n607) );
  IMUX40 U664 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n722), .S1(n714), .Q(n612) );
  IMUX40 U665 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n729), .S1(n714), .Q(n617) );
  IMUX40 U666 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n722), .S1(n715), .Q(n622) );
  IMUX40 U667 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n722), .S1(n715), .Q(n627) );
  IMUX40 U668 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n722), .S1(n716), .Q(n632) );
  IMUX40 U669 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n728), .S1(n716), .Q(n637) );
  IMUX40 U670 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n722), .S1(n715), .Q(n642) );
  IMUX40 U671 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n720), .S1(n716), .Q(n647) );
  IMUX40 U672 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n723), .S1(n715), .Q(n652) );
  IMUX40 U673 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n723), .S1(n718), .Q(n657) );
  IMUX40 U674 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n723), .S1(n718), .Q(n662) );
  IMUX40 U675 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n724), .S1(n718), .Q(n667) );
  IMUX40 U676 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n724), .S1(n716), .Q(n672) );
  IMUX40 U677 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n724), .S1(n716), .Q(n677) );
  IMUX40 U678 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n725), .S1(n712), .Q(n682) );
  IMUX40 U679 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n725), .S1(n717), .Q(n692) );
  IMUX40 U680 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n722), .S1(n716), .Q(n702) );
  BUF2 U681 ( .A(i_addr_Rt[3]), .Q(n366) );
  BUF2 U682 ( .A(i_addr_Rt[3]), .Q(n367) );
  BUF2 U683 ( .A(i_addr_Rs[3]), .Q(n709) );
  BUF2 U684 ( .A(i_addr_Rs[3]), .Q(n710) );
  INV3 U685 ( .A(i_addr_Rd[1]), .Q(n881) );
  INV3 U686 ( .A(i_addr_Rd[2]), .Q(n880) );
  INV3 U687 ( .A(i_addr_Rd[0]), .Q(n882) );
  INV3 U688 ( .A(i_con_RegWr), .Q(n883) );
  BUF2 U689 ( .A(i_addr_Rs[2]), .Q(n711) );
  INV3 U690 ( .A(i_addr_Rd[4]), .Q(n862) );
  INV3 U691 ( .A(i_addr_Rd[3]), .Q(n879) );
  MUX22 U692 ( .A(n404), .B(n399), .S(i_addr_Rs[4]), .Q(o_data_Rs[1]) );
  IMUX40 U693 ( .A(n405), .B(n406), .C(n407), .D(n408), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n404) );
  IMUX40 U694 ( .A(n400), .B(n401), .C(n402), .D(n403), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n399) );
  IMUX40 U695 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n726), .S1(n715), .Q(n405) );
  MUX22 U696 ( .A(n414), .B(n409), .S(i_addr_Rs[4]), .Q(o_data_Rs[2]) );
  IMUX40 U697 ( .A(n415), .B(n416), .C(n417), .D(n418), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n414) );
  IMUX40 U698 ( .A(n410), .B(n411), .C(n412), .D(n413), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n409) );
  IMUX40 U699 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n726), .S1(n718), .Q(n415) );
  MUX22 U700 ( .A(n424), .B(n419), .S(i_addr_Rs[4]), .Q(o_data_Rs[3]) );
  IMUX40 U701 ( .A(n425), .B(n426), .C(n427), .D(n428), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n424) );
  IMUX40 U702 ( .A(n420), .B(n421), .C(n422), .D(n423), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n419) );
  IMUX40 U703 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        i_addr_Rs[0]), .S1(n715), .Q(n425) );
  MUX22 U704 ( .A(n434), .B(n429), .S(i_addr_Rs[4]), .Q(o_data_Rs[4]) );
  IMUX40 U705 ( .A(n435), .B(n436), .C(n437), .D(n438), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n434) );
  IMUX40 U706 ( .A(n430), .B(n431), .C(n432), .D(n433), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n429) );
  IMUX40 U707 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n435) );
  MUX22 U708 ( .A(n444), .B(n439), .S(i_addr_Rs[4]), .Q(o_data_Rs[5]) );
  IMUX40 U709 ( .A(n445), .B(n446), .C(n447), .D(n448), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n444) );
  IMUX40 U710 ( .A(n440), .B(n441), .C(n442), .D(n443), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n439) );
  IMUX40 U711 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n727), .S1(i_addr_Rs[1]), .Q(n445) );
  MUX22 U712 ( .A(n454), .B(n449), .S(i_addr_Rs[4]), .Q(o_data_Rs[6]) );
  IMUX40 U713 ( .A(n455), .B(n456), .C(n457), .D(n458), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n454) );
  IMUX40 U714 ( .A(n450), .B(n451), .C(n452), .D(n453), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n449) );
  IMUX40 U715 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        i_addr_Rs[0]), .S1(n716), .Q(n455) );
  MUX22 U716 ( .A(n464), .B(n459), .S(i_addr_Rs[4]), .Q(o_data_Rs[7]) );
  IMUX40 U717 ( .A(n465), .B(n466), .C(n467), .D(n468), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n464) );
  IMUX40 U718 ( .A(n460), .B(n461), .C(n462), .D(n463), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n459) );
  IMUX40 U719 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        i_addr_Rs[0]), .S1(n718), .Q(n465) );
  MUX22 U720 ( .A(n474), .B(n469), .S(i_addr_Rs[4]), .Q(o_data_Rs[8]) );
  IMUX40 U721 ( .A(n475), .B(n476), .C(n477), .D(n478), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n474) );
  IMUX40 U722 ( .A(n470), .B(n471), .C(n472), .D(n473), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n469) );
  IMUX40 U723 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        i_addr_Rs[0]), .S1(n718), .Q(n475) );
  MUX22 U724 ( .A(n484), .B(n479), .S(i_addr_Rs[4]), .Q(o_data_Rs[9]) );
  IMUX40 U725 ( .A(n485), .B(n486), .C(n487), .D(n488), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n484) );
  IMUX40 U726 ( .A(n480), .B(n481), .C(n482), .D(n483), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n479) );
  IMUX40 U727 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n721), .S1(n718), .Q(n485) );
  MUX22 U728 ( .A(n494), .B(n489), .S(i_addr_Rs[4]), .Q(o_data_Rs[10]) );
  IMUX40 U729 ( .A(n495), .B(n496), .C(n497), .D(n498), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n494) );
  IMUX40 U730 ( .A(n490), .B(n491), .C(n492), .D(n493), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n489) );
  IMUX40 U731 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n728), .S1(n718), .Q(n495) );
  MUX22 U732 ( .A(n504), .B(n499), .S(i_addr_Rs[4]), .Q(o_data_Rs[11]) );
  IMUX40 U733 ( .A(n505), .B(n506), .C(n507), .D(n508), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n504) );
  IMUX40 U734 ( .A(n500), .B(n501), .C(n502), .D(n503), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n499) );
  IMUX40 U735 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n719), .S1(n712), .Q(n505) );
  MUX22 U736 ( .A(n514), .B(n509), .S(i_addr_Rs[4]), .Q(o_data_Rs[12]) );
  IMUX40 U737 ( .A(n515), .B(n516), .C(n517), .D(n518), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n514) );
  IMUX40 U738 ( .A(n510), .B(n511), .C(n512), .D(n513), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n509) );
  IMUX40 U739 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n729), .S1(i_addr_Rs[1]), .Q(n515) );
  MUX22 U740 ( .A(n524), .B(n519), .S(i_addr_Rs[4]), .Q(o_data_Rs[13]) );
  IMUX40 U741 ( .A(n525), .B(n526), .C(n527), .D(n528), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n524) );
  IMUX40 U742 ( .A(n520), .B(n521), .C(n522), .D(n523), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n519) );
  IMUX40 U743 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n730), .S1(n712), .Q(n525) );
  MUX22 U744 ( .A(n534), .B(n529), .S(i_addr_Rs[4]), .Q(o_data_Rs[14]) );
  IMUX40 U745 ( .A(n535), .B(n536), .C(n537), .D(n538), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n534) );
  IMUX40 U746 ( .A(n530), .B(n531), .C(n532), .D(n533), .S0(n710), .S1(n711), 
        .Q(n529) );
  IMUX40 U747 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n720), .S1(n716), .Q(n535) );
  MUX22 U748 ( .A(n544), .B(n539), .S(i_addr_Rs[4]), .Q(o_data_Rs[15]) );
  IMUX40 U749 ( .A(n545), .B(n546), .C(n547), .D(n548), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n544) );
  IMUX40 U750 ( .A(n540), .B(n541), .C(n542), .D(n543), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n539) );
  IMUX40 U751 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n721), .S1(n713), .Q(n545) );
  MUX22 U752 ( .A(n554), .B(n549), .S(i_addr_Rs[4]), .Q(o_data_Rs[16]) );
  IMUX40 U753 ( .A(n555), .B(n556), .C(n557), .D(n558), .S0(n710), .S1(n711), 
        .Q(n554) );
  IMUX40 U754 ( .A(n550), .B(n551), .C(n552), .D(n553), .S0(n710), .S1(n711), 
        .Q(n549) );
  IMUX40 U755 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n721), .S1(i_addr_Rs[1]), .Q(n555) );
  MUX22 U756 ( .A(n564), .B(n559), .S(i_addr_Rs[4]), .Q(o_data_Rs[17]) );
  IMUX40 U757 ( .A(n565), .B(n566), .C(n567), .D(n568), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n564) );
  IMUX40 U758 ( .A(n560), .B(n561), .C(n562), .D(n563), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n559) );
  IMUX40 U759 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n722), .S1(i_addr_Rs[1]), .Q(n565) );
  MUX22 U760 ( .A(n574), .B(n569), .S(i_addr_Rs[4]), .Q(o_data_Rs[18]) );
  IMUX40 U761 ( .A(n575), .B(n576), .C(n577), .D(n578), .S0(n710), .S1(n711), 
        .Q(n574) );
  IMUX40 U762 ( .A(n570), .B(n571), .C(n572), .D(n573), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n569) );
  IMUX40 U763 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n720), .S1(i_addr_Rs[1]), .Q(n575) );
  MUX22 U764 ( .A(n584), .B(n579), .S(i_addr_Rs[4]), .Q(o_data_Rs[19]) );
  IMUX40 U765 ( .A(n585), .B(n586), .C(n587), .D(n588), .S0(n710), .S1(n711), 
        .Q(n584) );
  IMUX40 U766 ( .A(n580), .B(n581), .C(n582), .D(n583), .S0(n710), .S1(n711), 
        .Q(n579) );
  IMUX40 U767 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n729), .S1(n718), .Q(n585) );
  MUX22 U768 ( .A(n594), .B(n589), .S(i_addr_Rs[4]), .Q(o_data_Rs[20]) );
  IMUX40 U769 ( .A(n595), .B(n596), .C(n597), .D(n598), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n594) );
  IMUX40 U770 ( .A(n590), .B(n591), .C(n592), .D(n593), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n589) );
  IMUX40 U771 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n730), .S1(i_addr_Rs[1]), .Q(n595) );
  MUX22 U772 ( .A(n604), .B(n599), .S(i_addr_Rs[4]), .Q(o_data_Rs[21]) );
  IMUX40 U773 ( .A(n605), .B(n606), .C(n607), .D(n608), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n604) );
  IMUX40 U774 ( .A(n600), .B(n601), .C(n602), .D(n603), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n599) );
  IMUX40 U775 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n728), .S1(n714), .Q(n605) );
  MUX22 U776 ( .A(n614), .B(n609), .S(i_addr_Rs[4]), .Q(o_data_Rs[22]) );
  IMUX40 U777 ( .A(n615), .B(n616), .C(n617), .D(n618), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n614) );
  IMUX40 U778 ( .A(n610), .B(n611), .C(n612), .D(n613), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n609) );
  IMUX40 U779 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n721), .S1(n714), .Q(n615) );
  MUX22 U780 ( .A(n624), .B(n619), .S(i_addr_Rs[4]), .Q(o_data_Rs[23]) );
  IMUX40 U781 ( .A(n625), .B(n626), .C(n627), .D(n628), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n624) );
  IMUX40 U782 ( .A(n620), .B(n621), .C(n622), .D(n623), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n619) );
  IMUX40 U783 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n722), .S1(n715), .Q(n625) );
  MUX22 U784 ( .A(n634), .B(n629), .S(i_addr_Rs[4]), .Q(o_data_Rs[24]) );
  IMUX40 U785 ( .A(n635), .B(n636), .C(n637), .D(n638), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n634) );
  IMUX40 U786 ( .A(n630), .B(n631), .C(n632), .D(n633), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n629) );
  IMUX40 U787 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n720), .S1(n716), .Q(n635) );
  MUX22 U788 ( .A(n644), .B(n639), .S(i_addr_Rs[4]), .Q(o_data_Rs[25]) );
  IMUX40 U789 ( .A(n645), .B(n646), .C(n647), .D(n648), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n644) );
  IMUX40 U790 ( .A(n640), .B(n641), .C(n642), .D(n643), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n639) );
  IMUX40 U791 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n721), .S1(n714), .Q(n645) );
  MUX22 U792 ( .A(n654), .B(n649), .S(i_addr_Rs[4]), .Q(o_data_Rs[26]) );
  IMUX40 U793 ( .A(n655), .B(n656), .C(n657), .D(n658), .S0(n709), .S1(n711), 
        .Q(n654) );
  IMUX40 U794 ( .A(n650), .B(n651), .C(n652), .D(n653), .S0(n709), .S1(n711), 
        .Q(n649) );
  IMUX40 U795 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n723), .S1(n716), .Q(n655) );
  MUX22 U796 ( .A(n664), .B(n659), .S(i_addr_Rs[4]), .Q(o_data_Rs[27]) );
  IMUX40 U797 ( .A(n665), .B(n666), .C(n667), .D(n668), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n664) );
  IMUX40 U798 ( .A(n660), .B(n661), .C(n662), .D(n663), .S0(n710), .S1(n711), 
        .Q(n659) );
  IMUX40 U799 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n724), .S1(n716), .Q(n665) );
  MUX22 U800 ( .A(n674), .B(n669), .S(i_addr_Rs[4]), .Q(o_data_Rs[28]) );
  IMUX40 U801 ( .A(n675), .B(n676), .C(n677), .D(n678), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n674) );
  IMUX40 U802 ( .A(n670), .B(n671), .C(n672), .D(n673), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n669) );
  IMUX40 U803 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n724), .S1(n716), .Q(n675) );
  MUX22 U804 ( .A(n684), .B(n679), .S(i_addr_Rs[4]), .Q(o_data_Rs[29]) );
  IMUX40 U805 ( .A(n685), .B(n686), .C(n687), .D(n688), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n684) );
  IMUX40 U806 ( .A(n680), .B(n681), .C(n682), .D(n683), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n679) );
  IMUX40 U807 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n725), .S1(n717), .Q(n687) );
  MUX22 U808 ( .A(n694), .B(n689), .S(i_addr_Rs[4]), .Q(o_data_Rs[30]) );
  IMUX40 U809 ( .A(n695), .B(n696), .C(n697), .D(n698), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n694) );
  IMUX40 U810 ( .A(n690), .B(n691), .C(n692), .D(n693), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n689) );
  IMUX40 U811 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n724), .S1(n717), .Q(n697) );
  MUX22 U812 ( .A(n704), .B(n699), .S(i_addr_Rs[4]), .Q(o_data_Rs[31]) );
  IMUX40 U813 ( .A(n705), .B(n706), .C(n707), .D(n708), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n704) );
  IMUX40 U814 ( .A(n700), .B(n701), .C(n702), .D(n703), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n699) );
  IMUX40 U815 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n721), .S1(n712), .Q(n707) );
  BUF2 U816 ( .A(n375), .Q(n369) );
  BUF2 U817 ( .A(i_addr_Rt[1]), .Q(n375) );
  BUF2 U818 ( .A(n718), .Q(n712) );
  BUF2 U819 ( .A(i_addr_Rs[1]), .Q(n718) );
  MUX22 U820 ( .A(n6), .B(n1), .S(i_addr_Rt[4]), .Q(o_data_Rt[0]) );
  IMUX40 U821 ( .A(n2), .B(n3), .C(n4), .D(n5), .S0(n365), .S1(i_addr_Rt[2]), 
        .Q(n1) );
  IMUX40 U822 ( .A(n7), .B(n8), .C(n9), .D(n10), .S0(n365), .S1(n368), .Q(n6)
         );
  MUX22 U823 ( .A(n16), .B(n11), .S(i_addr_Rt[4]), .Q(o_data_Rt[1]) );
  IMUX40 U824 ( .A(n17), .B(n18), .C(n19), .D(n20), .S0(n365), .S1(n368), .Q(
        n16) );
  IMUX40 U825 ( .A(n12), .B(n13), .C(n14), .D(n15), .S0(n365), .S1(n368), .Q(
        n11) );
  IMUX40 U826 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n379), .S1(n370), .Q(n17) );
  MUX22 U827 ( .A(n26), .B(n21), .S(i_addr_Rt[4]), .Q(o_data_Rt[2]) );
  IMUX40 U828 ( .A(n27), .B(n28), .C(n29), .D(n30), .S0(n366), .S1(n368), .Q(
        n26) );
  IMUX40 U829 ( .A(n22), .B(n23), .C(n24), .D(n25), .S0(n366), .S1(n368), .Q(
        n21) );
  IMUX40 U830 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n378), .S1(i_addr_Rt[1]), .Q(n27) );
  MUX22 U831 ( .A(n36), .B(n31), .S(i_addr_Rt[4]), .Q(o_data_Rt[3]) );
  IMUX40 U832 ( .A(n37), .B(n38), .C(n83), .D(n84), .S0(n366), .S1(n368), .Q(
        n36) );
  IMUX40 U833 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(n366), .S1(n368), .Q(
        n31) );
  IMUX40 U834 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n381), .S1(n369), .Q(n37) );
  MUX22 U835 ( .A(n90), .B(n85), .S(i_addr_Rt[4]), .Q(o_data_Rt[4]) );
  IMUX40 U836 ( .A(n91), .B(n92), .C(n93), .D(n94), .S0(n366), .S1(n368), .Q(
        n90) );
  IMUX40 U837 ( .A(n86), .B(n87), .C(n88), .D(n89), .S0(n366), .S1(n368), .Q(
        n85) );
  IMUX40 U838 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n376), .S1(i_addr_Rt[1]), .Q(n91) );
  MUX22 U839 ( .A(n100), .B(n95), .S(i_addr_Rt[4]), .Q(o_data_Rt[5]) );
  IMUX40 U840 ( .A(n101), .B(n102), .C(n103), .D(n104), .S0(n366), .S1(n368), 
        .Q(n100) );
  IMUX40 U841 ( .A(n96), .B(n97), .C(n98), .D(n99), .S0(n366), .S1(n368), .Q(
        n95) );
  IMUX40 U842 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n388), .S1(n375), .Q(n101) );
  MUX22 U843 ( .A(n110), .B(n105), .S(i_addr_Rt[4]), .Q(o_data_Rt[6]) );
  IMUX40 U844 ( .A(n111), .B(n112), .C(n113), .D(n114), .S0(n366), .S1(n368), 
        .Q(n110) );
  IMUX40 U845 ( .A(n106), .B(n107), .C(n108), .D(n109), .S0(n366), .S1(n368), 
        .Q(n105) );
  IMUX40 U846 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n386), .S1(i_addr_Rt[1]), .Q(n111) );
  MUX22 U847 ( .A(n120), .B(n115), .S(i_addr_Rt[4]), .Q(o_data_Rt[7]) );
  IMUX40 U848 ( .A(n121), .B(n122), .C(n123), .D(n124), .S0(n366), .S1(n368), 
        .Q(n120) );
  IMUX40 U849 ( .A(n116), .B(n117), .C(n118), .D(n119), .S0(n366), .S1(n368), 
        .Q(n115) );
  IMUX40 U850 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n386), .S1(n373), .Q(n121) );
  MUX22 U851 ( .A(n130), .B(n125), .S(i_addr_Rt[4]), .Q(o_data_Rt[8]) );
  IMUX40 U852 ( .A(n131), .B(n132), .C(n133), .D(n134), .S0(n367), .S1(n368), 
        .Q(n130) );
  IMUX40 U853 ( .A(n126), .B(n127), .C(n128), .D(n129), .S0(n367), .S1(n368), 
        .Q(n125) );
  IMUX40 U854 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n385), .S1(n375), .Q(n131) );
  MUX22 U855 ( .A(n140), .B(n135), .S(i_addr_Rt[4]), .Q(o_data_Rt[9]) );
  IMUX40 U856 ( .A(n141), .B(n142), .C(n143), .D(n144), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n140) );
  IMUX40 U857 ( .A(n136), .B(n137), .C(n138), .D(n139), .S0(n367), .S1(n368), 
        .Q(n135) );
  IMUX40 U858 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n388), .S1(i_addr_Rt[1]), .Q(n141) );
  MUX22 U859 ( .A(n150), .B(n145), .S(i_addr_Rt[4]), .Q(o_data_Rt[10]) );
  IMUX40 U860 ( .A(n151), .B(n152), .C(n153), .D(n154), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n150) );
  IMUX40 U861 ( .A(n146), .B(n147), .C(n148), .D(n149), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n145) );
  IMUX40 U862 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n385), .S1(i_addr_Rt[1]), .Q(n151) );
  MUX22 U863 ( .A(n160), .B(n155), .S(i_addr_Rt[4]), .Q(o_data_Rt[11]) );
  IMUX40 U864 ( .A(n161), .B(n162), .C(n163), .D(n164), .S0(n367), .S1(n368), 
        .Q(n160) );
  IMUX40 U865 ( .A(n156), .B(n157), .C(n158), .D(n159), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n155) );
  IMUX40 U866 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n376), .S1(n371), .Q(n161) );
  MUX22 U867 ( .A(n170), .B(n165), .S(i_addr_Rt[4]), .Q(o_data_Rt[12]) );
  IMUX40 U868 ( .A(n171), .B(n172), .C(n173), .D(n174), .S0(n367), .S1(n368), 
        .Q(n170) );
  IMUX40 U869 ( .A(n166), .B(n167), .C(n168), .D(n169), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n165) );
  IMUX40 U870 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n377), .S1(i_addr_Rt[1]), .Q(n171) );
  MUX22 U871 ( .A(n180), .B(n175), .S(i_addr_Rt[4]), .Q(o_data_Rt[13]) );
  IMUX40 U872 ( .A(n181), .B(n182), .C(n183), .D(n184), .S0(n367), .S1(n368), 
        .Q(n180) );
  IMUX40 U873 ( .A(n176), .B(n177), .C(n178), .D(n179), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n175) );
  IMUX40 U874 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n377), .S1(n375), .Q(n181) );
  MUX22 U875 ( .A(n190), .B(n185), .S(i_addr_Rt[4]), .Q(o_data_Rt[14]) );
  IMUX40 U876 ( .A(n191), .B(n192), .C(n193), .D(n194), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n190) );
  IMUX40 U877 ( .A(n186), .B(n187), .C(n188), .D(n189), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n185) );
  IMUX40 U878 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n378), .S1(n371), .Q(n191) );
  MUX22 U879 ( .A(n200), .B(n195), .S(i_addr_Rt[4]), .Q(o_data_Rt[15]) );
  IMUX40 U880 ( .A(n201), .B(n202), .C(n203), .D(n204), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n200) );
  IMUX40 U881 ( .A(n196), .B(n197), .C(n198), .D(n199), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n195) );
  IMUX40 U882 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n380), .S1(i_addr_Rt[1]), .Q(n201) );
  MUX22 U883 ( .A(n210), .B(n205), .S(i_addr_Rt[4]), .Q(o_data_Rt[16]) );
  IMUX40 U884 ( .A(n211), .B(n212), .C(n213), .D(n214), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n210) );
  IMUX40 U885 ( .A(n206), .B(n207), .C(n208), .D(n209), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n205) );
  IMUX40 U886 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n382), .S1(n372), .Q(n211) );
  MUX22 U887 ( .A(n220), .B(n215), .S(i_addr_Rt[4]), .Q(o_data_Rt[17]) );
  IMUX40 U888 ( .A(n221), .B(n222), .C(n223), .D(n224), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n220) );
  IMUX40 U889 ( .A(n216), .B(n217), .C(n218), .D(n219), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n215) );
  IMUX40 U890 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n384), .S1(n370), .Q(n221) );
  MUX22 U891 ( .A(n230), .B(n225), .S(i_addr_Rt[4]), .Q(o_data_Rt[18]) );
  IMUX40 U892 ( .A(n231), .B(n232), .C(n233), .D(n234), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n230) );
  IMUX40 U893 ( .A(n226), .B(n227), .C(n228), .D(n229), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n225) );
  IMUX40 U894 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n379), .S1(n370), .Q(n231) );
  MUX22 U895 ( .A(n240), .B(n235), .S(i_addr_Rt[4]), .Q(o_data_Rt[19]) );
  IMUX40 U896 ( .A(n241), .B(n242), .C(n243), .D(n244), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n240) );
  IMUX40 U897 ( .A(n236), .B(n237), .C(n238), .D(n239), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n235) );
  IMUX40 U898 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n379), .S1(i_addr_Rt[1]), .Q(n241) );
  MUX22 U899 ( .A(n250), .B(n245), .S(i_addr_Rt[4]), .Q(o_data_Rt[20]) );
  IMUX40 U900 ( .A(n251), .B(n252), .C(n253), .D(n254), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n250) );
  IMUX40 U901 ( .A(n246), .B(n247), .C(n248), .D(n249), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n245) );
  IMUX40 U902 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n380), .S1(i_addr_Rt[1]), .Q(n251) );
  MUX22 U903 ( .A(n260), .B(n255), .S(i_addr_Rt[4]), .Q(o_data_Rt[21]) );
  IMUX40 U904 ( .A(n261), .B(n262), .C(n263), .D(n264), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n260) );
  IMUX40 U905 ( .A(n256), .B(n257), .C(n258), .D(n259), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n255) );
  IMUX40 U906 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n377), .S1(n371), .Q(n261) );
  MUX22 U907 ( .A(n270), .B(n265), .S(i_addr_Rt[4]), .Q(o_data_Rt[22]) );
  IMUX40 U908 ( .A(n271), .B(n272), .C(n273), .D(n274), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n270) );
  IMUX40 U909 ( .A(n266), .B(n267), .C(n268), .D(n269), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n265) );
  IMUX40 U910 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n378), .S1(n371), .Q(n271) );
  MUX22 U911 ( .A(n280), .B(n275), .S(i_addr_Rt[4]), .Q(o_data_Rt[23]) );
  IMUX40 U912 ( .A(n281), .B(n282), .C(n283), .D(n284), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n280) );
  IMUX40 U913 ( .A(n276), .B(n277), .C(n278), .D(n279), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n275) );
  IMUX40 U914 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n381), .S1(n373), .Q(n281) );
  MUX22 U915 ( .A(n290), .B(n285), .S(i_addr_Rt[4]), .Q(o_data_Rt[24]) );
  IMUX40 U916 ( .A(n291), .B(n292), .C(n293), .D(n294), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n290) );
  IMUX40 U917 ( .A(n286), .B(n287), .C(n288), .D(n289), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n285) );
  IMUX40 U918 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n382), .S1(n374), .Q(n291) );
  MUX22 U919 ( .A(n300), .B(n295), .S(i_addr_Rt[4]), .Q(o_data_Rt[25]) );
  IMUX40 U920 ( .A(n301), .B(n302), .C(n303), .D(n304), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n300) );
  IMUX40 U921 ( .A(n296), .B(n297), .C(n298), .D(n299), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n295) );
  IMUX40 U922 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n382), .S1(n369), .Q(n301) );
  MUX22 U923 ( .A(n310), .B(n305), .S(i_addr_Rt[4]), .Q(o_data_Rt[26]) );
  IMUX40 U924 ( .A(n311), .B(n312), .C(n313), .D(n314), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n310) );
  IMUX40 U925 ( .A(n306), .B(n307), .C(n308), .D(n309), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n305) );
  IMUX40 U926 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n382), .S1(n372), .Q(n311) );
  MUX22 U927 ( .A(n320), .B(n315), .S(i_addr_Rt[4]), .Q(o_data_Rt[27]) );
  IMUX40 U928 ( .A(n321), .B(n322), .C(n323), .D(n324), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n320) );
  IMUX40 U929 ( .A(n316), .B(n317), .C(n318), .D(n319), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n315) );
  IMUX40 U930 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n383), .S1(n374), .Q(n321) );
  MUX22 U931 ( .A(n330), .B(n325), .S(i_addr_Rt[4]), .Q(o_data_Rt[28]) );
  IMUX40 U932 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n330) );
  IMUX40 U933 ( .A(n326), .B(n327), .C(n328), .D(n329), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n325) );
  IMUX40 U934 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n383), .S1(n372), .Q(n331) );
  MUX22 U935 ( .A(n340), .B(n335), .S(i_addr_Rt[4]), .Q(o_data_Rt[29]) );
  IMUX40 U936 ( .A(n341), .B(n342), .C(n343), .D(n344), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n340) );
  IMUX40 U937 ( .A(n336), .B(n337), .C(n338), .D(n339), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n335) );
  IMUX40 U938 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n384), .S1(n373), .Q(n341) );
  MUX22 U939 ( .A(n350), .B(n345), .S(i_addr_Rt[4]), .Q(o_data_Rt[30]) );
  IMUX40 U940 ( .A(n351), .B(n352), .C(n353), .D(n354), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n350) );
  IMUX40 U941 ( .A(n346), .B(n347), .C(n348), .D(n349), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n345) );
  IMUX40 U942 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        i_addr_Rt[0]), .S1(n374), .Q(n351) );
  MUX22 U943 ( .A(n360), .B(n355), .S(i_addr_Rt[4]), .Q(o_data_Rt[31]) );
  IMUX40 U944 ( .A(n361), .B(n362), .C(n363), .D(n364), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n360) );
  IMUX40 U945 ( .A(n356), .B(n357), .C(n358), .D(n359), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n355) );
  IMUX40 U946 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n381), .S1(n374), .Q(n361) );
  BUF2 U947 ( .A(i_addr_Rt[2]), .Q(n368) );
  BUF2 U948 ( .A(i_addr_Rt[3]), .Q(n365) );
endmodule


module D_shiftleft ( i_data_immE, o_data_immshiftl );
  input [15:0] i_data_immE;
  output [31:0] o_data_immshiftl;
  wire   n1;
  assign o_data_immshiftl[0] = o_data_immshiftl[1];
  assign o_data_immshiftl[19] = o_data_immshiftl[30];
  assign o_data_immshiftl[29] = o_data_immshiftl[30];
  assign o_data_immshiftl[25] = o_data_immshiftl[30];
  assign o_data_immshiftl[21] = o_data_immshiftl[30];
  assign o_data_immshiftl[31] = o_data_immshiftl[30];
  assign o_data_immshiftl[20] = o_data_immshiftl[30];
  assign o_data_immshiftl[27] = o_data_immshiftl[30];
  assign o_data_immshiftl[26] = o_data_immshiftl[30];
  assign o_data_immshiftl[22] = o_data_immshiftl[30];
  assign o_data_immshiftl[24] = i_data_immE[15];
  assign o_data_immshiftl[28] = i_data_immE[15];
  assign o_data_immshiftl[17] = i_data_immE[15];
  assign o_data_immshiftl[18] = i_data_immE[15];
  assign o_data_immshiftl[23] = i_data_immE[15];
  assign o_data_immshiftl[16] = i_data_immE[14];
  assign o_data_immshiftl[15] = i_data_immE[13];
  assign o_data_immshiftl[14] = i_data_immE[12];
  assign o_data_immshiftl[13] = i_data_immE[11];
  assign o_data_immshiftl[12] = i_data_immE[10];
  assign o_data_immshiftl[11] = i_data_immE[9];
  assign o_data_immshiftl[10] = i_data_immE[8];
  assign o_data_immshiftl[9] = i_data_immE[7];
  assign o_data_immshiftl[8] = i_data_immE[6];
  assign o_data_immshiftl[7] = i_data_immE[5];
  assign o_data_immshiftl[6] = i_data_immE[4];
  assign o_data_immshiftl[5] = i_data_immE[3];
  assign o_data_immshiftl[4] = i_data_immE[2];
  assign o_data_immshiftl[3] = i_data_immE[1];
  assign o_data_immshiftl[2] = i_data_immE[0];

  INV3 U2 ( .A(n1), .Q(o_data_immshiftl[30]) );
  INV3 U3 ( .A(i_data_immE[15]), .Q(n1) );
  LOGIC0 U4 ( .Q(o_data_immshiftl[1]) );
endmodule


module D_sign_extend ( i_data_immD, i_con_signext, o_data_immD );
  input [15:0] i_data_immD;
  output [31:0] o_data_immD;
  input i_con_signext;
  wire   n2;
  assign o_data_immD[15] = i_data_immD[15];
  assign o_data_immD[14] = i_data_immD[14];
  assign o_data_immD[13] = i_data_immD[13];
  assign o_data_immD[12] = i_data_immD[12];
  assign o_data_immD[11] = i_data_immD[11];
  assign o_data_immD[10] = i_data_immD[10];
  assign o_data_immD[9] = i_data_immD[9];
  assign o_data_immD[8] = i_data_immD[8];
  assign o_data_immD[7] = i_data_immD[7];
  assign o_data_immD[6] = i_data_immD[6];
  assign o_data_immD[5] = i_data_immD[5];
  assign o_data_immD[4] = i_data_immD[4];
  assign o_data_immD[3] = i_data_immD[3];
  assign o_data_immD[2] = i_data_immD[2];
  assign o_data_immD[1] = i_data_immD[1];
  assign o_data_immD[0] = i_data_immD[0];
  assign o_data_immD[16] = o_data_immD[31];
  assign o_data_immD[17] = o_data_immD[31];
  assign o_data_immD[18] = o_data_immD[31];
  assign o_data_immD[19] = o_data_immD[31];
  assign o_data_immD[20] = o_data_immD[31];
  assign o_data_immD[21] = o_data_immD[31];
  assign o_data_immD[22] = o_data_immD[31];
  assign o_data_immD[23] = o_data_immD[31];
  assign o_data_immD[24] = o_data_immD[31];
  assign o_data_immD[25] = o_data_immD[31];
  assign o_data_immD[26] = o_data_immD[31];
  assign o_data_immD[27] = o_data_immD[31];
  assign o_data_immD[28] = o_data_immD[31];
  assign o_data_immD[29] = o_data_immD[31];
  assign o_data_immD[30] = o_data_immD[31];

  INV3 U2 ( .A(n2), .Q(o_data_immD[31]) );
  NAND22 U3 ( .A(i_con_signext), .B(i_data_immD[15]), .Q(n2) );
endmodule


module D_jump_ext ( i_addr_j, i_PC4_j, o_addr_j );
  input [25:0] i_addr_j;
  input [3:0] i_PC4_j;
  output [31:0] o_addr_j;

  assign o_addr_j[0] = o_addr_j[1];
  assign o_addr_j[31] = i_PC4_j[3];
  assign o_addr_j[30] = i_PC4_j[2];
  assign o_addr_j[29] = i_PC4_j[1];
  assign o_addr_j[28] = i_PC4_j[0];
  assign o_addr_j[27] = i_addr_j[25];
  assign o_addr_j[26] = i_addr_j[24];
  assign o_addr_j[25] = i_addr_j[23];
  assign o_addr_j[24] = i_addr_j[22];
  assign o_addr_j[23] = i_addr_j[21];
  assign o_addr_j[22] = i_addr_j[20];
  assign o_addr_j[21] = i_addr_j[19];
  assign o_addr_j[20] = i_addr_j[18];
  assign o_addr_j[19] = i_addr_j[17];
  assign o_addr_j[18] = i_addr_j[16];
  assign o_addr_j[17] = i_addr_j[15];
  assign o_addr_j[16] = i_addr_j[14];
  assign o_addr_j[15] = i_addr_j[13];
  assign o_addr_j[14] = i_addr_j[12];
  assign o_addr_j[13] = i_addr_j[11];
  assign o_addr_j[12] = i_addr_j[10];
  assign o_addr_j[11] = i_addr_j[9];
  assign o_addr_j[10] = i_addr_j[8];
  assign o_addr_j[9] = i_addr_j[7];
  assign o_addr_j[8] = i_addr_j[6];
  assign o_addr_j[7] = i_addr_j[5];
  assign o_addr_j[6] = i_addr_j[4];
  assign o_addr_j[5] = i_addr_j[3];
  assign o_addr_j[4] = i_addr_j[2];
  assign o_addr_j[3] = i_addr_j[1];
  assign o_addr_j[2] = i_addr_j[0];

  LOGIC0 U2 ( .Q(o_addr_j[1]) );
endmodule


module E_forward ( i_addr_rs, i_addr_rt, i_addr_rdM, i_addr_rdW, i_addr_rtM, 
        i_addr_rtW, i_con_regwriteM, i_con_regwriteW, i_con_memreadM, 
        i_con_memreadW, o_con_fa, o_con_fb, o_con_cmpalu, o_con_cmpmem );
  input [4:0] i_addr_rs;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rdM;
  input [4:0] i_addr_rdW;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  output [2:0] o_con_fa;
  output [2:0] o_con_fb;
  input i_con_regwriteM, i_con_regwriteW, i_con_memreadM, i_con_memreadW;
  output o_con_cmpalu, o_con_cmpmem;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82;

  OAI310 U1 ( .A(n1), .B(n2), .C(n3), .D(n4), .Q(o_con_fb[2]) );
  OAI210 U2 ( .A(n5), .B(n6), .C(n4), .Q(o_con_fb[0]) );
  NAND30 U3 ( .A(n7), .B(n8), .C(i_con_memreadW), .Q(n4) );
  CLKIN0 U4 ( .A(n9), .Q(n7) );
  NAND40 U5 ( .A(n10), .B(n11), .C(n12), .D(n13), .Q(n6) );
  XNR20 U6 ( .A(i_addr_rt[1]), .B(i_addr_rdW[1]), .Q(n13) );
  XNR20 U7 ( .A(i_addr_rt[2]), .B(i_addr_rdW[2]), .Q(n12) );
  XNR20 U8 ( .A(i_addr_rt[3]), .B(i_addr_rdW[3]), .Q(n11) );
  XNR20 U9 ( .A(i_addr_rt[4]), .B(i_addr_rdW[4]), .Q(n10) );
  NAND40 U10 ( .A(n14), .B(i_con_regwriteW), .C(n15), .D(n16), .Q(n5) );
  CLKIN0 U11 ( .A(n17), .Q(n15) );
  XNR20 U12 ( .A(i_addr_rt[0]), .B(i_addr_rdW[0]), .Q(n14) );
  NOR20 U13 ( .A(o_con_fa[2]), .B(n18), .Q(o_con_fa[1]) );
  CLKIN0 U14 ( .A(n19), .Q(n18) );
  OAI210 U15 ( .A(o_con_cmpmem), .B(n20), .C(n21), .Q(o_con_fa[0]) );
  NAND20 U16 ( .A(n22), .B(n23), .Q(n21) );
  NOR40 U17 ( .A(o_con_fa[2]), .B(n19), .C(n24), .D(n25), .Q(n23) );
  XOR20 U18 ( .A(i_addr_rdW[0]), .B(i_addr_rs[0]), .Q(n25) );
  CLKIN0 U19 ( .A(i_con_regwriteW), .Q(n24) );
  NOR40 U20 ( .A(n26), .B(n27), .C(n28), .D(n29), .Q(n19) );
  OAI310 U21 ( .A(i_addr_rdM[0]), .B(i_addr_rdM[1]), .C(n30), .D(
        i_con_regwriteM), .Q(n28) );
  CLKIN0 U22 ( .A(n31), .Q(n30) );
  NOR30 U23 ( .A(i_addr_rdM[2]), .B(i_addr_rdM[4]), .C(i_addr_rdM[3]), .Q(n31)
         );
  NAND20 U24 ( .A(n32), .B(n20), .Q(o_con_fa[2]) );
  NOR40 U25 ( .A(n33), .B(n34), .C(n35), .D(n36), .Q(n22) );
  IMUX20 U26 ( .A(n37), .B(i_addr_rs[4]), .S(i_addr_rdW[4]), .Q(n36) );
  NOR20 U27 ( .A(n38), .B(i_addr_rs[4]), .Q(n37) );
  NOR40 U28 ( .A(i_addr_rdW[3]), .B(i_addr_rdW[2]), .C(i_addr_rdW[1]), .D(
        i_addr_rdW[0]), .Q(n38) );
  XOR20 U29 ( .A(i_addr_rdW[3]), .B(i_addr_rs[3]), .Q(n35) );
  XOR20 U30 ( .A(i_addr_rdW[2]), .B(i_addr_rs[2]), .Q(n34) );
  XOR20 U31 ( .A(i_addr_rdW[1]), .B(i_addr_rs[1]), .Q(n33) );
  NAND40 U32 ( .A(n39), .B(n40), .C(n41), .D(n42), .Q(n20) );
  NOR40 U33 ( .A(n43), .B(n44), .C(n45), .D(n46), .Q(n42) );
  XNR20 U34 ( .A(n47), .B(i_addr_rs[1]), .Q(n46) );
  XOR20 U35 ( .A(i_addr_rtW[0]), .B(i_addr_rs[0]), .Q(n45) );
  XNR20 U36 ( .A(i_addr_rtW[3]), .B(i_addr_rs[3]), .Q(n41) );
  XNR20 U37 ( .A(i_addr_rtW[4]), .B(i_addr_rs[4]), .Q(n40) );
  XNR20 U38 ( .A(i_addr_rtW[2]), .B(i_addr_rs[2]), .Q(n39) );
  NOR20 U39 ( .A(n17), .B(n16), .Q(o_con_fb[1]) );
  NAND40 U40 ( .A(n48), .B(i_con_regwriteM), .C(n49), .D(n50), .Q(n16) );
  NOR30 U41 ( .A(n51), .B(n52), .C(n53), .Q(n50) );
  XOR20 U42 ( .A(i_addr_rdM[2]), .B(i_addr_rt[2]), .Q(n53) );
  XOR20 U43 ( .A(i_addr_rdM[4]), .B(i_addr_rt[4]), .Q(n52) );
  XOR20 U44 ( .A(i_addr_rdM[3]), .B(i_addr_rt[3]), .Q(n51) );
  XNR20 U45 ( .A(i_addr_rt[0]), .B(i_addr_rdM[0]), .Q(n49) );
  XNR20 U46 ( .A(i_addr_rt[1]), .B(i_addr_rdM[1]), .Q(n48) );
  OAI210 U47 ( .A(n9), .B(n44), .C(n8), .Q(n17) );
  AOI210 U48 ( .A(n54), .B(i_con_memreadM), .C(n2), .Q(n8) );
  NOR30 U49 ( .A(i_addr_rt[0]), .B(i_addr_rt[1]), .C(n55), .Q(n2) );
  CLKIN0 U50 ( .A(n56), .Q(n55) );
  NOR30 U51 ( .A(i_addr_rt[2]), .B(i_addr_rt[4]), .C(i_addr_rt[3]), .Q(n56) );
  CLKIN0 U52 ( .A(n3), .Q(n54) );
  NAND40 U53 ( .A(n57), .B(n58), .C(n59), .D(n60), .Q(n3) );
  XNR20 U54 ( .A(i_addr_rt[0]), .B(i_addr_rtM[0]), .Q(n60) );
  NOR20 U55 ( .A(n61), .B(n62), .Q(n59) );
  XOR20 U56 ( .A(i_addr_rtM[3]), .B(i_addr_rt[3]), .Q(n62) );
  XNR20 U57 ( .A(n63), .B(i_addr_rt[1]), .Q(n61) );
  XNR20 U58 ( .A(i_addr_rt[2]), .B(i_addr_rtM[2]), .Q(n58) );
  XNR20 U59 ( .A(i_addr_rt[4]), .B(i_addr_rtM[4]), .Q(n57) );
  CLKIN0 U60 ( .A(i_con_memreadW), .Q(n44) );
  NAND40 U61 ( .A(n64), .B(n65), .C(n66), .D(n67), .Q(n9) );
  XNR20 U62 ( .A(i_addr_rt[0]), .B(i_addr_rtW[0]), .Q(n67) );
  NOR20 U63 ( .A(n68), .B(n69), .Q(n66) );
  XOR20 U64 ( .A(i_addr_rtW[3]), .B(i_addr_rt[3]), .Q(n69) );
  XNR20 U65 ( .A(n47), .B(i_addr_rt[1]), .Q(n68) );
  CLKIN0 U66 ( .A(i_addr_rtW[1]), .Q(n47) );
  XNR20 U67 ( .A(i_addr_rt[2]), .B(i_addr_rtW[2]), .Q(n65) );
  XNR20 U68 ( .A(i_addr_rt[4]), .B(i_addr_rtW[4]), .Q(n64) );
  CLKIN0 U69 ( .A(n32), .Q(o_con_cmpmem) );
  NAND40 U70 ( .A(n70), .B(n71), .C(n72), .D(n73), .Q(n32) );
  NOR40 U71 ( .A(n43), .B(n1), .C(n74), .D(n75), .Q(n73) );
  XNR20 U72 ( .A(n63), .B(i_addr_rs[1]), .Q(n75) );
  CLKIN0 U73 ( .A(i_addr_rtM[1]), .Q(n63) );
  XOR20 U74 ( .A(i_addr_rtM[0]), .B(i_addr_rs[0]), .Q(n74) );
  CLKIN0 U75 ( .A(i_con_memreadM), .Q(n1) );
  XNR20 U76 ( .A(i_addr_rtM[3]), .B(i_addr_rs[3]), .Q(n72) );
  XNR20 U77 ( .A(i_addr_rtM[4]), .B(i_addr_rs[4]), .Q(n71) );
  XNR20 U78 ( .A(i_addr_rtM[2]), .B(i_addr_rs[2]), .Q(n70) );
  NOR40 U79 ( .A(n29), .B(n76), .C(n27), .D(n26), .Q(o_con_cmpalu) );
  XOR20 U80 ( .A(i_addr_rs[4]), .B(i_addr_rdM[4]), .Q(n26) );
  NAND30 U81 ( .A(n77), .B(n78), .C(n79), .Q(n27) );
  XNR20 U82 ( .A(i_addr_rs[1]), .B(i_addr_rdM[1]), .Q(n79) );
  XNR20 U83 ( .A(i_addr_rs[2]), .B(i_addr_rdM[2]), .Q(n78) );
  XNR20 U84 ( .A(i_addr_rs[0]), .B(i_addr_rdM[0]), .Q(n77) );
  NAND20 U85 ( .A(i_con_regwriteM), .B(n80), .Q(n76) );
  CLKIN0 U86 ( .A(n43), .Q(n80) );
  NOR30 U87 ( .A(i_addr_rs[0]), .B(i_addr_rs[1]), .C(n81), .Q(n43) );
  CLKIN0 U88 ( .A(n82), .Q(n81) );
  NOR30 U89 ( .A(i_addr_rs[2]), .B(i_addr_rs[4]), .C(i_addr_rs[3]), .Q(n82) );
  XOR20 U90 ( .A(i_addr_rs[3]), .B(i_addr_rdM[3]), .Q(n29) );
endmodule


module decode ( i_clk, i_nrst, i_addr_pc4, i_data_instr, i_con_Wregwrite, 
        i_data_Wregwrite, i_addr_Wregwrite, i_addr_Erd, i_addr_Mrd, 
        i_con_Eregwrite, i_con_Mregwrite, i_addr_rtM, i_addr_rtW, 
        i_con_memreadM, i_con_memreadW, o_data_rs, o_data_rt, o_addr_rd, 
        o_addr_rt, o_data_jr, o_con_jump, o_addr_pc4, o_addr_branch, 
        o_addr_jump, o_con_Ealuop, o_con_Ealusrc, o_con_Eregdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Wloadmux, o_con_Walupc8, 
        o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall, o_con_Ebop, 
        o_data_signext, o_con_Efamux, o_con_Efbmux, o_data_Fmemout );
  input [31:0] i_addr_pc4;
  input [31:0] i_data_instr;
  input [31:0] i_data_Wregwrite;
  input [4:0] i_addr_Wregwrite;
  input [4:0] i_addr_Erd;
  input [4:0] i_addr_Mrd;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  output [31:0] o_data_rs;
  output [31:0] o_data_rt;
  output [4:0] o_addr_rd;
  output [4:0] o_addr_rt;
  output [31:0] o_data_jr;
  output [1:0] o_con_jump;
  output [31:0] o_addr_pc4;
  output [31:0] o_addr_branch;
  output [31:0] o_addr_jump;
  output [5:0] o_con_Ealuop;
  output [1:0] o_con_Wloadmux;
  output [2:0] o_con_Ebop;
  output [31:0] o_data_signext;
  output [2:0] o_con_Efamux;
  output [2:0] o_con_Efbmux;
  output [31:0] o_data_Fmemout;
  input i_clk, i_nrst, i_con_Wregwrite, i_con_Eregwrite, i_con_Mregwrite,
         i_con_memreadM, i_con_memreadW;
  output o_con_Ealusrc, o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite,
         o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall;
  wire   control_o_con_alusrc, control_o_con_regdst, jbcon_o_con_aluPC4,
         control_o_con_memread, control_o_con_memwrite, control_o_con_memtoreg,
         control_o_con_regwrite, signext_i_con_signext, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;
  wire   [31:0] regbank_o_data_Rt;
  wire   [5:0] control_o_con_aluop;
  wire   [1:0] control_o_con_loadsig;
  wire   [31:0] signext_o_data_immD;
  wire   [2:0] for_o_con_fa;
  wire   [2:0] for_o_con_fb;
  wire   [31:0] pcadd_o_addr_pcbranchE;
  wire   [2:0] jbcon_o_con_bop;
  wire   [31:2] pcadd_i_data_immshiftl;
  assign o_addr_jump[1] = o_addr_jump[0];

  DFC3 pipe_bop_reg_2_ ( .D(jbcon_o_con_bop[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[2]) );
  DFC3 pipe_bop_reg_1_ ( .D(jbcon_o_con_bop[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[1]) );
  DFC3 pipe_bop_reg_0_ ( .D(jbcon_o_con_bop[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[0]) );
  DFC3 pipe_data_rs_reg_31_ ( .D(o_data_jr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[31]) );
  DFC3 pipe_data_rs_reg_30_ ( .D(o_data_jr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[30]) );
  DFC3 pipe_data_rs_reg_29_ ( .D(o_data_jr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[29]) );
  DFC3 pipe_data_rs_reg_28_ ( .D(o_data_jr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[28]) );
  DFC3 pipe_data_rs_reg_27_ ( .D(o_data_jr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[27]) );
  DFC3 pipe_data_rs_reg_26_ ( .D(o_data_jr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[26]) );
  DFC3 pipe_data_rs_reg_25_ ( .D(o_data_jr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[25]) );
  DFC3 pipe_data_rs_reg_24_ ( .D(o_data_jr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[24]) );
  DFC3 pipe_data_rs_reg_23_ ( .D(o_data_jr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[23]) );
  DFC3 pipe_data_rs_reg_22_ ( .D(o_data_jr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[22]) );
  DFC3 pipe_data_rs_reg_21_ ( .D(o_data_jr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[21]) );
  DFC3 pipe_data_rs_reg_20_ ( .D(o_data_jr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[20]) );
  DFC3 pipe_data_rs_reg_19_ ( .D(o_data_jr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[19]) );
  DFC3 pipe_data_rs_reg_18_ ( .D(o_data_jr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[18]) );
  DFC3 pipe_data_rs_reg_17_ ( .D(o_data_jr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[17]) );
  DFC3 pipe_data_rs_reg_16_ ( .D(o_data_jr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[16]) );
  DFC3 pipe_data_rs_reg_15_ ( .D(o_data_jr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[15]) );
  DFC3 pipe_data_rs_reg_14_ ( .D(o_data_jr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[14]) );
  DFC3 pipe_data_rs_reg_13_ ( .D(o_data_jr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[13]) );
  DFC3 pipe_data_rs_reg_12_ ( .D(o_data_jr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[12]) );
  DFC3 pipe_data_rs_reg_11_ ( .D(o_data_jr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[11]) );
  DFC3 pipe_data_rs_reg_10_ ( .D(o_data_jr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[10]) );
  DFC3 pipe_data_rs_reg_9_ ( .D(o_data_jr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[9]) );
  DFC3 pipe_data_rs_reg_8_ ( .D(o_data_jr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[8]) );
  DFC3 pipe_data_rs_reg_7_ ( .D(o_data_jr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[7]) );
  DFC3 pipe_data_rs_reg_6_ ( .D(o_data_jr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[6]) );
  DFC3 pipe_data_rs_reg_5_ ( .D(o_data_jr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[5]) );
  DFC3 pipe_data_rs_reg_4_ ( .D(o_data_jr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[4]) );
  DFC3 pipe_data_rs_reg_3_ ( .D(o_data_jr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[3]) );
  DFC3 pipe_data_rs_reg_2_ ( .D(o_data_jr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[2]) );
  DFC3 pipe_data_rs_reg_1_ ( .D(o_data_jr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[1]) );
  DFC3 pipe_data_rs_reg_0_ ( .D(o_data_jr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[0]) );
  DFC3 pipe_data_rt_reg_31_ ( .D(regbank_o_data_Rt[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[31]) );
  DFC3 pipe_data_rt_reg_30_ ( .D(regbank_o_data_Rt[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC3 pipe_data_rt_reg_29_ ( .D(regbank_o_data_Rt[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[29]) );
  DFC3 pipe_data_rt_reg_28_ ( .D(regbank_o_data_Rt[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28]) );
  DFC3 pipe_data_rt_reg_27_ ( .D(regbank_o_data_Rt[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27]) );
  DFC3 pipe_data_rt_reg_26_ ( .D(regbank_o_data_Rt[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26]) );
  DFC3 pipe_data_rt_reg_25_ ( .D(regbank_o_data_Rt[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25]) );
  DFC3 pipe_data_rt_reg_24_ ( .D(regbank_o_data_Rt[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24]) );
  DFC3 pipe_data_rt_reg_23_ ( .D(regbank_o_data_Rt[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23]) );
  DFC3 pipe_data_rt_reg_22_ ( .D(regbank_o_data_Rt[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC3 pipe_data_rt_reg_21_ ( .D(regbank_o_data_Rt[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21]) );
  DFC3 pipe_data_rt_reg_20_ ( .D(regbank_o_data_Rt[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20]) );
  DFC3 pipe_data_rt_reg_19_ ( .D(regbank_o_data_Rt[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19]) );
  DFC3 pipe_data_rt_reg_18_ ( .D(regbank_o_data_Rt[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18]) );
  DFC3 pipe_data_rt_reg_17_ ( .D(regbank_o_data_Rt[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17]) );
  DFC3 pipe_data_rt_reg_16_ ( .D(regbank_o_data_Rt[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC3 pipe_data_rt_reg_15_ ( .D(regbank_o_data_Rt[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15]) );
  DFC3 pipe_data_rt_reg_14_ ( .D(regbank_o_data_Rt[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14]) );
  DFC3 pipe_data_rt_reg_13_ ( .D(regbank_o_data_Rt[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC3 pipe_data_rt_reg_12_ ( .D(regbank_o_data_Rt[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12]) );
  DFC3 pipe_data_rt_reg_11_ ( .D(regbank_o_data_Rt[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11]) );
  DFC3 pipe_data_rt_reg_10_ ( .D(regbank_o_data_Rt[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC3 pipe_data_rt_reg_9_ ( .D(regbank_o_data_Rt[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[9]) );
  DFC3 pipe_data_rt_reg_8_ ( .D(regbank_o_data_Rt[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[8]) );
  DFC3 pipe_data_rt_reg_7_ ( .D(regbank_o_data_Rt[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[7]) );
  DFC3 pipe_data_rt_reg_6_ ( .D(regbank_o_data_Rt[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[6]) );
  DFC3 pipe_data_rt_reg_5_ ( .D(regbank_o_data_Rt[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[5]) );
  DFC3 pipe_data_rt_reg_4_ ( .D(regbank_o_data_Rt[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[4]) );
  DFC3 pipe_data_rt_reg_3_ ( .D(regbank_o_data_Rt[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[3]) );
  DFC3 pipe_data_rt_reg_2_ ( .D(regbank_o_data_Rt[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[2]) );
  DFC3 pipe_data_rt_reg_1_ ( .D(regbank_o_data_Rt[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[1]) );
  DFC3 pipe_data_rt_reg_0_ ( .D(regbank_o_data_Rt[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[0]) );
  DFC3 pipe_addr_rd_reg_4_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[4]) );
  DFC3 pipe_addr_rd_reg_3_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[3]) );
  DFC3 pipe_addr_rd_reg_2_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[2]) );
  DFC3 pipe_addr_rd_reg_1_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[1]) );
  DFC3 pipe_addr_rd_reg_0_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[0]) );
  DFC3 pipe_addr_rt_reg_4_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[0]) );
  DFC3 pipe_addr_pc4_reg_31_ ( .D(i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_addr_pc4_reg_30_ ( .D(i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_addr_pc4_reg_29_ ( .D(i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_addr_pc4_reg_28_ ( .D(i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_addr_pc4_reg_27_ ( .D(i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_addr_pc4_reg_26_ ( .D(i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_addr_pc4_reg_25_ ( .D(i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_addr_pc4_reg_24_ ( .D(i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_addr_pc4_reg_23_ ( .D(i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_addr_pc4_reg_22_ ( .D(i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_addr_pc4_reg_21_ ( .D(i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_addr_pc4_reg_20_ ( .D(i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_addr_pc4_reg_19_ ( .D(i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_addr_pc4_reg_18_ ( .D(i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_addr_pc4_reg_17_ ( .D(i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_addr_pc4_reg_16_ ( .D(i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_addr_pc4_reg_15_ ( .D(i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_addr_pc4_reg_14_ ( .D(i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_addr_pc4_reg_13_ ( .D(i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_addr_pc4_reg_12_ ( .D(i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_addr_pc4_reg_11_ ( .D(i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_addr_pc4_reg_10_ ( .D(i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_addr_pc4_reg_9_ ( .D(i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_addr_pc4_reg_8_ ( .D(i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_addr_pc4_reg_7_ ( .D(i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_addr_pc4_reg_6_ ( .D(i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_addr_pc4_reg_5_ ( .D(i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_addr_pc4_reg_4_ ( .D(i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_addr_pc4_reg_3_ ( .D(i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_addr_pc4_reg_2_ ( .D(i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_addr_pc4_reg_1_ ( .D(i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_addr_pc4_reg_0_ ( .D(i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  DFC3 pipe_con_Ealuop_reg_5_ ( .D(control_o_con_aluop[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[5]) );
  DFC3 pipe_con_Ealuop_reg_4_ ( .D(control_o_con_aluop[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[4]) );
  DFC3 pipe_con_Ealuop_reg_3_ ( .D(control_o_con_aluop[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[3]) );
  DFC3 pipe_con_Ealuop_reg_2_ ( .D(control_o_con_aluop[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[2]) );
  DFC3 pipe_con_Ealuop_reg_1_ ( .D(control_o_con_aluop[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[1]) );
  DFC3 pipe_con_Ealuop_reg_0_ ( .D(control_o_con_aluop[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[0]) );
  DFC3 pipe_con_Ealusrc_reg ( .D(control_o_con_alusrc), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Ealusrc) );
  DFC3 pipe_con_Eregdst_reg ( .D(control_o_con_regdst), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Eregdst) );
  DFC3 pipe_con_EaluPC4_reg ( .D(jbcon_o_con_aluPC4), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Walupc8) );
  DFC3 pipe_con_Mmemread_reg ( .D(control_o_con_memread), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(control_o_con_memwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wloadmux_reg_1_ ( .D(control_o_con_loadsig[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_con_Wloadmux[1]) );
  DFC3 pipe_con_Wloadmux_reg_0_ ( .D(control_o_con_loadsig[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_con_Wloadmux[0]) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(control_o_con_memtoreg), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(control_o_con_regwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wregwrite) );
  DFC3 pipe_signext_o_data_immD_reg_31_ ( .D(signext_o_data_immD[31]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[31]) );
  DFC3 pipe_signext_o_data_immD_reg_30_ ( .D(signext_o_data_immD[30]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[30]) );
  DFC3 pipe_signext_o_data_immD_reg_29_ ( .D(signext_o_data_immD[29]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[29]) );
  DFC3 pipe_signext_o_data_immD_reg_28_ ( .D(signext_o_data_immD[28]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[28]) );
  DFC3 pipe_signext_o_data_immD_reg_27_ ( .D(signext_o_data_immD[27]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[27]) );
  DFC3 pipe_signext_o_data_immD_reg_26_ ( .D(signext_o_data_immD[26]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[26]) );
  DFC3 pipe_signext_o_data_immD_reg_25_ ( .D(signext_o_data_immD[25]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[25]) );
  DFC3 pipe_signext_o_data_immD_reg_24_ ( .D(signext_o_data_immD[24]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[24]) );
  DFC3 pipe_signext_o_data_immD_reg_23_ ( .D(signext_o_data_immD[23]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[23]) );
  DFC3 pipe_signext_o_data_immD_reg_22_ ( .D(signext_o_data_immD[22]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[22]) );
  DFC3 pipe_signext_o_data_immD_reg_21_ ( .D(signext_o_data_immD[21]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[21]) );
  DFC3 pipe_signext_o_data_immD_reg_20_ ( .D(signext_o_data_immD[20]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[20]) );
  DFC3 pipe_signext_o_data_immD_reg_19_ ( .D(signext_o_data_immD[19]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[19]) );
  DFC3 pipe_signext_o_data_immD_reg_18_ ( .D(signext_o_data_immD[18]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[18]) );
  DFC3 pipe_signext_o_data_immD_reg_17_ ( .D(signext_o_data_immD[17]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[17]) );
  DFC3 pipe_signext_o_data_immD_reg_16_ ( .D(signext_o_data_immD[16]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[16]) );
  DFC3 pipe_signext_o_data_immD_reg_15_ ( .D(signext_o_data_immD[15]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[15]) );
  DFC3 pipe_signext_o_data_immD_reg_14_ ( .D(signext_o_data_immD[14]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[14]) );
  DFC3 pipe_signext_o_data_immD_reg_13_ ( .D(signext_o_data_immD[13]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[13]) );
  DFC3 pipe_signext_o_data_immD_reg_12_ ( .D(signext_o_data_immD[12]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[12]) );
  DFC3 pipe_signext_o_data_immD_reg_11_ ( .D(signext_o_data_immD[11]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[11]) );
  DFC3 pipe_signext_o_data_immD_reg_10_ ( .D(signext_o_data_immD[10]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[10]) );
  DFC3 pipe_signext_o_data_immD_reg_9_ ( .D(signext_o_data_immD[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[9]) );
  DFC3 pipe_signext_o_data_immD_reg_8_ ( .D(signext_o_data_immD[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[8]) );
  DFC3 pipe_signext_o_data_immD_reg_7_ ( .D(signext_o_data_immD[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[7]) );
  DFC3 pipe_signext_o_data_immD_reg_6_ ( .D(signext_o_data_immD[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[6]) );
  DFC3 pipe_signext_o_data_immD_reg_5_ ( .D(signext_o_data_immD[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[5]) );
  DFC3 pipe_signext_o_data_immD_reg_4_ ( .D(signext_o_data_immD[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[4]) );
  DFC3 pipe_signext_o_data_immD_reg_3_ ( .D(signext_o_data_immD[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[3]) );
  DFC3 pipe_signext_o_data_immD_reg_2_ ( .D(signext_o_data_immD[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[2]) );
  DFC3 pipe_signext_o_data_immD_reg_1_ ( .D(signext_o_data_immD[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[1]) );
  DFC3 pipe_signext_o_data_immD_reg_0_ ( .D(signext_o_data_immD[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[0]) );
  DFC3 pipe_con_Efamux_reg_2_ ( .D(for_o_con_fa[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[2]) );
  DFC3 pipe_con_Efamux_reg_1_ ( .D(for_o_con_fa[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[1]) );
  DFC3 pipe_con_Efamux_reg_0_ ( .D(for_o_con_fa[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[0]) );
  DFC3 pipe_con_Efbmux_reg_2_ ( .D(for_o_con_fb[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[2]) );
  DFC3 pipe_con_Efbmux_reg_1_ ( .D(for_o_con_fb[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[1]) );
  DFC3 pipe_con_Efbmux_reg_0_ ( .D(for_o_con_fb[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[0]) );
  DFC3 pipe_memout_reg_31_ ( .D(i_data_Wregwrite[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[31]) );
  DFC3 pipe_memout_reg_30_ ( .D(i_data_Wregwrite[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[30]) );
  DFC3 pipe_memout_reg_29_ ( .D(i_data_Wregwrite[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[29]) );
  DFC3 pipe_memout_reg_28_ ( .D(i_data_Wregwrite[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[28]) );
  DFC3 pipe_memout_reg_27_ ( .D(i_data_Wregwrite[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[27]) );
  DFC3 pipe_memout_reg_26_ ( .D(i_data_Wregwrite[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[26]) );
  DFC3 pipe_memout_reg_25_ ( .D(i_data_Wregwrite[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[25]) );
  DFC3 pipe_memout_reg_24_ ( .D(i_data_Wregwrite[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[24]) );
  DFC3 pipe_memout_reg_23_ ( .D(i_data_Wregwrite[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[23]) );
  DFC3 pipe_memout_reg_22_ ( .D(i_data_Wregwrite[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[22]) );
  DFC3 pipe_memout_reg_20_ ( .D(i_data_Wregwrite[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[20]) );
  DFC3 pipe_memout_reg_19_ ( .D(i_data_Wregwrite[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[19]) );
  DFC3 pipe_memout_reg_18_ ( .D(i_data_Wregwrite[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[18]) );
  DFC3 pipe_memout_reg_16_ ( .D(i_data_Wregwrite[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[16]) );
  DFC3 pipe_memout_reg_15_ ( .D(i_data_Wregwrite[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[15]) );
  DFC3 pipe_memout_reg_14_ ( .D(i_data_Wregwrite[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[14]) );
  DFC3 pipe_memout_reg_13_ ( .D(i_data_Wregwrite[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[13]) );
  DFC3 pipe_memout_reg_12_ ( .D(i_data_Wregwrite[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[12]) );
  DFC3 pipe_memout_reg_11_ ( .D(i_data_Wregwrite[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[11]) );
  DFC3 pipe_memout_reg_10_ ( .D(i_data_Wregwrite[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[10]) );
  DFC3 pipe_memout_reg_8_ ( .D(i_data_Wregwrite[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[8]) );
  DFC3 pipe_memout_reg_4_ ( .D(i_data_Wregwrite[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[4]) );
  DFC3 pipe_memout_reg_3_ ( .D(i_data_Wregwrite[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[3]) );
  DFC3 pipe_memout_reg_0_ ( .D(i_data_Wregwrite[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[0]) );
  DFC3 pipe_addr_branch_reg_31_ ( .D(pcadd_o_addr_pcbranchE[31]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[31]) );
  DFC3 pipe_addr_branch_reg_30_ ( .D(pcadd_o_addr_pcbranchE[30]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[30]) );
  DFC3 pipe_addr_branch_reg_29_ ( .D(pcadd_o_addr_pcbranchE[29]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[29]) );
  DFC3 pipe_addr_branch_reg_28_ ( .D(pcadd_o_addr_pcbranchE[28]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[28]) );
  DFC3 pipe_addr_branch_reg_27_ ( .D(pcadd_o_addr_pcbranchE[27]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[27]) );
  DFC3 pipe_addr_branch_reg_26_ ( .D(pcadd_o_addr_pcbranchE[26]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[26]) );
  DFC3 pipe_addr_branch_reg_25_ ( .D(pcadd_o_addr_pcbranchE[25]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[25]) );
  DFC3 pipe_addr_branch_reg_24_ ( .D(pcadd_o_addr_pcbranchE[24]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[24]) );
  DFC3 pipe_addr_branch_reg_23_ ( .D(pcadd_o_addr_pcbranchE[23]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[23]) );
  DFC3 pipe_addr_branch_reg_22_ ( .D(pcadd_o_addr_pcbranchE[22]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[22]) );
  DFC3 pipe_addr_branch_reg_21_ ( .D(pcadd_o_addr_pcbranchE[21]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[21]) );
  DFC3 pipe_addr_branch_reg_20_ ( .D(pcadd_o_addr_pcbranchE[20]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[20]) );
  DFC3 pipe_addr_branch_reg_19_ ( .D(pcadd_o_addr_pcbranchE[19]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[19]) );
  DFC3 pipe_addr_branch_reg_18_ ( .D(pcadd_o_addr_pcbranchE[18]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[18]) );
  DFC3 pipe_addr_branch_reg_17_ ( .D(pcadd_o_addr_pcbranchE[17]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[17]) );
  DFC3 pipe_addr_branch_reg_16_ ( .D(pcadd_o_addr_pcbranchE[16]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[16]) );
  DFC3 pipe_addr_branch_reg_15_ ( .D(pcadd_o_addr_pcbranchE[15]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[15]) );
  DFC3 pipe_addr_branch_reg_14_ ( .D(pcadd_o_addr_pcbranchE[14]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[14]) );
  DFC3 pipe_addr_branch_reg_13_ ( .D(pcadd_o_addr_pcbranchE[13]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[13]) );
  DFC3 pipe_addr_branch_reg_12_ ( .D(pcadd_o_addr_pcbranchE[12]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[12]) );
  DFC3 pipe_addr_branch_reg_11_ ( .D(pcadd_o_addr_pcbranchE[11]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[11]) );
  DFC3 pipe_addr_branch_reg_10_ ( .D(pcadd_o_addr_pcbranchE[10]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[10]) );
  DFC3 pipe_addr_branch_reg_9_ ( .D(pcadd_o_addr_pcbranchE[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[9]) );
  DFC3 pipe_addr_branch_reg_8_ ( .D(pcadd_o_addr_pcbranchE[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[8]) );
  DFC3 pipe_addr_branch_reg_7_ ( .D(pcadd_o_addr_pcbranchE[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[7]) );
  DFC3 pipe_addr_branch_reg_6_ ( .D(pcadd_o_addr_pcbranchE[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[6]) );
  DFC3 pipe_addr_branch_reg_5_ ( .D(pcadd_o_addr_pcbranchE[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[5]) );
  DFC3 pipe_addr_branch_reg_4_ ( .D(pcadd_o_addr_pcbranchE[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[4]) );
  DFC3 pipe_addr_branch_reg_3_ ( .D(pcadd_o_addr_pcbranchE[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[3]) );
  DFC3 pipe_addr_branch_reg_2_ ( .D(pcadd_o_addr_pcbranchE[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[2]) );
  DFC3 pipe_addr_branch_reg_1_ ( .D(pcadd_o_addr_pcbranchE[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[1]) );
  DFC3 pipe_addr_branch_reg_0_ ( .D(pcadd_o_addr_pcbranchE[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[0]) );
  D_control u_control ( .o_con_regdst(control_o_con_regdst), .o_con_memread(
        control_o_con_memread), .o_con_memtoreg(control_o_con_memtoreg), 
        .o_con_memwrite(control_o_con_memwrite), .o_con_alusrc(
        control_o_con_alusrc), .o_con_regwrite(control_o_con_regwrite), 
        .o_con_ifsign(signext_i_con_signext), .o_con_loadsig(
        control_o_con_loadsig), .o_con_aluop(control_o_con_aluop), 
        .i_con_instru(i_data_instr[31:26]) );
  D_jb_control u_jb_control ( .o_con_jump(o_con_jump), .o_con_bop(
        jbcon_o_con_bop), .o_con_aluPC4(jbcon_o_con_aluPC4), .o_con_ifstall(
        o_con_ifstall), .i_con_instru(i_data_instr[31:26]), .i_con_func(
        i_data_instr[5:0]), .i_con_rt(i_data_instr[16]) );
  D_pcadd u_pcadd ( .i_addr_pcadd4E(i_addr_pc4), .i_data_immshiftl({
        pcadd_i_data_immshiftl, o_addr_jump[0], o_addr_jump[0]}), 
        .o_addr_pcbranchE(pcadd_o_addr_pcbranchE) );
  D_register_bank u_regbank ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_addr_Rs(
        i_data_instr[25:21]), .i_addr_Rt(i_data_instr[20:16]), .i_con_RegWr(
        i_con_Wregwrite), .i_addr_Rd(i_addr_Wregwrite), .i_data_Rd(
        i_data_Wregwrite), .o_data_Rs(o_data_jr), .o_data_Rt(regbank_o_data_Rt) );
  D_shiftleft u_sl ( .i_data_immE(i_data_instr[15:0]), .o_data_immshiftl({
        pcadd_i_data_immshiftl, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}) );
  D_sign_extend u_signext ( .i_data_immD(i_data_instr[15:0]), .i_con_signext(
        signext_i_con_signext), .o_data_immD(signext_o_data_immD) );
  D_jump_ext u_jump_ext ( .i_addr_j(i_data_instr[25:0]), .i_PC4_j(
        i_addr_pc4[31:28]), .o_addr_j({o_addr_jump[31:2], 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4}) );
  E_forward u_forward ( .i_addr_rs(i_data_instr[25:21]), .i_addr_rt(
        i_data_instr[20:16]), .i_addr_rdM(i_addr_Erd), .i_addr_rdW(i_addr_Mrd), 
        .i_addr_rtM(i_addr_rtM), .i_addr_rtW(i_addr_rtW), .i_con_regwriteM(
        i_con_Eregwrite), .i_con_regwriteW(i_con_Mregwrite), .i_con_memreadM(
        i_con_memreadM), .i_con_memreadW(i_con_memreadW), .o_con_fa(
        for_o_con_fa), .o_con_fb(for_o_con_fb) );
  DFC1 pipe_memout_reg_21_ ( .D(i_data_Wregwrite[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[21]) );
  DFC1 pipe_memout_reg_6_ ( .D(i_data_Wregwrite[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[6]) );
  DFC1 pipe_memout_reg_5_ ( .D(i_data_Wregwrite[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[5]) );
  DFC1 pipe_memout_reg_2_ ( .D(i_data_Wregwrite[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[2]) );
  DFC1 pipe_memout_reg_7_ ( .D(i_data_Wregwrite[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[7]) );
  DFC1 pipe_memout_reg_9_ ( .D(i_data_Wregwrite[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[9]) );
  DFC1 pipe_memout_reg_1_ ( .D(i_data_Wregwrite[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[1]) );
  DFC1 pipe_memout_reg_17_ ( .D(i_data_Wregwrite[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[17]) );
  LOGIC0 U3 ( .Q(o_addr_jump[0]) );
endmodule


module E_alu_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   ML_int_1__31_, ML_int_1__30_, ML_int_1__29_, ML_int_1__28_,
         ML_int_1__27_, ML_int_1__26_, ML_int_1__25_, ML_int_1__24_,
         ML_int_1__23_, ML_int_1__22_, ML_int_1__21_, ML_int_1__20_,
         ML_int_1__19_, ML_int_1__18_, ML_int_1__17_, ML_int_1__16_,
         ML_int_1__15_, ML_int_1__14_, ML_int_1__13_, ML_int_1__12_,
         ML_int_1__11_, ML_int_1__10_, ML_int_1__9_, ML_int_1__8_,
         ML_int_1__7_, ML_int_1__6_, ML_int_1__5_, ML_int_1__4_, ML_int_1__3_,
         ML_int_1__2_, ML_int_1__1_, ML_int_1__0_, ML_int_2__31_,
         ML_int_2__30_, ML_int_2__29_, ML_int_2__28_, ML_int_2__27_,
         ML_int_2__26_, ML_int_2__25_, ML_int_2__24_, ML_int_2__23_,
         ML_int_2__22_, ML_int_2__21_, ML_int_2__20_, ML_int_2__19_,
         ML_int_2__18_, ML_int_2__17_, ML_int_2__16_, ML_int_2__15_,
         ML_int_2__14_, ML_int_2__13_, ML_int_2__12_, ML_int_2__11_,
         ML_int_2__10_, ML_int_2__9_, ML_int_2__8_, ML_int_2__7_, ML_int_2__6_,
         ML_int_2__5_, ML_int_2__4_, ML_int_2__3_, ML_int_2__2_, ML_int_3__31_,
         ML_int_3__30_, ML_int_3__29_, ML_int_3__28_, ML_int_3__27_,
         ML_int_3__26_, ML_int_3__25_, ML_int_3__24_, ML_int_3__23_,
         ML_int_3__22_, ML_int_3__21_, ML_int_3__20_, ML_int_3__19_,
         ML_int_3__18_, ML_int_3__17_, ML_int_3__16_, ML_int_3__15_,
         ML_int_3__14_, ML_int_3__13_, ML_int_3__12_, ML_int_3__11_,
         ML_int_3__10_, ML_int_3__9_, ML_int_3__8_, ML_int_3__7_, ML_int_3__6_,
         ML_int_3__5_, ML_int_3__4_, ML_int_3__1_, ML_int_3__0_, ML_int_4__31_,
         ML_int_4__30_, ML_int_4__29_, ML_int_4__28_, ML_int_4__27_,
         ML_int_4__26_, ML_int_4__25_, ML_int_4__24_, ML_int_4__15_,
         ML_int_4__14_, ML_int_4__13_, ML_int_4__12_, ML_int_4__11_,
         ML_int_4__10_, ML_int_4__9_, ML_int_4__8_, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36;

  MUX21 U3 ( .A(A[12]), .B(A[11]), .S(SH[0]), .Q(ML_int_1__12_) );
  MUX21 U4 ( .A(A[6]), .B(A[5]), .S(SH[0]), .Q(ML_int_1__6_) );
  MUX21 U5 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Q(ML_int_1__2_) );
  MUX21 U6 ( .A(A[11]), .B(A[10]), .S(SH[0]), .Q(ML_int_1__11_) );
  MUX21 U7 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Q(ML_int_1__8_) );
  MUX21 U8 ( .A(A[9]), .B(A[8]), .S(SH[0]), .Q(ML_int_1__9_) );
  MUX21 U9 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Q(ML_int_1__10_) );
  MUX21 U10 ( .A(A[4]), .B(A[3]), .S(SH[0]), .Q(ML_int_1__4_) );
  MUX21 U11 ( .A(A[3]), .B(A[2]), .S(SH[0]), .Q(ML_int_1__3_) );
  MUX21 U12 ( .A(A[5]), .B(A[4]), .S(SH[0]), .Q(ML_int_1__5_) );
  MUX21 U13 ( .A(A[20]), .B(A[19]), .S(SH[0]), .Q(ML_int_1__20_) );
  MUX21 U14 ( .A(A[21]), .B(A[20]), .S(SH[0]), .Q(ML_int_1__21_) );
  MUX21 U15 ( .A(A[22]), .B(A[21]), .S(SH[0]), .Q(ML_int_1__22_) );
  MUX21 U16 ( .A(A[18]), .B(A[17]), .S(SH[0]), .Q(ML_int_1__18_) );
  MUX21 U17 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Q(ML_int_1__1_) );
  INV0 U18 ( .A(A[0]), .Q(n24) );
  MUX22 U19 ( .A(ML_int_3__8_), .B(ML_int_3__0_), .S(SH[3]), .Q(ML_int_4__8_)
         );
  MUX22 U20 ( .A(ML_int_3__9_), .B(ML_int_3__1_), .S(SH[3]), .Q(ML_int_4__9_)
         );
  MUX22 U21 ( .A(ML_int_1__8_), .B(ML_int_1__6_), .S(SH[1]), .Q(ML_int_2__8_)
         );
  MUX22 U22 ( .A(ML_int_1__10_), .B(ML_int_1__8_), .S(SH[1]), .Q(ML_int_2__10_) );
  MUX22 U23 ( .A(ML_int_1__9_), .B(ML_int_1__7_), .S(SH[1]), .Q(ML_int_2__9_)
         );
  MUX22 U24 ( .A(ML_int_1__7_), .B(ML_int_1__5_), .S(SH[1]), .Q(ML_int_2__7_)
         );
  MUX22 U25 ( .A(ML_int_1__4_), .B(ML_int_1__2_), .S(SH[1]), .Q(ML_int_2__4_)
         );
  MUX22 U26 ( .A(ML_int_1__6_), .B(ML_int_1__4_), .S(SH[1]), .Q(ML_int_2__6_)
         );
  MUX22 U27 ( .A(ML_int_1__5_), .B(ML_int_1__3_), .S(SH[1]), .Q(ML_int_2__5_)
         );
  MUX22 U28 ( .A(ML_int_2__8_), .B(ML_int_2__4_), .S(SH[2]), .Q(ML_int_3__8_)
         );
  MUX22 U29 ( .A(ML_int_2__9_), .B(ML_int_2__5_), .S(SH[2]), .Q(ML_int_3__9_)
         );
  MUX22 U30 ( .A(ML_int_2__10_), .B(ML_int_2__6_), .S(SH[2]), .Q(ML_int_3__10_) );
  MUX22 U31 ( .A(ML_int_2__11_), .B(ML_int_2__7_), .S(SH[2]), .Q(ML_int_3__11_) );
  MUX22 U32 ( .A(ML_int_2__12_), .B(ML_int_2__8_), .S(SH[2]), .Q(ML_int_3__12_) );
  MUX22 U33 ( .A(ML_int_2__13_), .B(ML_int_2__9_), .S(SH[2]), .Q(ML_int_3__13_) );
  MUX22 U34 ( .A(ML_int_2__14_), .B(ML_int_2__10_), .S(SH[2]), .Q(
        ML_int_3__14_) );
  MUX22 U35 ( .A(ML_int_3__10_), .B(n21), .S(SH[3]), .Q(ML_int_4__10_) );
  MUX22 U36 ( .A(ML_int_3__11_), .B(n20), .S(SH[3]), .Q(ML_int_4__11_) );
  MUX22 U37 ( .A(ML_int_3__12_), .B(ML_int_3__4_), .S(SH[3]), .Q(ML_int_4__12_) );
  MUX22 U38 ( .A(ML_int_3__13_), .B(ML_int_3__5_), .S(SH[3]), .Q(ML_int_4__13_) );
  MUX22 U39 ( .A(ML_int_3__14_), .B(ML_int_3__6_), .S(SH[3]), .Q(ML_int_4__14_) );
  MUX22 U40 ( .A(ML_int_1__2_), .B(ML_int_1__0_), .S(SH[1]), .Q(ML_int_2__2_)
         );
  MUX22 U41 ( .A(ML_int_1__3_), .B(ML_int_1__1_), .S(SH[1]), .Q(ML_int_2__3_)
         );
  MUX22 U42 ( .A(ML_int_2__4_), .B(n23), .S(SH[2]), .Q(ML_int_3__4_) );
  INV3 U43 ( .A(n36), .Q(n23) );
  MUX22 U44 ( .A(ML_int_2__5_), .B(n22), .S(SH[2]), .Q(ML_int_3__5_) );
  INV3 U45 ( .A(n35), .Q(n22) );
  MUX22 U46 ( .A(ML_int_2__7_), .B(ML_int_2__3_), .S(SH[2]), .Q(ML_int_3__7_)
         );
  MUX22 U47 ( .A(ML_int_2__6_), .B(ML_int_2__2_), .S(SH[2]), .Q(ML_int_3__6_)
         );
  MUX22 U48 ( .A(ML_int_1__16_), .B(ML_int_1__14_), .S(SH[1]), .Q(
        ML_int_2__16_) );
  MUX22 U49 ( .A(ML_int_1__17_), .B(ML_int_1__15_), .S(SH[1]), .Q(
        ML_int_2__17_) );
  MUX22 U50 ( .A(ML_int_1__18_), .B(ML_int_1__16_), .S(SH[1]), .Q(
        ML_int_2__18_) );
  MUX22 U51 ( .A(ML_int_1__11_), .B(ML_int_1__9_), .S(SH[1]), .Q(ML_int_2__11_) );
  MUX22 U52 ( .A(ML_int_2__16_), .B(ML_int_2__12_), .S(SH[2]), .Q(
        ML_int_3__16_) );
  MUX22 U53 ( .A(ML_int_2__17_), .B(ML_int_2__13_), .S(SH[2]), .Q(
        ML_int_3__17_) );
  MUX22 U54 ( .A(ML_int_1__12_), .B(ML_int_1__10_), .S(SH[1]), .Q(
        ML_int_2__12_) );
  MUX22 U55 ( .A(ML_int_1__13_), .B(ML_int_1__11_), .S(SH[1]), .Q(
        ML_int_2__13_) );
  MUX22 U56 ( .A(ML_int_1__14_), .B(ML_int_1__12_), .S(SH[1]), .Q(
        ML_int_2__14_) );
  MUX22 U57 ( .A(ML_int_2__18_), .B(ML_int_2__14_), .S(SH[2]), .Q(
        ML_int_3__18_) );
  MUX22 U58 ( .A(ML_int_2__19_), .B(ML_int_2__15_), .S(SH[2]), .Q(
        ML_int_3__19_) );
  MUX22 U59 ( .A(ML_int_1__15_), .B(ML_int_1__13_), .S(SH[1]), .Q(
        ML_int_2__15_) );
  MUX22 U60 ( .A(ML_int_2__15_), .B(ML_int_2__11_), .S(SH[2]), .Q(
        ML_int_3__15_) );
  MUX22 U61 ( .A(ML_int_2__20_), .B(ML_int_2__16_), .S(SH[2]), .Q(
        ML_int_3__20_) );
  MUX22 U62 ( .A(ML_int_2__21_), .B(ML_int_2__17_), .S(SH[2]), .Q(
        ML_int_3__21_) );
  MUX22 U63 ( .A(ML_int_2__22_), .B(ML_int_2__18_), .S(SH[2]), .Q(
        ML_int_3__22_) );
  MUX22 U64 ( .A(ML_int_3__15_), .B(ML_int_3__7_), .S(SH[3]), .Q(ML_int_4__15_) );
  MUX22 U65 ( .A(ML_int_1__19_), .B(ML_int_1__17_), .S(SH[1]), .Q(
        ML_int_2__19_) );
  MUX22 U66 ( .A(ML_int_1__24_), .B(ML_int_1__22_), .S(SH[1]), .Q(
        ML_int_2__24_) );
  MUX22 U67 ( .A(ML_int_1__20_), .B(ML_int_1__18_), .S(SH[1]), .Q(
        ML_int_2__20_) );
  MUX22 U68 ( .A(ML_int_1__21_), .B(ML_int_1__19_), .S(SH[1]), .Q(
        ML_int_2__21_) );
  MUX22 U69 ( .A(ML_int_1__25_), .B(ML_int_1__23_), .S(SH[1]), .Q(
        ML_int_2__25_) );
  MUX22 U70 ( .A(ML_int_1__22_), .B(ML_int_1__20_), .S(SH[1]), .Q(
        ML_int_2__22_) );
  MUX22 U71 ( .A(ML_int_1__26_), .B(ML_int_1__24_), .S(SH[1]), .Q(
        ML_int_2__26_) );
  MUX22 U72 ( .A(ML_int_1__23_), .B(ML_int_1__21_), .S(SH[1]), .Q(
        ML_int_2__23_) );
  MUX22 U73 ( .A(ML_int_1__27_), .B(ML_int_1__25_), .S(SH[1]), .Q(
        ML_int_2__27_) );
  MUX22 U74 ( .A(ML_int_2__23_), .B(ML_int_2__19_), .S(SH[2]), .Q(
        ML_int_3__23_) );
  MUX22 U75 ( .A(ML_int_4__30_), .B(ML_int_4__14_), .S(SH[4]), .Q(B[30]) );
  INV3 U76 ( .A(ML_int_4__8_), .Q(n19) );
  INV3 U77 ( .A(ML_int_4__10_), .Q(n17) );
  INV3 U78 ( .A(ML_int_4__11_), .Q(n16) );
  INV3 U79 ( .A(ML_int_4__12_), .Q(n15) );
  INV3 U80 ( .A(ML_int_4__13_), .Q(n14) );
  INV3 U81 ( .A(ML_int_4__14_), .Q(n13) );
  INV3 U82 ( .A(n34), .Q(n21) );
  INV3 U83 ( .A(n33), .Q(n20) );
  MUX22 U84 ( .A(A[7]), .B(A[6]), .S(SH[0]), .Q(ML_int_1__7_) );
  IMUX21 U85 ( .A(n1), .B(n32), .S(SH[4]), .Q(B[16]) );
  IMUX21 U86 ( .A(ML_int_3__16_), .B(ML_int_3__8_), .S(SH[3]), .Q(n1) );
  IMUX21 U87 ( .A(n2), .B(n31), .S(SH[4]), .Q(B[17]) );
  IMUX21 U88 ( .A(ML_int_3__17_), .B(ML_int_3__9_), .S(SH[3]), .Q(n2) );
  MUX22 U89 ( .A(ML_int_4__24_), .B(ML_int_4__8_), .S(SH[4]), .Q(B[24]) );
  MUX22 U90 ( .A(ML_int_3__24_), .B(ML_int_3__16_), .S(SH[3]), .Q(
        ML_int_4__24_) );
  MUX22 U91 ( .A(ML_int_2__24_), .B(ML_int_2__20_), .S(SH[2]), .Q(
        ML_int_3__24_) );
  MUX22 U92 ( .A(ML_int_4__25_), .B(ML_int_4__9_), .S(SH[4]), .Q(B[25]) );
  MUX22 U93 ( .A(ML_int_3__25_), .B(ML_int_3__17_), .S(SH[3]), .Q(
        ML_int_4__25_) );
  MUX22 U94 ( .A(ML_int_2__25_), .B(ML_int_2__21_), .S(SH[2]), .Q(
        ML_int_3__25_) );
  IMUX21 U95 ( .A(n3), .B(n30), .S(SH[4]), .Q(B[18]) );
  IMUX21 U96 ( .A(ML_int_3__18_), .B(ML_int_3__10_), .S(SH[3]), .Q(n3) );
  IMUX21 U97 ( .A(n4), .B(n29), .S(SH[4]), .Q(B[19]) );
  IMUX21 U98 ( .A(ML_int_3__19_), .B(ML_int_3__11_), .S(SH[3]), .Q(n4) );
  IMUX21 U99 ( .A(n5), .B(n28), .S(SH[4]), .Q(B[20]) );
  IMUX21 U100 ( .A(ML_int_3__20_), .B(ML_int_3__12_), .S(SH[3]), .Q(n5) );
  IMUX21 U101 ( .A(n6), .B(n27), .S(SH[4]), .Q(B[21]) );
  IMUX21 U102 ( .A(ML_int_3__21_), .B(ML_int_3__13_), .S(SH[3]), .Q(n6) );
  IMUX21 U103 ( .A(n7), .B(n26), .S(SH[4]), .Q(B[22]) );
  IMUX21 U104 ( .A(ML_int_3__22_), .B(ML_int_3__14_), .S(SH[3]), .Q(n7) );
  MUX22 U105 ( .A(ML_int_4__26_), .B(ML_int_4__10_), .S(SH[4]), .Q(B[26]) );
  MUX22 U106 ( .A(ML_int_3__26_), .B(ML_int_3__18_), .S(SH[3]), .Q(
        ML_int_4__26_) );
  MUX22 U107 ( .A(ML_int_2__26_), .B(ML_int_2__22_), .S(SH[2]), .Q(
        ML_int_3__26_) );
  MUX22 U108 ( .A(ML_int_4__28_), .B(ML_int_4__12_), .S(SH[4]), .Q(B[28]) );
  MUX22 U109 ( .A(ML_int_3__28_), .B(ML_int_3__20_), .S(SH[3]), .Q(
        ML_int_4__28_) );
  MUX22 U110 ( .A(ML_int_2__28_), .B(ML_int_2__24_), .S(SH[2]), .Q(
        ML_int_3__28_) );
  MUX22 U111 ( .A(ML_int_1__28_), .B(ML_int_1__26_), .S(SH[1]), .Q(
        ML_int_2__28_) );
  INV3 U112 ( .A(ML_int_4__9_), .Q(n18) );
  INV3 U113 ( .A(ML_int_4__15_), .Q(n12) );
  MUX22 U114 ( .A(A[14]), .B(A[13]), .S(SH[0]), .Q(ML_int_1__14_) );
  MUX22 U115 ( .A(A[13]), .B(A[12]), .S(SH[0]), .Q(ML_int_1__13_) );
  MUX22 U116 ( .A(A[15]), .B(A[14]), .S(SH[0]), .Q(ML_int_1__15_) );
  MUX22 U117 ( .A(ML_int_3__30_), .B(ML_int_3__22_), .S(SH[3]), .Q(
        ML_int_4__30_) );
  MUX22 U118 ( .A(ML_int_2__30_), .B(ML_int_2__26_), .S(SH[2]), .Q(
        ML_int_3__30_) );
  MUX22 U119 ( .A(ML_int_1__30_), .B(ML_int_1__28_), .S(SH[1]), .Q(
        ML_int_2__30_) );
  MUX22 U120 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Q(ML_int_1__30_) );
  IMUX21 U121 ( .A(n8), .B(n25), .S(SH[4]), .Q(B[23]) );
  IMUX21 U122 ( .A(ML_int_3__23_), .B(ML_int_3__15_), .S(SH[3]), .Q(n8) );
  MUX22 U123 ( .A(ML_int_4__27_), .B(ML_int_4__11_), .S(SH[4]), .Q(B[27]) );
  MUX22 U124 ( .A(ML_int_3__27_), .B(ML_int_3__19_), .S(SH[3]), .Q(
        ML_int_4__27_) );
  MUX22 U125 ( .A(ML_int_2__27_), .B(ML_int_2__23_), .S(SH[2]), .Q(
        ML_int_3__27_) );
  MUX22 U126 ( .A(ML_int_4__29_), .B(ML_int_4__13_), .S(SH[4]), .Q(B[29]) );
  MUX22 U127 ( .A(ML_int_3__29_), .B(ML_int_3__21_), .S(SH[3]), .Q(
        ML_int_4__29_) );
  MUX22 U128 ( .A(ML_int_2__29_), .B(ML_int_2__25_), .S(SH[2]), .Q(
        ML_int_3__29_) );
  MUX22 U129 ( .A(ML_int_1__29_), .B(ML_int_1__27_), .S(SH[1]), .Q(
        ML_int_2__29_) );
  MUX22 U130 ( .A(ML_int_4__31_), .B(ML_int_4__15_), .S(SH[4]), .Q(B[31]) );
  MUX22 U131 ( .A(ML_int_3__31_), .B(ML_int_3__23_), .S(SH[3]), .Q(
        ML_int_4__31_) );
  MUX22 U132 ( .A(ML_int_2__31_), .B(ML_int_2__27_), .S(SH[2]), .Q(
        ML_int_3__31_) );
  MUX22 U133 ( .A(ML_int_1__31_), .B(ML_int_1__29_), .S(SH[1]), .Q(
        ML_int_2__31_) );
  MUX22 U134 ( .A(A[24]), .B(A[23]), .S(SH[0]), .Q(ML_int_1__24_) );
  MUX22 U135 ( .A(A[19]), .B(A[18]), .S(SH[0]), .Q(ML_int_1__19_) );
  MUX22 U136 ( .A(A[25]), .B(A[24]), .S(SH[0]), .Q(ML_int_1__25_) );
  MUX22 U137 ( .A(A[29]), .B(A[28]), .S(SH[0]), .Q(ML_int_1__29_) );
  MUX22 U138 ( .A(A[26]), .B(A[25]), .S(SH[0]), .Q(ML_int_1__26_) );
  MUX22 U139 ( .A(A[28]), .B(A[27]), .S(SH[0]), .Q(ML_int_1__28_) );
  MUX22 U140 ( .A(A[23]), .B(A[22]), .S(SH[0]), .Q(ML_int_1__23_) );
  MUX22 U141 ( .A(A[27]), .B(A[26]), .S(SH[0]), .Q(ML_int_1__27_) );
  MUX22 U142 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Q(ML_int_1__31_) );
  INV3 U143 ( .A(SH[2]), .Q(n10) );
  INV3 U144 ( .A(SH[1]), .Q(n9) );
  INV3 U145 ( .A(SH[3]), .Q(n11) );
  MUX21 U146 ( .A(A[16]), .B(A[15]), .S(SH[0]), .Q(ML_int_1__16_) );
  MUX21 U147 ( .A(A[17]), .B(A[16]), .S(SH[0]), .Q(ML_int_1__17_) );
  NOR20 U148 ( .A(SH[4]), .B(n18), .Q(B[9]) );
  NOR20 U149 ( .A(SH[4]), .B(n19), .Q(B[8]) );
  NOR20 U150 ( .A(SH[4]), .B(n25), .Q(B[7]) );
  NOR20 U151 ( .A(SH[4]), .B(n26), .Q(B[6]) );
  NOR20 U152 ( .A(SH[4]), .B(n27), .Q(B[5]) );
  NOR20 U153 ( .A(SH[4]), .B(n28), .Q(B[4]) );
  NOR20 U154 ( .A(SH[4]), .B(n29), .Q(B[3]) );
  NOR20 U155 ( .A(SH[4]), .B(n30), .Q(B[2]) );
  NOR20 U156 ( .A(SH[4]), .B(n31), .Q(B[1]) );
  NOR20 U157 ( .A(SH[4]), .B(n12), .Q(B[15]) );
  NOR20 U158 ( .A(SH[4]), .B(n13), .Q(B[14]) );
  NOR20 U159 ( .A(SH[4]), .B(n14), .Q(B[13]) );
  NOR20 U160 ( .A(SH[4]), .B(n15), .Q(B[12]) );
  NOR20 U161 ( .A(SH[4]), .B(n16), .Q(B[11]) );
  NOR20 U162 ( .A(SH[4]), .B(n17), .Q(B[10]) );
  NOR20 U163 ( .A(SH[4]), .B(n32), .Q(B[0]) );
  NAND20 U164 ( .A(ML_int_3__7_), .B(n11), .Q(n25) );
  NAND20 U165 ( .A(ML_int_3__6_), .B(n11), .Q(n26) );
  NAND20 U166 ( .A(ML_int_3__5_), .B(n11), .Q(n27) );
  NAND20 U167 ( .A(ML_int_3__4_), .B(n11), .Q(n28) );
  NAND20 U168 ( .A(n20), .B(n11), .Q(n29) );
  NAND20 U169 ( .A(n21), .B(n11), .Q(n30) );
  NAND20 U170 ( .A(ML_int_3__1_), .B(n11), .Q(n31) );
  NAND20 U171 ( .A(ML_int_3__0_), .B(n11), .Q(n32) );
  NAND20 U172 ( .A(ML_int_2__3_), .B(n10), .Q(n33) );
  NAND20 U173 ( .A(ML_int_2__2_), .B(n10), .Q(n34) );
  NOR20 U174 ( .A(n35), .B(SH[2]), .Q(ML_int_3__1_) );
  NOR20 U175 ( .A(n36), .B(SH[2]), .Q(ML_int_3__0_) );
  NAND20 U176 ( .A(ML_int_1__1_), .B(n9), .Q(n35) );
  NAND20 U177 ( .A(ML_int_1__0_), .B(n9), .Q(n36) );
  NOR20 U178 ( .A(n24), .B(SH[0]), .Q(ML_int_1__0_) );
endmodule


module E_alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [15:1] carry;

  ADD32 U2_14 ( .A(A[14]), .B(n12), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADD32 U2_12 ( .A(A[12]), .B(n14), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADD32 U2_11 ( .A(A[11]), .B(n15), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADD32 U2_10 ( .A(A[10]), .B(n16), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADD32 U2_9 ( .A(A[9]), .B(n17), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADD32 U2_7 ( .A(A[7]), .B(n19), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADD32 U2_6 ( .A(A[6]), .B(n20), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADD32 U2_5 ( .A(A[5]), .B(n21), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADD32 U2_3 ( .A(A[3]), .B(n23), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADD32 U2_2 ( .A(A[2]), .B(n24), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADD32 U2_1 ( .A(A[1]), .B(n25), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NAND22 U1 ( .A(carry[4]), .B(A[4]), .Q(n1) );
  NAND22 U2 ( .A(carry[4]), .B(n22), .Q(n2) );
  NAND22 U3 ( .A(carry[8]), .B(n18), .Q(n5) );
  NAND22 U4 ( .A(carry[8]), .B(A[8]), .Q(n4) );
  NAND33 U5 ( .A(n8), .B(n9), .C(n10), .Q(carry[14]) );
  NAND22 U6 ( .A(A[13]), .B(n13), .Q(n10) );
  INV3 U7 ( .A(B[8]), .Q(n18) );
  INV3 U8 ( .A(B[0]), .Q(n26) );
  NAND33 U9 ( .A(n1), .B(n2), .C(n3), .Q(carry[5]) );
  NAND22 U10 ( .A(A[4]), .B(n22), .Q(n3) );
  NAND22 U11 ( .A(carry[13]), .B(A[13]), .Q(n8) );
  NAND22 U12 ( .A(carry[13]), .B(n13), .Q(n9) );
  NAND33 U13 ( .A(n4), .B(n5), .C(n6), .Q(carry[9]) );
  INV3 U14 ( .A(B[13]), .Q(n13) );
  NAND20 U15 ( .A(A[8]), .B(n18), .Q(n6) );
  INV2 U16 ( .A(B[4]), .Q(n22) );
  XOR30 U17 ( .A(carry[4]), .B(A[4]), .C(n22), .Q(DIFF[4]) );
  XOR30 U18 ( .A(carry[8]), .B(A[8]), .C(n18), .Q(DIFF[8]) );
  XOR20 U19 ( .A(A[13]), .B(n13), .Q(n7) );
  XOR21 U20 ( .A(carry[13]), .B(n7), .Q(DIFF[13]) );
  XOR20 U21 ( .A(A[0]), .B(n26), .Q(DIFF[0]) );
  INV3 U22 ( .A(B[10]), .Q(n16) );
  INV3 U23 ( .A(B[11]), .Q(n15) );
  INV3 U24 ( .A(B[12]), .Q(n14) );
  INV3 U25 ( .A(B[5]), .Q(n21) );
  INV3 U26 ( .A(B[9]), .Q(n17) );
  INV3 U27 ( .A(B[2]), .Q(n24) );
  INV3 U28 ( .A(B[3]), .Q(n23) );
  INV3 U29 ( .A(B[6]), .Q(n20) );
  INV3 U30 ( .A(B[7]), .Q(n19) );
  INV3 U31 ( .A(B[14]), .Q(n12) );
  XNR31 U32 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Q(DIFF[15]) );
  INV3 U33 ( .A(n11), .Q(carry[1]) );
  INV3 U34 ( .A(B[1]), .Q(n25) );
  NAND22 U35 ( .A(A[0]), .B(n26), .Q(n11) );
endmodule


module E_alu_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  wire   [15:1] carry;

  ADD32 U2_14 ( .A(A[14]), .B(n4), .CI(carry[14]), .CO(carry[15]), .S(DIFF[14]) );
  ADD32 U2_13 ( .A(A[13]), .B(n5), .CI(carry[13]), .CO(carry[14]), .S(DIFF[13]) );
  ADD32 U2_12 ( .A(A[12]), .B(n6), .CI(carry[12]), .CO(carry[13]), .S(DIFF[12]) );
  ADD32 U2_11 ( .A(A[11]), .B(n7), .CI(carry[11]), .CO(carry[12]), .S(DIFF[11]) );
  ADD32 U2_10 ( .A(A[10]), .B(n8), .CI(carry[10]), .CO(carry[11]), .S(DIFF[10]) );
  ADD32 U2_9 ( .A(A[9]), .B(n9), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9]) );
  ADD32 U2_8 ( .A(A[8]), .B(n10), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADD32 U2_7 ( .A(A[7]), .B(n11), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADD32 U2_6 ( .A(A[6]), .B(n12), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADD32 U2_5 ( .A(A[5]), .B(n13), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADD32 U2_4 ( .A(A[4]), .B(n14), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADD32 U2_3 ( .A(A[3]), .B(n15), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADD32 U2_2 ( .A(A[2]), .B(n16), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADD32 U2_1 ( .A(A[1]), .B(n17), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  NOR21 U1 ( .A(n18), .B(A[0]), .Q(n1) );
  INV3 U2 ( .A(B[4]), .Q(n14) );
  XNR20 U3 ( .A(A[0]), .B(n18), .Q(DIFF[0]) );
  INV3 U4 ( .A(A[15]), .Q(n2) );
  INV3 U5 ( .A(B[8]), .Q(n10) );
  INV3 U6 ( .A(B[9]), .Q(n9) );
  INV3 U7 ( .A(B[10]), .Q(n8) );
  INV3 U8 ( .A(B[11]), .Q(n7) );
  INV3 U9 ( .A(B[12]), .Q(n6) );
  INV3 U10 ( .A(B[13]), .Q(n5) );
  INV3 U11 ( .A(B[5]), .Q(n13) );
  INV3 U12 ( .A(B[2]), .Q(n16) );
  INV3 U13 ( .A(B[3]), .Q(n15) );
  INV3 U14 ( .A(B[6]), .Q(n12) );
  INV3 U15 ( .A(B[7]), .Q(n11) );
  INV3 U16 ( .A(B[14]), .Q(n4) );
  INV3 U17 ( .A(n1), .Q(carry[1]) );
  INV3 U18 ( .A(B[1]), .Q(n17) );
  INV3 U19 ( .A(B[0]), .Q(n18) );
  INV3 U20 ( .A(B[15]), .Q(n3) );
  XNR31 U21 ( .A(n2), .B(n3), .C(carry[15]), .Q(DIFF[15]) );
endmodule


module E_alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR31 U1 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Q(SUM[7]) );
  INV3 U2 ( .A(n1), .Q(carry[1]) );
  NOR21 U3 ( .A(B[0]), .B(A[0]), .Q(n1) );
  XNR21 U4 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
endmodule


module E_alu_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR21 U1 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  XOR31 U2 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Q(SUM[7]) );
  INV3 U3 ( .A(n1), .Q(carry[1]) );
  NAND22 U4 ( .A(A[0]), .B(B[0]), .Q(n1) );
endmodule


module E_alu_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  ADD31 U1 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  NOR20 U2 ( .A(B[0]), .B(A[0]), .Q(n1) );
  CLKIN3 U3 ( .A(n1), .Q(carry[1]) );
  XNR20 U4 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
endmodule


module E_alu_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  ADD31 U1 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  XOR20 U2 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  NAND20 U3 ( .A(A[0]), .B(B[0]), .Q(n1) );
  ADD31 U4 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV3 U5 ( .A(n1), .Q(carry[1]) );
endmodule


module E_alu_DW01_add_4 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  XNR20 U1 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  CLKIN3 U2 ( .A(n1), .Q(carry[1]) );
  NOR21 U3 ( .A(B[0]), .B(A[0]), .Q(n1) );
endmodule


module E_alu_DW01_add_5 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKIN3 U1 ( .A(n1), .Q(carry[1]) );
  NAND20 U2 ( .A(A[0]), .B(B[0]), .Q(n1) );
  XOR20 U3 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
endmodule


module E_alu_DW01_add_6 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND22 U1 ( .A(A[0]), .B(B[0]), .Q(n1) );
  CLKIN3 U2 ( .A(n1), .Q(carry[1]) );
  XOR20 U3 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
endmodule


module E_alu_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211;

  INV3 U3 ( .A(n126), .Q(n29) );
  INV3 U4 ( .A(n103), .Q(n24) );
  INV3 U5 ( .A(n113), .Q(n15) );
  INV3 U6 ( .A(n138), .Q(n34) );
  INV3 U7 ( .A(n116), .Q(n32) );
  INV3 U8 ( .A(n142), .Q(n31) );
  INV3 U9 ( .A(n164), .Q(n33) );
  INV3 U10 ( .A(n70), .Q(n37) );
  INV3 U11 ( .A(n102), .Q(n21) );
  INV3 U12 ( .A(n91), .Q(n46) );
  INV3 U13 ( .A(n92), .Q(n19) );
  INV3 U14 ( .A(n69), .Q(n20) );
  INV3 U15 ( .A(n63), .Q(n28) );
  INV3 U16 ( .A(n129), .Q(n13) );
  INV3 U17 ( .A(n106), .Q(n23) );
  INV3 U18 ( .A(A[18]), .Q(n38) );
  INV3 U19 ( .A(A[19]), .Q(n36) );
  INV3 U20 ( .A(n78), .Q(n35) );
  INV3 U21 ( .A(n159), .Q(n17) );
  INV3 U22 ( .A(n145), .Q(n26) );
  INV3 U23 ( .A(n110), .Q(n43) );
  INV3 U24 ( .A(n87), .Q(n27) );
  INV3 U25 ( .A(n82), .Q(n16) );
  INV3 U26 ( .A(n118), .Q(n49) );
  INV3 U27 ( .A(n88), .Q(n41) );
  INV3 U28 ( .A(n83), .Q(n40) );
  INV3 U29 ( .A(n77), .Q(n39) );
  BUF2 U30 ( .A(n95), .Q(n2) );
  INV3 U31 ( .A(n58), .Q(n47) );
  NOR21 U32 ( .A(n49), .B(n11), .Q(n91) );
  INV3 U33 ( .A(n123), .Q(n48) );
  INV3 U34 ( .A(n6), .Q(n5) );
  INV3 U35 ( .A(n53), .Q(n1) );
  NOR21 U36 ( .A(n50), .B(n11), .Q(n53) );
  INV3 U37 ( .A(n170), .Q(n18) );
  INV3 U38 ( .A(n120), .Q(n30) );
  INV3 U39 ( .A(n55), .Q(n14) );
  INV3 U40 ( .A(n54), .Q(n44) );
  INV3 U41 ( .A(n62), .Q(n45) );
  INV3 U42 ( .A(n76), .Q(n25) );
  INV3 U43 ( .A(n72), .Q(n42) );
  INV3 U44 ( .A(n179), .Q(n22) );
  BUF2 U45 ( .A(n97), .Q(n4) );
  INV3 U46 ( .A(n117), .Q(n50) );
  INV3 U47 ( .A(n12), .Q(n11) );
  INV3 U48 ( .A(n98), .Q(n6) );
  INV3 U49 ( .A(SH[2]), .Q(n9) );
  INV3 U50 ( .A(SH[1]), .Q(n8) );
  INV3 U51 ( .A(SH[0]), .Q(n7) );
  BUF2 U52 ( .A(n96), .Q(n3) );
  INV3 U53 ( .A(SH[3]), .Q(n10) );
  NOR21 U54 ( .A(SH[2]), .B(SH[3]), .Q(n117) );
  INV3 U55 ( .A(SH[4]), .Q(n12) );
  NOR21 U56 ( .A(n207), .B(SH[2]), .Q(n56) );
  OAI2110 U57 ( .A(n40), .B(n46), .C(n51), .D(n52), .Q(B[9]) );
  AOI220 U58 ( .A(n53), .B(n54), .C(n11), .D(n14), .Q(n52) );
  AOI220 U59 ( .A(n56), .B(n57), .C(n58), .D(n59), .Q(n51) );
  OAI2110 U60 ( .A(n41), .B(n46), .C(n60), .D(n61), .Q(B[8]) );
  AOI220 U61 ( .A(n53), .B(n62), .C(n11), .D(n63), .Q(n61) );
  AOI220 U62 ( .A(n56), .B(n64), .C(n58), .D(n65), .Q(n60) );
  OAI2110 U63 ( .A(n42), .B(n46), .C(n66), .D(n67), .Q(B[7]) );
  AOI220 U64 ( .A(n53), .B(n68), .C(n11), .D(n69), .Q(n67) );
  AOI220 U65 ( .A(n56), .B(n70), .C(n58), .D(n71), .Q(n66) );
  OAI2110 U66 ( .A(n43), .B(n46), .C(n73), .D(n74), .Q(B[6]) );
  AOI220 U67 ( .A(n53), .B(n75), .C(n11), .D(n25), .Q(n74) );
  AOI220 U68 ( .A(n56), .B(n77), .C(n58), .D(n78), .Q(n73) );
  OAI2110 U69 ( .A(n44), .B(n46), .C(n79), .D(n80), .Q(B[5]) );
  AOI220 U70 ( .A(n53), .B(n81), .C(n11), .D(n16), .Q(n80) );
  AOI220 U71 ( .A(n56), .B(n83), .C(n58), .D(n57), .Q(n79) );
  OAI2110 U72 ( .A(n45), .B(n46), .C(n84), .D(n85), .Q(B[4]) );
  AOI220 U73 ( .A(n53), .B(n86), .C(n11), .D(n27), .Q(n85) );
  AOI220 U74 ( .A(n56), .B(n88), .C(n58), .D(n64), .Q(n84) );
  OAI2110 U75 ( .A(n37), .B(n47), .C(n89), .D(n90), .Q(B[3]) );
  AOI220 U76 ( .A(n91), .B(n68), .C(n11), .D(n92), .Q(n90) );
  NAND20 U77 ( .A(n93), .B(n94), .Q(n68) );
  AOI220 U78 ( .A(A[10]), .B(n2), .C(A[9]), .D(n3), .Q(n94) );
  AOI220 U79 ( .A(A[8]), .B(n97), .C(A[7]), .D(n5), .Q(n93) );
  AOI220 U80 ( .A(n53), .B(n99), .C(n56), .D(n72), .Q(n89) );
  NAND20 U81 ( .A(n100), .B(n101), .Q(n99) );
  AOI220 U82 ( .A(A[6]), .B(n2), .C(A[5]), .D(n96), .Q(n101) );
  AOI220 U83 ( .A(A[4]), .B(n97), .C(A[3]), .D(n5), .Q(n100) );
  NOR20 U84 ( .A(n1), .B(n102), .Q(B[31]) );
  NOR20 U85 ( .A(n103), .B(n1), .Q(B[30]) );
  OAI2110 U86 ( .A(n39), .B(n47), .C(n104), .D(n105), .Q(B[2]) );
  AOI220 U87 ( .A(n91), .B(n75), .C(n11), .D(n106), .Q(n105) );
  NAND20 U88 ( .A(n107), .B(n108), .Q(n75) );
  AOI220 U89 ( .A(A[9]), .B(n2), .C(A[8]), .D(n3), .Q(n108) );
  AOI220 U90 ( .A(A[7]), .B(n97), .C(A[6]), .D(n5), .Q(n107) );
  AOI220 U91 ( .A(n53), .B(n109), .C(n56), .D(n110), .Q(n104) );
  NAND20 U92 ( .A(n111), .B(n112), .Q(n109) );
  AOI220 U93 ( .A(A[5]), .B(n2), .C(A[4]), .D(n96), .Q(n112) );
  AOI220 U94 ( .A(A[3]), .B(n4), .C(A[2]), .D(n5), .Q(n111) );
  NOR20 U95 ( .A(n113), .B(n1), .Q(B[29]) );
  NOR20 U96 ( .A(n29), .B(n1), .Q(B[28]) );
  NOR30 U97 ( .A(n114), .B(n11), .C(SH[3]), .Q(B[27]) );
  NOR20 U98 ( .A(n11), .B(n115), .Q(B[26]) );
  NOR20 U99 ( .A(n11), .B(n55), .Q(B[25]) );
  AOI220 U100 ( .A(n116), .B(n117), .C(n15), .D(n118), .Q(n55) );
  NOR20 U101 ( .A(n11), .B(n28), .Q(B[24]) );
  OAI220 U102 ( .A(n33), .B(n50), .C(n29), .D(n49), .Q(n63) );
  NOR20 U103 ( .A(n11), .B(n20), .Q(B[23]) );
  OAI210 U104 ( .A(n34), .B(n50), .C(n119), .Q(n69) );
  AOI220 U105 ( .A(n48), .B(n21), .C(n118), .D(n120), .Q(n119) );
  NOR20 U106 ( .A(n11), .B(n76), .Q(B[22]) );
  AOI210 U107 ( .A(n121), .B(n117), .C(n122), .Q(n76) );
  OAI220 U108 ( .A(n123), .B(n103), .C(n49), .D(n31), .Q(n122) );
  NOR20 U109 ( .A(n11), .B(n82), .Q(B[21]) );
  AOI210 U110 ( .A(n59), .B(n117), .C(n124), .Q(n82) );
  OAI220 U111 ( .A(n123), .B(n113), .C(n49), .D(n32), .Q(n124) );
  NOR20 U112 ( .A(n11), .B(n87), .Q(B[20]) );
  AOI210 U113 ( .A(n65), .B(n117), .C(n125), .Q(n87) );
  OAI220 U114 ( .A(n123), .B(n29), .C(n49), .D(n33), .Q(n125) );
  OAI2110 U115 ( .A(n40), .B(n47), .C(n127), .D(n128), .Q(B[1]) );
  AOI220 U116 ( .A(n91), .B(n81), .C(n11), .D(n129), .Q(n128) );
  NAND20 U117 ( .A(n130), .B(n131), .Q(n81) );
  AOI220 U118 ( .A(A[8]), .B(n95), .C(A[7]), .D(n96), .Q(n131) );
  AOI220 U119 ( .A(A[6]), .B(n97), .C(A[5]), .D(n5), .Q(n130) );
  AOI220 U120 ( .A(n53), .B(n132), .C(n56), .D(n54), .Q(n127) );
  NAND20 U121 ( .A(n133), .B(n134), .Q(n54) );
  AOI220 U122 ( .A(A[12]), .B(n95), .C(A[11]), .D(n3), .Q(n134) );
  AOI220 U123 ( .A(A[10]), .B(n97), .C(A[9]), .D(n5), .Q(n133) );
  NAND20 U124 ( .A(n135), .B(n136), .Q(n132) );
  AOI220 U125 ( .A(A[4]), .B(n95), .C(A[3]), .D(n96), .Q(n136) );
  AOI220 U126 ( .A(A[2]), .B(n4), .C(A[1]), .D(n5), .Q(n135) );
  NOR20 U127 ( .A(n11), .B(n19), .Q(B[19]) );
  OAI210 U128 ( .A(n114), .B(n10), .C(n137), .Q(n92) );
  AOI220 U129 ( .A(n118), .B(n138), .C(n117), .D(n71), .Q(n137) );
  NOR20 U130 ( .A(n11), .B(n23), .Q(B[18]) );
  OAI2110 U131 ( .A(n35), .B(n50), .C(n139), .D(n140), .Q(n106) );
  AOI220 U132 ( .A(n141), .B(n24), .C(n48), .D(n142), .Q(n140) );
  NAND20 U133 ( .A(n118), .B(n121), .Q(n139) );
  NOR20 U134 ( .A(n11), .B(n13), .Q(B[17]) );
  NAND20 U135 ( .A(n143), .B(n144), .Q(n129) );
  AOI220 U136 ( .A(n141), .B(n15), .C(n48), .D(n116), .Q(n144) );
  AOI220 U137 ( .A(n118), .B(n59), .C(n117), .D(n57), .Q(n143) );
  NOR20 U138 ( .A(n11), .B(n26), .Q(B[16]) );
  OAI2110 U139 ( .A(n30), .B(n47), .C(n146), .D(n147), .Q(B[15]) );
  AOI220 U140 ( .A(n91), .B(n71), .C(n53), .D(n70), .Q(n147) );
  AOI220 U141 ( .A(n148), .B(n21), .C(n56), .D(n138), .Q(n146) );
  OAI2110 U142 ( .A(n31), .B(n47), .C(n149), .D(n150), .Q(B[14]) );
  AOI220 U143 ( .A(n91), .B(n78), .C(n53), .D(n77), .Q(n150) );
  AOI220 U144 ( .A(n148), .B(n24), .C(n56), .D(n121), .Q(n149) );
  OAI2110 U145 ( .A(n32), .B(n47), .C(n151), .D(n152), .Q(B[13]) );
  AOI220 U146 ( .A(n91), .B(n57), .C(n53), .D(n83), .Q(n152) );
  NAND20 U147 ( .A(n153), .B(n154), .Q(n83) );
  AOI220 U148 ( .A(A[16]), .B(n2), .C(A[15]), .D(n3), .Q(n154) );
  AOI220 U149 ( .A(A[14]), .B(n4), .C(A[13]), .D(n5), .Q(n153) );
  NAND20 U150 ( .A(n155), .B(n156), .Q(n57) );
  AOI220 U151 ( .A(A[20]), .B(n2), .C(A[19]), .D(n3), .Q(n156) );
  AOI220 U152 ( .A(A[18]), .B(n4), .C(A[17]), .D(n5), .Q(n155) );
  AOI220 U153 ( .A(n148), .B(n15), .C(n56), .D(n59), .Q(n151) );
  NAND20 U154 ( .A(n157), .B(n158), .Q(n59) );
  AOI220 U155 ( .A(A[24]), .B(n2), .C(A[23]), .D(n3), .Q(n158) );
  AOI220 U156 ( .A(A[22]), .B(n4), .C(A[21]), .D(n5), .Q(n157) );
  AOI210 U157 ( .A(n98), .B(A[29]), .C(n17), .Q(n113) );
  AOI220 U158 ( .A(A[31]), .B(n3), .C(A[30]), .D(n4), .Q(n159) );
  NAND20 U159 ( .A(n160), .B(n161), .Q(n116) );
  AOI220 U160 ( .A(A[28]), .B(n2), .C(A[27]), .D(n3), .Q(n161) );
  AOI220 U161 ( .A(A[26]), .B(n4), .C(A[25]), .D(n5), .Q(n160) );
  OAI2110 U162 ( .A(n33), .B(n47), .C(n162), .D(n163), .Q(B[12]) );
  AOI220 U163 ( .A(n91), .B(n64), .C(n53), .D(n88), .Q(n163) );
  AOI220 U164 ( .A(n148), .B(n126), .C(n56), .D(n65), .Q(n162) );
  NOR20 U165 ( .A(n12), .B(n50), .Q(n148) );
  OAI2110 U166 ( .A(n34), .B(n47), .C(n18), .D(n165), .Q(B[11]) );
  AOI220 U167 ( .A(n91), .B(n70), .C(n53), .D(n72), .Q(n165) );
  NAND20 U168 ( .A(n166), .B(n167), .Q(n72) );
  AOI220 U169 ( .A(A[14]), .B(n95), .C(A[13]), .D(n3), .Q(n167) );
  AOI220 U170 ( .A(A[12]), .B(n4), .C(A[11]), .D(n5), .Q(n166) );
  NAND20 U171 ( .A(n168), .B(n169), .Q(n70) );
  AOI220 U172 ( .A(A[18]), .B(n95), .C(A[17]), .D(n3), .Q(n169) );
  AOI220 U173 ( .A(A[16]), .B(n4), .C(A[15]), .D(n98), .Q(n168) );
  OAI310 U174 ( .A(n114), .B(SH[3]), .C(n12), .D(n171), .Q(n170) );
  NAND20 U175 ( .A(n71), .B(n56), .Q(n171) );
  OAI2110 U176 ( .A(n36), .B(n6), .C(n172), .D(n173), .Q(n71) );
  AOI220 U177 ( .A(A[22]), .B(n2), .C(A[21]), .D(n3), .Q(n173) );
  NAND20 U178 ( .A(n4), .B(A[20]), .Q(n172) );
  IMUX20 U179 ( .A(n21), .B(n120), .S(n9), .Q(n114) );
  NAND20 U180 ( .A(n174), .B(n175), .Q(n120) );
  AOI220 U181 ( .A(A[30]), .B(n2), .C(A[29]), .D(n3), .Q(n175) );
  AOI220 U182 ( .A(A[28]), .B(n4), .C(A[27]), .D(n5), .Q(n174) );
  NAND20 U183 ( .A(A[31]), .B(n98), .Q(n102) );
  NAND20 U184 ( .A(n176), .B(n177), .Q(n138) );
  AOI220 U185 ( .A(A[26]), .B(n95), .C(A[25]), .D(n3), .Q(n177) );
  AOI220 U186 ( .A(A[24]), .B(n97), .C(A[23]), .D(n98), .Q(n176) );
  OAI2110 U187 ( .A(n39), .B(n46), .C(n178), .D(n22), .Q(B[10]) );
  OAI220 U188 ( .A(n1), .B(n43), .C(n12), .D(n115), .Q(n179) );
  AOI220 U189 ( .A(n142), .B(n117), .C(n24), .D(n118), .Q(n115) );
  AOI220 U190 ( .A(n5), .B(A[30]), .C(n4), .D(A[31]), .Q(n103) );
  NAND20 U191 ( .A(n180), .B(n181), .Q(n142) );
  AOI220 U192 ( .A(A[29]), .B(n2), .C(A[28]), .D(n3), .Q(n181) );
  AOI220 U193 ( .A(A[27]), .B(n4), .C(A[26]), .D(n5), .Q(n180) );
  NAND20 U194 ( .A(n182), .B(n183), .Q(n110) );
  AOI220 U195 ( .A(A[13]), .B(n2), .C(A[12]), .D(n3), .Q(n183) );
  AOI220 U196 ( .A(A[11]), .B(n97), .C(A[10]), .D(n5), .Q(n182) );
  AOI220 U197 ( .A(n56), .B(n78), .C(n58), .D(n121), .Q(n178) );
  NAND20 U198 ( .A(n184), .B(n185), .Q(n121) );
  AOI220 U199 ( .A(A[25]), .B(n95), .C(A[24]), .D(n3), .Q(n185) );
  AOI220 U200 ( .A(A[23]), .B(n4), .C(A[22]), .D(n5), .Q(n184) );
  OAI2110 U201 ( .A(n38), .B(n6), .C(n186), .D(n187), .Q(n78) );
  AOI220 U202 ( .A(A[21]), .B(n2), .C(n96), .D(A[20]), .Q(n187) );
  NAND20 U203 ( .A(n4), .B(A[19]), .Q(n186) );
  NAND20 U204 ( .A(n188), .B(n189), .Q(n77) );
  AOI220 U205 ( .A(A[17]), .B(n95), .C(A[16]), .D(n96), .Q(n189) );
  AOI220 U206 ( .A(A[15]), .B(n4), .C(A[14]), .D(n5), .Q(n188) );
  OAI2110 U207 ( .A(n41), .B(n47), .C(n190), .D(n191), .Q(B[0]) );
  AOI220 U208 ( .A(n91), .B(n86), .C(n11), .D(n145), .Q(n191) );
  NAND20 U209 ( .A(n192), .B(n193), .Q(n145) );
  AOI220 U210 ( .A(n141), .B(n126), .C(n48), .D(n164), .Q(n193) );
  NAND20 U211 ( .A(n194), .B(n195), .Q(n164) );
  AOI220 U212 ( .A(A[27]), .B(n95), .C(A[26]), .D(n3), .Q(n195) );
  AOI220 U213 ( .A(A[25]), .B(n97), .C(A[24]), .D(n98), .Q(n194) );
  NAND20 U214 ( .A(SH[3]), .B(n9), .Q(n123) );
  NAND20 U215 ( .A(n196), .B(n197), .Q(n126) );
  AOI220 U216 ( .A(A[31]), .B(n2), .C(A[30]), .D(n3), .Q(n197) );
  AOI220 U217 ( .A(A[29]), .B(n4), .C(A[28]), .D(n98), .Q(n196) );
  NOR20 U218 ( .A(n9), .B(n10), .Q(n141) );
  AOI220 U219 ( .A(n118), .B(n65), .C(n117), .D(n64), .Q(n192) );
  NAND20 U220 ( .A(n198), .B(n199), .Q(n64) );
  AOI220 U221 ( .A(A[19]), .B(n2), .C(A[18]), .D(n3), .Q(n199) );
  AOI220 U222 ( .A(A[17]), .B(n4), .C(A[16]), .D(n98), .Q(n198) );
  NAND20 U223 ( .A(n200), .B(n201), .Q(n65) );
  AOI220 U224 ( .A(A[23]), .B(n2), .C(A[22]), .D(n3), .Q(n201) );
  AOI220 U225 ( .A(A[21]), .B(n4), .C(n98), .D(A[20]), .Q(n200) );
  NAND20 U226 ( .A(n202), .B(n203), .Q(n86) );
  AOI220 U227 ( .A(A[7]), .B(n2), .C(A[6]), .D(n96), .Q(n203) );
  AOI220 U228 ( .A(A[5]), .B(n4), .C(A[4]), .D(n5), .Q(n202) );
  NOR20 U229 ( .A(n9), .B(SH[3]), .Q(n118) );
  AOI220 U230 ( .A(n53), .B(n204), .C(n56), .D(n62), .Q(n190) );
  NAND20 U231 ( .A(n205), .B(n206), .Q(n62) );
  AOI220 U232 ( .A(A[11]), .B(n2), .C(A[10]), .D(n96), .Q(n206) );
  AOI220 U233 ( .A(A[9]), .B(n4), .C(A[8]), .D(n5), .Q(n205) );
  NAND20 U234 ( .A(n208), .B(n209), .Q(n204) );
  AOI220 U235 ( .A(A[3]), .B(n2), .C(A[2]), .D(n96), .Q(n209) );
  AOI220 U236 ( .A(A[1]), .B(n97), .C(A[0]), .D(n5), .Q(n208) );
  NOR20 U237 ( .A(n9), .B(n207), .Q(n58) );
  NAND20 U238 ( .A(SH[3]), .B(n12), .Q(n207) );
  NAND20 U239 ( .A(n210), .B(n211), .Q(n88) );
  AOI220 U240 ( .A(A[15]), .B(n2), .C(A[14]), .D(n3), .Q(n211) );
  NOR20 U241 ( .A(n8), .B(SH[0]), .Q(n96) );
  NOR20 U242 ( .A(n8), .B(n7), .Q(n95) );
  AOI220 U243 ( .A(A[13]), .B(n4), .C(A[12]), .D(n5), .Q(n210) );
  NOR20 U244 ( .A(SH[0]), .B(SH[1]), .Q(n98) );
  NOR20 U245 ( .A(n7), .B(SH[1]), .Q(n97) );
endmodule


module E_alu_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147;

  AOI220 U1 ( .A(B[22]), .B(n34), .C(B[21]), .D(n46), .Q(n38) );
  INV1 U2 ( .A(B[21]), .Q(n60) );
  NAND20 U3 ( .A(n47), .B(B[20]), .Q(n37) );
  INV0 U4 ( .A(B[20]), .Q(n59) );
  NOR20 U5 ( .A(B[11]), .B(n81), .Q(n76) );
  NAND20 U6 ( .A(B[5]), .B(n106), .Q(n128) );
  NOR20 U7 ( .A(B[5]), .B(n106), .Q(n105) );
  INV0 U8 ( .A(A[17]), .Q(n66) );
  INV0 U9 ( .A(A[18]), .Q(n56) );
  INV0 U10 ( .A(A[19]), .Q(n40) );
  AOI2110 U11 ( .A(A[1]), .B(n122), .C(n123), .D(n124), .Q(n121) );
  INV0 U12 ( .A(B[1]), .Q(n122) );
  NOR20 U13 ( .A(A[7]), .B(n92), .Q(n89) );
  AOI310 U14 ( .A(n115), .B(n126), .C(B[1]), .D(n107), .Q(n95) );
  NOR20 U15 ( .A(A[1]), .B(n130), .Q(n126) );
  NAND20 U16 ( .A(A[3]), .B(n118), .Q(n115) );
  AOI310 U17 ( .A(n115), .B(n116), .C(B[2]), .D(n117), .Q(n97) );
  NAND20 U18 ( .A(A[9]), .B(n112), .Q(n109) );
  INV0 U19 ( .A(B[9]), .Q(n112) );
  INV0 U20 ( .A(B[3]), .Q(n118) );
  NAND20 U21 ( .A(B[4]), .B(n108), .Q(n119) );
  NAND20 U22 ( .A(n93), .B(B[8]), .Q(n87) );
  INV0 U23 ( .A(B[8]), .Q(n111) );
  NAND20 U24 ( .A(A[2]), .B(n131), .Q(n120) );
  INV0 U25 ( .A(B[2]), .Q(n131) );
  INV0 U26 ( .A(A[6]), .Q(n129) );
  INV0 U27 ( .A(A[0]), .Q(n125) );
  INV0 U28 ( .A(A[5]), .Q(n106) );
  NAND20 U29 ( .A(A[7]), .B(n114), .Q(n99) );
  NAND20 U30 ( .A(A[6]), .B(n113), .Q(n100) );
  NOR20 U31 ( .A(B[4]), .B(n108), .Q(n103) );
  NOR20 U32 ( .A(B[10]), .B(n79), .Q(n78) );
  NAND20 U33 ( .A(B[9]), .B(n94), .Q(n85) );
  INV2 U34 ( .A(A[9]), .Q(n94) );
  NAND20 U35 ( .A(B[10]), .B(n79), .Q(n86) );
  INV0 U36 ( .A(A[4]), .Q(n108) );
  INV0 U37 ( .A(A[2]), .Q(n116) );
  INV0 U38 ( .A(B[0]), .Q(n123) );
  NOR20 U39 ( .A(B[0]), .B(n125), .Q(n124) );
  INV3 U40 ( .A(n24), .Q(n17) );
  OAI2111 U41 ( .A(n72), .B(n73), .C(n74), .D(n75), .Q(n49) );
  NOR31 U42 ( .A(n71), .B(n82), .C(n83), .Q(n74) );
  AOI221 U43 ( .A(n76), .B(n77), .C(n78), .D(n77), .Q(n75) );
  NAND41 U44 ( .A(n85), .B(n86), .C(n87), .D(n88), .Q(n73) );
  OAI2111 U45 ( .A(n25), .B(n26), .C(n27), .D(n28), .Q(n2) );
  AOI2111 U46 ( .A(A[25]), .B(n35), .C(n24), .D(n36), .Q(n27) );
  AOI221 U47 ( .A(n29), .B(n30), .C(n31), .D(n30), .Q(n28) );
  NAND31 U48 ( .A(n37), .B(n38), .C(n39), .Q(n26) );
  AOI311 U49 ( .A(n1), .B(n2), .C(n3), .D(n4), .Q(LT_LE) );
  AOI311 U50 ( .A(B[25]), .B(n16), .C(n17), .D(n10), .Q(n3) );
  AOI2111 U51 ( .A(n140), .B(B[26]), .C(n141), .D(n142), .Q(n1) );
  NOR21 U52 ( .A(A[14]), .B(n71), .Q(n132) );
  INV3 U53 ( .A(n92), .Q(n101) );
  INV3 U54 ( .A(B[15]), .Q(n139) );
  NAND22 U55 ( .A(n18), .B(n14), .Q(n10) );
  NOR21 U56 ( .A(n21), .B(n22), .Q(n18) );
  NOR21 U57 ( .A(A[30]), .B(n13), .Q(n22) );
  NOR21 U58 ( .A(A[29]), .B(n23), .Q(n21) );
  NAND22 U59 ( .A(n57), .B(n58), .Q(n45) );
  NAND22 U60 ( .A(A[21]), .B(n60), .Q(n57) );
  NAND22 U61 ( .A(A[20]), .B(n59), .Q(n58) );
  AOI221 U62 ( .A(n61), .B(n62), .C(n63), .D(n62), .Q(n52) );
  NOR21 U63 ( .A(B[17]), .B(n66), .Q(n61) );
  NOR31 U64 ( .A(n10), .B(B[29]), .C(n12), .Q(n8) );
  INV3 U65 ( .A(A[29]), .Q(n12) );
  NOR31 U66 ( .A(n10), .B(B[28]), .C(n11), .Q(n9) );
  INV3 U67 ( .A(A[28]), .Q(n11) );
  NOR31 U68 ( .A(n45), .B(n54), .C(n55), .Q(n53) );
  NOR21 U69 ( .A(B[19]), .B(n40), .Q(n55) );
  NOR21 U70 ( .A(B[18]), .B(n56), .Q(n54) );
  NAND22 U71 ( .A(n69), .B(n70), .Q(n65) );
  NAND22 U72 ( .A(B[17]), .B(n66), .Q(n70) );
  NAND22 U73 ( .A(B[18]), .B(n56), .Q(n69) );
  INV3 U74 ( .A(n19), .Q(n14) );
  NOR21 U75 ( .A(A[31]), .B(n20), .Q(n19) );
  INV3 U76 ( .A(B[31]), .Q(n20) );
  NAND22 U77 ( .A(n42), .B(n43), .Q(n33) );
  NAND22 U78 ( .A(B[24]), .B(n44), .Q(n42) );
  NAND22 U79 ( .A(B[23]), .B(n32), .Q(n43) );
  INV3 U80 ( .A(A[24]), .Q(n44) );
  NAND31 U81 ( .A(n5), .B(n6), .C(n7), .Q(n4) );
  NAND22 U82 ( .A(n14), .B(n15), .Q(n5) );
  NAND31 U83 ( .A(A[30]), .B(n13), .C(n14), .Q(n6) );
  NOR21 U84 ( .A(n8), .B(n9), .Q(n7) );
  INV3 U85 ( .A(A[11]), .Q(n81) );
  INV3 U86 ( .A(A[12]), .Q(n84) );
  INV3 U87 ( .A(A[10]), .Q(n79) );
  INV3 U88 ( .A(A[13]), .Q(n67) );
  AOI311 U89 ( .A(n40), .B(n41), .C(B[19]), .D(n33), .Q(n39) );
  NOR21 U90 ( .A(A[20]), .B(n45), .Q(n47) );
  INV3 U91 ( .A(B[30]), .Q(n13) );
  NOR21 U92 ( .A(A[15]), .B(n139), .Q(n134) );
  INV3 U93 ( .A(B[29]), .Q(n23) );
  XOR21 U94 ( .A(B[31]), .B(A[31]), .Q(n15) );
  INV3 U95 ( .A(A[21]), .Q(n46) );
  NOR21 U96 ( .A(A[16]), .B(n135), .Q(n133) );
  NAND22 U97 ( .A(n144), .B(n145), .Q(n24) );
  NAND22 U98 ( .A(A[27]), .B(n147), .Q(n144) );
  NAND22 U99 ( .A(A[26]), .B(n146), .Q(n145) );
  INV3 U100 ( .A(B[27]), .Q(n147) );
  INV3 U101 ( .A(A[23]), .Q(n32) );
  NOR21 U102 ( .A(A[26]), .B(n24), .Q(n140) );
  INV3 U103 ( .A(A[22]), .Q(n34) );
  NOR21 U104 ( .A(A[28]), .B(n143), .Q(n141) );
  INV3 U105 ( .A(B[28]), .Q(n143) );
  NOR21 U106 ( .A(B[24]), .B(n44), .Q(n36) );
  NOR21 U107 ( .A(A[27]), .B(n147), .Q(n142) );
  NOR21 U108 ( .A(B[23]), .B(n32), .Q(n31) );
  NOR21 U109 ( .A(B[22]), .B(n34), .Q(n29) );
  INV3 U110 ( .A(B[26]), .Q(n146) );
  INV3 U111 ( .A(B[25]), .Q(n35) );
  INV3 U112 ( .A(A[25]), .Q(n16) );
  INV3 U113 ( .A(A[16]), .Q(n64) );
  INV3 U114 ( .A(n120), .Q(n130) );
  NAND22 U115 ( .A(n109), .B(n110), .Q(n92) );
  NAND22 U116 ( .A(A[8]), .B(n111), .Q(n110) );
  INV3 U117 ( .A(B[7]), .Q(n114) );
  NAND22 U118 ( .A(n136), .B(n137), .Q(n71) );
  NAND22 U119 ( .A(A[14]), .B(n138), .Q(n137) );
  NAND22 U120 ( .A(A[15]), .B(n139), .Q(n136) );
  INV3 U121 ( .A(B[14]), .Q(n138) );
  AOI311 U122 ( .A(n48), .B(n49), .C(n50), .D(n51), .Q(n25) );
  NAND22 U123 ( .A(n52), .B(n53), .Q(n51) );
  AOI311 U124 ( .A(n67), .B(n68), .C(B[13]), .D(n65), .Q(n50) );
  AOI2111 U125 ( .A(n132), .B(B[14]), .C(n133), .D(n134), .Q(n48) );
  AOI311 U126 ( .A(n95), .B(n96), .C(n97), .D(n98), .Q(n72) );
  NAND41 U127 ( .A(n120), .B(n125), .C(n115), .D(n121), .Q(n96) );
  NAND41 U128 ( .A(n99), .B(n100), .C(n101), .D(n102), .Q(n98) );
  INV3 U129 ( .A(B[6]), .Q(n113) );
  AOI211 U130 ( .A(n89), .B(B[7]), .C(n80), .Q(n88) );
  AOI221 U131 ( .A(n103), .B(n104), .C(n105), .D(n104), .Q(n102) );
  NAND22 U132 ( .A(n127), .B(n128), .Q(n107) );
  NAND22 U133 ( .A(B[6]), .B(n129), .Q(n127) );
  NAND22 U134 ( .A(n90), .B(n91), .Q(n80) );
  NAND22 U135 ( .A(B[12]), .B(n84), .Q(n90) );
  NAND22 U136 ( .A(B[11]), .B(n81), .Q(n91) );
  NOR21 U137 ( .A(A[8]), .B(n92), .Q(n93) );
  NOR21 U138 ( .A(B[12]), .B(n84), .Q(n82) );
  NOR21 U139 ( .A(B[13]), .B(n67), .Q(n83) );
  INV0 U140 ( .A(B[16]), .Q(n135) );
  NOR20 U141 ( .A(B[16]), .B(n64), .Q(n63) );
  CLKIN3 U142 ( .A(n33), .Q(n30) );
  CLKIN3 U143 ( .A(n45), .Q(n41) );
  CLKIN3 U144 ( .A(n65), .Q(n62) );
  CLKIN3 U145 ( .A(n71), .Q(n68) );
  CLKIN3 U146 ( .A(n80), .Q(n77) );
  CLKIN3 U147 ( .A(n107), .Q(n104) );
  OAI212 U148 ( .A(A[3]), .B(n118), .C(n119), .Q(n117) );
endmodule


module E_alu_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150;

  NAND22 U3 ( .A(n89), .B(n97), .Q(n106) );
  NAND22 U4 ( .A(n58), .B(n61), .Q(n70) );
  NAND22 U5 ( .A(n42), .B(n39), .Q(n43) );
  NAND22 U6 ( .A(n35), .B(n37), .Q(n38) );
  NAND22 U7 ( .A(n21), .B(n18), .Q(n22) );
  NAND22 U8 ( .A(n14), .B(n16), .Q(n17) );
  INV3 U9 ( .A(B[4]), .Q(n26) );
  INV3 U10 ( .A(n56), .Q(n77) );
  INV3 U11 ( .A(B[0]), .Q(n46) );
  INV0 U12 ( .A(A[2]), .Q(n132) );
  INV3 U13 ( .A(B[1]), .Q(n128) );
  NAND20 U14 ( .A(n3), .B(n4), .Q(n1) );
  INV0 U15 ( .A(A[1]), .Q(n133) );
  NAND20 U16 ( .A(A[0]), .B(n46), .Q(n44) );
  NAND21 U17 ( .A(A[5]), .B(n144), .Q(n18) );
  NOR20 U18 ( .A(A[3]), .B(n121), .Q(n135) );
  XOR20 U19 ( .A(n75), .B(n72), .Q(DIFF[13]) );
  XNR20 U20 ( .A(n70), .B(n68), .Q(DIFF[14]) );
  OAI211 U21 ( .A(n77), .B(n78), .C(n79), .Q(n76) );
  AOI210 U22 ( .A(n34), .B(n35), .C(n36), .Q(n33) );
  NAND20 U23 ( .A(n41), .B(n42), .Q(n40) );
  NAND21 U24 ( .A(A[1]), .B(n128), .Q(n39) );
  NAND22 U25 ( .A(A[4]), .B(n26), .Q(n25) );
  AOI221 U26 ( .A(A[3]), .B(n121), .C(n129), .D(n130), .Q(n119) );
  IMUX20 U27 ( .A(n82), .B(n83), .S(n77), .Q(DIFF[12]) );
  NAND20 U28 ( .A(n112), .B(n7), .Q(n111) );
  INV0 U29 ( .A(n29), .Q(n23) );
  INV0 U30 ( .A(A[6]), .Q(n146) );
  NAND20 U31 ( .A(B[2]), .B(n132), .Q(n35) );
  NAND20 U32 ( .A(B[1]), .B(n133), .Q(n42) );
  INV0 U33 ( .A(A[5]), .Q(n145) );
  NAND21 U34 ( .A(A[6]), .B(n142), .Q(n16) );
  NAND20 U35 ( .A(A[2]), .B(n125), .Q(n37) );
  INV0 U36 ( .A(B[2]), .Q(n125) );
  INV0 U37 ( .A(B[8]), .Q(n10) );
  NAND20 U38 ( .A(A[9]), .B(n108), .Q(n4) );
  INV0 U39 ( .A(B[9]), .Q(n108) );
  INV0 U40 ( .A(B[3]), .Q(n121) );
  NOR20 U41 ( .A(A[0]), .B(n46), .Q(n134) );
  NOR20 U42 ( .A(A[7]), .B(n118), .Q(n147) );
  XNR20 U43 ( .A(B[3]), .B(A[3]), .Q(n32) );
  NAND20 U44 ( .A(B[10]), .B(n150), .Q(n89) );
  NAND20 U45 ( .A(B[9]), .B(n109), .Q(n3) );
  INV0 U46 ( .A(A[9]), .Q(n109) );
  INV0 U47 ( .A(B[10]), .Q(n149) );
  NOR20 U48 ( .A(A[4]), .B(n26), .Q(n24) );
  XOR20 U49 ( .A(B[4]), .B(A[4]), .Q(n28) );
  NOR20 U50 ( .A(A[4]), .B(n26), .Q(n30) );
  IMUX20 U51 ( .A(n5), .B(n6), .S(n7), .Q(DIFF[8]) );
  XOR20 U52 ( .A(B[8]), .B(A[8]), .Q(n5) );
  XNR20 U53 ( .A(B[7]), .B(A[7]), .Q(n11) );
  INV0 U54 ( .A(A[7]), .Q(n139) );
  NOR20 U55 ( .A(A[0]), .B(n46), .Q(n45) );
  AOI2111 U56 ( .A(n47), .B(n48), .C(n49), .D(n50), .Q(DIFF[16]) );
  NOR21 U57 ( .A(B[15]), .B(n51), .Q(n50) );
  INV3 U58 ( .A(n65), .Q(n47) );
  XNR21 U59 ( .A(n66), .B(n67), .Q(DIFF[15]) );
  XNR21 U60 ( .A(B[15]), .B(A[15]), .Q(n66) );
  AOI211 U61 ( .A(n68), .B(n58), .C(n69), .Q(n67) );
  AOI211 U62 ( .A(n31), .B(n21), .C(n143), .Q(n141) );
  NOR21 U63 ( .A(A[12]), .B(n55), .Q(n78) );
  AOI211 U64 ( .A(n126), .B(n42), .C(n127), .Q(n124) );
  NOR31 U65 ( .A(n52), .B(n77), .C(n53), .Q(n49) );
  NAND22 U66 ( .A(n57), .B(n58), .Q(n52) );
  NOR21 U67 ( .A(n131), .B(n123), .Q(n130) );
  AOI211 U68 ( .A(n9), .B(n3), .C(n98), .Q(n96) );
  NAND22 U69 ( .A(n99), .B(n111), .Q(n110) );
  INV3 U70 ( .A(n148), .Q(n112) );
  XNR21 U71 ( .A(n22), .B(n20), .Q(DIFF[5]) );
  XNR21 U72 ( .A(n17), .B(n13), .Q(DIFF[6]) );
  XOR21 U73 ( .A(n1), .B(n2), .Q(DIFF[9]) );
  NAND22 U74 ( .A(n57), .B(n64), .Q(n75) );
  NAND22 U75 ( .A(A[8]), .B(n10), .Q(n99) );
  NAND22 U76 ( .A(n18), .B(n19), .Q(n13) );
  NAND22 U77 ( .A(n20), .B(n21), .Q(n19) );
  XNR21 U78 ( .A(n106), .B(n104), .Q(DIFF[10]) );
  NOR21 U79 ( .A(n87), .B(n88), .Q(n86) );
  NAND22 U80 ( .A(n3), .B(n89), .Q(n88) );
  AOI211 U81 ( .A(n62), .B(n57), .C(n63), .Q(n60) );
  INV3 U82 ( .A(n64), .Q(n63) );
  XNR21 U83 ( .A(n43), .B(n41), .Q(DIFF[1]) );
  XNR21 U84 ( .A(n38), .B(n34), .Q(DIFF[2]) );
  NAND22 U85 ( .A(A[12]), .B(n55), .Q(n79) );
  NAND22 U86 ( .A(n39), .B(n40), .Q(n34) );
  NOR21 U87 ( .A(A[8]), .B(n10), .Q(n148) );
  NOR21 U88 ( .A(A[15]), .B(n54), .Q(n65) );
  INV3 U89 ( .A(B[15]), .Q(n54) );
  INV3 U90 ( .A(A[15]), .Q(n51) );
  INV3 U91 ( .A(A[11]), .Q(n94) );
  INV3 U92 ( .A(n100), .Q(n91) );
  NOR21 U93 ( .A(A[11]), .B(n90), .Q(n100) );
  NAND22 U94 ( .A(B[5]), .B(n145), .Q(n21) );
  NAND22 U95 ( .A(B[6]), .B(n146), .Q(n14) );
  NAND22 U96 ( .A(n113), .B(n114), .Q(n7) );
  AOI211 U97 ( .A(n136), .B(n137), .C(n138), .Q(n113) );
  NAND22 U98 ( .A(n29), .B(n115), .Q(n114) );
  NOR21 U99 ( .A(B[7]), .B(n139), .Q(n138) );
  NAND22 U100 ( .A(n119), .B(n120), .Q(n29) );
  NOR21 U101 ( .A(n134), .B(n135), .Q(n129) );
  NAND22 U102 ( .A(n84), .B(n85), .Q(n56) );
  AOI211 U103 ( .A(n91), .B(n92), .C(n93), .Q(n84) );
  NAND22 U104 ( .A(n7), .B(n86), .Q(n85) );
  NOR21 U105 ( .A(B[11]), .B(n94), .Q(n93) );
  INV3 U106 ( .A(B[6]), .Q(n142) );
  INV3 U107 ( .A(B[5]), .Q(n144) );
  XNR21 U108 ( .A(n32), .B(n33), .Q(DIFF[3]) );
  IMUX21 U109 ( .A(n27), .B(n28), .S(n23), .Q(DIFF[4]) );
  NOR21 U110 ( .A(n30), .B(n31), .Q(n27) );
  NOR21 U111 ( .A(n8), .B(n9), .Q(n6) );
  NOR21 U112 ( .A(A[8]), .B(n10), .Q(n8) );
  XOR21 U113 ( .A(B[12]), .B(A[12]), .Q(n83) );
  NOR21 U114 ( .A(n101), .B(n62), .Q(n82) );
  NOR21 U115 ( .A(A[12]), .B(n55), .Q(n101) );
  INV3 U116 ( .A(B[7]), .Q(n118) );
  XNR21 U117 ( .A(n11), .B(n12), .Q(DIFF[7]) );
  AOI211 U118 ( .A(n13), .B(n14), .C(n15), .Q(n12) );
  XNR21 U119 ( .A(n102), .B(n103), .Q(DIFF[11]) );
  XNR21 U120 ( .A(B[11]), .B(A[11]), .Q(n102) );
  AOI211 U121 ( .A(n104), .B(n89), .C(n105), .Q(n103) );
  NOR21 U122 ( .A(n116), .B(n117), .Q(n115) );
  NAND22 U123 ( .A(n21), .B(n14), .Q(n117) );
  INV3 U124 ( .A(n147), .Q(n136) );
  NAND22 U125 ( .A(B[14]), .B(n74), .Q(n58) );
  INV3 U126 ( .A(A[14]), .Q(n74) );
  INV3 U127 ( .A(A[10]), .Q(n150) );
  NAND22 U128 ( .A(B[13]), .B(n81), .Q(n57) );
  INV3 U129 ( .A(A[13]), .Q(n81) );
  NAND22 U130 ( .A(A[13]), .B(n80), .Q(n64) );
  INV3 U131 ( .A(B[13]), .Q(n80) );
  INV3 U132 ( .A(B[12]), .Q(n55) );
  NAND22 U133 ( .A(A[14]), .B(n73), .Q(n61) );
  INV3 U134 ( .A(B[14]), .Q(n73) );
  NAND22 U135 ( .A(n44), .B(n45), .Q(n41) );
  INV3 U136 ( .A(B[11]), .Q(n90) );
  NAND22 U137 ( .A(A[10]), .B(n149), .Q(n97) );
  CLKIN3 U138 ( .A(n16), .Q(n15) );
  OAI212 U139 ( .A(n23), .B(n24), .C(n25), .Q(n20) );
  CLKIN3 U140 ( .A(n37), .Q(n36) );
  OAI222 U141 ( .A(A[15]), .B(n54), .C(A[12]), .D(n55), .Q(n53) );
  OAI212 U142 ( .A(n59), .B(n60), .C(n61), .Q(n48) );
  CLKIN3 U143 ( .A(n58), .Q(n59) );
  CLKIN3 U144 ( .A(n61), .Q(n69) );
  OAI212 U145 ( .A(n71), .B(n72), .C(n64), .Q(n68) );
  CLKIN3 U146 ( .A(n57), .Q(n71) );
  CLKIN3 U147 ( .A(n76), .Q(n72) );
  OAI222 U148 ( .A(A[8]), .B(n10), .C(A[11]), .D(n90), .Q(n87) );
  OAI212 U149 ( .A(n95), .B(n96), .C(n97), .Q(n92) );
  CLKIN3 U150 ( .A(n4), .Q(n98) );
  CLKIN3 U151 ( .A(n99), .Q(n9) );
  CLKIN3 U152 ( .A(n89), .Q(n95) );
  CLKIN3 U153 ( .A(n79), .Q(n62) );
  CLKIN3 U154 ( .A(n97), .Q(n105) );
  OAI212 U155 ( .A(n2), .B(n107), .C(n4), .Q(n104) );
  CLKIN3 U156 ( .A(n3), .Q(n107) );
  CLKIN3 U157 ( .A(n110), .Q(n2) );
  OAI222 U158 ( .A(A[7]), .B(n118), .C(A[4]), .D(n26), .Q(n116) );
  OAI212 U159 ( .A(A[3]), .B(n121), .C(n122), .Q(n120) );
  OAI212 U160 ( .A(n123), .B(n124), .C(n37), .Q(n122) );
  CLKIN3 U161 ( .A(n39), .Q(n127) );
  CLKIN3 U162 ( .A(n35), .Q(n123) );
  CLKIN3 U163 ( .A(n42), .Q(n131) );
  OAI212 U164 ( .A(n140), .B(n141), .C(n16), .Q(n137) );
  CLKIN3 U165 ( .A(n18), .Q(n143) );
  CLKIN3 U166 ( .A(n25), .Q(n31) );
  CLKIN3 U167 ( .A(n14), .Q(n140) );
  OAI212 U168 ( .A(A[0]), .B(n46), .C(n44), .Q(DIFF[0]) );
  CLKIN3 U169 ( .A(n44), .Q(n126) );
endmodule


module E_alu ( o_data_AluRes, i_data_A, i_data_B, i_con_AluCtrl, i_data_shamt
 );
  output [31:0] o_data_AluRes;
  input [31:0] i_data_A;
  input [31:0] i_data_B;
  input [3:0] i_con_AluCtrl;
  input [4:0] i_data_shamt;
  wire   N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N306, n41, n42,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n426, n428, n429, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n144, n145, n146, n147, n162, n204, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n427, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440;
  wire   [8:0] sum_1;
  wire   [8:0] pre_sum_2a;
  wire   [8:0] pre_sum_2b;
  wire   [8:0] pre_sum_3a;
  wire   [8:0] pre_sum_3b;
  wire   [7:0] pre_sum_4a;
  wire   [7:0] pre_sum_4b;
  wire   [16:0] half_sub;
  wire   [15:0] pre_suba;
  wire   [15:0] pre_subb;

  OAI222 U28 ( .A(n439), .B(n417), .C(n32), .D(n74), .Q(n137) );
  OAI222 U36 ( .A(n72), .B(n419), .C(n31), .D(n139), .Q(n152) );
  OAI222 U46 ( .A(n72), .B(n421), .C(i_data_A[7]), .D(n139), .Q(n159) );
  OAI222 U54 ( .A(n72), .B(n423), .C(i_data_A[6]), .D(n139), .Q(n167) );
  OAI222 U62 ( .A(n72), .B(n425), .C(i_data_A[5]), .D(n139), .Q(n174) );
  OAI222 U70 ( .A(n72), .B(n430), .C(i_data_A[4]), .D(n74), .Q(n181) );
  OAI222 U78 ( .A(n72), .B(n432), .C(i_data_A[3]), .D(n139), .Q(n188) );
  OAI212 U85 ( .A(n109), .B(n71), .C(i_data_B[31]), .Q(n197) );
  OAI212 U87 ( .A(n199), .B(n108), .C(n200), .Q(n195) );
  OAI212 U95 ( .A(n440), .B(n129), .C(n211), .Q(n209) );
  OAI222 U102 ( .A(n439), .B(n110), .C(n64), .D(n139), .Q(n214) );
  OAI222 U107 ( .A(n439), .B(n434), .C(i_data_A[2]), .D(n139), .Q(n219) );
  OAI212 U114 ( .A(n440), .B(n131), .C(n228), .Q(n226) );
  OAI222 U121 ( .A(n439), .B(n111), .C(i_data_A[29]), .D(n139), .Q(n231) );
  OAI212 U125 ( .A(n440), .B(n144), .C(n238), .Q(n236) );
  OAI222 U132 ( .A(n439), .B(n112), .C(n61), .D(n139), .Q(n241) );
  OAI212 U136 ( .A(n440), .B(n146), .C(n248), .Q(n246) );
  OAI222 U143 ( .A(n439), .B(n113), .C(n59), .D(n139), .Q(n251) );
  OAI212 U147 ( .A(n440), .B(n162), .C(n258), .Q(n256) );
  OAI222 U154 ( .A(n72), .B(n114), .C(n57), .D(n139), .Q(n261) );
  OAI212 U158 ( .A(n416), .B(n440), .C(n268), .Q(n266) );
  OAI222 U165 ( .A(n72), .B(n115), .C(n55), .D(n139), .Q(n271) );
  OAI212 U169 ( .A(n418), .B(n440), .C(n278), .Q(n276) );
  OAI212 U183 ( .A(n420), .B(n440), .C(n291), .Q(n289) );
  OAI222 U190 ( .A(n439), .B(n117), .C(i_data_A[23]), .D(n74), .Q(n295) );
  OAI212 U194 ( .A(n422), .B(n440), .C(n303), .Q(n301) );
  OAI222 U201 ( .A(n439), .B(n118), .C(n50), .D(n74), .Q(n306) );
  OAI212 U205 ( .A(n424), .B(n440), .C(n313), .Q(n311) );
  OAI222 U212 ( .A(n439), .B(n119), .C(i_data_A[21]), .D(n74), .Q(n316) );
  OAI212 U216 ( .A(n427), .B(n440), .C(n323), .Q(n321) );
  OAI222 U223 ( .A(n439), .B(n120), .C(n48), .D(n74), .Q(n326) );
  OAI222 U228 ( .A(n72), .B(n436), .C(i_data_A[1]), .D(n74), .Q(n331) );
  OAI212 U235 ( .A(n431), .B(n440), .C(n340), .Q(n338) );
  OAI222 U242 ( .A(n439), .B(n121), .C(n46), .D(n74), .Q(n343) );
  OAI212 U246 ( .A(n440), .B(n433), .C(n350), .Q(n348) );
  OAI222 U253 ( .A(n72), .B(n123), .C(n44), .D(n74), .Q(n353) );
  OAI212 U257 ( .A(n440), .B(n435), .C(n360), .Q(n358) );
  OAI222 U264 ( .A(n72), .B(n125), .C(n43), .D(n74), .Q(n363) );
  OAI212 U268 ( .A(n440), .B(n437), .C(n370), .Q(n368) );
  OAI222 U281 ( .A(n439), .B(n127), .C(n40), .D(n74), .Q(n373) );
  OAI222 U284 ( .A(n72), .B(n128), .C(i_data_A[15]), .D(n74), .Q(n378) );
  OAI222 U292 ( .A(n72), .B(n130), .C(n38), .D(n74), .Q(n385) );
  OAI222 U300 ( .A(n439), .B(n132), .C(n36), .D(n74), .Q(n392) );
  OAI222 U308 ( .A(n72), .B(n145), .C(n35), .D(n74), .Q(n399) );
  OAI222 U316 ( .A(n72), .B(n147), .C(n34), .D(n74), .Q(n406) );
  OAI222 U325 ( .A(n72), .B(n204), .C(n33), .D(n139), .Q(n413) );
  E_alu_DW01_ash_0 sll_56 ( .A({i_data_B[31:20], n18, n15, n13, i_data_B[16:0]}), .DATA_TC(n42), .SH(i_data_shamt), .SH_TC(n42), .B({N224, N223, N222, N221, 
        N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, 
        N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, 
        N196, N195, N194, N193}) );
  E_alu_DW01_sub_0 sub_1_root_sub_35_2 ( .A({n66, n64, n62, n61, n59, n57, n55, 
        i_data_A[24], n52, n51, i_data_A[21], n48, n47, n45, n43, i_data_A[16]}), .B({i_data_B[31:23], n22, i_data_B[21:19], n16, n13, n12}), .CI(n41), 
        .DIFF(pre_subb) );
  E_alu_DW01_sub_1 sub_34 ( .A({n66, n63, i_data_A[29], n61, n59, n57, n54, 
        n53, n52, n50, n49, n48, n46, n45, i_data_A[17:16]}), .B({
        i_data_B[31:19], n16, n13, n12}), .CI(n42), .DIFF(pre_suba) );
  E_alu_DW01_add_0 add_1_root_add_31_2 ( .A({n65, n63, n62, n60, n58, n56, n54, 
        n53}), .B(i_data_B[31:24]), .CI(n41), .SUM(pre_sum_4b) );
  E_alu_DW01_add_1 add_30 ( .A({n65, n63, n62, n60, n58, n56, n54, n53}), .B(
        i_data_B[31:24]), .CI(n42), .SUM(pre_sum_4a) );
  E_alu_DW01_add_2 add_1_root_add_29_2 ( .A({n42, n52, n51, n49, n48, n47, n44, 
        n2, n40}), .B({n42, i_data_B[23], n22, i_data_B[21:19], n16, n13, n12}), .CI(n41), .SUM(pre_sum_3b) );
  E_alu_DW01_add_3 add_28 ( .A({n42, i_data_A[23], n50, n49, n48, n46, n44, n2, 
        n40}), .B({n42, i_data_B[23], n22, i_data_B[21:19], n16, n13, n12}), 
        .CI(n42), .SUM(pre_sum_3a) );
  E_alu_DW01_add_4 add_1_root_add_27_2 ( .A({n42, n39, n38, n36, n35, n34, n33, 
        n32, i_data_A[8]}), .B({n42, i_data_B[15:8]}), .CI(n41), .SUM(
        pre_sum_2b) );
  E_alu_DW01_add_5 add_26 ( .A({n42, n39, n37, n36, n35, n34, n33, n32, 
        i_data_A[8]}), .B({n42, i_data_B[15:8]}), .CI(n42), .SUM(pre_sum_2a)
         );
  E_alu_DW01_add_6 add_25 ( .A({n42, i_data_A[7:0]}), .B({n42, i_data_B[7:0]}), 
        .CI(n42), .SUM(sum_1) );
  E_alu_DW_rash_0 r130 ( .A({i_data_B[31:23], n22, i_data_B[21:20], n18, n15, 
        n13, n12, i_data_B[15:0]}), .DATA_TC(n42), .SH(i_data_shamt), .SH_TC(
        n42), .B({N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, 
        N234, N233, N232, N231, N230, N229, N228, N227, N226, N225}) );
  E_alu_DW01_cmp2_1 r131 ( .A({n65, n63, n62, n60, n58, n56, n54, n53, 
        i_data_A[23], n50, n49, n48, n46, n44, n2, n40, n39, n37, n36, n35, 
        n34, n33, n32, n31, i_data_A[7:0]}), .B({i_data_B[31:23], n22, 
        i_data_B[21:20], n18, n15, n13, n12, i_data_B[15:0]}), .LEQ(n42), .TC(
        n42), .LT_LE(N306) );
  E_alu_DW01_sub_3 sub_33 ( .A({n42, n39, n37, n36, n35, n34, n33, i_data_A[9], 
        n31, i_data_A[7:0]}), .B({n42, i_data_B[15:0]}), .CI(n42), .DIFF(
        half_sub) );
  BUF15 U3 ( .A(i_data_B[16]), .Q(n12) );
  BUF6 U4 ( .A(i_data_A[18]), .Q(n45) );
  INV8 U5 ( .A(n14), .Q(n16) );
  BUF6 U6 ( .A(n201), .Q(n3) );
  NAND22 U7 ( .A(n194), .B(n7), .Q(o_data_AluRes[31]) );
  AOI221 U8 ( .A(i_data_B[30]), .B(n212), .C(pre_suba[14]), .D(n69), .Q(n207)
         );
  AOI220 U9 ( .A(i_data_B[21]), .B(n314), .C(pre_suba[5]), .D(n69), .Q(n309)
         );
  INV1 U10 ( .A(i_data_A[29]), .Q(n111) );
  OAI220 U11 ( .A(n439), .B(n116), .C(i_data_A[24]), .D(n74), .Q(n282) );
  OAI2110 U12 ( .A(i_data_A[24]), .B(n72), .C(n70), .D(n280), .Q(n279) );
  NAND20 U13 ( .A(i_data_A[24]), .B(n67), .Q(n280) );
  INV0 U14 ( .A(i_data_A[24]), .Q(n116) );
  AOI220 U15 ( .A(i_data_B[20]), .B(n324), .C(pre_suba[4]), .D(n69), .Q(n319)
         );
  INV0 U16 ( .A(i_data_B[21]), .Q(n20) );
  INV0 U17 ( .A(i_data_B[20]), .Q(n19) );
  NOR21 U18 ( .A(n77), .B(half_sub[16]), .Q(n202) );
  BUF2 U19 ( .A(i_data_A[20]), .Q(n48) );
  NAND31 U20 ( .A(i_con_AluCtrl[0]), .B(n83), .C(n90), .Q(n438) );
  XOR21 U21 ( .A(i_data_B[31]), .B(n66), .Q(n1) );
  NOR20 U22 ( .A(n78), .B(n281), .Q(n201) );
  INV3 U23 ( .A(pre_subb[15]), .Q(n108) );
  INV3 U24 ( .A(n6), .Q(n7) );
  NAND31 U25 ( .A(n193), .B(n191), .C(n192), .Q(n6) );
  BUF2 U26 ( .A(i_data_A[17]), .Q(n43) );
  INV3 U27 ( .A(sum_1[8]), .Q(n106) );
  NOR21 U29 ( .A(n106), .B(n78), .Q(n140) );
  AOI2112 U30 ( .A(pre_sum_4a[7]), .B(n104), .C(n196), .D(n195), .Q(n194) );
  AOI2111 U31 ( .A(N223), .B(n99), .C(n209), .D(n210), .Q(n208) );
  AOI222 U32 ( .A(pre_sum_2a[8]), .B(n106), .C(pre_sum_2b[8]), .D(sum_1[8]), 
        .Q(n284) );
  BUF2 U33 ( .A(i_data_A[17]), .Q(n2) );
  CLKIN3 U34 ( .A(n68), .Q(n69) );
  NAND22 U35 ( .A(n208), .B(n5), .Q(o_data_AluRes[30]) );
  CLKIN0 U37 ( .A(n14), .Q(n15) );
  NAND31 U38 ( .A(n207), .B(n205), .C(n206), .Q(n4) );
  INV3 U39 ( .A(n4), .Q(n5) );
  AOI220 U40 ( .A(n214), .B(n30), .C(pre_sum_4a[6]), .D(n104), .Q(n205) );
  NAND20 U41 ( .A(pre_sum_4b[6]), .B(n201), .Q(n206) );
  CLKIN3 U42 ( .A(n199), .Q(n107) );
  AOI220 U43 ( .A(i_data_B[29]), .B(n229), .C(pre_suba[13]), .D(n69), .Q(n224)
         );
  NAND20 U44 ( .A(pre_sum_4b[5]), .B(n3), .Q(n223) );
  AOI220 U45 ( .A(i_data_B[28]), .B(n239), .C(pre_suba[12]), .D(n202), .Q(n234) );
  NAND20 U47 ( .A(pre_sum_4b[4]), .B(n3), .Q(n233) );
  BUF12 U48 ( .A(i_data_B[17]), .Q(n13) );
  AOI220 U49 ( .A(pre_sum_2b[7]), .B(n140), .C(i_data_B[15]), .D(n379), .Q(
        n376) );
  AOI220 U50 ( .A(i_data_B[27]), .B(n249), .C(pre_suba[11]), .D(n69), .Q(n244)
         );
  NAND20 U51 ( .A(pre_sum_4b[3]), .B(n3), .Q(n243) );
  AOI220 U52 ( .A(pre_sum_2b[3]), .B(n140), .C(i_data_B[11]), .D(n407), .Q(
        n404) );
  AOI220 U53 ( .A(pre_sum_2b[4]), .B(n140), .C(i_data_B[12]), .D(n400), .Q(
        n397) );
  AOI220 U55 ( .A(pre_sum_2b[5]), .B(n140), .C(i_data_B[13]), .D(n393), .Q(
        n390) );
  AOI220 U56 ( .A(pre_sum_2b[6]), .B(n140), .C(i_data_B[14]), .D(n386), .Q(
        n383) );
  INV0 U57 ( .A(i_data_B[5]), .Q(n424) );
  AOI222 U58 ( .A(pre_subb[14]), .B(n107), .C(N255), .D(n8), .Q(n211) );
  CLKIN1 U59 ( .A(n284), .Q(n105) );
  NOR20 U60 ( .A(n78), .B(n284), .Q(n294) );
  CLKIN3 U61 ( .A(n283), .Q(n104) );
  NAND20 U63 ( .A(n281), .B(n100), .Q(n283) );
  NAND20 U64 ( .A(pre_sum_3b[6]), .B(n294), .Q(n298) );
  NAND20 U65 ( .A(pre_sum_4b[0]), .B(n3), .Q(n273) );
  NAND20 U66 ( .A(pre_sum_4b[1]), .B(n3), .Q(n263) );
  NAND20 U67 ( .A(pre_sum_4b[2]), .B(n3), .Q(n253) );
  NAND20 U68 ( .A(pre_sum_3b[0]), .B(n294), .Q(n365) );
  NAND20 U69 ( .A(pre_sum_3b[1]), .B(n294), .Q(n355) );
  NAND20 U71 ( .A(pre_sum_3b[2]), .B(n294), .Q(n345) );
  NAND20 U72 ( .A(pre_sum_3b[3]), .B(n294), .Q(n335) );
  NAND20 U73 ( .A(pre_sum_3b[4]), .B(n294), .Q(n318) );
  NAND20 U74 ( .A(pre_sum_3b[7]), .B(n294), .Q(n286) );
  AOI220 U75 ( .A(N201), .B(n99), .C(n31), .D(n71), .Q(n148) );
  AOI220 U76 ( .A(n282), .B(n24), .C(pre_sum_4a[0]), .D(n104), .Q(n272) );
  AOI220 U77 ( .A(n271), .B(n25), .C(pre_sum_4a[1]), .D(n104), .Q(n262) );
  AOI220 U79 ( .A(n261), .B(n26), .C(pre_sum_4a[2]), .D(n104), .Q(n252) );
  AOI220 U80 ( .A(n251), .B(n27), .C(pre_sum_4a[3]), .D(n104), .Q(n242) );
  AOI220 U81 ( .A(n241), .B(n28), .C(pre_sum_4a[4]), .D(n104), .Q(n232) );
  AOI220 U82 ( .A(n231), .B(n29), .C(pre_sum_4a[5]), .D(n104), .Q(n222) );
  OAI2110 U83 ( .A(n2), .B(n439), .C(n438), .D(n362), .Q(n361) );
  NAND20 U84 ( .A(n2), .B(n143), .Q(n362) );
  OAI2110 U86 ( .A(n44), .B(n439), .C(n438), .D(n352), .Q(n351) );
  NAND20 U88 ( .A(n44), .B(n143), .Q(n352) );
  OAI2110 U89 ( .A(n46), .B(n439), .C(n438), .D(n342), .Q(n341) );
  NAND20 U90 ( .A(n47), .B(n143), .Q(n342) );
  OAI2110 U91 ( .A(n40), .B(n439), .C(n438), .D(n372), .Q(n371) );
  NAND20 U92 ( .A(n40), .B(n67), .Q(n372) );
  INV2 U93 ( .A(n32), .Q(n417) );
  INV0 U94 ( .A(n31), .Q(n419) );
  INV0 U96 ( .A(n40), .Q(n127) );
  INV0 U97 ( .A(n2), .Q(n125) );
  INV0 U98 ( .A(n44), .Q(n123) );
  INV0 U99 ( .A(n47), .Q(n121) );
  AOI220 U100 ( .A(pre_sum_2b[0]), .B(n140), .C(i_data_B[8]), .D(n153), .Q(
        n150) );
  OAI2110 U101 ( .A(n31), .B(n439), .C(n70), .D(n154), .Q(n153) );
  NAND20 U103 ( .A(n31), .B(n67), .Q(n154) );
  AOI220 U104 ( .A(pre_sum_2b[1]), .B(n140), .C(i_data_B[9]), .D(n141), .Q(
        n135) );
  OAI2110 U105 ( .A(i_data_A[9]), .B(n439), .C(n70), .D(n142), .Q(n141) );
  NAND20 U106 ( .A(n67), .B(i_data_A[9]), .Q(n142) );
  AOI220 U108 ( .A(pre_sum_2b[2]), .B(n140), .C(i_data_B[10]), .D(n414), .Q(
        n411) );
  AOI220 U109 ( .A(N193), .B(n99), .C(i_data_A[0]), .D(n71), .Q(n96) );
  NAND20 U110 ( .A(i_data_A[7]), .B(n71), .Q(n156) );
  NAND20 U111 ( .A(i_data_A[3]), .B(n71), .Q(n185) );
  AOI220 U112 ( .A(n188), .B(n431), .C(i_data_B[3]), .D(n189), .Q(n187) );
  NAND20 U113 ( .A(i_data_A[4]), .B(n71), .Q(n178) );
  AOI220 U115 ( .A(n181), .B(n427), .C(i_data_B[4]), .D(n182), .Q(n180) );
  NAND20 U116 ( .A(i_data_A[6]), .B(n71), .Q(n164) );
  NAND20 U117 ( .A(i_data_A[5]), .B(n71), .Q(n171) );
  NAND20 U118 ( .A(i_data_A[2]), .B(n71), .Q(n216) );
  AOI220 U119 ( .A(n219), .B(n433), .C(i_data_B[2]), .D(n220), .Q(n218) );
  NAND20 U120 ( .A(i_data_A[1]), .B(n71), .Q(n328) );
  AOI220 U122 ( .A(n331), .B(n435), .C(i_data_B[1]), .D(n332), .Q(n330) );
  INV0 U123 ( .A(n17), .Q(n18) );
  OAI2110 U124 ( .A(i_data_A[1]), .B(n439), .C(n438), .D(n333), .Q(n332) );
  NAND20 U126 ( .A(i_data_A[1]), .B(n67), .Q(n333) );
  OAI2110 U127 ( .A(i_data_A[2]), .B(n72), .C(n70), .D(n221), .Q(n220) );
  NAND20 U128 ( .A(i_data_A[2]), .B(n67), .Q(n221) );
  OAI2110 U129 ( .A(i_data_A[3]), .B(n72), .C(n70), .D(n190), .Q(n189) );
  NAND20 U130 ( .A(i_data_A[3]), .B(n67), .Q(n190) );
  OAI2110 U131 ( .A(i_data_A[4]), .B(n72), .C(n70), .D(n183), .Q(n182) );
  NAND20 U133 ( .A(i_data_A[4]), .B(n67), .Q(n183) );
  OAI2110 U134 ( .A(i_data_A[5]), .B(n439), .C(n70), .D(n176), .Q(n175) );
  NAND20 U135 ( .A(i_data_A[5]), .B(n67), .Q(n176) );
  OAI2110 U137 ( .A(i_data_A[6]), .B(n439), .C(n70), .D(n169), .Q(n168) );
  NAND20 U138 ( .A(i_data_A[6]), .B(n67), .Q(n169) );
  OAI2110 U139 ( .A(i_data_A[7]), .B(n439), .C(n70), .D(n161), .Q(n160) );
  NAND20 U140 ( .A(i_data_A[7]), .B(n67), .Q(n161) );
  OAI2110 U141 ( .A(i_data_A[0]), .B(n439), .C(n428), .D(n70), .Q(n93) );
  NAND20 U142 ( .A(i_data_A[0]), .B(n143), .Q(n428) );
  INV0 U144 ( .A(i_data_A[1]), .Q(n436) );
  INV0 U145 ( .A(i_data_A[2]), .Q(n434) );
  INV0 U146 ( .A(i_data_A[3]), .Q(n432) );
  INV0 U148 ( .A(i_data_A[4]), .Q(n430) );
  INV0 U149 ( .A(i_data_A[5]), .Q(n425) );
  INV0 U150 ( .A(i_data_A[6]), .Q(n423) );
  INV0 U151 ( .A(i_data_A[7]), .Q(n421) );
  INV0 U152 ( .A(i_data_B[2]), .Q(n433) );
  INV0 U153 ( .A(i_data_B[1]), .Q(n435) );
  INV0 U155 ( .A(i_data_B[8]), .Q(n418) );
  INV0 U156 ( .A(i_data_B[9]), .Q(n416) );
  INV0 U157 ( .A(i_data_B[10]), .Q(n162) );
  INV0 U159 ( .A(i_data_B[3]), .Q(n431) );
  INV0 U160 ( .A(i_data_B[4]), .Q(n427) );
  INV0 U161 ( .A(i_data_B[0]), .Q(n437) );
  NOR21 U162 ( .A(n105), .B(n78), .Q(n296) );
  AOI221 U163 ( .A(pre_sum_3a[8]), .B(n284), .C(pre_sum_3b[8]), .D(n105), .Q(
        n281) );
  NAND22 U164 ( .A(half_sub[16]), .B(n101), .Q(n199) );
  INV3 U166 ( .A(n202), .Q(n68) );
  INV3 U167 ( .A(n71), .Q(n70) );
  NOR21 U168 ( .A(n70), .B(n127), .Q(n369) );
  NOR21 U170 ( .A(n70), .B(n125), .Q(n359) );
  NOR21 U171 ( .A(n70), .B(n123), .Q(n349) );
  NOR21 U172 ( .A(n70), .B(n119), .Q(n312) );
  NOR21 U173 ( .A(n70), .B(n118), .Q(n302) );
  NOR21 U174 ( .A(n70), .B(n117), .Q(n290) );
  NOR21 U175 ( .A(n70), .B(n116), .Q(n277) );
  NOR21 U176 ( .A(n70), .B(n115), .Q(n267) );
  NOR21 U177 ( .A(n70), .B(n114), .Q(n257) );
  NOR21 U178 ( .A(n70), .B(n113), .Q(n247) );
  NOR21 U179 ( .A(n70), .B(n112), .Q(n237) );
  NOR21 U180 ( .A(n70), .B(n111), .Q(n227) );
  NOR21 U181 ( .A(n70), .B(n121), .Q(n339) );
  NOR21 U182 ( .A(n70), .B(n120), .Q(n322) );
  INV3 U184 ( .A(n75), .Q(n74) );
  INV3 U185 ( .A(n73), .Q(n72) );
  BUF2 U186 ( .A(n98), .Q(n10) );
  BUF2 U187 ( .A(n98), .Q(n9) );
  BUF2 U188 ( .A(n98), .Q(n8) );
  NAND22 U189 ( .A(i_data_B[15]), .B(n203), .Q(n192) );
  AOI221 U191 ( .A(N256), .B(n9), .C(n73), .D(n1), .Q(n191) );
  AOI221 U192 ( .A(N224), .B(n99), .C(n66), .D(n71), .Q(n193) );
  NAND41 U193 ( .A(n364), .B(n365), .C(n366), .D(n367), .Q(o_data_AluRes[16])
         );
  AOI2111 U195 ( .A(N209), .B(n99), .C(n368), .D(n369), .Q(n367) );
  NAND41 U196 ( .A(n354), .B(n355), .C(n356), .D(n357), .Q(o_data_AluRes[17])
         );
  AOI221 U197 ( .A(i_data_B[17]), .B(n361), .C(pre_suba[1]), .D(n69), .Q(n356)
         );
  AOI2111 U198 ( .A(N210), .B(n99), .C(n358), .D(n359), .Q(n357) );
  NAND41 U199 ( .A(n344), .B(n345), .C(n346), .D(n347), .Q(o_data_AluRes[18])
         );
  AOI221 U200 ( .A(n16), .B(n351), .C(pre_suba[2]), .D(n202), .Q(n346) );
  AOI2111 U202 ( .A(N211), .B(n99), .C(n348), .D(n349), .Q(n347) );
  NAND41 U203 ( .A(n334), .B(n335), .C(n336), .D(n337), .Q(o_data_AluRes[19])
         );
  AOI221 U204 ( .A(i_data_B[19]), .B(n341), .C(pre_suba[3]), .D(n69), .Q(n336)
         );
  AOI2111 U206 ( .A(N212), .B(n99), .C(n338), .D(n339), .Q(n337) );
  NAND41 U207 ( .A(n317), .B(n318), .C(n319), .D(n320), .Q(o_data_AluRes[20])
         );
  AOI2111 U208 ( .A(N213), .B(n99), .C(n321), .D(n322), .Q(n320) );
  NAND41 U209 ( .A(n307), .B(n308), .C(n309), .D(n310), .Q(o_data_AluRes[21])
         );
  AOI2111 U210 ( .A(N214), .B(n99), .C(n311), .D(n312), .Q(n310) );
  NAND22 U211 ( .A(pre_sum_3b[5]), .B(n294), .Q(n308) );
  NAND41 U213 ( .A(n297), .B(n298), .C(n299), .D(n300), .Q(o_data_AluRes[22])
         );
  AOI221 U214 ( .A(i_data_B[22]), .B(n304), .C(pre_suba[6]), .D(n202), .Q(n299) );
  AOI2111 U215 ( .A(N215), .B(n99), .C(n301), .D(n302), .Q(n300) );
  NAND41 U217 ( .A(n285), .B(n286), .C(n287), .D(n288), .Q(o_data_AluRes[23])
         );
  AOI221 U218 ( .A(i_data_B[23]), .B(n292), .C(pre_suba[7]), .D(n69), .Q(n287)
         );
  AOI2111 U219 ( .A(N216), .B(n99), .C(n289), .D(n290), .Q(n288) );
  NAND41 U220 ( .A(n272), .B(n273), .C(n274), .D(n275), .Q(o_data_AluRes[24])
         );
  AOI221 U221 ( .A(i_data_B[24]), .B(n279), .C(pre_suba[8]), .D(n202), .Q(n274) );
  AOI2111 U222 ( .A(N217), .B(n99), .C(n276), .D(n277), .Q(n275) );
  NAND41 U224 ( .A(n262), .B(n263), .C(n264), .D(n265), .Q(o_data_AluRes[25])
         );
  AOI221 U225 ( .A(i_data_B[25]), .B(n269), .C(pre_suba[9]), .D(n69), .Q(n264)
         );
  AOI2111 U226 ( .A(N218), .B(n99), .C(n266), .D(n267), .Q(n265) );
  NAND41 U227 ( .A(n252), .B(n253), .C(n254), .D(n255), .Q(o_data_AluRes[26])
         );
  AOI221 U229 ( .A(i_data_B[26]), .B(n259), .C(pre_suba[10]), .D(n202), .Q(
        n254) );
  AOI2111 U230 ( .A(N219), .B(n99), .C(n256), .D(n257), .Q(n255) );
  NAND41 U231 ( .A(n242), .B(n243), .C(n244), .D(n245), .Q(o_data_AluRes[27])
         );
  AOI2111 U232 ( .A(N220), .B(n99), .C(n246), .D(n247), .Q(n245) );
  NAND41 U233 ( .A(n232), .B(n233), .C(n234), .D(n235), .Q(o_data_AluRes[28])
         );
  AOI2111 U234 ( .A(N221), .B(n99), .C(n236), .D(n237), .Q(n235) );
  NAND41 U236 ( .A(n222), .B(n223), .C(n224), .D(n225), .Q(o_data_AluRes[29])
         );
  AOI2111 U237 ( .A(N222), .B(n99), .C(n226), .D(n227), .Q(n225) );
  AOI221 U238 ( .A(n373), .B(n126), .C(pre_sum_3a[0]), .D(n296), .Q(n364) );
  AOI221 U239 ( .A(n363), .B(n124), .C(pre_sum_3a[1]), .D(n296), .Q(n354) );
  INV3 U240 ( .A(i_data_B[17]), .Q(n124) );
  AOI221 U241 ( .A(n353), .B(n122), .C(pre_sum_3a[2]), .D(n296), .Q(n344) );
  INV3 U243 ( .A(n16), .Q(n122) );
  AOI221 U244 ( .A(n343), .B(n17), .C(pre_sum_3a[3]), .D(n296), .Q(n334) );
  AOI221 U245 ( .A(n326), .B(n19), .C(pre_sum_3a[4]), .D(n296), .Q(n317) );
  AOI221 U247 ( .A(n316), .B(n20), .C(pre_sum_3a[5]), .D(n296), .Q(n307) );
  AOI221 U248 ( .A(n306), .B(n21), .C(pre_sum_3a[6]), .D(n296), .Q(n297) );
  AOI221 U249 ( .A(n295), .B(n23), .C(pre_sum_3a[7]), .D(n296), .Q(n285) );
  AOI221 U250 ( .A(pre_subb[12]), .B(n107), .C(N253), .D(n8), .Q(n238) );
  AOI221 U251 ( .A(pre_subb[13]), .B(n107), .C(N254), .D(n8), .Q(n228) );
  OAI311 U252 ( .A(n139), .B(i_data_B[31]), .C(n66), .D(n197), .Q(n196) );
  AOI221 U254 ( .A(pre_sum_4b[7]), .B(n3), .C(pre_suba[15]), .D(n69), .Q(n200)
         );
  NOR21 U255 ( .A(n78), .B(sum_1[8]), .Q(n138) );
  NAND41 U256 ( .A(n148), .B(n149), .C(n150), .D(n151), .Q(o_data_AluRes[8])
         );
  AOI221 U258 ( .A(N233), .B(n9), .C(half_sub[8]), .D(n101), .Q(n149) );
  AOI221 U259 ( .A(n152), .B(n418), .C(pre_sum_2a[0]), .D(n138), .Q(n151) );
  NAND41 U260 ( .A(n133), .B(n134), .C(n135), .D(n136), .Q(o_data_AluRes[9])
         );
  AOI221 U261 ( .A(N202), .B(n99), .C(n71), .D(i_data_A[9]), .Q(n133) );
  AOI221 U262 ( .A(N234), .B(n10), .C(half_sub[9]), .D(n101), .Q(n134) );
  AOI221 U263 ( .A(n137), .B(n416), .C(pre_sum_2a[1]), .D(n138), .Q(n136) );
  NAND41 U265 ( .A(n409), .B(n410), .C(n411), .D(n412), .Q(o_data_AluRes[10])
         );
  AOI221 U266 ( .A(N203), .B(n99), .C(i_data_A[10]), .D(n71), .Q(n409) );
  AOI221 U267 ( .A(N235), .B(n9), .C(half_sub[10]), .D(n101), .Q(n410) );
  AOI221 U269 ( .A(n413), .B(n162), .C(pre_sum_2a[2]), .D(n138), .Q(n412) );
  NAND41 U270 ( .A(n402), .B(n403), .C(n404), .D(n405), .Q(o_data_AluRes[11])
         );
  AOI221 U271 ( .A(N204), .B(n99), .C(n34), .D(n71), .Q(n402) );
  AOI221 U272 ( .A(N236), .B(n10), .C(half_sub[11]), .D(n101), .Q(n403) );
  AOI221 U273 ( .A(n406), .B(n146), .C(pre_sum_2a[3]), .D(n138), .Q(n405) );
  NAND41 U274 ( .A(n395), .B(n396), .C(n397), .D(n398), .Q(o_data_AluRes[12])
         );
  AOI221 U275 ( .A(N237), .B(n9), .C(half_sub[12]), .D(n101), .Q(n396) );
  AOI221 U276 ( .A(N205), .B(n99), .C(n35), .D(n71), .Q(n395) );
  AOI221 U277 ( .A(n399), .B(n144), .C(pre_sum_2a[4]), .D(n138), .Q(n398) );
  NAND41 U278 ( .A(n388), .B(n389), .C(n390), .D(n391), .Q(o_data_AluRes[13])
         );
  AOI221 U279 ( .A(N206), .B(n99), .C(i_data_A[13]), .D(n71), .Q(n388) );
  AOI221 U280 ( .A(N238), .B(n10), .C(half_sub[13]), .D(n101), .Q(n389) );
  AOI221 U282 ( .A(n392), .B(n131), .C(pre_sum_2a[5]), .D(n138), .Q(n391) );
  NAND41 U283 ( .A(n381), .B(n382), .C(n383), .D(n384), .Q(o_data_AluRes[14])
         );
  AOI221 U285 ( .A(N207), .B(n99), .C(n38), .D(n71), .Q(n381) );
  AOI221 U286 ( .A(N239), .B(n9), .C(half_sub[14]), .D(n101), .Q(n382) );
  AOI221 U287 ( .A(n385), .B(n129), .C(pre_sum_2a[6]), .D(n138), .Q(n384) );
  NAND41 U288 ( .A(n374), .B(n375), .C(n376), .D(n377), .Q(o_data_AluRes[15])
         );
  AOI221 U289 ( .A(N208), .B(n99), .C(i_data_A[15]), .D(n71), .Q(n374) );
  AOI221 U290 ( .A(N240), .B(n10), .C(half_sub[15]), .D(n101), .Q(n375) );
  AOI221 U291 ( .A(n378), .B(n11), .C(pre_sum_2a[7]), .D(n138), .Q(n377) );
  AOI221 U293 ( .A(pre_subb[3]), .B(n107), .C(N244), .D(n9), .Q(n340) );
  AOI221 U294 ( .A(pre_subb[4]), .B(n107), .C(N245), .D(n10), .Q(n323) );
  AOI221 U295 ( .A(pre_subb[5]), .B(n107), .C(N246), .D(n8), .Q(n313) );
  AOI221 U296 ( .A(pre_subb[6]), .B(n107), .C(N247), .D(n8), .Q(n303) );
  AOI221 U297 ( .A(pre_subb[7]), .B(n107), .C(N248), .D(n8), .Q(n291) );
  AOI221 U298 ( .A(pre_subb[8]), .B(n107), .C(N249), .D(n8), .Q(n278) );
  AOI221 U299 ( .A(pre_subb[9]), .B(n107), .C(N250), .D(n8), .Q(n268) );
  AOI221 U301 ( .A(pre_subb[1]), .B(n107), .C(N242), .D(n9), .Q(n360) );
  AOI221 U302 ( .A(pre_subb[2]), .B(n107), .C(N243), .D(n10), .Q(n350) );
  AOI221 U303 ( .A(pre_subb[10]), .B(n107), .C(N251), .D(n8), .Q(n258) );
  AOI221 U304 ( .A(pre_subb[11]), .B(n107), .C(N252), .D(n8), .Q(n248) );
  OAI2111 U305 ( .A(i_data_A[15]), .B(n72), .C(n438), .D(n380), .Q(n379) );
  NAND22 U306 ( .A(i_data_A[15]), .B(n143), .Q(n380) );
  OAI2111 U307 ( .A(n48), .B(n439), .C(n438), .D(n325), .Q(n324) );
  NAND22 U309 ( .A(n48), .B(n143), .Q(n325) );
  OAI2111 U310 ( .A(i_data_A[21]), .B(n439), .C(n70), .D(n315), .Q(n314) );
  NAND22 U311 ( .A(n49), .B(n143), .Q(n315) );
  OAI2111 U312 ( .A(n50), .B(n439), .C(n70), .D(n305), .Q(n304) );
  NAND22 U313 ( .A(n51), .B(n143), .Q(n305) );
  OAI2111 U314 ( .A(i_data_A[23]), .B(n72), .C(n438), .D(n293), .Q(n292) );
  NAND22 U315 ( .A(n52), .B(n143), .Q(n293) );
  OAI2111 U317 ( .A(n55), .B(n439), .C(n70), .D(n270), .Q(n269) );
  NAND22 U318 ( .A(n55), .B(n67), .Q(n270) );
  OAI2111 U319 ( .A(n57), .B(n72), .C(n70), .D(n260), .Q(n259) );
  NAND22 U320 ( .A(n57), .B(n67), .Q(n260) );
  OAI2111 U321 ( .A(n59), .B(n72), .C(n438), .D(n250), .Q(n249) );
  NAND22 U322 ( .A(n59), .B(n67), .Q(n250) );
  OAI2111 U323 ( .A(n61), .B(n72), .C(n438), .D(n240), .Q(n239) );
  NAND22 U324 ( .A(n61), .B(n67), .Q(n240) );
  OAI2111 U326 ( .A(i_data_A[29]), .B(n72), .C(n438), .D(n230), .Q(n229) );
  NAND22 U327 ( .A(i_data_A[29]), .B(n67), .Q(n230) );
  OAI2111 U328 ( .A(n64), .B(n439), .C(n438), .D(n213), .Q(n212) );
  NAND22 U329 ( .A(n64), .B(n67), .Q(n213) );
  INV3 U330 ( .A(n438), .Q(n71) );
  NAND22 U331 ( .A(n102), .B(n103), .Q(n429) );
  INV3 U332 ( .A(n77), .Q(n101) );
  INV3 U333 ( .A(n139), .Q(n75) );
  BUF2 U334 ( .A(n143), .Q(n67) );
  INV3 U335 ( .A(n203), .Q(n440) );
  INV3 U336 ( .A(n34), .Q(n147) );
  INV3 U337 ( .A(n35), .Q(n145) );
  INV3 U338 ( .A(i_data_A[13]), .Q(n132) );
  INV3 U339 ( .A(n38), .Q(n130) );
  INV3 U340 ( .A(i_data_A[15]), .Q(n128) );
  INV3 U341 ( .A(i_data_A[10]), .Q(n204) );
  INV3 U342 ( .A(n198), .Q(n109) );
  NAND22 U343 ( .A(n67), .B(n66), .Q(n198) );
  INV3 U344 ( .A(n439), .Q(n73) );
  INV3 U345 ( .A(n92), .Q(n98) );
  INV3 U346 ( .A(n48), .Q(n120) );
  INV3 U347 ( .A(n57), .Q(n114) );
  INV3 U348 ( .A(n59), .Q(n113) );
  INV3 U349 ( .A(n61), .Q(n112) );
  INV3 U350 ( .A(n49), .Q(n119) );
  INV3 U351 ( .A(n55), .Q(n115) );
  INV3 U352 ( .A(n64), .Q(n110) );
  INV3 U353 ( .A(n51), .Q(n118) );
  INV3 U354 ( .A(n52), .Q(n117) );
  NOR21 U355 ( .A(n70), .B(n110), .Q(n210) );
  BUF2 U356 ( .A(i_data_A[18]), .Q(n44) );
  NAND41 U357 ( .A(n97), .B(n96), .C(n95), .D(n94), .Q(o_data_AluRes[0]) );
  IMUX30 U358 ( .A(n75), .B(n73), .C(n93), .S0(i_data_A[0]), .S1(i_data_B[0]), 
        .Q(n94) );
  AOI221 U359 ( .A(N225), .B(n9), .C(half_sub[0]), .D(n101), .Q(n95) );
  AOI221 U360 ( .A(i_con_AluCtrl[0]), .B(n89), .C(sum_1[0]), .D(n100), .Q(n97)
         );
  NAND41 U361 ( .A(n163), .B(n164), .C(n165), .D(n166), .Q(o_data_AluRes[6])
         );
  AOI221 U362 ( .A(n167), .B(n422), .C(i_data_B[6]), .D(n168), .Q(n166) );
  AOI221 U363 ( .A(N231), .B(n9), .C(half_sub[6]), .D(n101), .Q(n165) );
  NAND41 U364 ( .A(n155), .B(n156), .C(n157), .D(n158), .Q(o_data_AluRes[7])
         );
  AOI221 U365 ( .A(n159), .B(n420), .C(i_data_B[7]), .D(n160), .Q(n158) );
  AOI221 U366 ( .A(N232), .B(n10), .C(half_sub[7]), .D(n101), .Q(n157) );
  AOI221 U367 ( .A(N199), .B(n99), .C(sum_1[6]), .D(n100), .Q(n163) );
  AOI221 U368 ( .A(N200), .B(n99), .C(sum_1[7]), .D(n100), .Q(n155) );
  AOI221 U369 ( .A(pre_subb[0]), .B(n107), .C(N241), .D(n10), .Q(n370) );
  OAI2111 U370 ( .A(i_data_A[10]), .B(n72), .C(n438), .D(n415), .Q(n414) );
  NAND22 U371 ( .A(i_data_A[10]), .B(n143), .Q(n415) );
  OAI2111 U372 ( .A(n34), .B(n72), .C(n70), .D(n408), .Q(n407) );
  NAND22 U373 ( .A(n34), .B(n143), .Q(n408) );
  OAI2111 U374 ( .A(n35), .B(n72), .C(n438), .D(n401), .Q(n400) );
  NAND22 U375 ( .A(n35), .B(n143), .Q(n401) );
  OAI2111 U376 ( .A(i_data_A[13]), .B(n72), .C(n438), .D(n394), .Q(n393) );
  NAND22 U377 ( .A(i_data_A[13]), .B(n143), .Q(n394) );
  OAI2111 U378 ( .A(n38), .B(n72), .C(n438), .D(n387), .Q(n386) );
  NAND22 U379 ( .A(n38), .B(n143), .Q(n387) );
  BUF2 U380 ( .A(i_data_A[21]), .Q(n49) );
  BUF2 U381 ( .A(i_data_A[19]), .Q(n46) );
  INV3 U382 ( .A(n21), .Q(n22) );
  BUF2 U383 ( .A(i_data_A[9]), .Q(n32) );
  BUF2 U384 ( .A(i_data_A[10]), .Q(n33) );
  BUF2 U385 ( .A(i_data_A[19]), .Q(n47) );
  AOI221 U386 ( .A(N194), .B(n99), .C(sum_1[1]), .D(n100), .Q(n327) );
  AOI221 U387 ( .A(N195), .B(n99), .C(sum_1[2]), .D(n100), .Q(n215) );
  AOI221 U388 ( .A(N197), .B(n99), .C(sum_1[4]), .D(n100), .Q(n177) );
  NAND41 U389 ( .A(n327), .B(n328), .C(n329), .D(n330), .Q(o_data_AluRes[1])
         );
  AOI221 U390 ( .A(N226), .B(n9), .C(half_sub[1]), .D(n101), .Q(n329) );
  NAND41 U391 ( .A(n215), .B(n216), .C(n217), .D(n218), .Q(o_data_AluRes[2])
         );
  AOI221 U392 ( .A(N227), .B(n10), .C(half_sub[2]), .D(n101), .Q(n217) );
  NAND41 U393 ( .A(n184), .B(n185), .C(n186), .D(n187), .Q(o_data_AluRes[3])
         );
  AOI221 U394 ( .A(N196), .B(n99), .C(sum_1[3]), .D(n100), .Q(n184) );
  NAND41 U395 ( .A(n177), .B(n178), .C(n179), .D(n180), .Q(o_data_AluRes[4])
         );
  AOI221 U396 ( .A(N229), .B(n9), .C(half_sub[4]), .D(n101), .Q(n179) );
  NAND41 U397 ( .A(n170), .B(n171), .C(n172), .D(n173), .Q(o_data_AluRes[5])
         );
  AOI221 U398 ( .A(n174), .B(n424), .C(i_data_B[5]), .D(n175), .Q(n173) );
  AOI221 U399 ( .A(N230), .B(n10), .C(half_sub[5]), .D(n101), .Q(n172) );
  AOI221 U400 ( .A(N228), .B(n10), .C(half_sub[3]), .D(n101), .Q(n186) );
  AOI221 U401 ( .A(N198), .B(n99), .C(sum_1[5]), .D(n100), .Q(n170) );
  IMUX21 U402 ( .A(n87), .B(n82), .S(n1), .Q(n84) );
  BUF2 U403 ( .A(i_data_A[11]), .Q(n34) );
  BUF2 U404 ( .A(i_data_A[12]), .Q(n35) );
  BUF2 U405 ( .A(i_data_A[25]), .Q(n54) );
  BUF2 U406 ( .A(i_data_A[16]), .Q(n40) );
  BUF2 U407 ( .A(i_data_A[24]), .Q(n53) );
  BUF2 U408 ( .A(i_data_A[22]), .Q(n50) );
  BUF2 U409 ( .A(i_data_A[13]), .Q(n36) );
  BUF2 U410 ( .A(i_data_A[22]), .Q(n51) );
  BUF2 U411 ( .A(i_data_A[23]), .Q(n52) );
  INV3 U412 ( .A(n78), .Q(n100) );
  NAND31 U413 ( .A(i_con_AluCtrl[1]), .B(n80), .C(n90), .Q(n78) );
  BUF2 U414 ( .A(i_data_A[8]), .Q(n31) );
  BUF2 U415 ( .A(i_data_A[26]), .Q(n57) );
  BUF2 U416 ( .A(i_data_A[27]), .Q(n59) );
  BUF2 U417 ( .A(i_data_A[15]), .Q(n39) );
  BUF2 U418 ( .A(i_data_A[14]), .Q(n38) );
  BUF2 U419 ( .A(i_data_A[14]), .Q(n37) );
  BUF2 U420 ( .A(i_data_A[26]), .Q(n56) );
  BUF2 U421 ( .A(i_data_A[27]), .Q(n58) );
  BUF2 U422 ( .A(i_data_A[25]), .Q(n55) );
  NOR40 U423 ( .A(n102), .B(i_con_AluCtrl[0]), .C(i_con_AluCtrl[1]), .D(
        i_con_AluCtrl[2]), .Q(n203) );
  NAND31 U424 ( .A(i_con_AluCtrl[1]), .B(i_con_AluCtrl[2]), .C(n102), .Q(n88)
         );
  NAND31 U425 ( .A(i_con_AluCtrl[0]), .B(i_con_AluCtrl[1]), .C(n90), .Q(n91)
         );
  NOR21 U426 ( .A(n429), .B(i_con_AluCtrl[1]), .Q(n143) );
  NOR21 U427 ( .A(n103), .B(i_con_AluCtrl[1]), .Q(n426) );
  INV3 U428 ( .A(i_data_B[11]), .Q(n146) );
  BUF2 U429 ( .A(i_data_A[31]), .Q(n66) );
  INV3 U430 ( .A(i_data_B[12]), .Q(n144) );
  INV3 U431 ( .A(i_data_B[7]), .Q(n420) );
  INV3 U432 ( .A(i_data_B[14]), .Q(n129) );
  INV3 U433 ( .A(i_data_B[13]), .Q(n131) );
  BUF2 U434 ( .A(i_data_A[28]), .Q(n61) );
  BUF2 U435 ( .A(i_data_A[30]), .Q(n63) );
  INV3 U436 ( .A(i_data_B[6]), .Q(n422) );
  BUF2 U437 ( .A(i_data_A[31]), .Q(n65) );
  BUF2 U438 ( .A(i_data_A[29]), .Q(n62) );
  BUF2 U439 ( .A(i_data_A[28]), .Q(n60) );
  BUF2 U440 ( .A(i_data_A[30]), .Q(n64) );
  INV3 U441 ( .A(i_data_B[18]), .Q(n14) );
  INV3 U442 ( .A(i_data_B[19]), .Q(n17) );
  INV3 U443 ( .A(i_data_B[22]), .Q(n21) );
  INV3 U444 ( .A(i_data_B[28]), .Q(n28) );
  INV3 U445 ( .A(i_data_B[27]), .Q(n27) );
  INV3 U446 ( .A(i_data_B[26]), .Q(n26) );
  INV3 U447 ( .A(i_data_B[25]), .Q(n25) );
  INV3 U448 ( .A(i_data_B[29]), .Q(n29) );
  INV3 U449 ( .A(i_data_B[30]), .Q(n30) );
  INV3 U450 ( .A(i_data_B[23]), .Q(n23) );
  INV3 U451 ( .A(i_data_B[24]), .Q(n24) );
  INV3 U452 ( .A(i_data_B[15]), .Q(n11) );
  LOGIC0 U453 ( .Q(n42) );
  LOGIC1 U454 ( .Q(n41) );
  INV0 U455 ( .A(n12), .Q(n126) );
  AOI220 U456 ( .A(n12), .B(n371), .C(pre_suba[0]), .D(n69), .Q(n366) );
  CLKIN3 U457 ( .A(i_con_AluCtrl[3]), .Q(n102) );
  CLKIN3 U458 ( .A(n88), .Q(n76) );
  CLKIN3 U459 ( .A(i_con_AluCtrl[0]), .Q(n80) );
  NAND22 U460 ( .A(n76), .B(n80), .Q(n77) );
  CLKIN3 U461 ( .A(n429), .Q(n90) );
  CLKIN3 U462 ( .A(i_con_AluCtrl[1]), .Q(n83) );
  NAND22 U463 ( .A(n426), .B(i_con_AluCtrl[3]), .Q(n79) );
  CLKIN3 U464 ( .A(n79), .Q(n81) );
  NAND22 U465 ( .A(n81), .B(n80), .Q(n139) );
  NAND22 U466 ( .A(n81), .B(i_con_AluCtrl[0]), .Q(n439) );
  CLKIN3 U467 ( .A(N306), .Q(n87) );
  CLKIN3 U468 ( .A(n66), .Q(n82) );
  NAND22 U469 ( .A(n84), .B(n83), .Q(n86) );
  CLKIN3 U470 ( .A(i_con_AluCtrl[2]), .Q(n103) );
  NAND22 U471 ( .A(i_con_AluCtrl[3]), .B(n103), .Q(n85) );
  OAI222 U472 ( .A(n88), .B(n87), .C(n86), .D(n85), .Q(n89) );
  CLKIN3 U473 ( .A(n91), .Q(n99) );
  NAND22 U474 ( .A(n426), .B(n102), .Q(n92) );
endmodule


module E_alu_control ( o_con_AluCtrl, i_con_AluOp, i_con_FuncCode );
  output [3:0] o_con_AluCtrl;
  input [5:0] i_con_AluOp;
  input [5:0] i_con_FuncCode;
  wire   n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;

  OAI212 U5 ( .A(n21), .B(n22), .C(n5), .Q(n18) );
  OAI212 U11 ( .A(n30), .B(n32), .C(n5), .Q(n31) );
  OAI222 U17 ( .A(n38), .B(n6), .C(i_con_AluOp[1]), .D(n6), .Q(n34) );
  OAI2111 U3 ( .A(n23), .B(n24), .C(n25), .D(n20), .Q(o_con_AluCtrl[2]) );
  NOR40 U4 ( .A(n8), .B(n26), .C(n12), .D(n22), .Q(n23) );
  INV3 U6 ( .A(n28), .Q(n12) );
  INV3 U7 ( .A(n29), .Q(n8) );
  OAI2111 U8 ( .A(n16), .B(n27), .C(n7), .D(n14), .Q(n22) );
  NAND31 U9 ( .A(n17), .B(n16), .C(n39), .Q(n41) );
  NOR21 U10 ( .A(n17), .B(n10), .Q(n26) );
  INV3 U12 ( .A(n42), .Q(n7) );
  NOR40 U13 ( .A(n21), .B(n30), .C(n26), .D(n43), .Q(n42) );
  NAND31 U14 ( .A(n41), .B(n27), .C(n28), .Q(n43) );
  NAND41 U15 ( .A(n41), .B(n9), .C(n7), .D(n14), .Q(n32) );
  INV3 U16 ( .A(n26), .Q(n9) );
  INV3 U18 ( .A(n24), .Q(n5) );
  NAND31 U19 ( .A(i_con_FuncCode[5]), .B(n15), .C(i_con_FuncCode[2]), .Q(n27)
         );
  NOR31 U20 ( .A(i_con_FuncCode[3]), .B(i_con_FuncCode[5]), .C(
        i_con_FuncCode[2]), .Q(n39) );
  NAND31 U21 ( .A(n18), .B(n19), .C(n20), .Q(o_con_AluCtrl[3]) );
  NAND31 U22 ( .A(i_con_AluOp[0]), .B(i_con_AluOp[3]), .C(i_con_AluOp[2]), .Q(
        n19) );
  NOR21 U23 ( .A(n10), .B(i_con_FuncCode[0]), .Q(n21) );
  NAND22 U24 ( .A(n39), .B(i_con_FuncCode[1]), .Q(n28) );
  INV3 U25 ( .A(i_con_FuncCode[1]), .Q(n16) );
  INV3 U26 ( .A(n45), .Q(n10) );
  NOR40 U27 ( .A(n11), .B(n15), .C(n16), .D(i_con_FuncCode[2]), .Q(n45) );
  INV3 U28 ( .A(i_con_FuncCode[5]), .Q(n11) );
  INV3 U29 ( .A(i_con_FuncCode[3]), .Q(n15) );
  OAI2111 U30 ( .A(n35), .B(n24), .C(n36), .D(n20), .Q(o_con_AluCtrl[0]) );
  NAND31 U31 ( .A(i_con_AluOp[3]), .B(n4), .C(i_con_AluOp[0]), .Q(n36) );
  AOI2111 U32 ( .A(n39), .B(i_con_FuncCode[0]), .C(n40), .D(n32), .Q(n35) );
  OAI311 U33 ( .A(n27), .B(i_con_FuncCode[1]), .C(n17), .D(n44), .Q(n40) );
  NAND41 U34 ( .A(n1), .B(i_con_AluOp[1]), .C(n2), .D(n31), .Q(
        o_con_AluCtrl[1]) );
  INV3 U35 ( .A(n33), .Q(n2) );
  INV3 U36 ( .A(n34), .Q(n1) );
  AOI211 U37 ( .A(n3), .B(i_con_AluOp[4]), .C(i_con_AluOp[5]), .Q(n38) );
  NOR31 U38 ( .A(i_con_FuncCode[2]), .B(i_con_FuncCode[3]), .C(n11), .Q(n30)
         );
  INV3 U39 ( .A(i_con_AluOp[0]), .Q(n6) );
  NOR21 U40 ( .A(n34), .B(n37), .Q(n20) );
  NOR40 U41 ( .A(n4), .B(n6), .C(n3), .D(i_con_AluOp[4]), .Q(n37) );
  AOI311 U42 ( .A(i_con_FuncCode[1]), .B(n17), .C(n13), .D(n21), .Q(n44) );
  INV3 U43 ( .A(n27), .Q(n13) );
  INV3 U44 ( .A(i_con_FuncCode[0]), .Q(n17) );
  NAND22 U45 ( .A(i_con_FuncCode[1]), .B(n30), .Q(n29) );
  INV3 U46 ( .A(i_con_AluOp[2]), .Q(n4) );
  INV3 U47 ( .A(i_con_AluOp[3]), .Q(n3) );
  INV3 U48 ( .A(i_con_FuncCode[4]), .Q(n14) );
  OAI311 U49 ( .A(i_con_AluOp[2]), .B(i_con_AluOp[3]), .C(n6), .D(n25), .Q(n33) );
  NAND31 U50 ( .A(i_con_AluOp[4]), .B(n4), .C(i_con_AluOp[0]), .Q(n25) );
  NAND22 U51 ( .A(i_con_AluOp[1]), .B(n6), .Q(n24) );
endmodule


module E_famux5 ( i_data_rs, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fa, o_data_alusra );
  input [31:0] i_data_rs;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fa;
  output [31:0] o_data_alusra;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV3 U1 ( .A(n13), .Q(n112) );
  INV3 U2 ( .A(i_con_fa[2]), .Q(n12) );
  INV3 U3 ( .A(i_con_fa[0]), .Q(n14) );
  AOI221 U4 ( .A(i_data_lwM[16]), .B(n114), .C(i_data_lwW[16]), .D(n9), .Q(n66) );
  AOI220 U5 ( .A(i_data_rs[16]), .B(n5), .C(i_data_writeres[16]), .D(n7), .Q(
        n68) );
  AOI221 U6 ( .A(i_data_lwM[7]), .B(n114), .C(i_data_lwW[7]), .D(n9), .Q(n39)
         );
  AOI221 U7 ( .A(i_data_rs[7]), .B(n4), .C(i_data_writeres[7]), .D(n6), .Q(n41) );
  NAND22 U8 ( .A(n14), .B(n2), .Q(n13) );
  NAND20 U9 ( .A(n12), .B(i_con_fa[1]), .Q(n1) );
  INV2 U10 ( .A(n1), .Q(n2) );
  NAND33 U11 ( .A(n68), .B(n67), .C(n66), .Q(o_data_alusra[16]) );
  NAND33 U12 ( .A(n71), .B(n70), .C(n69), .Q(o_data_alusra[17]) );
  AOI221 U13 ( .A(i_data_rs[17]), .B(n5), .C(i_data_writeres[17]), .D(n6), .Q(
        n71) );
  AOI220 U14 ( .A(i_data_lwM[0]), .B(n114), .C(i_data_lwW[0]), .D(n9), .Q(n18)
         );
  AOI220 U15 ( .A(i_data_rs[0]), .B(n4), .C(i_data_writeres[0]), .D(n6), .Q(
        n20) );
  AOI220 U16 ( .A(i_data_lwM[17]), .B(n114), .C(i_data_lwW[17]), .D(n8), .Q(
        n69) );
  AOI220 U17 ( .A(i_data_rs[23]), .B(n5), .C(i_data_writeres[23]), .D(n111), 
        .Q(n89) );
  AOI220 U18 ( .A(i_data_lwM[23]), .B(n114), .C(i_data_lwW[23]), .D(n8), .Q(
        n87) );
  AOI220 U19 ( .A(i_data_rs[12]), .B(n4), .C(i_data_writeres[12]), .D(n7), .Q(
        n56) );
  AOI220 U20 ( .A(i_data_lwM[12]), .B(n114), .C(i_data_lwW[12]), .D(n9), .Q(
        n54) );
  AOI220 U21 ( .A(i_data_rs[13]), .B(n4), .C(i_data_writeres[13]), .D(n111), 
        .Q(n59) );
  AOI220 U22 ( .A(i_data_lwM[13]), .B(n114), .C(i_data_lwW[13]), .D(n8), .Q(
        n57) );
  AOI220 U23 ( .A(i_data_rs[20]), .B(n5), .C(i_data_writeres[20]), .D(n7), .Q(
        n80) );
  AOI220 U24 ( .A(i_data_lwM[20]), .B(n114), .C(i_data_lwW[20]), .D(n9), .Q(
        n78) );
  AOI220 U25 ( .A(i_data_lwM[8]), .B(n114), .C(i_data_lwW[8]), .D(n9), .Q(n42)
         );
  AOI220 U26 ( .A(i_data_rs[18]), .B(n5), .C(i_data_writeres[18]), .D(n7), .Q(
        n74) );
  AOI220 U27 ( .A(i_data_lwM[18]), .B(n114), .C(i_data_lwW[18]), .D(n9), .Q(
        n72) );
  AOI220 U28 ( .A(i_data_rs[21]), .B(n5), .C(i_data_writeres[21]), .D(n6), .Q(
        n83) );
  AOI220 U29 ( .A(i_data_lwM[21]), .B(n114), .C(i_data_lwW[21]), .D(n8), .Q(
        n81) );
  AOI220 U30 ( .A(i_data_rs[19]), .B(n5), .C(i_data_writeres[19]), .D(n6), .Q(
        n77) );
  AOI220 U31 ( .A(i_data_lwM[19]), .B(n114), .C(i_data_lwW[19]), .D(n8), .Q(
        n75) );
  AOI220 U32 ( .A(i_data_rs[9]), .B(n4), .C(i_data_writeres[9]), .D(n6), .Q(
        n47) );
  AOI220 U33 ( .A(i_data_lwM[9]), .B(n114), .C(i_data_lwW[9]), .D(n9), .Q(n45)
         );
  AOI220 U34 ( .A(i_data_rs[15]), .B(n4), .C(i_data_writeres[15]), .D(n111), 
        .Q(n65) );
  AOI220 U35 ( .A(i_data_lwM[15]), .B(n114), .C(i_data_lwW[15]), .D(n8), .Q(
        n63) );
  AOI220 U36 ( .A(i_data_rs[22]), .B(n5), .C(i_data_writeres[22]), .D(n7), .Q(
        n86) );
  AOI220 U37 ( .A(i_data_lwM[22]), .B(n114), .C(i_data_lwW[22]), .D(n9), .Q(
        n84) );
  AOI220 U38 ( .A(i_data_rs[1]), .B(n4), .C(i_data_writeres[1]), .D(n6), .Q(
        n23) );
  AOI220 U39 ( .A(i_data_lwM[1]), .B(n114), .C(i_data_lwW[1]), .D(n9), .Q(n21)
         );
  AOI220 U40 ( .A(i_data_rs[2]), .B(n4), .C(i_data_writeres[2]), .D(n6), .Q(
        n26) );
  AOI220 U41 ( .A(i_data_lwM[2]), .B(n114), .C(i_data_lwW[2]), .D(n9), .Q(n24)
         );
  AOI220 U42 ( .A(i_data_lwM[5]), .B(n114), .C(i_data_lwW[5]), .D(n113), .Q(
        n33) );
  AOI220 U43 ( .A(i_data_rs[14]), .B(n4), .C(i_data_writeres[14]), .D(n7), .Q(
        n62) );
  AOI220 U44 ( .A(i_data_lwM[14]), .B(n114), .C(i_data_lwW[14]), .D(n9), .Q(
        n60) );
  NAND30 U45 ( .A(i_con_fa[2]), .B(i_con_fa[0]), .C(n16), .Q(n17) );
  NAND30 U46 ( .A(i_con_fa[0]), .B(n12), .C(n16), .Q(n11) );
  AOI220 U47 ( .A(i_data_rs[27]), .B(n5), .C(i_data_writeres[27]), .D(n111), 
        .Q(n101) );
  AOI220 U48 ( .A(i_data_lwM[27]), .B(n114), .C(i_data_lwW[27]), .D(n8), .Q(
        n99) );
  AOI220 U49 ( .A(i_data_rs[28]), .B(n5), .C(i_data_writeres[28]), .D(n7), .Q(
        n104) );
  AOI220 U50 ( .A(i_data_lwM[28]), .B(n114), .C(i_data_lwW[28]), .D(n9), .Q(
        n102) );
  AOI220 U51 ( .A(i_data_rs[24]), .B(n5), .C(i_data_writeres[24]), .D(n7), .Q(
        n92) );
  AOI220 U52 ( .A(i_data_lwM[24]), .B(n114), .C(i_data_lwW[24]), .D(n9), .Q(
        n90) );
  AOI220 U53 ( .A(i_data_rs[29]), .B(n5), .C(i_data_writeres[29]), .D(n7), .Q(
        n107) );
  AOI220 U54 ( .A(i_data_lwM[29]), .B(n114), .C(i_data_lwW[29]), .D(n8), .Q(
        n105) );
  AOI220 U55 ( .A(i_data_rs[25]), .B(n5), .C(i_data_writeres[25]), .D(n111), 
        .Q(n95) );
  AOI220 U56 ( .A(i_data_lwM[25]), .B(n114), .C(i_data_lwW[25]), .D(n8), .Q(
        n93) );
  AOI220 U57 ( .A(i_data_rs[26]), .B(n5), .C(i_data_writeres[26]), .D(n7), .Q(
        n98) );
  AOI220 U58 ( .A(i_data_lwM[26]), .B(n114), .C(i_data_lwW[26]), .D(n9), .Q(
        n96) );
  AOI220 U59 ( .A(i_data_rs[31]), .B(n5), .C(i_data_writeres[31]), .D(n111), 
        .Q(n117) );
  AOI220 U60 ( .A(i_data_lwM[31]), .B(n114), .C(i_data_lwW[31]), .D(n8), .Q(
        n115) );
  AOI220 U61 ( .A(i_data_rs[30]), .B(n5), .C(i_data_writeres[30]), .D(n7), .Q(
        n110) );
  AOI220 U62 ( .A(i_data_lwM[30]), .B(n114), .C(i_data_lwW[30]), .D(n9), .Q(
        n108) );
  BUF2 U63 ( .A(n3), .Q(n5) );
  BUF2 U64 ( .A(n3), .Q(n4) );
  XOR21 U65 ( .A(n16), .B(n10), .Q(n3) );
  BUF2 U66 ( .A(n113), .Q(n8) );
  BUF2 U67 ( .A(n111), .Q(n7) );
  BUF2 U68 ( .A(n113), .Q(n9) );
  BUF2 U69 ( .A(n111), .Q(n6) );
  AOI221 U70 ( .A(i_data_lwM[4]), .B(n114), .C(i_data_lwW[4]), .D(n8), .Q(n30)
         );
  AOI221 U71 ( .A(i_data_rs[4]), .B(n4), .C(i_data_writeres[4]), .D(n6), .Q(
        n32) );
  AOI221 U72 ( .A(i_data_lwM[6]), .B(n114), .C(i_data_lwW[6]), .D(n113), .Q(
        n36) );
  AOI221 U73 ( .A(i_data_rs[6]), .B(n4), .C(i_data_writeres[6]), .D(n6), .Q(
        n38) );
  INV3 U74 ( .A(n15), .Q(n114) );
  NAND31 U75 ( .A(i_con_fa[2]), .B(n14), .C(n16), .Q(n15) );
  NAND31 U76 ( .A(n74), .B(n73), .C(n72), .Q(o_data_alusra[18]) );
  AOI221 U77 ( .A(i_data_lwM[3]), .B(n114), .C(i_data_lwW[3]), .D(n9), .Q(n27)
         );
  AOI221 U78 ( .A(i_data_rs[3]), .B(n4), .C(i_data_writeres[3]), .D(n6), .Q(
        n29) );
  AOI221 U79 ( .A(i_data_rs[5]), .B(n4), .C(i_data_writeres[5]), .D(n6), .Q(
        n35) );
  INV3 U80 ( .A(n11), .Q(n111) );
  INV3 U81 ( .A(n17), .Q(n113) );
  NAND31 U82 ( .A(n53), .B(n52), .C(n51), .Q(o_data_alusra[11]) );
  AOI221 U83 ( .A(i_data_lwM[11]), .B(n114), .C(i_data_lwW[11]), .D(n8), .Q(
        n51) );
  AOI221 U84 ( .A(i_data_rs[11]), .B(n4), .C(i_data_writeres[11]), .D(n111), 
        .Q(n53) );
  NAND31 U85 ( .A(n44), .B(n43), .C(n42), .Q(o_data_alusra[8]) );
  AOI221 U86 ( .A(i_data_rs[8]), .B(n4), .C(i_data_writeres[8]), .D(n6), .Q(
        n44) );
  NAND31 U87 ( .A(n62), .B(n61), .C(n60), .Q(o_data_alusra[14]) );
  NAND31 U88 ( .A(n83), .B(n82), .C(n81), .Q(o_data_alusra[21]) );
  NAND31 U89 ( .A(n65), .B(n64), .C(n63), .Q(o_data_alusra[15]) );
  NAND31 U90 ( .A(n77), .B(n76), .C(n75), .Q(o_data_alusra[19]) );
  NAND31 U91 ( .A(n80), .B(n79), .C(n78), .Q(o_data_alusra[20]) );
  NAND31 U92 ( .A(n47), .B(n46), .C(n45), .Q(o_data_alusra[9]) );
  NAND31 U93 ( .A(n50), .B(n49), .C(n48), .Q(o_data_alusra[10]) );
  AOI221 U94 ( .A(i_data_lwM[10]), .B(n114), .C(i_data_lwW[10]), .D(n9), .Q(
        n48) );
  AOI221 U95 ( .A(i_data_rs[10]), .B(n4), .C(i_data_writeres[10]), .D(n6), .Q(
        n50) );
  NAND31 U96 ( .A(n56), .B(n55), .C(n54), .Q(o_data_alusra[12]) );
  NAND31 U97 ( .A(n59), .B(n58), .C(n57), .Q(o_data_alusra[13]) );
  NAND31 U98 ( .A(n117), .B(n116), .C(n115), .Q(o_data_alusra[31]) );
  NAND31 U99 ( .A(n107), .B(n106), .C(n105), .Q(o_data_alusra[29]) );
  NAND31 U100 ( .A(n95), .B(n94), .C(n93), .Q(o_data_alusra[25]) );
  NAND31 U101 ( .A(n86), .B(n85), .C(n84), .Q(o_data_alusra[22]) );
  NAND31 U102 ( .A(n101), .B(n100), .C(n99), .Q(o_data_alusra[27]) );
  NAND31 U103 ( .A(n104), .B(n103), .C(n102), .Q(o_data_alusra[28]) );
  NAND31 U104 ( .A(n89), .B(n88), .C(n87), .Q(o_data_alusra[23]) );
  NAND31 U105 ( .A(n92), .B(n91), .C(n90), .Q(o_data_alusra[24]) );
  NAND31 U106 ( .A(n98), .B(n97), .C(n96), .Q(o_data_alusra[26]) );
  NAND31 U107 ( .A(n110), .B(n109), .C(n108), .Q(o_data_alusra[30]) );
  CLKIN3 U108 ( .A(i_con_fa[1]), .Q(n16) );
  NAND22 U109 ( .A(n12), .B(n14), .Q(n10) );
  NAND22 U110 ( .A(i_data_alures[0]), .B(n112), .Q(n19) );
  NAND33 U111 ( .A(n20), .B(n19), .C(n18), .Q(o_data_alusra[0]) );
  NAND22 U112 ( .A(i_data_alures[1]), .B(n112), .Q(n22) );
  NAND33 U113 ( .A(n23), .B(n22), .C(n21), .Q(o_data_alusra[1]) );
  NAND22 U114 ( .A(i_data_alures[2]), .B(n112), .Q(n25) );
  NAND33 U115 ( .A(n26), .B(n25), .C(n24), .Q(o_data_alusra[2]) );
  NAND22 U116 ( .A(i_data_alures[3]), .B(n112), .Q(n28) );
  NAND33 U117 ( .A(n29), .B(n28), .C(n27), .Q(o_data_alusra[3]) );
  NAND22 U118 ( .A(i_data_alures[4]), .B(n112), .Q(n31) );
  NAND33 U119 ( .A(n32), .B(n31), .C(n30), .Q(o_data_alusra[4]) );
  NAND22 U120 ( .A(i_data_alures[5]), .B(n112), .Q(n34) );
  NAND33 U121 ( .A(n35), .B(n34), .C(n33), .Q(o_data_alusra[5]) );
  NAND22 U122 ( .A(i_data_alures[6]), .B(n112), .Q(n37) );
  NAND33 U123 ( .A(n38), .B(n37), .C(n36), .Q(o_data_alusra[6]) );
  NAND22 U124 ( .A(i_data_alures[7]), .B(n112), .Q(n40) );
  NAND33 U125 ( .A(n41), .B(n40), .C(n39), .Q(o_data_alusra[7]) );
  NAND22 U126 ( .A(i_data_alures[8]), .B(n112), .Q(n43) );
  NAND22 U127 ( .A(i_data_alures[9]), .B(n112), .Q(n46) );
  NAND22 U128 ( .A(i_data_alures[10]), .B(n112), .Q(n49) );
  NAND22 U129 ( .A(i_data_alures[11]), .B(n112), .Q(n52) );
  NAND22 U130 ( .A(i_data_alures[12]), .B(n112), .Q(n55) );
  NAND22 U131 ( .A(i_data_alures[13]), .B(n112), .Q(n58) );
  NAND22 U132 ( .A(i_data_alures[14]), .B(n112), .Q(n61) );
  NAND22 U133 ( .A(i_data_alures[15]), .B(n112), .Q(n64) );
  NAND22 U134 ( .A(i_data_alures[16]), .B(n112), .Q(n67) );
  NAND22 U135 ( .A(i_data_alures[17]), .B(n112), .Q(n70) );
  NAND22 U136 ( .A(i_data_alures[18]), .B(n112), .Q(n73) );
  NAND22 U137 ( .A(i_data_alures[19]), .B(n112), .Q(n76) );
  NAND22 U138 ( .A(i_data_alures[20]), .B(n112), .Q(n79) );
  NAND22 U139 ( .A(i_data_alures[21]), .B(n112), .Q(n82) );
  NAND22 U140 ( .A(i_data_alures[22]), .B(n112), .Q(n85) );
  NAND22 U141 ( .A(i_data_alures[23]), .B(n112), .Q(n88) );
  NAND22 U142 ( .A(i_data_alures[24]), .B(n112), .Q(n91) );
  NAND22 U143 ( .A(i_data_alures[25]), .B(n112), .Q(n94) );
  NAND22 U144 ( .A(i_data_alures[26]), .B(n112), .Q(n97) );
  NAND22 U145 ( .A(i_data_alures[27]), .B(n112), .Q(n100) );
  NAND22 U146 ( .A(i_data_alures[28]), .B(n112), .Q(n103) );
  NAND22 U147 ( .A(i_data_alures[29]), .B(n112), .Q(n106) );
  NAND22 U148 ( .A(i_data_alures[30]), .B(n112), .Q(n109) );
  NAND22 U149 ( .A(i_data_alures[31]), .B(n112), .Q(n116) );
endmodule


module E_fbmux5 ( i_data_rt, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fb, o_data_alusrb );
  input [31:0] i_data_rt;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fb;
  output [31:0] o_data_alusrb;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119;

  INV3 U1 ( .A(n1), .Q(n2) );
  NAND22 U2 ( .A(n71), .B(n72), .Q(n1) );
  NAND26 U3 ( .A(n67), .B(n8), .Q(o_data_alusrb[16]) );
  NAND33 U4 ( .A(n69), .B(n70), .C(n68), .Q(n7) );
  INV3 U5 ( .A(i_con_fb[1]), .Q(n17) );
  AOI221 U6 ( .A(i_data_lwW[16]), .B(n115), .C(i_data_lwM[16]), .D(n116), .Q(
        n70) );
  NAND22 U7 ( .A(i_data_rt[16]), .B(n9), .Q(n68) );
  NAND31 U8 ( .A(n24), .B(n23), .C(n22), .Q(o_data_alusrb[1]) );
  NAND22 U9 ( .A(n17), .B(n5), .Q(n18) );
  INV6 U10 ( .A(n18), .Q(n115) );
  NAND20 U11 ( .A(i_data_alures[14]), .B(n6), .Q(n62) );
  NAND20 U12 ( .A(i_data_alures[13]), .B(n6), .Q(n59) );
  NAND20 U13 ( .A(i_data_alures[28]), .B(n6), .Q(n105) );
  NAND20 U14 ( .A(i_data_alures[25]), .B(n6), .Q(n96) );
  NAND20 U15 ( .A(i_data_alures[30]), .B(n6), .Q(n111) );
  NAND20 U16 ( .A(i_data_alures[27]), .B(n6), .Q(n102) );
  NAND21 U17 ( .A(i_data_alures[26]), .B(n6), .Q(n99) );
  AOI221 U18 ( .A(i_data_lwM[17]), .B(n116), .C(i_data_lwW[17]), .D(n115), .Q(
        n71) );
  NAND26 U19 ( .A(n73), .B(n2), .Q(o_data_alusrb[17]) );
  INV6 U20 ( .A(n12), .Q(n113) );
  NAND30 U21 ( .A(i_con_fb[0]), .B(n13), .C(n17), .Q(n12) );
  NAND24 U22 ( .A(i_data_writeres[16]), .B(n113), .Q(n67) );
  CLKIN3 U23 ( .A(n16), .Q(n3) );
  CLKIN3 U24 ( .A(n16), .Q(n116) );
  NAND30 U25 ( .A(i_con_fb[2]), .B(n15), .C(n17), .Q(n16) );
  CLKIN3 U26 ( .A(n14), .Q(n6) );
  NAND22 U27 ( .A(i_data_alures[16]), .B(n114), .Q(n69) );
  INV2 U28 ( .A(n4), .Q(n5) );
  INV6 U29 ( .A(n7), .Q(n8) );
  NAND20 U30 ( .A(i_con_fb[0]), .B(i_con_fb[2]), .Q(n4) );
  NAND30 U31 ( .A(i_con_fb[1]), .B(n13), .C(n15), .Q(n14) );
  AOI220 U32 ( .A(i_data_rt[2]), .B(n10), .C(i_data_writeres[2]), .D(n113), 
        .Q(n27) );
  AOI220 U33 ( .A(i_data_rt[9]), .B(n10), .C(i_data_writeres[9]), .D(n113), 
        .Q(n48) );
  BUF6 U34 ( .A(n9), .Q(n10) );
  AOI220 U35 ( .A(i_data_lwM[1]), .B(n3), .C(i_data_lwW[1]), .D(n115), .Q(n22)
         );
  AOI220 U36 ( .A(i_data_lwM[18]), .B(n116), .C(i_data_lwW[18]), .D(n115), .Q(
        n74) );
  NAND33 U37 ( .A(n76), .B(n75), .C(n74), .Q(o_data_alusrb[18]) );
  NAND31 U38 ( .A(n21), .B(n20), .C(n19), .Q(o_data_alusrb[0]) );
  AOI220 U39 ( .A(i_data_lwM[0]), .B(n3), .C(i_data_lwW[0]), .D(n115), .Q(n19)
         );
  AOI220 U40 ( .A(i_data_rt[0]), .B(n10), .C(i_data_writeres[0]), .D(n113), 
        .Q(n21) );
  AOI220 U41 ( .A(i_data_lwM[9]), .B(n3), .C(i_data_lwW[9]), .D(n115), .Q(n46)
         );
  AOI220 U42 ( .A(i_data_rt[10]), .B(n10), .C(i_data_writeres[10]), .D(n113), 
        .Q(n51) );
  AOI220 U43 ( .A(i_data_lwM[10]), .B(n3), .C(i_data_lwW[10]), .D(n115), .Q(
        n49) );
  AOI220 U44 ( .A(i_data_rt[6]), .B(n10), .C(i_data_writeres[6]), .D(n113), 
        .Q(n39) );
  AOI220 U45 ( .A(i_data_lwM[6]), .B(n3), .C(i_data_lwW[6]), .D(n115), .Q(n37)
         );
  AOI220 U46 ( .A(i_data_rt[11]), .B(n10), .C(i_data_writeres[11]), .D(n113), 
        .Q(n54) );
  AOI220 U47 ( .A(i_data_lwM[11]), .B(n3), .C(i_data_lwW[11]), .D(n115), .Q(
        n52) );
  AOI220 U48 ( .A(i_data_rt[12]), .B(n10), .C(i_data_writeres[12]), .D(n113), 
        .Q(n57) );
  AOI220 U49 ( .A(i_data_lwM[12]), .B(n3), .C(i_data_lwW[12]), .D(n115), .Q(
        n55) );
  AOI220 U50 ( .A(i_data_rt[13]), .B(n10), .C(i_data_writeres[13]), .D(n113), 
        .Q(n60) );
  AOI220 U51 ( .A(i_data_lwM[13]), .B(n3), .C(i_data_lwW[13]), .D(n115), .Q(
        n58) );
  AOI220 U52 ( .A(i_data_rt[15]), .B(n10), .C(i_data_writeres[15]), .D(n113), 
        .Q(n66) );
  AOI220 U53 ( .A(i_data_lwM[15]), .B(n3), .C(i_data_lwW[15]), .D(n115), .Q(
        n64) );
  AOI220 U54 ( .A(i_data_lwM[19]), .B(n3), .C(i_data_lwW[19]), .D(n115), .Q(
        n77) );
  AOI220 U55 ( .A(i_data_lwM[20]), .B(n3), .C(i_data_lwW[20]), .D(n115), .Q(
        n80) );
  AOI220 U56 ( .A(i_data_lwM[21]), .B(n3), .C(i_data_lwW[21]), .D(n115), .Q(
        n83) );
  AOI220 U57 ( .A(i_data_lwM[22]), .B(n3), .C(i_data_lwW[22]), .D(n115), .Q(
        n86) );
  AOI220 U58 ( .A(i_data_lwM[23]), .B(n3), .C(i_data_lwW[23]), .D(n115), .Q(
        n89) );
  AOI220 U59 ( .A(i_data_lwM[2]), .B(n3), .C(i_data_lwW[2]), .D(n115), .Q(n25)
         );
  AOI220 U60 ( .A(i_data_rt[5]), .B(n10), .C(i_data_writeres[5]), .D(n113), 
        .Q(n36) );
  AOI220 U61 ( .A(i_data_lwM[5]), .B(n3), .C(i_data_lwW[5]), .D(n115), .Q(n34)
         );
  AOI220 U62 ( .A(i_data_rt[7]), .B(n10), .C(i_data_writeres[7]), .D(n113), 
        .Q(n42) );
  AOI220 U63 ( .A(i_data_lwM[7]), .B(n3), .C(i_data_lwW[7]), .D(n115), .Q(n40)
         );
  AOI220 U64 ( .A(i_data_rt[14]), .B(n10), .C(i_data_writeres[14]), .D(n113), 
        .Q(n63) );
  AOI220 U65 ( .A(i_data_lwM[14]), .B(n3), .C(i_data_lwW[14]), .D(n115), .Q(
        n61) );
  AOI220 U66 ( .A(i_data_lwM[24]), .B(n3), .C(i_data_lwW[24]), .D(n115), .Q(
        n92) );
  AOI220 U67 ( .A(i_data_lwM[25]), .B(n3), .C(i_data_lwW[25]), .D(n115), .Q(
        n95) );
  AOI220 U68 ( .A(i_data_lwM[26]), .B(n3), .C(i_data_lwW[26]), .D(n115), .Q(
        n98) );
  AOI220 U69 ( .A(i_data_lwM[27]), .B(n3), .C(i_data_lwW[27]), .D(n115), .Q(
        n101) );
  AOI220 U70 ( .A(i_data_lwM[28]), .B(n3), .C(i_data_lwW[28]), .D(n115), .Q(
        n104) );
  AOI220 U71 ( .A(i_data_lwM[29]), .B(n3), .C(i_data_lwW[29]), .D(n115), .Q(
        n107) );
  AOI220 U72 ( .A(i_data_lwM[30]), .B(n3), .C(i_data_lwW[30]), .D(n115), .Q(
        n110) );
  AOI220 U73 ( .A(i_data_lwM[31]), .B(n3), .C(i_data_lwW[31]), .D(n115), .Q(
        n117) );
  XOR21 U74 ( .A(n17), .B(n11), .Q(n9) );
  CLKIN3 U75 ( .A(n14), .Q(n114) );
  AOI221 U76 ( .A(i_data_rt[1]), .B(n10), .C(i_data_writeres[1]), .D(n113), 
        .Q(n24) );
  NAND31 U77 ( .A(n79), .B(n78), .C(n77), .Q(o_data_alusrb[19]) );
  NAND31 U78 ( .A(n82), .B(n81), .C(n80), .Q(o_data_alusrb[20]) );
  NAND31 U79 ( .A(n27), .B(n26), .C(n25), .Q(o_data_alusrb[2]) );
  NAND31 U80 ( .A(n42), .B(n41), .C(n40), .Q(o_data_alusrb[7]) );
  NAND31 U81 ( .A(n66), .B(n65), .C(n64), .Q(o_data_alusrb[15]) );
  NAND31 U82 ( .A(n85), .B(n84), .C(n83), .Q(o_data_alusrb[21]) );
  NAND31 U83 ( .A(n88), .B(n87), .C(n86), .Q(o_data_alusrb[22]) );
  NAND31 U84 ( .A(n30), .B(n29), .C(n28), .Q(o_data_alusrb[3]) );
  AOI221 U85 ( .A(i_data_lwM[3]), .B(n3), .C(i_data_lwW[3]), .D(n115), .Q(n28)
         );
  AOI221 U86 ( .A(i_data_rt[3]), .B(n10), .C(i_data_writeres[3]), .D(n113), 
        .Q(n30) );
  NAND31 U87 ( .A(n33), .B(n32), .C(n31), .Q(o_data_alusrb[4]) );
  AOI221 U88 ( .A(i_data_lwM[4]), .B(n3), .C(i_data_lwW[4]), .D(n115), .Q(n31)
         );
  AOI221 U89 ( .A(i_data_rt[4]), .B(n10), .C(i_data_writeres[4]), .D(n113), 
        .Q(n33) );
  NAND31 U90 ( .A(n36), .B(n35), .C(n34), .Q(o_data_alusrb[5]) );
  NAND31 U91 ( .A(n39), .B(n38), .C(n37), .Q(o_data_alusrb[6]) );
  NAND31 U92 ( .A(n45), .B(n44), .C(n43), .Q(o_data_alusrb[8]) );
  AOI221 U93 ( .A(i_data_lwM[8]), .B(n3), .C(i_data_lwW[8]), .D(n115), .Q(n43)
         );
  AOI221 U94 ( .A(i_data_rt[8]), .B(n10), .C(i_data_writeres[8]), .D(n113), 
        .Q(n45) );
  NAND31 U95 ( .A(n48), .B(n47), .C(n46), .Q(o_data_alusrb[9]) );
  NAND31 U96 ( .A(n51), .B(n50), .C(n49), .Q(o_data_alusrb[10]) );
  NAND31 U97 ( .A(n54), .B(n53), .C(n52), .Q(o_data_alusrb[11]) );
  NAND31 U98 ( .A(n57), .B(n56), .C(n55), .Q(o_data_alusrb[12]) );
  NAND31 U99 ( .A(n60), .B(n59), .C(n58), .Q(o_data_alusrb[13]) );
  NAND31 U100 ( .A(n63), .B(n62), .C(n61), .Q(o_data_alusrb[14]) );
  NAND31 U101 ( .A(n91), .B(n90), .C(n89), .Q(o_data_alusrb[23]) );
  NAND31 U102 ( .A(n94), .B(n93), .C(n92), .Q(o_data_alusrb[24]) );
  NAND31 U103 ( .A(n97), .B(n96), .C(n95), .Q(o_data_alusrb[25]) );
  NAND31 U104 ( .A(n100), .B(n99), .C(n98), .Q(o_data_alusrb[26]) );
  NAND31 U105 ( .A(n103), .B(n102), .C(n101), .Q(o_data_alusrb[27]) );
  NAND31 U106 ( .A(n106), .B(n105), .C(n104), .Q(o_data_alusrb[28]) );
  NAND31 U107 ( .A(n109), .B(n108), .C(n107), .Q(o_data_alusrb[29]) );
  NAND31 U108 ( .A(n112), .B(n111), .C(n110), .Q(o_data_alusrb[30]) );
  NAND31 U109 ( .A(n119), .B(n118), .C(n117), .Q(o_data_alusrb[31]) );
  AOI220 U110 ( .A(i_data_rt[30]), .B(n10), .C(i_data_writeres[30]), .D(n113), 
        .Q(n112) );
  AOI220 U111 ( .A(i_data_rt[29]), .B(n10), .C(i_data_writeres[29]), .D(n113), 
        .Q(n109) );
  AOI220 U112 ( .A(i_data_rt[26]), .B(n10), .C(i_data_writeres[26]), .D(n113), 
        .Q(n100) );
  AOI220 U113 ( .A(i_data_rt[28]), .B(n10), .C(i_data_writeres[28]), .D(n113), 
        .Q(n106) );
  AOI220 U114 ( .A(i_data_rt[25]), .B(n10), .C(i_data_writeres[25]), .D(n113), 
        .Q(n97) );
  AOI220 U115 ( .A(i_data_rt[27]), .B(n10), .C(i_data_writeres[27]), .D(n113), 
        .Q(n103) );
  AOI220 U116 ( .A(i_data_rt[31]), .B(n10), .C(i_data_writeres[31]), .D(n113), 
        .Q(n119) );
  AOI220 U117 ( .A(i_data_rt[24]), .B(n10), .C(i_data_writeres[24]), .D(n113), 
        .Q(n94) );
  AOI220 U118 ( .A(i_data_rt[23]), .B(n10), .C(i_data_writeres[23]), .D(n113), 
        .Q(n91) );
  AOI220 U119 ( .A(i_data_rt[22]), .B(n10), .C(i_data_writeres[22]), .D(n113), 
        .Q(n88) );
  AOI220 U120 ( .A(i_data_rt[21]), .B(n10), .C(i_data_writeres[21]), .D(n113), 
        .Q(n85) );
  AOI220 U121 ( .A(i_data_rt[20]), .B(n10), .C(i_data_writeres[20]), .D(n113), 
        .Q(n82) );
  AOI220 U122 ( .A(i_data_rt[19]), .B(n10), .C(i_data_writeres[19]), .D(n113), 
        .Q(n79) );
  AOI220 U123 ( .A(i_data_rt[18]), .B(n10), .C(i_data_writeres[18]), .D(n113), 
        .Q(n76) );
  CLKIN3 U124 ( .A(i_con_fb[2]), .Q(n13) );
  CLKIN3 U125 ( .A(i_con_fb[0]), .Q(n15) );
  NAND22 U126 ( .A(n13), .B(n15), .Q(n11) );
  NAND22 U127 ( .A(i_data_alures[0]), .B(n6), .Q(n20) );
  NAND22 U128 ( .A(i_data_alures[1]), .B(n6), .Q(n23) );
  NAND22 U129 ( .A(i_data_alures[2]), .B(n6), .Q(n26) );
  NAND22 U130 ( .A(i_data_alures[3]), .B(n6), .Q(n29) );
  NAND22 U131 ( .A(i_data_alures[4]), .B(n6), .Q(n32) );
  NAND22 U132 ( .A(i_data_alures[5]), .B(n6), .Q(n35) );
  NAND22 U133 ( .A(i_data_alures[6]), .B(n6), .Q(n38) );
  NAND22 U134 ( .A(i_data_alures[7]), .B(n6), .Q(n41) );
  NAND22 U135 ( .A(i_data_alures[8]), .B(n114), .Q(n44) );
  NAND22 U136 ( .A(i_data_alures[9]), .B(n6), .Q(n47) );
  NAND22 U137 ( .A(i_data_alures[10]), .B(n6), .Q(n50) );
  NAND22 U138 ( .A(i_data_alures[11]), .B(n6), .Q(n53) );
  NAND22 U139 ( .A(i_data_alures[12]), .B(n6), .Q(n56) );
  NAND22 U140 ( .A(i_data_alures[15]), .B(n6), .Q(n65) );
  AOI222 U141 ( .A(i_data_rt[17]), .B(n10), .C(i_data_writeres[17]), .D(n113), 
        .Q(n73) );
  NAND22 U142 ( .A(i_data_alures[17]), .B(n114), .Q(n72) );
  NAND22 U143 ( .A(i_data_alures[18]), .B(n6), .Q(n75) );
  NAND22 U144 ( .A(i_data_alures[19]), .B(n6), .Q(n78) );
  NAND22 U145 ( .A(i_data_alures[20]), .B(n6), .Q(n81) );
  NAND22 U146 ( .A(i_data_alures[21]), .B(n6), .Q(n84) );
  NAND22 U147 ( .A(i_data_alures[22]), .B(n6), .Q(n87) );
  NAND22 U148 ( .A(i_data_alures[23]), .B(n6), .Q(n90) );
  NAND22 U149 ( .A(i_data_alures[24]), .B(n6), .Q(n93) );
  NAND22 U150 ( .A(i_data_alures[29]), .B(n6), .Q(n108) );
  NAND22 U151 ( .A(i_data_alures[31]), .B(n6), .Q(n118) );
endmodule


module E_alubmux ( i_data_fb, i_data_imm, i_con_imm, o_data_alub );
  input [31:0] i_data_fb;
  input [31:0] i_data_imm;
  output [31:0] o_data_alub;
  input i_con_imm;
  wire   n1, n2, n3, n4, n5, n6;

  CLKIN3 U1 ( .A(n5), .Q(o_data_alub[16]) );
  MUX26 U2 ( .A(i_data_fb[20]), .B(i_data_imm[20]), .S(n3), .Q(o_data_alub[20]) );
  NAND22 U3 ( .A(n1), .B(n2), .Q(o_data_alub[0]) );
  INV3 U4 ( .A(n6), .Q(o_data_alub[17]) );
  MUX22 U5 ( .A(i_data_fb[8]), .B(i_data_imm[8]), .S(i_con_imm), .Q(
        o_data_alub[8]) );
  NAND22 U6 ( .A(i_data_fb[0]), .B(n4), .Q(n1) );
  MUX22 U7 ( .A(i_data_fb[1]), .B(i_data_imm[1]), .S(i_con_imm), .Q(
        o_data_alub[1]) );
  NAND22 U8 ( .A(i_data_imm[0]), .B(n3), .Q(n2) );
  CLKIN3 U9 ( .A(n4), .Q(n3) );
  AOI222 U10 ( .A(i_data_fb[16]), .B(n4), .C(i_data_imm[16]), .D(i_con_imm), 
        .Q(n5) );
  MUX22 U11 ( .A(i_data_fb[2]), .B(i_data_imm[2]), .S(n3), .Q(o_data_alub[2])
         );
  MUX22 U12 ( .A(i_data_fb[18]), .B(i_data_imm[18]), .S(i_con_imm), .Q(
        o_data_alub[18]) );
  MUX22 U13 ( .A(i_data_fb[19]), .B(i_data_imm[19]), .S(n3), .Q(
        o_data_alub[19]) );
  MUX22 U14 ( .A(i_data_fb[11]), .B(i_data_imm[11]), .S(i_con_imm), .Q(
        o_data_alub[11]) );
  MUX22 U15 ( .A(i_data_fb[10]), .B(i_data_imm[10]), .S(i_con_imm), .Q(
        o_data_alub[10]) );
  MUX22 U16 ( .A(i_data_fb[9]), .B(i_data_imm[9]), .S(i_con_imm), .Q(
        o_data_alub[9]) );
  MUX22 U17 ( .A(i_data_fb[3]), .B(i_data_imm[3]), .S(n3), .Q(o_data_alub[3])
         );
  MUX22 U18 ( .A(i_data_fb[4]), .B(i_data_imm[4]), .S(i_con_imm), .Q(
        o_data_alub[4]) );
  MUX22 U19 ( .A(i_data_fb[5]), .B(i_data_imm[5]), .S(i_con_imm), .Q(
        o_data_alub[5]) );
  MUX22 U20 ( .A(i_data_fb[21]), .B(i_data_imm[21]), .S(n3), .Q(
        o_data_alub[21]) );
  MUX22 U21 ( .A(i_data_fb[22]), .B(i_data_imm[22]), .S(n3), .Q(
        o_data_alub[22]) );
  INV3 U22 ( .A(i_con_imm), .Q(n4) );
  MUX22 U23 ( .A(i_data_fb[12]), .B(i_data_imm[12]), .S(i_con_imm), .Q(
        o_data_alub[12]) );
  MUX22 U24 ( .A(i_data_fb[7]), .B(i_data_imm[7]), .S(i_con_imm), .Q(
        o_data_alub[7]) );
  MUX22 U25 ( .A(i_data_fb[14]), .B(i_data_imm[14]), .S(i_con_imm), .Q(
        o_data_alub[14]) );
  MUX22 U26 ( .A(i_data_fb[13]), .B(i_data_imm[13]), .S(i_con_imm), .Q(
        o_data_alub[13]) );
  MUX22 U27 ( .A(i_data_fb[6]), .B(i_data_imm[6]), .S(i_con_imm), .Q(
        o_data_alub[6]) );
  MUX22 U28 ( .A(i_data_fb[28]), .B(i_data_imm[28]), .S(n3), .Q(
        o_data_alub[28]) );
  MUX22 U29 ( .A(i_data_fb[27]), .B(i_data_imm[27]), .S(n3), .Q(
        o_data_alub[27]) );
  MUX22 U30 ( .A(i_data_fb[26]), .B(i_data_imm[26]), .S(n3), .Q(
        o_data_alub[26]) );
  MUX22 U31 ( .A(i_data_fb[25]), .B(i_data_imm[25]), .S(n3), .Q(
        o_data_alub[25]) );
  MUX22 U32 ( .A(i_data_fb[29]), .B(i_data_imm[29]), .S(n3), .Q(
        o_data_alub[29]) );
  MUX22 U33 ( .A(i_data_fb[30]), .B(i_data_imm[30]), .S(n3), .Q(
        o_data_alub[30]) );
  MUX22 U34 ( .A(i_data_fb[23]), .B(i_data_imm[23]), .S(n3), .Q(
        o_data_alub[23]) );
  MUX22 U35 ( .A(i_data_fb[24]), .B(i_data_imm[24]), .S(n3), .Q(
        o_data_alub[24]) );
  MUX22 U36 ( .A(i_data_fb[31]), .B(i_data_imm[31]), .S(i_con_imm), .Q(
        o_data_alub[31]) );
  MUX22 U37 ( .A(i_data_fb[15]), .B(i_data_imm[15]), .S(i_con_imm), .Q(
        o_data_alub[15]) );
  AOI222 U38 ( .A(i_data_fb[17]), .B(n4), .C(i_data_imm[17]), .D(i_con_imm), 
        .Q(n6) );
endmodule


module E_rdmux ( i_data_rtE, i_data_rdE, i_con_regdst, i_con_aluPC4, 
        o_data_writeE );
  input [4:0] i_data_rtE;
  input [4:0] i_data_rdE;
  output [4:0] o_data_writeE;
  input i_con_regdst, i_con_aluPC4;
  wire   n7, n8, n9, n10, n11, n1, n2, n3, n4, n5, n6;

  OAI2111 U2 ( .A(i_con_regdst), .B(n4), .C(n6), .D(n10), .Q(o_data_writeE[1])
         );
  INV3 U3 ( .A(i_data_rtE[1]), .Q(n4) );
  NAND22 U4 ( .A(i_data_rdE[1]), .B(i_con_regdst), .Q(n10) );
  OAI2111 U5 ( .A(i_con_regdst), .B(n5), .C(n6), .D(n11), .Q(o_data_writeE[0])
         );
  INV3 U6 ( .A(i_data_rtE[0]), .Q(n5) );
  NAND22 U7 ( .A(i_data_rdE[0]), .B(i_con_regdst), .Q(n11) );
  OAI2111 U8 ( .A(i_con_regdst), .B(n1), .C(n6), .D(n7), .Q(o_data_writeE[4])
         );
  INV3 U9 ( .A(i_data_rtE[4]), .Q(n1) );
  NAND22 U10 ( .A(i_data_rdE[4]), .B(i_con_regdst), .Q(n7) );
  OAI2111 U11 ( .A(i_con_regdst), .B(n3), .C(n6), .D(n9), .Q(o_data_writeE[2])
         );
  INV3 U12 ( .A(i_data_rtE[2]), .Q(n3) );
  NAND22 U13 ( .A(i_data_rdE[2]), .B(i_con_regdst), .Q(n9) );
  OAI2111 U14 ( .A(i_con_regdst), .B(n2), .C(n6), .D(n8), .Q(o_data_writeE[3])
         );
  INV3 U15 ( .A(i_data_rtE[3]), .Q(n2) );
  NAND22 U16 ( .A(i_data_rdE[3]), .B(i_con_regdst), .Q(n8) );
  INV3 U17 ( .A(i_con_aluPC4), .Q(n6) );
endmodule


module D_compare_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  NAND21 U1 ( .A(A[0]), .B(n4), .Q(n28) );
  INV2 U2 ( .A(n27), .Q(n2) );
  INV0 U3 ( .A(A[1]), .Q(n3) );
  INV2 U4 ( .A(NE), .Q(EQ) );
  INV3 U5 ( .A(B[0]), .Q(n4) );
  NAND20 U6 ( .A(n5), .B(n6), .Q(NE) );
  NOR40 U7 ( .A(n7), .B(n8), .C(n9), .D(n10), .Q(n6) );
  NAND40 U8 ( .A(n11), .B(n12), .C(n13), .D(n14), .Q(n10) );
  XNR20 U9 ( .A(B[11]), .B(A[11]), .Q(n14) );
  XNR20 U10 ( .A(B[12]), .B(A[12]), .Q(n13) );
  XNR20 U11 ( .A(B[13]), .B(A[13]), .Q(n12) );
  XNR20 U12 ( .A(B[14]), .B(A[14]), .Q(n11) );
  NAND40 U13 ( .A(n15), .B(n16), .C(n17), .D(n18), .Q(n9) );
  XNR20 U14 ( .A(B[7]), .B(A[7]), .Q(n18) );
  XNR20 U15 ( .A(B[8]), .B(A[8]), .Q(n17) );
  XNR20 U16 ( .A(B[9]), .B(A[9]), .Q(n16) );
  XNR20 U17 ( .A(B[10]), .B(A[10]), .Q(n15) );
  NAND40 U18 ( .A(n19), .B(n20), .C(n21), .D(n22), .Q(n8) );
  XNR20 U19 ( .A(B[3]), .B(A[3]), .Q(n22) );
  XNR20 U20 ( .A(B[4]), .B(A[4]), .Q(n21) );
  XNR20 U21 ( .A(B[5]), .B(A[5]), .Q(n20) );
  XNR20 U22 ( .A(B[6]), .B(A[6]), .Q(n19) );
  NAND40 U23 ( .A(n23), .B(n24), .C(n2), .D(n25), .Q(n7) );
  OAI220 U24 ( .A(n26), .B(n3), .C(B[1]), .D(n26), .Q(n25) );
  NOR20 U25 ( .A(n4), .B(A[0]), .Q(n26) );
  AOI220 U26 ( .A(n3), .B(n28), .C(n28), .D(B[1]), .Q(n27) );
  XNR20 U27 ( .A(B[31]), .B(A[31]), .Q(n24) );
  XNR20 U28 ( .A(B[2]), .B(A[2]), .Q(n23) );
  NOR40 U29 ( .A(n29), .B(n30), .C(n31), .D(n32), .Q(n5) );
  NAND40 U30 ( .A(n33), .B(n34), .C(n35), .D(n36), .Q(n32) );
  XNR20 U31 ( .A(B[27]), .B(A[27]), .Q(n36) );
  XNR20 U32 ( .A(B[28]), .B(A[28]), .Q(n35) );
  XNR20 U33 ( .A(B[29]), .B(A[29]), .Q(n34) );
  XNR20 U34 ( .A(B[30]), .B(A[30]), .Q(n33) );
  NAND40 U35 ( .A(n37), .B(n38), .C(n39), .D(n40), .Q(n31) );
  XNR20 U36 ( .A(B[23]), .B(A[23]), .Q(n40) );
  XNR20 U37 ( .A(B[24]), .B(A[24]), .Q(n39) );
  XNR20 U38 ( .A(B[25]), .B(A[25]), .Q(n38) );
  XNR20 U39 ( .A(B[26]), .B(A[26]), .Q(n37) );
  NAND40 U40 ( .A(n41), .B(n42), .C(n43), .D(n44), .Q(n30) );
  XNR20 U41 ( .A(B[19]), .B(A[19]), .Q(n44) );
  XNR20 U42 ( .A(B[20]), .B(A[20]), .Q(n43) );
  XNR20 U43 ( .A(B[21]), .B(A[21]), .Q(n42) );
  XNR20 U44 ( .A(B[22]), .B(A[22]), .Q(n41) );
  NAND40 U45 ( .A(n45), .B(n46), .C(n47), .D(n48), .Q(n29) );
  XNR20 U46 ( .A(B[15]), .B(A[15]), .Q(n48) );
  XNR20 U47 ( .A(B[16]), .B(A[16]), .Q(n47) );
  XNR20 U48 ( .A(B[17]), .B(A[17]), .Q(n46) );
  XNR20 U49 ( .A(B[18]), .B(A[18]), .Q(n45) );
endmodule


module D_compare ( o_con_ifbranch, i_data_rs, i_data_rt, i_con_bop );
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [2:0] i_con_bop;
  output o_con_ifbranch;
  wire   N32, N33, n4, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n1, n2, n3, n5, n6;

  AOI222 U7 ( .A(N32), .B(n3), .C(i_data_rs[31]), .D(i_con_bop[2]), .Q(n14) );
  D_compare_DW01_cmp6_0 r49 ( .A(i_data_rs), .B(i_data_rt), .TC(n4), .EQ(N32), 
        .NE(N33) );
  AOI211 U2 ( .A(N33), .B(n6), .C(n16), .Q(n10) );
  OAI311 U3 ( .A(n5), .B(i_con_bop[2]), .C(n10), .D(n11), .Q(o_con_ifbranch)
         );
  INV0 U4 ( .A(i_data_rs[31]), .Q(n1) );
  NOR30 U5 ( .A(i_data_rs[0]), .B(i_data_rs[11]), .C(i_data_rs[10]), .Q(n19)
         );
  AOI312 U6 ( .A(n6), .B(n1), .C(n12), .D(n13), .Q(n11) );
  INV3 U8 ( .A(n15), .Q(n2) );
  NOR40 U9 ( .A(i_data_rs[2]), .B(i_data_rs[29]), .C(i_data_rs[28]), .D(
        i_data_rs[27]), .Q(n24) );
  NOR40 U10 ( .A(i_data_rs[5]), .B(i_data_rs[4]), .C(i_data_rs[3]), .D(
        i_data_rs[30]), .Q(n25) );
  NOR40 U11 ( .A(i_data_rs[9]), .B(i_data_rs[8]), .C(i_data_rs[7]), .D(
        i_data_rs[6]), .Q(n26) );
  AOI211 U12 ( .A(n15), .B(n5), .C(n3), .Q(n12) );
  NOR21 U13 ( .A(n17), .B(n18), .Q(n15) );
  NAND41 U14 ( .A(n19), .B(n20), .C(n21), .D(n22), .Q(n18) );
  NAND41 U15 ( .A(n23), .B(n24), .C(n25), .D(n26), .Q(n17) );
  NOR40 U16 ( .A(i_data_rs[19]), .B(i_data_rs[18]), .C(i_data_rs[17]), .D(
        i_data_rs[16]), .Q(n21) );
  NOR40 U17 ( .A(i_data_rs[22]), .B(i_data_rs[21]), .C(i_data_rs[20]), .D(
        i_data_rs[1]), .Q(n22) );
  NOR40 U18 ( .A(i_data_rs[15]), .B(i_data_rs[14]), .C(i_data_rs[13]), .D(
        i_data_rs[12]), .Q(n20) );
  NOR40 U19 ( .A(i_data_rs[26]), .B(i_data_rs[25]), .C(i_data_rs[24]), .D(
        i_data_rs[23]), .Q(n23) );
  AOI211 U20 ( .A(n1), .B(n2), .C(n6), .Q(n16) );
  NOR32 U21 ( .A(n6), .B(i_con_bop[1]), .C(n14), .Q(n13) );
  INV3 U22 ( .A(i_con_bop[0]), .Q(n6) );
  INV3 U23 ( .A(i_con_bop[1]), .Q(n5) );
  INV3 U24 ( .A(i_con_bop[2]), .Q(n3) );
  LOGIC0 U25 ( .Q(n4) );
endmodule


module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Ealuop, i_con_Ealusrc, 
        i_con_Eregdst, i_con_Mmemread, i_con_Mmemwrite, i_con_Wloadmux, 
        i_con_Walupc8, i_con_Wmemtoreg, i_con_Wregwrite, i_con_Efamux, 
        i_con_Efbmux, i_con_bop, o_data_pc4, o_data_alures, o_data_rt, 
        o_addr_regdst, o_con_Mmemread, o_con_Mmemwrite, o_con_Wloadmux, 
        o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_addr_Erd, 
        o_addr_Mrt, o_con_ifbranch );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [5:0] i_con_Ealuop;
  input [1:0] i_con_Wloadmux;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [2:0] i_con_bop;
  output [31:0] o_data_pc4;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [1:0] o_con_Wloadmux;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Walupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Walupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch;

  wire   [31:0] alu_o_data_AluRes;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;

  DFC3 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[0]) );
  DFC3 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC3 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC3 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC3 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC3 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC3 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC3 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC3 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC3 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC3 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC3 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC3 pipe_rt_reg_28_ ( .D(compare_i_data_rt[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[28]) );
  DFC3 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  DFC3 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC3 pipe_rt_reg_25_ ( .D(compare_i_data_rt[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[25]) );
  DFC3 pipe_rt_reg_24_ ( .D(compare_i_data_rt[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[24]) );
  DFC3 pipe_rt_reg_23_ ( .D(compare_i_data_rt[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[23]) );
  DFC3 pipe_rt_reg_22_ ( .D(compare_i_data_rt[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[22]) );
  DFC3 pipe_rt_reg_18_ ( .D(compare_i_data_rt[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[18]) );
  DFC3 pipe_rt_reg_15_ ( .D(compare_i_data_rt[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[15]) );
  DFC3 pipe_rt_reg_14_ ( .D(compare_i_data_rt[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[14]) );
  DFC3 pipe_rt_reg_13_ ( .D(compare_i_data_rt[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[13]) );
  DFC3 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC3 pipe_rt_reg_11_ ( .D(compare_i_data_rt[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[11]) );
  DFC3 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC3 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC3 pipe_rt_reg_0_ ( .D(compare_i_data_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[0]) );
  DFC3 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC3 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC3 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC3 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC3 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC3 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wloadmux_reg_1_ ( .D(i_con_Wloadmux[1]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[1]) );
  DFC3 pipe_con_Wloadmux_reg_0_ ( .D(i_con_Wloadmux[0]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[0]) );
  DFC3 pipe_con_Walupc8_reg ( .D(i_con_Walupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Walupc8) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  E_alu u_alu ( .o_data_AluRes(alu_o_data_AluRes), .i_data_A(compare_i_data_rs), .i_data_B(alu_i_data_B), .i_con_AluCtrl(alu_i_con_AluCtrl), .i_data_shamt(
        i_data_immext[10:6]) );
  E_alu_control u_alu_control ( .o_con_AluCtrl(alu_i_con_AluCtrl), 
        .i_con_AluOp(i_con_Ealuop), .i_con_FuncCode(i_data_immext[5:0]) );
  E_famux5 u_famux5 ( .i_data_rs(i_data_rs), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fa(i_con_Efamux), .o_data_alusra(
        compare_i_data_rs) );
  E_fbmux5 u_fbmux ( .i_data_rt(i_data_rt), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fb(i_con_Efbmux), .o_data_alusrb(
        compare_i_data_rt) );
  E_alubmux u_alubmux ( .i_data_fb(compare_i_data_rt), .i_data_imm(
        i_data_immext), .i_con_imm(i_con_Ealusrc), .o_data_alub(alu_i_data_B)
         );
  E_rdmux u_rdmux ( .i_data_rtE(i_addr_rt), .i_data_rdE(i_addr_rd), 
        .i_con_regdst(i_con_Eregdst), .i_con_aluPC4(i_con_Walupc8), 
        .o_data_writeE(o_addr_Erd) );
  D_compare u_compare ( .o_con_ifbranch(o_con_ifbranch), .i_data_rs(
        compare_i_data_rs), .i_data_rt(compare_i_data_rt), .i_con_bop(
        i_con_bop) );
  DFC1 pipe_rt_reg_16_ ( .D(compare_i_data_rt[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[16]) );
  DFC1 pipe_rt_reg_21_ ( .D(compare_i_data_rt[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[21]) );
  DFC1 pipe_rt_reg_20_ ( .D(compare_i_data_rt[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[20]) );
  DFC1 pipe_rt_reg_19_ ( .D(compare_i_data_rt[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[19]) );
  DFC1 pipe_rt_reg_10_ ( .D(compare_i_data_rt[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[10]) );
  DFC1 pipe_rt_reg_9_ ( .D(compare_i_data_rt[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[9]) );
  DFC1 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC1 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC1 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC1 pipe_rt_reg_2_ ( .D(compare_i_data_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[2]) );
  DFC1 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  DFC1 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC1 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC1 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC1 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC1 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC1 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC1 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC1 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC1 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC1 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC1 pipe_rt_reg_5_ ( .D(compare_i_data_rt[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[5]) );
  DFC1 pipe_alures_reg_15_ ( .D(alu_o_data_AluRes[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[15]) );
  DFC1 pipe_alures_reg_14_ ( .D(alu_o_data_AluRes[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[14]) );
  DFC1 pipe_alures_reg_13_ ( .D(alu_o_data_AluRes[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[13]) );
  DFC1 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC1 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC1 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC1 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC1 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_rt_reg_17_ ( .D(compare_i_data_rt[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[17]) );
endmodule


module mem_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  NOR21 U2 ( .A(n81), .B(n82), .Q(n80) );
  INV3 U3 ( .A(n83), .Q(n81) );
  NOR31 U4 ( .A(n10), .B(n84), .C(n7), .Q(n83) );
  NAND22 U5 ( .A(n34), .B(n35), .Q(n33) );
  NOR31 U6 ( .A(n38), .B(n36), .C(n37), .Q(n35) );
  NOR21 U7 ( .A(n22), .B(n33), .Q(n21) );
  INV3 U8 ( .A(n23), .Q(n22) );
  NOR31 U9 ( .A(n26), .B(n24), .C(n25), .Q(n23) );
  NOR21 U10 ( .A(n50), .B(n54), .Q(n53) );
  NOR21 U11 ( .A(n38), .B(n42), .Q(n41) );
  NOR21 U12 ( .A(n26), .B(n30), .Q(n29) );
  XNR21 U13 ( .A(n31), .B(n26), .Q(SUM[25]) );
  XNR21 U14 ( .A(n53), .B(n49), .Q(SUM[18]) );
  XNR21 U15 ( .A(n41), .B(n37), .Q(SUM[22]) );
  XNR21 U16 ( .A(n29), .B(n25), .Q(SUM[26]) );
  INV3 U17 ( .A(n57), .Q(n46) );
  NAND31 U18 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  NOR21 U19 ( .A(n62), .B(n63), .Q(n58) );
  INV3 U20 ( .A(n61), .Q(n59) );
  NOR21 U21 ( .A(n78), .B(n2), .Q(n77) );
  NOR21 U22 ( .A(n63), .B(n67), .Q(n66) );
  XNR21 U23 ( .A(n1), .B(n2), .Q(SUM[9]) );
  XNR21 U24 ( .A(n68), .B(n63), .Q(SUM[13]) );
  XNR21 U25 ( .A(n55), .B(n50), .Q(SUM[17]) );
  XNR21 U26 ( .A(n43), .B(n38), .Q(SUM[21]) );
  XNR21 U27 ( .A(n66), .B(n62), .Q(SUM[14]) );
  XNR21 U28 ( .A(n77), .B(n74), .Q(SUM[10]) );
  XNR21 U29 ( .A(n6), .B(n7), .Q(SUM[6]) );
  INV3 U30 ( .A(n8), .Q(n6) );
  NAND22 U31 ( .A(n9), .B(A[5]), .Q(n8) );
  XNR21 U32 ( .A(n9), .B(n10), .Q(SUM[5]) );
  NAND22 U33 ( .A(A[3]), .B(A[2]), .Q(n82) );
  NOR21 U34 ( .A(n19), .B(n20), .Q(n18) );
  INV3 U35 ( .A(A[28]), .Q(n20) );
  NOR21 U36 ( .A(n71), .B(n3), .Q(n60) );
  INV3 U37 ( .A(n72), .Q(n71) );
  NOR31 U38 ( .A(n2), .B(n73), .C(n74), .Q(n72) );
  NAND22 U39 ( .A(A[11]), .B(A[8]), .Q(n73) );
  NOR21 U40 ( .A(n33), .B(n32), .Q(n31) );
  INV3 U41 ( .A(A[24]), .Q(n32) );
  INV3 U42 ( .A(A[9]), .Q(n2) );
  INV3 U43 ( .A(A[5]), .Q(n10) );
  NOR21 U44 ( .A(n15), .B(n16), .Q(n14) );
  INV3 U45 ( .A(A[29]), .Q(n16) );
  NOR21 U46 ( .A(n57), .B(n56), .Q(n55) );
  INV3 U47 ( .A(A[16]), .Q(n56) );
  NOR21 U48 ( .A(n45), .B(n44), .Q(n43) );
  INV3 U49 ( .A(A[20]), .Q(n44) );
  INV3 U50 ( .A(A[6]), .Q(n7) );
  INV3 U51 ( .A(A[10]), .Q(n74) );
  XNR21 U52 ( .A(A[24]), .B(n33), .Q(SUM[24]) );
  XNR21 U53 ( .A(A[28]), .B(n19), .Q(SUM[28]) );
  XNR21 U54 ( .A(A[29]), .B(n15), .Q(SUM[29]) );
  XOR21 U55 ( .A(A[30]), .B(n14), .Q(SUM[30]) );
  XOR21 U56 ( .A(n51), .B(n52), .Q(SUM[19]) );
  INV3 U57 ( .A(A[19]), .Q(n51) );
  NAND22 U58 ( .A(n53), .B(A[18]), .Q(n52) );
  XOR21 U59 ( .A(n39), .B(n40), .Q(SUM[23]) );
  INV3 U60 ( .A(A[23]), .Q(n39) );
  NAND22 U61 ( .A(n41), .B(A[22]), .Q(n40) );
  XOR21 U62 ( .A(n27), .B(n28), .Q(SUM[27]) );
  INV3 U63 ( .A(A[27]), .Q(n27) );
  NAND22 U64 ( .A(n29), .B(A[26]), .Q(n28) );
  XOR21 U65 ( .A(n12), .B(n13), .Q(SUM[31]) );
  INV3 U66 ( .A(A[31]), .Q(n12) );
  NAND22 U67 ( .A(A[30]), .B(n14), .Q(n13) );
  NAND22 U68 ( .A(A[7]), .B(A[4]), .Q(n84) );
  INV3 U69 ( .A(A[2]), .Q(SUM[2]) );
  INV3 U70 ( .A(n45), .Q(n34) );
  NAND22 U71 ( .A(n46), .B(n47), .Q(n45) );
  NOR31 U72 ( .A(n50), .B(n48), .C(n49), .Q(n47) );
  NAND22 U73 ( .A(A[19]), .B(A[16]), .Q(n48) );
  NOR21 U74 ( .A(n82), .B(n11), .Q(n9) );
  INV3 U75 ( .A(A[4]), .Q(n11) );
  NOR21 U76 ( .A(n3), .B(n79), .Q(n1) );
  INV3 U77 ( .A(A[8]), .Q(n79) );
  INV3 U78 ( .A(A[17]), .Q(n50) );
  INV3 U79 ( .A(A[21]), .Q(n38) );
  INV3 U80 ( .A(A[25]), .Q(n26) );
  INV3 U81 ( .A(A[13]), .Q(n63) );
  NOR21 U82 ( .A(n69), .B(n70), .Q(n68) );
  INV3 U83 ( .A(A[12]), .Q(n70) );
  INV3 U84 ( .A(A[14]), .Q(n62) );
  INV3 U85 ( .A(A[18]), .Q(n49) );
  INV3 U86 ( .A(A[22]), .Q(n37) );
  INV3 U87 ( .A(A[26]), .Q(n25) );
  XNR21 U88 ( .A(A[8]), .B(n3), .Q(SUM[8]) );
  XNR21 U89 ( .A(A[12]), .B(n69), .Q(SUM[12]) );
  XNR21 U90 ( .A(A[16]), .B(n57), .Q(SUM[16]) );
  XNR21 U91 ( .A(A[20]), .B(n45), .Q(SUM[20]) );
  XOR21 U92 ( .A(n4), .B(n5), .Q(SUM[7]) );
  INV3 U93 ( .A(A[7]), .Q(n4) );
  NAND22 U94 ( .A(n6), .B(A[6]), .Q(n5) );
  XOR21 U95 ( .A(n75), .B(n76), .Q(SUM[11]) );
  INV3 U96 ( .A(A[11]), .Q(n75) );
  NAND22 U97 ( .A(n77), .B(A[10]), .Q(n76) );
  XOR21 U98 ( .A(n64), .B(n65), .Q(SUM[15]) );
  INV3 U99 ( .A(A[15]), .Q(n64) );
  NAND22 U100 ( .A(n66), .B(A[14]), .Q(n65) );
  NAND22 U101 ( .A(A[23]), .B(A[20]), .Q(n36) );
  NAND22 U102 ( .A(A[27]), .B(A[24]), .Q(n24) );
  NAND22 U103 ( .A(A[15]), .B(A[12]), .Q(n61) );
  XNR21 U104 ( .A(A[4]), .B(n82), .Q(SUM[4]) );
  XOR21 U105 ( .A(A[3]), .B(A[2]), .Q(SUM[3]) );
  CLKIN3 U106 ( .A(n18), .Q(n15) );
  CLKIN3 U107 ( .A(n21), .Q(n19) );
  CLKIN3 U108 ( .A(n31), .Q(n30) );
  CLKIN3 U109 ( .A(n43), .Q(n42) );
  CLKIN3 U110 ( .A(n55), .Q(n54) );
  CLKIN3 U111 ( .A(n68), .Q(n67) );
  CLKIN3 U112 ( .A(n60), .Q(n69) );
  CLKIN3 U113 ( .A(n1), .Q(n78) );
  CLKIN3 U114 ( .A(n80), .Q(n3) );
endmodule


module mem ( i_clk, i_nrst, i_data_pc4, i_data_alures, i_data_memout, 
        i_addr_regdst, i_con_Wloadmux, i_con_Walupc8, i_con_Wmemtoreg, 
        i_con_Wregwrite, i_con_FWmemread, i_addr_Mrt, o_data_pc8, 
        o_data_alures, o_data_memout, o_addr_regdst, o_con_Wloadmux, 
        o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread, 
        o_addr_Wrt );
  input [31:0] i_data_pc4;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [4:0] i_addr_regdst;
  input [1:0] i_con_Wloadmux;
  input [4:0] i_addr_Mrt;
  output [31:0] o_data_pc8;
  output [31:0] o_data_alures;
  output [31:0] o_data_memout;
  output [4:0] o_addr_regdst;
  output [1:0] o_con_Wloadmux;
  output [4:0] o_addr_Wrt;
  input i_clk, i_nrst, i_con_Walupc8, i_con_Wmemtoreg, i_con_Wregwrite,
         i_con_FWmemread;
  output o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread;
  wire   n_Logic1_, n_Logic0_;
  wire   [31:0] pc8;

  DFC3 pipe_rt_reg_4_ ( .D(i_addr_Mrt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(i_addr_Mrt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(i_addr_Mrt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[2]) );
  DFC3 pipe_rt_reg_1_ ( .D(i_addr_Mrt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[1]) );
  DFC3 pipe_rt_reg_0_ ( .D(i_addr_Mrt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[0]) );
  DFC3 pipe_data_pc8_reg_31_ ( .D(pc8[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[31]) );
  DFC3 pipe_data_pc8_reg_30_ ( .D(pc8[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[30]) );
  DFC3 pipe_data_pc8_reg_29_ ( .D(pc8[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[29]) );
  DFC3 pipe_data_pc8_reg_28_ ( .D(pc8[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[28]) );
  DFC3 pipe_data_pc8_reg_27_ ( .D(pc8[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[27]) );
  DFC3 pipe_data_pc8_reg_26_ ( .D(pc8[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[26]) );
  DFC3 pipe_data_pc8_reg_25_ ( .D(pc8[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[25]) );
  DFC3 pipe_data_pc8_reg_24_ ( .D(pc8[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[24]) );
  DFC3 pipe_data_pc8_reg_23_ ( .D(pc8[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[23]) );
  DFC3 pipe_data_pc8_reg_22_ ( .D(pc8[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[22]) );
  DFC3 pipe_data_pc8_reg_21_ ( .D(pc8[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[21]) );
  DFC3 pipe_data_pc8_reg_20_ ( .D(pc8[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[20]) );
  DFC3 pipe_data_pc8_reg_19_ ( .D(pc8[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[19]) );
  DFC3 pipe_data_pc8_reg_18_ ( .D(pc8[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[18]) );
  DFC3 pipe_data_pc8_reg_17_ ( .D(pc8[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[17]) );
  DFC3 pipe_data_pc8_reg_16_ ( .D(pc8[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[16]) );
  DFC3 pipe_data_pc8_reg_15_ ( .D(pc8[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[15]) );
  DFC3 pipe_data_pc8_reg_14_ ( .D(pc8[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[14]) );
  DFC3 pipe_data_pc8_reg_13_ ( .D(pc8[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[13]) );
  DFC3 pipe_data_pc8_reg_12_ ( .D(pc8[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[12]) );
  DFC3 pipe_data_pc8_reg_11_ ( .D(pc8[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[11]) );
  DFC3 pipe_data_pc8_reg_10_ ( .D(pc8[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[10]) );
  DFC3 pipe_data_pc8_reg_9_ ( .D(pc8[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[9]) );
  DFC3 pipe_data_pc8_reg_8_ ( .D(pc8[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[8]) );
  DFC3 pipe_data_pc8_reg_7_ ( .D(pc8[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[7]) );
  DFC3 pipe_data_pc8_reg_6_ ( .D(pc8[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[6]) );
  DFC3 pipe_data_pc8_reg_5_ ( .D(pc8[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[5]) );
  DFC3 pipe_data_pc8_reg_4_ ( .D(pc8[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[4]) );
  DFC3 pipe_data_pc8_reg_3_ ( .D(pc8[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[3]) );
  DFC3 pipe_data_pc8_reg_2_ ( .D(pc8[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[2]) );
  DFC3 pipe_data_pc8_reg_1_ ( .D(pc8[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[1]) );
  DFC3 pipe_data_pc8_reg_0_ ( .D(pc8[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[0]) );
  DFC3 pipe_data_alures_reg_31_ ( .D(i_data_alures[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[31]) );
  DFC3 pipe_data_alures_reg_30_ ( .D(i_data_alures[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[30]) );
  DFC3 pipe_data_alures_reg_29_ ( .D(i_data_alures[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[29]) );
  DFC3 pipe_data_alures_reg_28_ ( .D(i_data_alures[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[28]) );
  DFC3 pipe_data_alures_reg_27_ ( .D(i_data_alures[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[27]) );
  DFC3 pipe_data_alures_reg_26_ ( .D(i_data_alures[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[26]) );
  DFC3 pipe_data_alures_reg_25_ ( .D(i_data_alures[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[25]) );
  DFC3 pipe_data_alures_reg_24_ ( .D(i_data_alures[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[24]) );
  DFC3 pipe_data_alures_reg_23_ ( .D(i_data_alures[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[23]) );
  DFC3 pipe_data_alures_reg_22_ ( .D(i_data_alures[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[22]) );
  DFC3 pipe_data_alures_reg_21_ ( .D(i_data_alures[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[21]) );
  DFC3 pipe_data_alures_reg_20_ ( .D(i_data_alures[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[20]) );
  DFC3 pipe_data_alures_reg_19_ ( .D(i_data_alures[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[19]) );
  DFC3 pipe_data_alures_reg_18_ ( .D(i_data_alures[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[18]) );
  DFC3 pipe_data_alures_reg_17_ ( .D(i_data_alures[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[17]) );
  DFC3 pipe_data_alures_reg_16_ ( .D(i_data_alures[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[16]) );
  DFC3 pipe_data_alures_reg_15_ ( .D(i_data_alures[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[15]) );
  DFC3 pipe_data_alures_reg_14_ ( .D(i_data_alures[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[14]) );
  DFC3 pipe_data_alures_reg_13_ ( .D(i_data_alures[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[13]) );
  DFC3 pipe_data_alures_reg_12_ ( .D(i_data_alures[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[12]) );
  DFC3 pipe_data_alures_reg_11_ ( .D(i_data_alures[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[11]) );
  DFC3 pipe_data_alures_reg_10_ ( .D(i_data_alures[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[10]) );
  DFC3 pipe_data_alures_reg_9_ ( .D(i_data_alures[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC3 pipe_data_alures_reg_8_ ( .D(i_data_alures[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC3 pipe_data_alures_reg_7_ ( .D(i_data_alures[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC3 pipe_data_alures_reg_6_ ( .D(i_data_alures[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC3 pipe_data_alures_reg_5_ ( .D(i_data_alures[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC3 pipe_data_alures_reg_4_ ( .D(i_data_alures[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC3 pipe_data_alures_reg_3_ ( .D(i_data_alures[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC3 pipe_data_alures_reg_2_ ( .D(i_data_alures[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC3 pipe_data_alures_reg_1_ ( .D(i_data_alures[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC3 pipe_data_alures_reg_0_ ( .D(i_data_alures[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC3 pipe_data_memout_reg_31_ ( .D(i_data_memout[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[31]) );
  DFC3 pipe_data_memout_reg_30_ ( .D(i_data_memout[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[30]) );
  DFC3 pipe_data_memout_reg_29_ ( .D(i_data_memout[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[29]) );
  DFC3 pipe_data_memout_reg_28_ ( .D(i_data_memout[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[28]) );
  DFC3 pipe_data_memout_reg_27_ ( .D(i_data_memout[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[27]) );
  DFC3 pipe_data_memout_reg_26_ ( .D(i_data_memout[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[26]) );
  DFC3 pipe_data_memout_reg_25_ ( .D(i_data_memout[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[25]) );
  DFC3 pipe_data_memout_reg_24_ ( .D(i_data_memout[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[24]) );
  DFC3 pipe_data_memout_reg_23_ ( .D(i_data_memout[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[23]) );
  DFC3 pipe_data_memout_reg_22_ ( .D(i_data_memout[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[22]) );
  DFC3 pipe_data_memout_reg_21_ ( .D(i_data_memout[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[21]) );
  DFC3 pipe_data_memout_reg_20_ ( .D(i_data_memout[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[20]) );
  DFC3 pipe_data_memout_reg_19_ ( .D(i_data_memout[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[19]) );
  DFC3 pipe_data_memout_reg_18_ ( .D(i_data_memout[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[18]) );
  DFC3 pipe_data_memout_reg_17_ ( .D(i_data_memout[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[17]) );
  DFC3 pipe_data_memout_reg_16_ ( .D(i_data_memout[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[16]) );
  DFC3 pipe_data_memout_reg_15_ ( .D(i_data_memout[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[15]) );
  DFC3 pipe_data_memout_reg_14_ ( .D(i_data_memout[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[14]) );
  DFC3 pipe_data_memout_reg_13_ ( .D(i_data_memout[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[13]) );
  DFC3 pipe_data_memout_reg_12_ ( .D(i_data_memout[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[12]) );
  DFC3 pipe_data_memout_reg_11_ ( .D(i_data_memout[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[11]) );
  DFC3 pipe_data_memout_reg_10_ ( .D(i_data_memout[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[10]) );
  DFC3 pipe_data_memout_reg_9_ ( .D(i_data_memout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[9]) );
  DFC3 pipe_data_memout_reg_8_ ( .D(i_data_memout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[8]) );
  DFC3 pipe_data_memout_reg_7_ ( .D(i_data_memout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[7]) );
  DFC3 pipe_data_memout_reg_6_ ( .D(i_data_memout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[6]) );
  DFC3 pipe_data_memout_reg_5_ ( .D(i_data_memout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[5]) );
  DFC3 pipe_data_memout_reg_4_ ( .D(i_data_memout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[4]) );
  DFC3 pipe_data_memout_reg_3_ ( .D(i_data_memout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[3]) );
  DFC3 pipe_data_memout_reg_2_ ( .D(i_data_memout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[2]) );
  DFC3 pipe_data_memout_reg_1_ ( .D(i_data_memout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[1]) );
  DFC3 pipe_data_memout_reg_0_ ( .D(i_data_memout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[0]) );
  DFC3 pipe_addr_regdst_reg_4_ ( .D(i_addr_regdst[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[4]) );
  DFC3 pipe_addr_regdst_reg_3_ ( .D(i_addr_regdst[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[3]) );
  DFC3 pipe_addr_regdst_reg_2_ ( .D(i_addr_regdst[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[2]) );
  DFC3 pipe_addr_regdst_reg_1_ ( .D(i_addr_regdst[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[1]) );
  DFC3 pipe_addr_regdst_reg_0_ ( .D(i_addr_regdst[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[0]) );
  DFC3 pipe_con_Wloadmux_reg_1_ ( .D(i_con_Wloadmux[1]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[1]) );
  DFC3 pipe_con_Wloadmux_reg_0_ ( .D(i_con_Wloadmux[0]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[0]) );
  DFC3 pipe_con_Walupc8_reg ( .D(i_con_Walupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Walupc8) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_con_FWmemread_reg ( .D(i_con_FWmemread), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_FWmemread) );
  mem_DW01_add_1 add_31 ( .A(i_data_pc4), .B({n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic1_, n_Logic0_, n_Logic0_}), .CI(n_Logic0_), .SUM(pc8) );
  LOGIC0 U3 ( .Q(n_Logic0_) );
  LOGIC1 U4 ( .Q(n_Logic1_) );
endmodule


module W_resmux ( i_data_alures, i_data_pc8, i_con_pc8, o_data_alu );
  input [31:0] i_data_alures;
  input [31:0] i_data_pc8;
  output [31:0] o_data_alu;
  input i_con_pc8;
  wire   n1, n2;

  MUX22 U1 ( .A(i_data_alures[7]), .B(i_data_pc8[7]), .S(n1), .Q(o_data_alu[7]) );
  MUX21 U2 ( .A(i_data_alures[16]), .B(i_data_pc8[16]), .S(i_con_pc8), .Q(
        o_data_alu[16]) );
  MUX21 U3 ( .A(i_data_alures[15]), .B(i_data_pc8[15]), .S(i_con_pc8), .Q(
        o_data_alu[15]) );
  MUX21 U4 ( .A(i_data_alures[13]), .B(i_data_pc8[13]), .S(i_con_pc8), .Q(
        o_data_alu[13]) );
  MUX21 U5 ( .A(i_data_alures[14]), .B(i_data_pc8[14]), .S(i_con_pc8), .Q(
        o_data_alu[14]) );
  MUX21 U6 ( .A(i_data_alures[22]), .B(i_data_pc8[22]), .S(n2), .Q(
        o_data_alu[22]) );
  MUX21 U7 ( .A(i_data_alures[19]), .B(i_data_pc8[19]), .S(i_con_pc8), .Q(
        o_data_alu[19]) );
  MUX21 U8 ( .A(i_data_alures[23]), .B(i_data_pc8[23]), .S(i_con_pc8), .Q(
        o_data_alu[23]) );
  MUX21 U9 ( .A(i_data_alures[24]), .B(i_data_pc8[24]), .S(n2), .Q(
        o_data_alu[24]) );
  MUX21 U10 ( .A(i_data_alures[25]), .B(i_data_pc8[25]), .S(i_con_pc8), .Q(
        o_data_alu[25]) );
  MUX21 U11 ( .A(i_data_alures[0]), .B(i_data_pc8[0]), .S(n1), .Q(
        o_data_alu[0]) );
  MUX21 U12 ( .A(i_data_alures[1]), .B(i_data_pc8[1]), .S(n1), .Q(
        o_data_alu[1]) );
  MUX21 U13 ( .A(i_data_alures[8]), .B(i_data_pc8[8]), .S(n1), .Q(
        o_data_alu[8]) );
  MUX21 U14 ( .A(i_data_alures[11]), .B(i_data_pc8[11]), .S(n1), .Q(
        o_data_alu[11]) );
  MUX21 U15 ( .A(i_data_alures[12]), .B(i_data_pc8[12]), .S(n1), .Q(
        o_data_alu[12]) );
  MUX21 U16 ( .A(i_data_alures[3]), .B(i_data_pc8[3]), .S(n1), .Q(
        o_data_alu[3]) );
  MUX21 U17 ( .A(i_data_alures[4]), .B(i_data_pc8[4]), .S(n1), .Q(
        o_data_alu[4]) );
  MUX21 U18 ( .A(i_data_alures[2]), .B(i_data_pc8[2]), .S(n1), .Q(
        o_data_alu[2]) );
  MUX21 U19 ( .A(i_data_alures[5]), .B(i_data_pc8[5]), .S(n1), .Q(
        o_data_alu[5]) );
  MUX21 U20 ( .A(i_data_alures[6]), .B(i_data_pc8[6]), .S(n1), .Q(
        o_data_alu[6]) );
  MUX22 U21 ( .A(i_data_alures[17]), .B(i_data_pc8[17]), .S(i_con_pc8), .Q(
        o_data_alu[17]) );
  MUX22 U22 ( .A(i_data_alures[18]), .B(i_data_pc8[18]), .S(i_con_pc8), .Q(
        o_data_alu[18]) );
  MUX22 U23 ( .A(i_data_alures[20]), .B(i_data_pc8[20]), .S(n2), .Q(
        o_data_alu[20]) );
  BUF2 U24 ( .A(i_con_pc8), .Q(n1) );
  MUX22 U25 ( .A(i_data_alures[21]), .B(i_data_pc8[21]), .S(n2), .Q(
        o_data_alu[21]) );
  MUX22 U26 ( .A(i_data_alures[9]), .B(i_data_pc8[9]), .S(n1), .Q(
        o_data_alu[9]) );
  MUX22 U27 ( .A(i_data_alures[10]), .B(i_data_pc8[10]), .S(n1), .Q(
        o_data_alu[10]) );
  BUF2 U28 ( .A(i_con_pc8), .Q(n2) );
  MUX22 U29 ( .A(i_data_alures[26]), .B(i_data_pc8[26]), .S(n2), .Q(
        o_data_alu[26]) );
  MUX22 U30 ( .A(i_data_alures[27]), .B(i_data_pc8[27]), .S(n2), .Q(
        o_data_alu[27]) );
  MUX22 U31 ( .A(i_data_alures[28]), .B(i_data_pc8[28]), .S(n2), .Q(
        o_data_alu[28]) );
  MUX22 U32 ( .A(i_data_alures[29]), .B(i_data_pc8[29]), .S(n2), .Q(
        o_data_alu[29]) );
  MUX22 U33 ( .A(i_data_alures[30]), .B(i_data_pc8[30]), .S(n2), .Q(
        o_data_alu[30]) );
  MUX22 U34 ( .A(i_data_alures[31]), .B(i_data_pc8[31]), .S(n2), .Q(
        o_data_alu[31]) );
endmodule


module W_loadmux3 ( i_data_Rdata, i_con_loadsig, o_data_Wdata );
  input [31:0] i_data_Rdata;
  input [1:0] i_con_loadsig;
  output [31:0] o_data_Wdata;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50;

  NAND20 U2 ( .A(n50), .B(n47), .Q(o_data_Wdata[30]) );
  NAND20 U3 ( .A(n50), .B(n43), .Q(o_data_Wdata[26]) );
  NAND20 U4 ( .A(n50), .B(n45), .Q(o_data_Wdata[28]) );
  NAND20 U5 ( .A(n50), .B(n42), .Q(o_data_Wdata[25]) );
  NAND20 U6 ( .A(n50), .B(n44), .Q(o_data_Wdata[27]) );
  NAND20 U7 ( .A(n50), .B(n49), .Q(o_data_Wdata[31]) );
  NAND20 U8 ( .A(n50), .B(n40), .Q(o_data_Wdata[23]) );
  NAND20 U9 ( .A(n50), .B(n39), .Q(o_data_Wdata[22]) );
  NAND20 U10 ( .A(n50), .B(n37), .Q(o_data_Wdata[20]) );
  NAND20 U11 ( .A(n50), .B(n46), .Q(o_data_Wdata[29]) );
  NAND20 U12 ( .A(n50), .B(n38), .Q(o_data_Wdata[21]) );
  NAND20 U13 ( .A(n50), .B(n41), .Q(o_data_Wdata[24]) );
  INV3 U14 ( .A(n1), .Q(n2) );
  INV6 U15 ( .A(n26), .Q(n3) );
  INV6 U16 ( .A(n33), .Q(n50) );
  INV3 U17 ( .A(i_con_loadsig[1]), .Q(n5) );
  NAND22 U18 ( .A(n26), .B(n27), .Q(n4) );
  NAND22 U19 ( .A(i_data_Rdata[15]), .B(n28), .Q(n32) );
  INV3 U20 ( .A(n27), .Q(n28) );
  NAND22 U21 ( .A(n50), .B(n34), .Q(o_data_Wdata[17]) );
  NOR21 U22 ( .A(n15), .B(n14), .Q(o_data_Wdata[7]) );
  CLKIN3 U23 ( .A(n26), .Q(n48) );
  NAND22 U24 ( .A(n25), .B(i_con_loadsig[0]), .Q(n13) );
  NAND21 U25 ( .A(i_con_loadsig[1]), .B(i_data_Rdata[7]), .Q(n1) );
  NAND22 U26 ( .A(n32), .B(n31), .Q(n33) );
  NAND22 U27 ( .A(n31), .B(n30), .Q(o_data_Wdata[16]) );
  NAND23 U28 ( .A(n16), .B(n2), .Q(n31) );
  NAND22 U29 ( .A(n5), .B(n16), .Q(n26) );
  NAND20 U30 ( .A(n31), .B(n22), .Q(o_data_Wdata[13]) );
  NAND20 U31 ( .A(n31), .B(n19), .Q(o_data_Wdata[10]) );
  NAND20 U32 ( .A(n31), .B(n17), .Q(o_data_Wdata[8]) );
  NAND20 U33 ( .A(n31), .B(n23), .Q(o_data_Wdata[14]) );
  NAND20 U34 ( .A(n31), .B(n21), .Q(o_data_Wdata[12]) );
  NAND20 U35 ( .A(n31), .B(n20), .Q(o_data_Wdata[11]) );
  NAND20 U36 ( .A(n31), .B(n18), .Q(o_data_Wdata[9]) );
  NAND22 U37 ( .A(i_con_loadsig[0]), .B(n5), .Q(n27) );
  AOI212 U38 ( .A(i_data_Rdata[16]), .B(n48), .C(n29), .Q(n30) );
  INV0 U39 ( .A(i_data_Rdata[7]), .Q(n14) );
  INV0 U40 ( .A(i_data_Rdata[15]), .Q(n24) );
  INV3 U41 ( .A(n32), .Q(n29) );
  CLKIN6 U42 ( .A(i_con_loadsig[0]), .Q(n16) );
  NAND21 U43 ( .A(i_data_Rdata[30]), .B(n3), .Q(n47) );
  NAND21 U44 ( .A(i_data_Rdata[29]), .B(n3), .Q(n46) );
  NAND21 U45 ( .A(i_data_Rdata[26]), .B(n3), .Q(n43) );
  NAND21 U46 ( .A(i_data_Rdata[28]), .B(n3), .Q(n45) );
  NAND21 U47 ( .A(i_data_Rdata[25]), .B(n3), .Q(n42) );
  NAND21 U48 ( .A(i_data_Rdata[27]), .B(n3), .Q(n44) );
  NAND21 U49 ( .A(i_data_Rdata[31]), .B(n3), .Q(n49) );
  NAND21 U50 ( .A(i_data_Rdata[24]), .B(n3), .Q(n41) );
  NAND21 U51 ( .A(i_data_Rdata[23]), .B(n3), .Q(n40) );
  NAND21 U52 ( .A(i_data_Rdata[22]), .B(n3), .Q(n39) );
  NAND21 U53 ( .A(i_data_Rdata[21]), .B(n3), .Q(n38) );
  NAND21 U54 ( .A(i_data_Rdata[20]), .B(n3), .Q(n37) );
  NAND21 U55 ( .A(i_data_Rdata[19]), .B(n3), .Q(n36) );
  NAND21 U56 ( .A(i_data_Rdata[18]), .B(n3), .Q(n35) );
  NAND21 U57 ( .A(i_data_Rdata[17]), .B(n3), .Q(n34) );
  OAI210 U58 ( .A(n25), .B(n24), .C(n31), .Q(o_data_Wdata[15]) );
  NAND21 U59 ( .A(n50), .B(n36), .Q(o_data_Wdata[19]) );
  NAND21 U60 ( .A(n50), .B(n35), .Q(o_data_Wdata[18]) );
  CLKIN3 U61 ( .A(n4), .Q(n25) );
  NAND22 U62 ( .A(i_data_Rdata[0]), .B(n13), .Q(n6) );
  CLKIN3 U63 ( .A(n6), .Q(o_data_Wdata[0]) );
  NAND22 U64 ( .A(i_data_Rdata[1]), .B(n13), .Q(n7) );
  CLKIN3 U65 ( .A(n7), .Q(o_data_Wdata[1]) );
  NAND22 U66 ( .A(i_data_Rdata[2]), .B(n13), .Q(n8) );
  CLKIN3 U67 ( .A(n8), .Q(o_data_Wdata[2]) );
  NAND22 U68 ( .A(i_data_Rdata[3]), .B(n13), .Q(n9) );
  CLKIN3 U69 ( .A(n9), .Q(o_data_Wdata[3]) );
  NAND22 U70 ( .A(i_data_Rdata[4]), .B(n13), .Q(n10) );
  CLKIN3 U71 ( .A(n10), .Q(o_data_Wdata[4]) );
  NAND22 U72 ( .A(i_data_Rdata[5]), .B(n13), .Q(n11) );
  CLKIN3 U73 ( .A(n11), .Q(o_data_Wdata[5]) );
  NAND22 U74 ( .A(i_data_Rdata[6]), .B(n13), .Q(n12) );
  CLKIN3 U75 ( .A(n12), .Q(o_data_Wdata[6]) );
  CLKIN3 U76 ( .A(n13), .Q(n15) );
  NAND22 U77 ( .A(i_data_Rdata[8]), .B(n4), .Q(n17) );
  NAND22 U78 ( .A(i_data_Rdata[9]), .B(n4), .Q(n18) );
  NAND22 U79 ( .A(i_data_Rdata[10]), .B(n4), .Q(n19) );
  NAND22 U80 ( .A(i_data_Rdata[11]), .B(n4), .Q(n20) );
  NAND22 U81 ( .A(i_data_Rdata[12]), .B(n4), .Q(n21) );
  NAND22 U82 ( .A(i_data_Rdata[13]), .B(n4), .Q(n22) );
  NAND22 U83 ( .A(i_data_Rdata[14]), .B(n4), .Q(n23) );
endmodule


module W_datamux ( i_data_alu, i_data_load, i_con_memtoreg, o_data_toreg );
  input [31:0] i_data_alu;
  input [31:0] i_data_load;
  output [31:0] o_data_toreg;
  input i_con_memtoreg;
  wire   n1, n2, n3, n4, n5, n6;

  MUX22 U1 ( .A(i_data_alu[24]), .B(i_data_load[24]), .S(n1), .Q(
        o_data_toreg[24]) );
  MUX22 U2 ( .A(i_data_alu[23]), .B(i_data_load[23]), .S(n1), .Q(
        o_data_toreg[23]) );
  MUX22 U3 ( .A(i_data_alu[28]), .B(i_data_load[28]), .S(n1), .Q(
        o_data_toreg[28]) );
  MUX22 U4 ( .A(i_data_alu[7]), .B(i_data_load[7]), .S(n1), .Q(o_data_toreg[7]) );
  AOI221 U5 ( .A(i_data_load[16]), .B(n2), .C(i_data_alu[16]), .D(n3), .Q(n4)
         );
  INV3 U6 ( .A(i_con_memtoreg), .Q(n3) );
  CLKIN3 U7 ( .A(n3), .Q(n2) );
  MUX22 U8 ( .A(i_data_alu[4]), .B(i_data_load[4]), .S(n2), .Q(o_data_toreg[4]) );
  MUX21 U9 ( .A(i_data_alu[3]), .B(i_data_load[3]), .S(n2), .Q(o_data_toreg[3]) );
  MUX22 U10 ( .A(i_data_alu[2]), .B(i_data_load[2]), .S(n2), .Q(
        o_data_toreg[2]) );
  AOI221 U11 ( .A(i_data_load[18]), .B(n2), .C(i_data_alu[18]), .D(n3), .Q(n6)
         );
  MUX22 U12 ( .A(i_data_alu[0]), .B(i_data_load[0]), .S(n1), .Q(
        o_data_toreg[0]) );
  MUX21 U13 ( .A(i_data_alu[15]), .B(i_data_load[15]), .S(n2), .Q(
        o_data_toreg[15]) );
  MUX21 U14 ( .A(i_data_alu[11]), .B(i_data_load[11]), .S(n2), .Q(
        o_data_toreg[11]) );
  MUX21 U15 ( .A(i_data_alu[12]), .B(i_data_load[12]), .S(n2), .Q(
        o_data_toreg[12]) );
  MUX21 U16 ( .A(i_data_alu[13]), .B(i_data_load[13]), .S(n2), .Q(
        o_data_toreg[13]) );
  MUX21 U17 ( .A(i_data_alu[14]), .B(i_data_load[14]), .S(i_con_memtoreg), .Q(
        o_data_toreg[14]) );
  MUX21 U18 ( .A(i_data_alu[22]), .B(i_data_load[22]), .S(n1), .Q(
        o_data_toreg[22]) );
  MUX21 U19 ( .A(i_data_alu[20]), .B(i_data_load[20]), .S(n1), .Q(
        o_data_toreg[20]) );
  MUX21 U20 ( .A(i_data_alu[5]), .B(i_data_load[5]), .S(n2), .Q(
        o_data_toreg[5]) );
  MUX21 U21 ( .A(i_data_alu[6]), .B(i_data_load[6]), .S(n1), .Q(
        o_data_toreg[6]) );
  MUX21 U22 ( .A(i_data_alu[25]), .B(i_data_load[25]), .S(n1), .Q(
        o_data_toreg[25]) );
  MUX21 U23 ( .A(i_data_alu[26]), .B(i_data_load[26]), .S(n1), .Q(
        o_data_toreg[26]) );
  MUX21 U24 ( .A(i_data_alu[27]), .B(i_data_load[27]), .S(n1), .Q(
        o_data_toreg[27]) );
  MUX21 U25 ( .A(i_data_alu[29]), .B(i_data_load[29]), .S(n1), .Q(
        o_data_toreg[29]) );
  MUX21 U26 ( .A(i_data_alu[30]), .B(i_data_load[30]), .S(n1), .Q(
        o_data_toreg[30]) );
  MUX21 U27 ( .A(i_data_alu[31]), .B(i_data_load[31]), .S(n1), .Q(
        o_data_toreg[31]) );
  INV3 U28 ( .A(n3), .Q(n1) );
  INV3 U29 ( .A(n4), .Q(o_data_toreg[16]) );
  MUX22 U30 ( .A(i_data_alu[1]), .B(i_data_load[1]), .S(n1), .Q(
        o_data_toreg[1]) );
  MUX22 U31 ( .A(i_data_alu[19]), .B(i_data_load[19]), .S(n1), .Q(
        o_data_toreg[19]) );
  MUX22 U32 ( .A(i_data_alu[8]), .B(i_data_load[8]), .S(n2), .Q(
        o_data_toreg[8]) );
  MUX22 U33 ( .A(i_data_alu[21]), .B(i_data_load[21]), .S(n1), .Q(
        o_data_toreg[21]) );
  MUX22 U34 ( .A(i_data_alu[9]), .B(i_data_load[9]), .S(n2), .Q(
        o_data_toreg[9]) );
  MUX22 U35 ( .A(i_data_alu[10]), .B(i_data_load[10]), .S(n2), .Q(
        o_data_toreg[10]) );
  AOI222 U36 ( .A(i_data_load[17]), .B(n2), .C(i_data_alu[17]), .D(n3), .Q(n5)
         );
  CLKIN3 U37 ( .A(n5), .Q(o_data_toreg[17]) );
  CLKIN3 U38 ( .A(n6), .Q(o_data_toreg[18]) );
endmodule


module writeback ( i_data_pc8, i_data_alures, i_data_memout, i_con_Wloadmux, 
        i_con_Walupc8, i_con_Wmemtoreg, o_data_regwrite );
  input [31:0] i_data_pc8;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [1:0] i_con_Wloadmux;
  output [31:0] o_data_regwrite;
  input i_con_Walupc8, i_con_Wmemtoreg;

  wire   [31:0] datamux_i_data_alu;
  wire   [31:0] datamux_i_data_load;

  W_resmux u_resmux ( .i_data_alures(i_data_alures), .i_data_pc8(i_data_pc8), 
        .i_con_pc8(i_con_Walupc8), .o_data_alu(datamux_i_data_alu) );
  W_loadmux3 u_loadmux ( .i_data_Rdata(i_data_memout), .i_con_loadsig(
        i_con_Wloadmux), .o_data_Wdata(datamux_i_data_load) );
  W_datamux u_datamux ( .i_data_alu(datamux_i_data_alu), .i_data_load(
        datamux_i_data_load), .i_con_memtoreg(i_con_Wmemtoreg), .o_data_toreg(
        o_data_regwrite) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Mmemread, ex_con_Mmemwrite, ex_con_Walupc8, ex_con_Wmemtoreg,
         mem_con_Walupc8, mem_con_Wmemtoreg, wb_con_Walupc8, wb_con_Wmemtoreg,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2;
  wire   [31:0] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [31:0] id_addr_pc4;
  wire   [31:0] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [1:0] ex_con_Wloadmux;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] wb_data_memout;
  wire   [31:0] mem_data_pc4;
  wire   [1:0] mem_con_Wloadmux;
  wire   [31:0] wb_data_pc8;
  wire   [31:0] mem_data_alures;
  wire   [1:0] wb_con_Wloadmux;

  fetch u_fetch ( .i_clk(clk), .i_nrst(rst_n), .i_addr_b(if_addr_b), 
        .i_addr_j({if_addr_j, n1, n1}), .i_addr_jr(id_data_jr), .i_con_b(
        if_con_b), .i_con_j(if_con_j), .i_data_instr(read_instruction), 
        .i_con_ifstall(if_con_ifstall), .o_addr_pc(instruction_address), 
        .o_addr_pc4(id_addr_pc4), .o_data_instr(id_data_instr) );
  decode u_decode ( .i_clk(clk), .i_nrst(rst_n), .i_addr_pc4(id_addr_pc4), 
        .i_data_instr(id_data_instr), .i_con_Wregwrite(id_con_Wregwrite), 
        .i_data_Wregwrite({n16, n15, n14, id_data_Wregwrite[28:27], n13, n12, 
        id_data_Wregwrite[24:23], n11, id_data_Wregwrite[21], n10, n9, n8, 
        id_data_Wregwrite[17:15], n7, n6, id_data_Wregwrite[12], n5, 
        id_data_Wregwrite[10:9], n4, id_data_Wregwrite[7], n3, n2, 
        id_data_Wregwrite[4:0]}), .i_addr_Wregwrite(id_addr_Wregwrite), 
        .i_addr_Erd(for_o_addr_Erd), .i_addr_Mrd(mem_addr_regdst), 
        .i_con_Eregwrite(ex_con_Wregwrite), .i_con_Mregwrite(mem_con_Wregwrite), .i_addr_rtM(for_addr_rtM), .i_addr_rtW(for_addr_rtW), .i_con_memreadM(
        mem_read), .i_con_memreadW(for_FWmemread), .o_data_rs(id_data_rs), 
        .o_data_rt(ex_data_rt), .o_addr_rd(ex_addr_rd), .o_addr_rt(ex_addr_rt), 
        .o_data_jr(id_data_jr), .o_con_jump(if_con_j), .o_addr_pc4(ex_data_pc4), .o_addr_branch(if_addr_b), .o_addr_jump({if_addr_j, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .o_con_Ealuop(ex_con_Ealuop), 
        .o_con_Ealusrc(ex_con_Ealusrc), .o_con_Eregdst(ex_con_Eregdst), 
        .o_con_Mmemread(ex_con_Mmemread), .o_con_Mmemwrite(ex_con_Mmemwrite), 
        .o_con_Wloadmux(ex_con_Wloadmux), .o_con_Walupc8(ex_con_Walupc8), 
        .o_con_Wmemtoreg(ex_con_Wmemtoreg), .o_con_Wregwrite(ex_con_Wregwrite), 
        .o_con_ifstall(if_con_ifstall), .o_con_Ebop(ex_con_bop), 
        .o_data_signext(ex_data_immext), .o_con_Efamux(for_o_con_Efamux), 
        .o_con_Efbmux(for_o_con_Efbmux), .o_data_Fmemout(for_memout) );
  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext(
        ex_data_immext), .i_addr_rt(ex_addr_rt), .i_addr_rd(ex_addr_rd), 
        .i_data_FEalures(data_address), .i_data_FMalures({n16, n15, n14, 
        id_data_Wregwrite[28:27], n13, n12, id_data_Wregwrite[24:23], n11, 
        id_data_Wregwrite[21], n10, n9, n8, id_data_Wregwrite[17:15], n7, n6, 
        id_data_Wregwrite[12], n5, id_data_Wregwrite[10:9], n4, 
        id_data_Wregwrite[7], n3, n2, id_data_Wregwrite[4:0]}), 
        .i_data_FMmemout(wb_data_memout), .i_data_FWmemout(for_memout), 
        .i_con_Ealuop(ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), 
        .i_con_Mmemwrite(ex_con_Mmemwrite), .i_con_Wloadmux(ex_con_Wloadmux), 
        .i_con_Walupc8(ex_con_Walupc8), .i_con_Wmemtoreg(ex_con_Wmemtoreg), 
        .i_con_Wregwrite(ex_con_Wregwrite), .i_con_Efamux(for_o_con_Efamux), 
        .i_con_Efbmux(for_o_con_Efbmux), .i_con_bop(ex_con_bop), .o_data_pc4(
        mem_data_pc4), .o_data_alures(data_address), .o_data_rt(write_data), 
        .o_addr_regdst(mem_addr_regdst), .o_con_Mmemread(mem_read), 
        .o_con_Mmemwrite(mem_write), .o_con_Wloadmux(mem_con_Wloadmux), 
        .o_con_Walupc8(mem_con_Walupc8), .o_con_Wmemtoreg(mem_con_Wmemtoreg), 
        .o_con_Wregwrite(mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), 
        .o_addr_Mrt(for_addr_rtM), .o_con_ifbranch(if_con_b) );
  mem u_mem ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(mem_data_pc4), 
        .i_data_alures(data_address), .i_data_memout(read_data), 
        .i_addr_regdst(mem_addr_regdst), .i_con_Wloadmux(mem_con_Wloadmux), 
        .i_con_Walupc8(mem_con_Walupc8), .i_con_Wmemtoreg(mem_con_Wmemtoreg), 
        .i_con_Wregwrite(mem_con_Wregwrite), .i_con_FWmemread(ex_con_Mmemread), 
        .i_addr_Mrt(for_addr_rtM), .o_data_pc8(wb_data_pc8), .o_data_alures(
        mem_data_alures), .o_data_memout(wb_data_memout), .o_addr_regdst(
        id_addr_Wregwrite), .o_con_Wloadmux(wb_con_Wloadmux), .o_con_Walupc8(
        wb_con_Walupc8), .o_con_Wmemtoreg(wb_con_Wmemtoreg), .o_con_Wregwrite(
        id_con_Wregwrite), .o_con_FWmemread(for_FWmemread), .o_addr_Wrt(
        for_addr_rtW) );
  writeback u_writeback ( .i_data_pc8(wb_data_pc8), .i_data_alures(
        mem_data_alures), .i_data_memout(wb_data_memout), .i_con_Wloadmux(
        wb_con_Wloadmux), .i_con_Walupc8(wb_con_Walupc8), .i_con_Wmemtoreg(
        wb_con_Wmemtoreg), .o_data_regwrite(id_data_Wregwrite) );
  BUF8 U1 ( .A(id_data_Wregwrite[18]), .Q(n8) );
  BUF6 U2 ( .A(id_data_Wregwrite[8]), .Q(n4) );
  BUF6 U3 ( .A(id_data_Wregwrite[19]), .Q(n9) );
  BUF6 U4 ( .A(id_data_Wregwrite[20]), .Q(n10) );
  BUF2 U5 ( .A(id_data_Wregwrite[5]), .Q(n2) );
  BUF2 U6 ( .A(id_data_Wregwrite[6]), .Q(n3) );
  BUF2 U7 ( .A(id_data_Wregwrite[22]), .Q(n11) );
  BUF2 U8 ( .A(id_data_Wregwrite[11]), .Q(n5) );
  BUF2 U9 ( .A(id_data_Wregwrite[13]), .Q(n6) );
  BUF2 U10 ( .A(id_data_Wregwrite[14]), .Q(n7) );
  BUF2 U11 ( .A(id_data_Wregwrite[25]), .Q(n12) );
  BUF2 U12 ( .A(id_data_Wregwrite[26]), .Q(n13) );
  BUF2 U13 ( .A(id_data_Wregwrite[29]), .Q(n14) );
  BUF2 U14 ( .A(id_data_Wregwrite[30]), .Q(n15) );
  BUF2 U15 ( .A(id_data_Wregwrite[31]), .Q(n16) );
  LOGIC0 U16 ( .Q(n1) );
endmodule

