`timescale 1ns / 1ps
module D_compare