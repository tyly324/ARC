`timescale 1ns / 1ps
module D_unsign_extend