module decode();