
module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Efamux, i_con_Efbmux, 
        i_con_Ealuop, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread, 
        i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_bop, o_data_pc4, o_data_alures, o_data_rt, o_addr_regdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_addr_Erd, o_addr_Mrt, o_con_ifbranch );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [5:0] i_con_Ealuop;
  input [2:0] i_con_bop;
  output [31:0] o_data_pc4;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch;
  wire   u_alu_N306, u_alu_DP_OP_83J3_124_3384_n154,
         u_alu_DP_OP_84J3_125_2615_n145, u_alu_DP_OP_84J3_125_2615_n140,
         u_alu_DP_OP_84J3_125_2615_n137, u_alu_DP_OP_84J3_125_2615_n136,
         u_alu_DP_OP_84J3_125_2615_n134, u_alu_DP_OP_84J3_125_2615_n111,
         u_alu_DP_OP_84J3_125_2615_n109, u_alu_DP_OP_84J3_125_2615_n108,
         u_alu_DP_OP_84J3_125_2615_n95, u_alu_DP_OP_84J3_125_2615_n92,
         u_alu_DP_OP_84J3_125_2615_n91, u_alu_DP_OP_84J3_125_2615_n90,
         u_alu_DP_OP_84J3_125_2615_n89, u_alu_DP_OP_84J3_125_2615_n86,
         u_alu_DP_OP_84J3_125_2615_n81, u_alu_DP_OP_84J3_125_2615_n80,
         u_alu_DP_OP_84J3_125_2615_n77, u_alu_DP_OP_84J3_125_2615_n73,
         u_alu_DP_OP_84J3_125_2615_n70, u_alu_DP_OP_84J3_125_2615_n68,
         u_alu_DP_OP_84J3_125_2615_n50, u_alu_DP_OP_84J3_125_2615_n49,
         u_alu_DP_OP_84J3_125_2615_n48, u_alu_DP_OP_84J3_125_2615_n46,
         u_alu_DP_OP_84J3_125_2615_n45, u_alu_DP_OP_84J3_125_2615_n40,
         u_alu_DP_OP_84J3_125_2615_n39, u_alu_DP_OP_84J3_125_2615_n37,
         u_alu_DP_OP_84J3_125_2615_n36, u_alu_DP_OP_84J3_125_2615_n33,
         u_alu_DP_OP_84J3_125_2615_n32, u_alu_DP_OP_84J3_125_2615_n31,
         u_alu_DP_OP_84J3_125_2615_n30, u_alu_DP_OP_84J3_125_2615_n23,
         u_alu_DP_OP_84J3_125_2615_n22, u_alu_DP_OP_84J3_125_2615_n18,
         u_alu_DP_OP_84J3_125_2615_n17, u_alu_DP_OP_84J3_125_2615_n16,
         u_alu_DP_OP_84J3_125_2615_n15, u_alu_DP_OP_84J3_125_2615_n14,
         u_alu_DP_OP_84J3_125_2615_n11, u_alu_DP_OP_84J3_125_2615_n7,
         u_alu_DP_OP_84J3_125_2615_n6, u_alu_DP_OP_84J3_125_2615_n5,
         u_alu_DP_OP_84J3_125_2615_n4, u_alu_DP_OP_84J3_125_2615_n3,
         u_alu_DP_OP_84J3_125_2615_n2, u_alu_DP_OP_84J3_125_2615_n1,
         u_alu_lt_x_11_A_23_, u_alu_lt_x_11_A_12_, u_alu_lt_x_11_A_10_,
         u_alu_lt_x_11_A_5_, u_alu_lt_x_11_A_3_, u_alu_lt_x_11_A_2_,
         u_alu_lt_x_11_A_0_, u_alu_lt_x_11_B_22_, u_alu_lt_x_11_B_21_,
         u_alu_lt_x_11_B_20_, u_alu_lt_x_11_B_19_, u_alu_lt_x_11_B_18_,
         u_alu_lt_x_11_B_17_, u_alu_lt_x_11_B_16_, u_alu_lt_x_11_B_15_,
         u_alu_lt_x_11_B_14_, u_alu_lt_x_11_B_13_, u_alu_lt_x_11_B_9_,
         u_alu_lt_x_11_B_8_, u_alu_lt_x_11_B_5_, u_alu_lt_x_11_B_1_,
         u_alu_lt_x_11_B_0_, u_alu_lt_x_11_n172, u_alu_lt_x_11_n171,
         u_alu_lt_x_11_n159, u_alu_lt_x_11_n143, u_alu_lt_x_11_n142,
         u_alu_lt_x_11_n140, u_alu_lt_x_11_n139, u_alu_lt_x_11_n138,
         u_alu_lt_x_11_n137, u_alu_lt_x_11_n136, u_alu_lt_x_11_n135,
         u_alu_lt_x_11_n134, u_alu_lt_x_11_n133, u_alu_lt_x_11_n131,
         u_alu_lt_x_11_n130, u_alu_lt_x_11_n129, u_alu_lt_x_11_n127,
         u_alu_lt_x_11_n126, u_alu_lt_x_11_n125, u_alu_lt_x_11_n124,
         u_alu_lt_x_11_n123, u_alu_lt_x_11_n122, u_alu_lt_x_11_n120,
         u_alu_lt_x_11_n119, u_alu_lt_x_11_n118, u_alu_lt_x_11_n117,
         u_alu_lt_x_11_n116, u_alu_lt_x_11_n115, u_alu_lt_x_11_n113,
         u_alu_lt_x_11_n112, u_alu_lt_x_11_n111, u_alu_lt_x_11_n110,
         u_alu_lt_x_11_n109, u_alu_lt_x_11_n108, u_alu_lt_x_11_n107,
         u_alu_lt_x_11_n106, u_alu_lt_x_11_n105, u_alu_lt_x_11_n104,
         u_alu_lt_x_11_n103, u_alu_lt_x_11_n101, u_alu_lt_x_11_n100,
         u_alu_lt_x_11_n99, u_alu_lt_x_11_n98, u_alu_lt_x_11_n97,
         u_alu_lt_x_11_n96, u_alu_lt_x_11_n94, u_alu_lt_x_11_n92,
         u_alu_lt_x_11_n91, u_alu_lt_x_11_n90, u_alu_lt_x_11_n87,
         u_alu_lt_x_11_n86, u_alu_lt_x_11_n85, u_alu_lt_x_11_n84,
         u_alu_lt_x_11_n83, u_alu_lt_x_11_n82, u_alu_lt_x_11_n81,
         u_alu_lt_x_11_n80, u_alu_lt_x_11_n79, u_alu_lt_x_11_n78,
         u_alu_lt_x_11_n77, u_alu_lt_x_11_n76, u_alu_lt_x_11_n75,
         u_alu_lt_x_11_n74, u_alu_lt_x_11_n73, u_alu_lt_x_11_n72,
         u_alu_lt_x_11_n71, u_alu_lt_x_11_n70, u_alu_lt_x_11_n69,
         u_alu_lt_x_11_n68, u_alu_lt_x_11_n67, u_alu_lt_x_11_n66,
         u_alu_lt_x_11_n65, u_alu_lt_x_11_n64, u_alu_lt_x_11_n63,
         u_alu_lt_x_11_n62, u_alu_lt_x_11_n61, u_alu_lt_x_11_n60,
         u_alu_lt_x_11_n59, u_alu_lt_x_11_n58, u_alu_lt_x_11_n57,
         u_alu_lt_x_11_n56, u_alu_lt_x_11_n55, u_alu_lt_x_11_n54,
         u_alu_lt_x_11_n52, u_alu_lt_x_11_n50, u_alu_lt_x_11_n49,
         u_alu_lt_x_11_n48, u_alu_lt_x_11_n47, u_alu_lt_x_11_n46,
         u_alu_lt_x_11_n45, u_alu_lt_x_11_n44, u_alu_lt_x_11_n43,
         u_alu_lt_x_11_n42, u_alu_lt_x_11_n41, u_alu_lt_x_11_n40,
         u_alu_lt_x_11_n39, u_alu_lt_x_11_n38, u_alu_lt_x_11_n37,
         u_alu_lt_x_11_n36, u_alu_lt_x_11_n35, u_alu_lt_x_11_n33,
         u_alu_lt_x_11_n31, u_alu_lt_x_11_n30, u_alu_lt_x_11_n29,
         u_alu_lt_x_11_n28, u_alu_lt_x_11_n27, u_alu_lt_x_11_n26,
         u_alu_lt_x_11_n24, u_alu_lt_x_11_n22, u_alu_lt_x_11_n21,
         u_alu_lt_x_11_n20, u_alu_lt_x_11_n19, u_alu_lt_x_11_n18,
         u_alu_lt_x_11_n17, u_alu_lt_x_11_n16, u_alu_lt_x_11_n15,
         u_alu_lt_x_11_n14, u_alu_lt_x_11_n13, u_alu_lt_x_11_n12,
         u_alu_lt_x_11_n11, u_alu_lt_x_11_n10, u_alu_lt_x_11_n9,
         u_alu_lt_x_11_n8, u_alu_lt_x_11_n7, u_alu_lt_x_11_n6,
         u_alu_lt_x_11_n5, u_alu_lt_x_11_n4, u_alu_lt_x_11_n3,
         u_alu_lt_x_11_n2, u_alu_lt_x_11_n1, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203;
  wire   [31:0] alu_o_data_AluRes;
  wire   [31:13] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:7] alu_i_data_B;
  wire   [7:1] u_alu_pre_sum_4b;
  wire   [7:0] u_alu_pre_sum_4a;

  DFC1 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC1 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC1 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC1 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC1 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC1 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[31]) );
  DFC1 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[30]) );
  DFC1 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[29]) );
  DFC1 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[28]) );
  DFC1 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[27]) );
  DFC1 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[26]) );
  DFC1 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[25]) );
  DFC1 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[24]) );
  DFC1 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[23]) );
  DFC1 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[22]) );
  DFC1 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[21]) );
  DFC1 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[20]) );
  DFC1 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[19]) );
  DFC1 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[18]) );
  DFC1 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[17]) );
  DFC1 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[16]) );
  DFC1 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[15]) );
  DFC1 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[14]) );
  DFC1 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[13]) );
  DFC1 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[12]) );
  DFC1 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[11]) );
  DFC1 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[10]) );
  DFC1 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[9]) );
  DFC1 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[8]) );
  DFC1 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[7]) );
  DFC1 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[6]) );
  DFC1 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[5]) );
  DFC1 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[4]) );
  DFC1 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[3]) );
  DFC1 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[2]) );
  DFC1 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[1]) );
  DFC1 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[0]) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  DFC1 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC1 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC1 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC1 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC1 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC1 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC1 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC1 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC1 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC1 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC1 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC1 pipe_alures_reg_15_ ( .D(n3196), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[15]) );
  DFC1 pipe_alures_reg_14_ ( .D(n3195), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[14]) );
  DFC1 pipe_alures_reg_13_ ( .D(n3194), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[13]) );
  DFC1 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC1 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC1 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC1 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC1 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC1 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC1 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC1 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC1 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC1 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC1 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC1 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC1 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC1 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC1 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC1 pipe_rt_reg_28_ ( .D(n1019), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28])
         );
  DFC1 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  DFC1 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC1 pipe_rt_reg_25_ ( .D(n565), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25])
         );
  DFC1 pipe_rt_reg_24_ ( .D(n3186), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24])
         );
  DFC1 pipe_rt_reg_23_ ( .D(n3183), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23])
         );
  DFC1 pipe_rt_reg_22_ ( .D(n3187), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22])
         );
  DFC1 pipe_rt_reg_21_ ( .D(n3190), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21])
         );
  DFC1 pipe_rt_reg_20_ ( .D(n3189), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20])
         );
  DFC1 pipe_rt_reg_19_ ( .D(n1325), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19])
         );
  DFC1 pipe_rt_reg_18_ ( .D(n3182), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18])
         );
  DFC1 pipe_rt_reg_17_ ( .D(n3180), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17])
         );
  DFC1 pipe_rt_reg_16_ ( .D(compare_i_data_rt[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[16]) );
  DFC1 pipe_rt_reg_15_ ( .D(n133), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15])
         );
  DFC1 pipe_rt_reg_14_ ( .D(n3193), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14])
         );
  DFC1 pipe_rt_reg_13_ ( .D(compare_i_data_rt[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[13]) );
  DFC1 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC1 pipe_rt_reg_11_ ( .D(n366), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11])
         );
  DFC1 pipe_rt_reg_10_ ( .D(compare_i_data_rt[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[10]) );
  DFC1 pipe_rt_reg_9_ ( .D(n3181), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[9]) );
  DFC1 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC1 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC1 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC1 pipe_rt_reg_5_ ( .D(n3188), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[5]) );
  DFC1 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC1 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC1 pipe_rt_reg_2_ ( .D(n3191), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[2]) );
  DFC1 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC1 pipe_rt_reg_0_ ( .D(compare_i_data_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[0]) );
  DFC1 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC1 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC1 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC1 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC1 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC1 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC1 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC1 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC1 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U102 ( .A(u_alu_DP_OP_84J3_125_2615_n5), .B(
        u_alu_DP_OP_84J3_125_2615_n95), .Q(u_alu_pre_sum_4b[3]) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U24 ( .A(u_alu_DP_OP_84J3_125_2615_n4), .B(
        u_alu_DP_OP_84J3_125_2615_n32), .Q(u_alu_pre_sum_4a[4]) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U90 ( .A(u_alu_DP_OP_84J3_125_2615_n4), .B(
        u_alu_DP_OP_84J3_125_2615_n89), .Q(u_alu_pre_sum_4b[4]) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U72 ( .A(u_alu_DP_OP_84J3_125_2615_n2), .B(
        u_alu_DP_OP_84J3_125_2615_n73), .Q(u_alu_pre_sum_4b[6]) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U6 ( .A(u_alu_DP_OP_84J3_125_2615_n2), .B(
        u_alu_DP_OP_84J3_125_2615_n16), .Q(u_alu_pre_sum_4a[6]) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U23 ( .A(n3054), .B(compare_i_data_rs[29]), 
        .Q(u_alu_DP_OP_84J3_125_2615_n22) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U20 ( .A(u_alu_DP_OP_84J3_125_2615_n109), 
        .B(u_alu_DP_OP_84J3_125_2615_n22), .Q(u_alu_DP_OP_84J3_125_2615_n3) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U54 ( .A(u_alu_DP_OP_84J3_125_2615_n136), 
        .B(n356), .Q(u_alu_DP_OP_84J3_125_2615_n40) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U44 ( .A(u_alu_DP_OP_84J3_125_2615_n137), 
        .B(u_alu_DP_OP_84J3_125_2615_n145), .Q(u_alu_DP_OP_84J3_125_2615_n37)
         );
  NAND22 u_alu_DP_OP_84J3_125_2615_U41 ( .A(u_alu_DP_OP_84J3_125_2615_n111), 
        .B(u_alu_DP_OP_84J3_125_2615_n37), .Q(u_alu_DP_OP_84J3_125_2615_n5) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U32 ( .A(u_alu_DP_OP_84J3_125_2615_n81), 
        .B(u_alu_DP_OP_84J3_125_2615_n31), .Q(u_alu_DP_OP_84J3_125_2615_n4) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U16 ( .A(u_alu_DP_OP_84J3_125_2615_n81), 
        .B(u_alu_DP_OP_84J3_125_2615_n109), .Q(u_alu_DP_OP_84J3_125_2615_n17)
         );
  AOI211 u_alu_DP_OP_84J3_125_2615_U17 ( .A(u_alu_DP_OP_84J3_125_2615_n109), 
        .B(u_alu_DP_OP_84J3_125_2615_n86), .C(u_alu_DP_OP_84J3_125_2615_n77), 
        .Q(u_alu_DP_OP_84J3_125_2615_n18) );
  OAI212 u_alu_DP_OP_84J3_125_2615_U15 ( .A(u_alu_DP_OP_84J3_125_2615_n17), 
        .B(u_alu_DP_OP_84J3_125_2615_n33), .C(u_alu_DP_OP_84J3_125_2615_n18), 
        .Q(u_alu_DP_OP_84J3_125_2615_n16) );
  NOR21 u_alu_DP_OP_84J3_125_2615_U12 ( .A(compare_i_data_rs[30]), .B(n384), 
        .Q(u_alu_DP_OP_84J3_125_2615_n14) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U13 ( .A(n384), .B(compare_i_data_rs[30]), 
        .Q(u_alu_DP_OP_84J3_125_2615_n15) );
  XOR21 u_alu_DP_OP_84J3_125_2615_U1 ( .A(u_alu_DP_OP_84J3_125_2615_n1), .B(
        u_alu_DP_OP_84J3_125_2615_n11), .Q(u_alu_pre_sum_4a[7]) );
  AOI211 u_alu_DP_OP_84J3_125_2615_U73 ( .A(u_alu_DP_OP_84J3_125_2615_n73), 
        .B(u_alu_DP_OP_84J3_125_2615_n108), .C(u_alu_DP_OP_84J3_125_2615_n70), 
        .Q(u_alu_DP_OP_84J3_125_2615_n68) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U10 ( .A(u_alu_DP_OP_84J3_125_2615_n108), 
        .B(u_alu_DP_OP_84J3_125_2615_n15), .Q(u_alu_DP_OP_84J3_125_2615_n2) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U51 ( .A(n427), .B(
        u_alu_DP_OP_84J3_125_2615_n40), .Q(u_alu_DP_OP_84J3_125_2615_n6) );
  XOR21 u_alu_DP_OP_84J3_125_2615_U45 ( .A(u_alu_DP_OP_84J3_125_2615_n6), .B(
        u_alu_DP_OP_84J3_125_2615_n45), .Q(u_alu_pre_sum_4a[2]) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U58 ( .A(n756), .B(
        u_alu_DP_OP_84J3_125_2615_n48), .Q(u_alu_DP_OP_84J3_125_2615_n7) );
  XOR21 u_alu_DP_OP_84J3_125_2615_U121 ( .A(u_alu_DP_OP_84J3_125_2615_n49), 
        .B(u_alu_DP_OP_84J3_125_2615_n7), .Q(u_alu_pre_sum_4b[1]) );
  NAND20 u_alu_lt_x_11_U45 ( .A(u_alu_lt_x_11_B_22_), .B(n451), .Q(
        u_alu_lt_x_11_n44) );
  NOR20 u_alu_lt_x_11_U132 ( .A(n1775), .B(n628), .Q(u_alu_lt_x_11_n131) );
  OAI212 u_alu_lt_x_11_U1 ( .A(u_alu_lt_x_11_n1), .B(u_alu_lt_x_11_n55), .C(
        u_alu_lt_x_11_n2), .Q(u_alu_N306) );
  AOI211 u_alu_lt_x_11_U13 ( .A(u_alu_lt_x_11_n20), .B(u_alu_lt_x_11_n13), .C(
        u_alu_lt_x_11_n14), .Q(u_alu_lt_x_11_n12) );
  AOI211 u_alu_lt_x_11_U23 ( .A(n566), .B(u_alu_lt_x_11_n28), .C(
        u_alu_lt_x_11_n24), .Q(u_alu_lt_x_11_n22) );
  AOI211 u_alu_lt_x_11_U47 ( .A(u_alu_lt_x_11_n47), .B(u_alu_lt_x_11_n52), .C(
        u_alu_lt_x_11_n48), .Q(u_alu_lt_x_11_n46) );
  AOI211 u_alu_lt_x_11_U60 ( .A(u_alu_lt_x_11_n67), .B(u_alu_lt_x_11_n60), .C(
        u_alu_lt_x_11_n61), .Q(u_alu_lt_x_11_n59) );
  AOI211 u_alu_lt_x_11_U70 ( .A(u_alu_lt_x_11_n70), .B(u_alu_lt_x_11_n75), .C(
        u_alu_lt_x_11_n71), .Q(u_alu_lt_x_11_n69) );
  AOI211 u_alu_lt_x_11_U82 ( .A(u_alu_lt_x_11_n82), .B(u_alu_lt_x_11_n97), .C(
        u_alu_lt_x_11_n83), .Q(u_alu_lt_x_11_n81) );
  AOI211 u_alu_lt_x_11_U100 ( .A(u_alu_lt_x_11_n100), .B(u_alu_lt_x_11_n105), 
        .C(u_alu_lt_x_11_n101), .Q(u_alu_lt_x_11_n99) );
  NAND22 u_alu_lt_x_11_U69 ( .A(u_alu_lt_x_11_n74), .B(u_alu_lt_x_11_n70), .Q(
        u_alu_lt_x_11_n68) );
  NAND22 u_alu_lt_x_11_U81 ( .A(u_alu_lt_x_11_n82), .B(u_alu_lt_x_11_n96), .Q(
        u_alu_lt_x_11_n80) );
  NOR21 u_alu_lt_x_11_U97 ( .A(u_alu_lt_x_11_n108), .B(u_alu_lt_x_11_n98), .Q(
        u_alu_lt_x_11_n96) );
  NOR21 u_alu_lt_x_11_U83 ( .A(u_alu_lt_x_11_n84), .B(u_alu_lt_x_11_n86), .Q(
        u_alu_lt_x_11_n82) );
  NAND22 u_alu_lt_x_11_U87 ( .A(n1003), .B(u_alu_lt_x_11_n92), .Q(
        u_alu_lt_x_11_n86) );
  OAI212 u_alu_lt_x_11_U111 ( .A(u_alu_lt_x_11_n111), .B(u_alu_lt_x_11_n133), 
        .C(u_alu_lt_x_11_n112), .Q(u_alu_lt_x_11_n110) );
  AOI211 u_alu_lt_x_11_U134 ( .A(u_alu_lt_x_11_n140), .B(u_alu_lt_x_11_n134), 
        .C(u_alu_lt_x_11_n135), .Q(u_alu_lt_x_11_n133) );
  NOR21 u_alu_lt_x_11_U135 ( .A(u_alu_lt_x_11_n138), .B(u_alu_lt_x_11_n136), 
        .Q(u_alu_lt_x_11_n134) );
  NAND22 u_alu_lt_x_11_U112 ( .A(u_alu_lt_x_11_n113), .B(u_alu_lt_x_11_n127), 
        .Q(u_alu_lt_x_11_n111) );
  NAND22 u_alu_lt_x_11_U118 ( .A(u_alu_lt_x_11_n123), .B(u_alu_lt_x_11_n119), 
        .Q(u_alu_lt_x_11_n117) );
  NAND22 u_alu_lt_x_11_U2 ( .A(u_alu_lt_x_11_n9), .B(u_alu_lt_x_11_n3), .Q(
        u_alu_lt_x_11_n1) );
  NOR21 u_alu_lt_x_11_U10 ( .A(u_alu_lt_x_11_n33), .B(u_alu_lt_x_11_n11), .Q(
        u_alu_lt_x_11_n9) );
  NAND22 u_alu_lt_x_11_U12 ( .A(u_alu_lt_x_11_n19), .B(u_alu_lt_x_11_n13), .Q(
        u_alu_lt_x_11_n11) );
  NOR21 u_alu_lt_x_11_U14 ( .A(u_alu_lt_x_11_n17), .B(u_alu_lt_x_11_n15), .Q(
        u_alu_lt_x_11_n13) );
  NOR21 u_alu_lt_x_11_U20 ( .A(u_alu_lt_x_11_n31), .B(u_alu_lt_x_11_n21), .Q(
        u_alu_lt_x_11_n19) );
  NAND22 u_alu_lt_x_11_U22 ( .A(u_alu_lt_x_11_n27), .B(n566), .Q(
        u_alu_lt_x_11_n21) );
  NAND22 u_alu_lt_x_11_U34 ( .A(u_alu_lt_x_11_n35), .B(u_alu_lt_x_11_n41), .Q(
        u_alu_lt_x_11_n33) );
  NOR21 u_alu_lt_x_11_U42 ( .A(u_alu_lt_x_11_n43), .B(u_alu_lt_x_11_n45), .Q(
        u_alu_lt_x_11_n41) );
  NOR21 u_alu_lt_x_11_U44 ( .A(n451), .B(u_alu_lt_x_11_B_22_), .Q(
        u_alu_lt_x_11_n43) );
  NOR21 u_alu_lt_x_11_U36 ( .A(u_alu_lt_x_11_n39), .B(u_alu_lt_x_11_n37), .Q(
        u_alu_lt_x_11_n35) );
  NAND20 u_alu_lt_x_11_U17 ( .A(n3054), .B(n444), .Q(u_alu_lt_x_11_n16) );
  NAND20 u_alu_lt_x_11_U19 ( .A(n680), .B(u_alu_lt_x_11_n172), .Q(
        u_alu_lt_x_11_n18) );
  NAND20 u_alu_lt_x_11_U27 ( .A(u_alu_DP_OP_84J3_125_2615_n137), .B(
        u_alu_lt_x_11_n171), .Q(u_alu_lt_x_11_n26) );
  NAND20 u_alu_lt_x_11_U39 ( .A(u_alu_DP_OP_84J3_125_2615_n134), .B(n433), .Q(
        u_alu_lt_x_11_n38) );
  NAND20 u_alu_lt_x_11_U55 ( .A(u_alu_lt_x_11_B_20_), .B(n452), .Q(
        u_alu_lt_x_11_n54) );
  NAND20 u_alu_lt_x_11_U64 ( .A(u_alu_lt_x_11_B_19_), .B(n443), .Q(
        u_alu_lt_x_11_n63) );
  NAND20 u_alu_lt_x_11_U66 ( .A(n2636), .B(u_alu_lt_x_11_B_18_), .Q(
        u_alu_lt_x_11_n65) );
  NAND20 u_alu_lt_x_11_U78 ( .A(n432), .B(u_alu_lt_x_11_B_16_), .Q(
        u_alu_lt_x_11_n77) );
  NAND20 u_alu_lt_x_11_U86 ( .A(u_alu_lt_x_11_B_14_), .B(n403), .Q(
        u_alu_lt_x_11_n85) );
  NAND20 u_alu_lt_x_11_U92 ( .A(u_alu_lt_x_11_B_13_), .B(n417), .Q(
        u_alu_lt_x_11_n91) );
  NAND20 u_alu_lt_x_11_U104 ( .A(n471), .B(n406), .Q(u_alu_lt_x_11_n103) );
  NAND20 u_alu_lt_x_11_U108 ( .A(n440), .B(n2027), .Q(u_alu_lt_x_11_n107) );
  NOR20 u_alu_lt_x_11_U77 ( .A(u_alu_lt_x_11_B_16_), .B(n432), .Q(
        u_alu_lt_x_11_n76) );
  NAND20 u_alu_lt_x_11_U123 ( .A(alu_i_data_B[7]), .B(n357), .Q(
        u_alu_lt_x_11_n122) );
  NAND20 u_alu_lt_x_11_U144 ( .A(u_alu_lt_x_11_B_0_), .B(n419), .Q(
        u_alu_lt_x_11_n143) );
  NOR21 u_alu_lt_x_11_U137 ( .A(n418), .B(n369), .Q(u_alu_lt_x_11_n136) );
  OAI211 u_alu_lt_x_11_U136 ( .A(u_alu_lt_x_11_n139), .B(u_alu_lt_x_11_n136), 
        .C(u_alu_lt_x_11_n137), .Q(u_alu_lt_x_11_n135) );
  OAI211 u_alu_lt_x_11_U37 ( .A(u_alu_lt_x_11_n40), .B(u_alu_lt_x_11_n37), .C(
        u_alu_lt_x_11_n38), .Q(u_alu_lt_x_11_n36) );
  OAI211 u_alu_lt_x_11_U5 ( .A(u_alu_lt_x_11_n8), .B(u_alu_lt_x_11_n5), .C(
        u_alu_lt_x_11_n6), .Q(u_alu_lt_x_11_n4) );
  OAI211 u_alu_lt_x_11_U68 ( .A(u_alu_lt_x_11_n79), .B(u_alu_lt_x_11_n68), .C(
        u_alu_lt_x_11_n69), .Q(u_alu_lt_x_11_n67) );
  NOR21 u_alu_lt_x_11_U61 ( .A(u_alu_lt_x_11_n64), .B(u_alu_lt_x_11_n62), .Q(
        u_alu_lt_x_11_n60) );
  NAND22 u_alu_lt_x_11_U59 ( .A(u_alu_lt_x_11_n60), .B(u_alu_lt_x_11_n66), .Q(
        u_alu_lt_x_11_n58) );
  AOI211 u_alu_DP_OP_84J3_125_2615_U25 ( .A(u_alu_DP_OP_84J3_125_2615_n32), 
        .B(u_alu_DP_OP_84J3_125_2615_n81), .C(u_alu_DP_OP_84J3_125_2615_n86), 
        .Q(u_alu_DP_OP_84J3_125_2615_n23) );
  NOR21 u_alu_lt_x_11_U8 ( .A(n447), .B(n384), .Q(u_alu_lt_x_11_n7) );
  OAI210 u_alu_lt_x_11_U141 ( .A(n2413), .B(u_alu_lt_x_11_n143), .C(
        u_alu_lt_x_11_n142), .Q(u_alu_lt_x_11_n140) );
  NOR21 u_alu_lt_x_11_U63 ( .A(n443), .B(u_alu_lt_x_11_B_19_), .Q(
        u_alu_lt_x_11_n62) );
  NOR21 u_alu_lt_x_11_U38 ( .A(n433), .B(u_alu_DP_OP_84J3_125_2615_n134), .Q(
        u_alu_lt_x_11_n37) );
  NOR21 u_alu_lt_x_11_U67 ( .A(u_alu_lt_x_11_n68), .B(u_alu_lt_x_11_n78), .Q(
        u_alu_lt_x_11_n66) );
  NOR21 u_alu_lt_x_11_U128 ( .A(u_alu_lt_x_11_n131), .B(u_alu_lt_x_11_n129), 
        .Q(u_alu_lt_x_11_n127) );
  OAI211 u_alu_lt_x_11_U15 ( .A(u_alu_lt_x_11_n18), .B(u_alu_lt_x_11_n15), .C(
        u_alu_lt_x_11_n16), .Q(u_alu_lt_x_11_n14) );
  NOR20 u_alu_lt_x_11_U30 ( .A(n355), .B(u_alu_DP_OP_84J3_125_2615_n136), .Q(
        u_alu_lt_x_11_n29) );
  NAND20 u_alu_lt_x_11_U31 ( .A(u_alu_DP_OP_84J3_125_2615_n136), .B(n355), .Q(
        u_alu_lt_x_11_n30) );
  NOR21 u_alu_DP_OP_84J3_125_2615_U34 ( .A(compare_i_data_rs[28]), .B(n680), 
        .Q(u_alu_DP_OP_84J3_125_2615_n30) );
  NOR21 u_alu_lt_x_11_U4 ( .A(u_alu_lt_x_11_n7), .B(u_alu_lt_x_11_n5), .Q(
        u_alu_lt_x_11_n3) );
  NOR20 u_alu_lt_x_11_U65 ( .A(u_alu_lt_x_11_B_18_), .B(n2636), .Q(
        u_alu_lt_x_11_n64) );
  AOI211 u_alu_DP_OP_84J3_125_2615_U91 ( .A(u_alu_DP_OP_84J3_125_2615_n89), 
        .B(u_alu_DP_OP_84J3_125_2615_n81), .C(u_alu_DP_OP_84J3_125_2615_n86), 
        .Q(u_alu_DP_OP_84J3_125_2615_n80) );
  NOR20 u_alu_lt_x_11_U18 ( .A(u_alu_lt_x_11_n172), .B(n680), .Q(
        u_alu_lt_x_11_n17) );
  OAI211 u_alu_lt_x_11_U43 ( .A(u_alu_lt_x_11_n43), .B(u_alu_lt_x_11_n46), .C(
        u_alu_lt_x_11_n44), .Q(u_alu_lt_x_11_n42) );
  OAI211 u_alu_lt_x_11_U62 ( .A(u_alu_lt_x_11_n65), .B(u_alu_lt_x_11_n62), .C(
        u_alu_lt_x_11_n63), .Q(u_alu_lt_x_11_n61) );
  OAI212 u_alu_lt_x_11_U98 ( .A(u_alu_lt_x_11_n109), .B(u_alu_lt_x_11_n98), 
        .C(u_alu_lt_x_11_n99), .Q(u_alu_lt_x_11_n97) );
  OAI212 u_alu_lt_x_11_U58 ( .A(u_alu_lt_x_11_n58), .B(u_alu_lt_x_11_n81), .C(
        u_alu_lt_x_11_n59), .Q(u_alu_lt_x_11_n57) );
  AOI211 u_alu_lt_x_11_U3 ( .A(u_alu_lt_x_11_n10), .B(u_alu_lt_x_11_n3), .C(
        u_alu_lt_x_11_n4), .Q(u_alu_lt_x_11_n2) );
  OAI211 u_alu_lt_x_11_U21 ( .A(n3010), .B(u_alu_lt_x_11_n21), .C(
        u_alu_lt_x_11_n22), .Q(u_alu_lt_x_11_n20) );
  DFC1 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC3 pipe_con_Malupc8_reg ( .D(i_con_Malupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Malupc8) );
  NAND24 U3 ( .A(n9), .B(i_data_FMalures[25]), .Q(n1435) );
  NOR23 U4 ( .A(n2848), .B(n2847), .Q(n2885) );
  INV15 U5 ( .A(n1166), .Q(n401) );
  AOI222 U6 ( .A(n3067), .B(u_alu_lt_x_11_B_15_), .C(n2308), .D(n410), .Q(
        n2600) );
  AOI212 U7 ( .A(n2099), .B(n458), .C(n78), .Q(n2056) );
  NAND26 U8 ( .A(n435), .B(compare_i_data_rs[28]), .Q(n3081) );
  NAND26 U9 ( .A(n1045), .B(n1930), .Q(n1946) );
  AOI211 U10 ( .A(n860), .B(n410), .C(n2264), .Q(n2520) );
  INV3 U11 ( .A(n311), .Q(n310) );
  NAND24 U12 ( .A(n382), .B(i_data_rt[13]), .Q(n2165) );
  NOR23 U13 ( .A(n252), .B(n2010), .Q(n2434) );
  NOR22 U14 ( .A(n2010), .B(n2423), .Q(n2011) );
  NAND26 U15 ( .A(n438), .B(n1039), .Q(n2010) );
  NOR22 U16 ( .A(n1171), .B(n1946), .Q(n3144) );
  NAND33 U17 ( .A(n3114), .B(n3113), .C(n1155), .Q(n3125) );
  AOI212 U18 ( .A(n3039), .B(n378), .C(n3038), .Q(n3040) );
  INV12 U19 ( .A(n1150), .Q(n343) );
  NAND31 U20 ( .A(n1171), .B(n386), .C(u_alu_lt_x_11_B_19_), .Q(n55) );
  NAND23 U21 ( .A(n390), .B(i_data_rt[18]), .Q(n1128) );
  NAND24 U22 ( .A(n2822), .B(n1), .Q(n2825) );
  CLKIN6 U23 ( .A(n2821), .Q(n1) );
  NAND24 U24 ( .A(n2819), .B(n2818), .Q(n2821) );
  NOR24 U25 ( .A(n2723), .B(n2724), .Q(n2818) );
  NAND24 U26 ( .A(n4), .B(n2), .Q(n2822) );
  OAI212 U27 ( .A(n2623), .B(n2622), .C(n3), .Q(n2) );
  CLKIN3 U28 ( .A(n2657), .Q(n3) );
  NOR24 U29 ( .A(n2514), .B(n2513), .Q(n2622) );
  CLKIN6 U30 ( .A(n2658), .Q(n2623) );
  CLKIN6 U31 ( .A(n2660), .Q(n4) );
  NAND24 U32 ( .A(n978), .B(n2624), .Q(n2660) );
  NOR24 U33 ( .A(n1167), .B(n2309), .Q(n2310) );
  NAND24 U34 ( .A(n2598), .B(n186), .Q(n2309) );
  CLKIN6 U35 ( .A(n5), .Q(n2598) );
  NAND24 U36 ( .A(n471), .B(n132), .Q(n5) );
  INV12 U37 ( .A(n6), .Q(n7) );
  NAND34 U38 ( .A(n1548), .B(n1546), .C(n259), .Q(n1681) );
  NAND23 U39 ( .A(n928), .B(n2966), .Q(n1027) );
  NAND26 U40 ( .A(n2669), .B(n2668), .Q(u_alu_lt_x_11_B_21_) );
  NAND24 U41 ( .A(n1489), .B(n139), .Q(n2669) );
  INV6 U42 ( .A(n967), .Q(n6) );
  NOR22 U43 ( .A(n628), .B(n1775), .Q(n627) );
  NAND24 U44 ( .A(n728), .B(n726), .Q(n1942) );
  NAND23 U45 ( .A(n2204), .B(n400), .Q(n885) );
  NOR22 U46 ( .A(n1565), .B(n1564), .Q(n1570) );
  INV6 U47 ( .A(i_data_immext[0]), .Q(n1565) );
  NAND26 U48 ( .A(i_data_immext[3]), .B(i_data_immext[5]), .Q(n1564) );
  INV12 U49 ( .A(n3161), .Q(n1153) );
  NOR23 U50 ( .A(n332), .B(n1631), .Q(n3161) );
  NAND26 U51 ( .A(n1060), .B(n330), .Q(n1152) );
  NAND26 U52 ( .A(n172), .B(n171), .Q(n2393) );
  NAND24 U53 ( .A(n1364), .B(n759), .Q(compare_i_data_rt[3]) );
  NAND33 U54 ( .A(n1739), .B(n1738), .C(n1737), .Q(n2595) );
  NAND26 U55 ( .A(u_alu_lt_x_11_n40), .B(n2836), .Q(n2843) );
  NOR22 U56 ( .A(n765), .B(n1448), .Q(n762) );
  NAND23 U57 ( .A(n1136), .B(i_data_FMmemout[15]), .Q(n1216) );
  NAND26 U58 ( .A(n501), .B(n499), .Q(n894) );
  INV15 U59 ( .A(n312), .Q(n2636) );
  NAND28 U60 ( .A(n585), .B(n584), .Q(n594) );
  CLKIN4 U61 ( .A(n604), .Q(n584) );
  AOI212 U62 ( .A(n2855), .B(n2854), .C(n823), .Q(n2662) );
  NOR23 U63 ( .A(n364), .B(n241), .Q(n240) );
  NOR23 U64 ( .A(n241), .B(n786), .Q(n785) );
  NAND23 U65 ( .A(n2243), .B(n2242), .Q(n3193) );
  AOI212 U66 ( .A(n3024), .B(n3025), .C(n386), .Q(n3108) );
  NAND20 U67 ( .A(n3032), .B(n400), .Q(n2978) );
  NAND26 U68 ( .A(u_alu_lt_x_11_B_16_), .B(n1171), .Q(n267) );
  NAND26 U69 ( .A(n825), .B(n2394), .Q(u_alu_lt_x_11_B_16_) );
  NOR23 U70 ( .A(n401), .B(n2057), .Q(n505) );
  CLKIN4 U71 ( .A(n873), .Q(n3033) );
  NAND26 U72 ( .A(n876), .B(n1953), .Q(n3192) );
  INV8 U73 ( .A(n3192), .Q(n875) );
  NAND24 U74 ( .A(n1137), .B(i_data_FMmemout[11]), .Q(n595) );
  NAND23 U75 ( .A(n1137), .B(i_data_FMmemout[24]), .Q(n1055) );
  BUF15 U76 ( .A(n1437), .Q(n8) );
  NOR24 U77 ( .A(n699), .B(n565), .Q(n698) );
  NOR24 U78 ( .A(n1389), .B(n352), .Q(n1437) );
  AOI212 U79 ( .A(n9), .B(i_data_FMalures[9]), .C(n238), .Q(n48) );
  NOR23 U80 ( .A(n1356), .B(n351), .Q(n238) );
  NAND24 U81 ( .A(n1038), .B(n117), .Q(n3191) );
  NOR23 U82 ( .A(n203), .B(n649), .Q(n648) );
  XOR22 U83 ( .A(u_alu_DP_OP_84J3_125_2615_n3), .B(
        u_alu_DP_OP_84J3_125_2615_n23), .Q(u_alu_pre_sum_4a[5]) );
  NAND26 U84 ( .A(u_alu_lt_x_11_B_18_), .B(n1171), .Q(n2714) );
  NOR23 U85 ( .A(n458), .B(n3029), .Q(n3030) );
  NAND24 U86 ( .A(n338), .B(i_data_FWmemout[1]), .Q(n1679) );
  NAND24 U87 ( .A(n338), .B(i_data_FWmemout[13]), .Q(n2191) );
  INV15 U88 ( .A(n350), .Q(n352) );
  INV12 U89 ( .A(n381), .Q(n383) );
  NAND26 U90 ( .A(n1609), .B(n377), .Q(n3009) );
  NOR32 U91 ( .A(n1496), .B(n1124), .C(n1497), .Q(n548) );
  INV12 U92 ( .A(n471), .Q(n2374) );
  NOR23 U93 ( .A(n203), .B(n2585), .Q(n2586) );
  CLKBU15 U94 ( .A(n594), .Q(n347) );
  NAND34 U95 ( .A(n208), .B(n207), .C(n206), .Q(n205) );
  NOR33 U96 ( .A(n2635), .B(n2636), .C(u_alu_lt_x_11_B_18_), .Q(n878) );
  AOI212 U97 ( .A(n3047), .B(n1053), .C(n3046), .Q(n3048) );
  NOR22 U98 ( .A(n2654), .B(n2333), .Q(n2282) );
  NOR22 U99 ( .A(n1504), .B(n347), .Q(n1291) );
  NOR23 U100 ( .A(n1438), .B(n8), .Q(n702) );
  NOR33 U101 ( .A(n2013), .B(n1140), .C(n2012), .Q(n2124) );
  AOI212 U102 ( .A(n2321), .B(n2208), .C(n2207), .Q(n2225) );
  CLKIN4 U103 ( .A(n1345), .Q(n1348) );
  NOR24 U104 ( .A(n458), .B(n1906), .Q(n1831) );
  NOR23 U105 ( .A(n420), .B(n2139), .Q(n2487) );
  NAND26 U106 ( .A(n446), .B(u_alu_lt_x_11_A_12_), .Q(n2198) );
  NAND23 U107 ( .A(n842), .B(n841), .Q(n840) );
  NAND23 U108 ( .A(n3126), .B(n2958), .Q(n1057) );
  NAND43 U109 ( .A(n1240), .B(n1241), .C(n1243), .D(n249), .Q(n250) );
  INV6 U110 ( .A(n94), .Q(n249) );
  INV12 U111 ( .A(n1111), .Q(n9) );
  INV12 U112 ( .A(n1111), .Q(n456) );
  NOR24 U113 ( .A(n394), .B(n3109), .Q(n3110) );
  INV12 U114 ( .A(n2202), .Q(n2300) );
  NOR22 U115 ( .A(u_alu_lt_x_11_B_8_), .B(n1039), .Q(n1095) );
  NAND23 U116 ( .A(u_alu_lt_x_11_B_8_), .B(n1171), .Q(n187) );
  INV12 U117 ( .A(u_alu_lt_x_11_B_8_), .Q(n438) );
  AOI212 U118 ( .A(n2673), .B(n410), .C(n2672), .Q(n2674) );
  NAND24 U119 ( .A(n454), .B(i_data_FEalures[21]), .Q(n1110) );
  NAND26 U120 ( .A(n3197), .B(n139), .Q(n2286) );
  NAND26 U121 ( .A(n2971), .B(n2441), .Q(n1149) );
  NAND26 U122 ( .A(n155), .B(n154), .Q(n3187) );
  AOI212 U123 ( .A(n1836), .B(n2907), .C(n1835), .Q(n1837) );
  NAND24 U124 ( .A(n365), .B(n401), .Q(n1526) );
  INV3 U125 ( .A(n2555), .Q(n2556) );
  INV3 U126 ( .A(n1205), .Q(n215) );
  NOR21 U127 ( .A(n1171), .B(n2593), .Q(n2594) );
  NOR21 U128 ( .A(n1170), .B(n1168), .Q(n837) );
  NAND23 U129 ( .A(n2442), .B(n1473), .Q(n288) );
  NAND22 U130 ( .A(n1296), .B(n461), .Q(n1297) );
  NOR21 U131 ( .A(n1295), .B(n351), .Q(n1298) );
  NAND22 U132 ( .A(n1617), .B(n1616), .Q(n1864) );
  NAND22 U133 ( .A(n142), .B(i_data_FMmemout[14]), .Q(n211) );
  NAND22 U134 ( .A(n398), .B(i_data_rs[27]), .Q(n262) );
  NAND22 U135 ( .A(n143), .B(i_data_FMmemout[27]), .Q(n1427) );
  NOR21 U136 ( .A(n386), .B(n1617), .Q(n2930) );
  INV3 U137 ( .A(n2933), .Q(n175) );
  INV3 U138 ( .A(i_data_immext[4]), .Q(n719) );
  INV6 U139 ( .A(n725), .Q(n473) );
  INV3 U140 ( .A(n360), .Q(n134) );
  INV3 U141 ( .A(n287), .Q(n286) );
  NOR32 U142 ( .A(n288), .B(n496), .C(compare_i_data_rt[16]), .Q(n287) );
  NAND22 U143 ( .A(compare_i_data_rt[16]), .B(n288), .Q(n285) );
  NAND22 U144 ( .A(compare_i_data_rt[16]), .B(n496), .Q(n284) );
  NOR22 U145 ( .A(n1875), .B(n886), .Q(n2416) );
  NAND26 U146 ( .A(n1121), .B(n406), .Q(n2108) );
  NAND22 U147 ( .A(n2164), .B(n365), .Q(n2429) );
  NAND33 U148 ( .A(n2168), .B(n2188), .C(n391), .Q(n2248) );
  NAND22 U149 ( .A(n2963), .B(n1171), .Q(n2981) );
  NAND22 U150 ( .A(n2304), .B(n2376), .Q(n530) );
  INV3 U151 ( .A(n2349), .Q(n2359) );
  NAND22 U152 ( .A(n2474), .B(n2462), .Q(n2463) );
  BUF6 U153 ( .A(n2835), .Q(u_alu_lt_x_11_B_22_) );
  NAND22 U154 ( .A(u_alu_lt_x_11_B_18_), .B(n2636), .Q(n2830) );
  NAND26 U155 ( .A(n1440), .B(n563), .Q(compare_i_data_rs[25]) );
  NAND22 U156 ( .A(u_alu_lt_x_11_B_17_), .B(n2897), .Q(n1043) );
  NAND22 U157 ( .A(n2981), .B(n707), .Q(n3147) );
  NAND22 U158 ( .A(n471), .B(n420), .Q(n707) );
  INV3 U159 ( .A(n2421), .Q(n881) );
  NAND22 U160 ( .A(n958), .B(n957), .Q(n882) );
  NOR32 U161 ( .A(n638), .B(n1416), .C(n607), .Q(n606) );
  NAND22 U162 ( .A(n1418), .B(n608), .Q(n607) );
  NOR21 U163 ( .A(n1286), .B(n1158), .Q(n1239) );
  NOR21 U164 ( .A(n1167), .B(n1712), .Q(n311) );
  INV3 U165 ( .A(n798), .Q(n218) );
  NOR23 U166 ( .A(n2382), .B(n2381), .Q(n2383) );
  INV3 U167 ( .A(n630), .Q(n2392) );
  NOR22 U168 ( .A(n407), .B(n438), .Q(n2031) );
  NAND22 U169 ( .A(n2156), .B(n2350), .Q(n225) );
  INV6 U170 ( .A(n618), .Q(n2362) );
  AOI221 U171 ( .A(n2489), .B(n401), .C(n2590), .D(n397), .Q(n2527) );
  NAND22 U172 ( .A(n2552), .B(n2559), .Q(n2557) );
  NOR21 U173 ( .A(n2636), .B(u_alu_lt_x_11_B_18_), .Q(n2580) );
  NAND26 U174 ( .A(n199), .B(n198), .Q(n1632) );
  INV3 U175 ( .A(n1601), .Q(n198) );
  INV6 U176 ( .A(n1602), .Q(n199) );
  INV3 U177 ( .A(n2520), .Q(n2524) );
  NAND22 U178 ( .A(n3097), .B(n2611), .Q(n2522) );
  NAND23 U179 ( .A(n1493), .B(n139), .Q(n2618) );
  INV3 U180 ( .A(n2838), .Q(n2764) );
  NAND22 U181 ( .A(n2770), .B(n2818), .Q(n2782) );
  NAND24 U182 ( .A(n2451), .B(n2450), .Q(n3167) );
  NAND23 U183 ( .A(n405), .B(n414), .Q(n756) );
  INV12 U184 ( .A(n1388), .Q(n350) );
  NAND26 U185 ( .A(n1457), .B(n1456), .Q(compare_i_data_rs[21]) );
  INV3 U186 ( .A(u_alu_lt_x_11_A_5_), .Q(n437) );
  NAND24 U187 ( .A(n907), .B(n874), .Q(n897) );
  INV12 U188 ( .A(u_alu_lt_x_11_A_3_), .Q(n418) );
  NAND22 U189 ( .A(n1137), .B(i_data_FMmemout[4]), .Q(n1201) );
  NAND23 U190 ( .A(n338), .B(i_data_FWmemout[19]), .Q(n206) );
  INV3 U191 ( .A(n2390), .Q(n1958) );
  INV3 U192 ( .A(n1155), .Q(n303) );
  NAND23 U193 ( .A(n336), .B(u_alu_lt_x_11_B_14_), .Q(n2358) );
  NAND24 U194 ( .A(n170), .B(n168), .Q(n167) );
  INV3 U195 ( .A(n2456), .Q(n2315) );
  NAND22 U196 ( .A(n2296), .B(n458), .Q(n275) );
  NOR22 U197 ( .A(n1164), .B(n379), .Q(n849) );
  NAND23 U198 ( .A(u_alu_DP_OP_83J3_124_3384_n154), .B(u_alu_lt_x_11_B_16_), 
        .Q(n2514) );
  XNR21 U199 ( .A(n2757), .B(n214), .Q(n2758) );
  NOR21 U200 ( .A(n2812), .B(n2815), .Q(n2783) );
  INV12 U201 ( .A(n1044), .Q(n421) );
  NAND24 U202 ( .A(n3158), .B(n400), .Q(n3074) );
  NOR22 U203 ( .A(n3131), .B(n3135), .Q(n3141) );
  INV3 U204 ( .A(n977), .Q(n3138) );
  INV12 U205 ( .A(n402), .Q(n381) );
  NAND33 U206 ( .A(n831), .B(n1468), .C(n2559), .Q(compare_i_data_rs[19]) );
  NAND22 U207 ( .A(n970), .B(n364), .Q(n510) );
  INV12 U208 ( .A(n1160), .Q(n1158) );
  NOR21 U209 ( .A(n1346), .B(n1158), .Q(n1347) );
  INV8 U210 ( .A(i_data_immext[6]), .Q(n1164) );
  NOR22 U211 ( .A(n683), .B(n1443), .Q(n682) );
  NAND22 U212 ( .A(n2189), .B(n2188), .Q(n316) );
  NOR23 U213 ( .A(n1352), .B(n347), .Q(n237) );
  INV3 U214 ( .A(n264), .Q(n323) );
  BUF6 U215 ( .A(n399), .Q(n361) );
  NAND22 U216 ( .A(n2595), .B(n2594), .Q(n2596) );
  INV3 U217 ( .A(n939), .Q(n2521) );
  NAND22 U218 ( .A(n398), .B(i_data_rs[25]), .Q(n1439) );
  INV3 U219 ( .A(n836), .Q(n2975) );
  NAND22 U220 ( .A(n384), .B(n837), .Q(n836) );
  NAND23 U221 ( .A(n680), .B(n1171), .Q(n3027) );
  NAND22 U222 ( .A(n410), .B(n1167), .Q(n184) );
  NAND22 U223 ( .A(alu_i_data_B[31]), .B(n837), .Q(n873) );
  NAND22 U224 ( .A(u_alu_lt_x_11_B_21_), .B(n837), .Q(n271) );
  INV3 U225 ( .A(i_con_Ealuop[5]), .Q(n1555) );
  INV6 U226 ( .A(n1039), .Q(n235) );
  INV3 U227 ( .A(compare_i_data_rt[12]), .Q(n230) );
  NOR20 U228 ( .A(n2027), .B(n440), .Q(u_alu_lt_x_11_n106) );
  NAND23 U229 ( .A(n2027), .B(n1171), .Q(n939) );
  BUF6 U230 ( .A(u_alu_lt_x_11_B_15_), .Q(n193) );
  NAND22 U231 ( .A(n940), .B(n939), .Q(n937) );
  NOR32 U232 ( .A(n1236), .B(n1237), .C(n1235), .Q(n771) );
  NAND22 U233 ( .A(n343), .B(i_data_rs[7]), .Q(n1238) );
  NOR22 U234 ( .A(n1683), .B(n804), .Q(n1922) );
  NAND23 U235 ( .A(u_alu_lt_x_11_B_9_), .B(n436), .Q(u_alu_lt_x_11_n109) );
  NAND26 U236 ( .A(n800), .B(n1475), .Q(n3185) );
  NAND22 U237 ( .A(n2139), .B(n436), .Q(n2370) );
  NAND22 U238 ( .A(n187), .B(n186), .Q(n185) );
  NAND22 U239 ( .A(n141), .B(i_data_FMmemout[13]), .Q(n1250) );
  NOR21 U240 ( .A(n164), .B(n3185), .Q(n2130) );
  INV3 U241 ( .A(n211), .Q(n210) );
  INV3 U242 ( .A(u_alu_lt_x_11_n90), .Q(n1003) );
  AOI211 U243 ( .A(n2500), .B(n410), .C(n1988), .Q(n2175) );
  NOR21 U244 ( .A(n1168), .B(n267), .Q(n1988) );
  NOR22 U245 ( .A(n420), .B(n2763), .Q(n2612) );
  INV3 U246 ( .A(n662), .Q(n2552) );
  INV3 U247 ( .A(n2517), .Q(n2513) );
  INV6 U248 ( .A(n2933), .Q(n2793) );
  NAND22 U249 ( .A(n306), .B(n385), .Q(n2740) );
  NOR23 U250 ( .A(n1340), .B(n347), .Q(n153) );
  NOR32 U251 ( .A(n491), .B(n490), .C(n486), .Q(n489) );
  INV3 U252 ( .A(n1119), .Q(n512) );
  NAND22 U253 ( .A(n2521), .B(n410), .Q(n2716) );
  NAND22 U254 ( .A(n371), .B(n1170), .Q(n2715) );
  NAND22 U255 ( .A(n2930), .B(n1167), .Q(n319) );
  NOR32 U256 ( .A(n2396), .B(n1171), .C(n2395), .Q(n2869) );
  NOR21 U257 ( .A(n2952), .B(n3167), .Q(n966) );
  NOR22 U258 ( .A(n537), .B(n536), .Q(n2937) );
  NOR22 U259 ( .A(n394), .B(n2889), .Q(n2976) );
  NAND24 U260 ( .A(n668), .B(n377), .Q(u_alu_DP_OP_84J3_125_2615_n136) );
  NAND22 U261 ( .A(n213), .B(n363), .Q(n212) );
  INV3 U262 ( .A(n1196), .Q(n213) );
  NOR23 U263 ( .A(n1428), .B(n1122), .Q(n1070) );
  INV3 U264 ( .A(n262), .Q(n1428) );
  NAND22 U265 ( .A(n2930), .B(n394), .Q(n2931) );
  NAND22 U266 ( .A(n174), .B(n180), .Q(n179) );
  NOR21 U267 ( .A(n615), .B(n362), .Q(n180) );
  NAND23 U268 ( .A(n3015), .B(n3014), .Q(n986) );
  NAND31 U269 ( .A(n182), .B(n181), .C(n386), .Q(n3099) );
  NAND22 U270 ( .A(n175), .B(n2952), .Q(n181) );
  INV6 U271 ( .A(n3129), .Q(n3130) );
  INV3 U272 ( .A(n3012), .Q(n3007) );
  NAND22 U273 ( .A(n1409), .B(n472), .Q(n1410) );
  INV3 U274 ( .A(n1413), .Q(n190) );
  NAND22 U275 ( .A(n398), .B(i_data_rs[30]), .Q(n1413) );
  NOR21 U276 ( .A(n1370), .B(n292), .Q(n1412) );
  NOR21 U277 ( .A(i_data_immext[3]), .B(i_data_immext[4]), .Q(n1563) );
  NAND22 U278 ( .A(n360), .B(u_alu_lt_x_11_A_0_), .Q(n136) );
  AOI211 U279 ( .A(n1726), .B(n1741), .C(n1722), .Q(n1723) );
  INV3 U280 ( .A(n1922), .Q(n855) );
  NAND23 U281 ( .A(n1378), .B(n1377), .Q(compare_i_data_rs[31]) );
  NOR32 U282 ( .A(n1376), .B(n1375), .C(n1374), .Q(n1378) );
  NAND23 U283 ( .A(n1692), .B(n1691), .Q(u_alu_lt_x_11_A_2_) );
  AOI211 U284 ( .A(n1690), .B(n1689), .C(n2384), .Q(n1727) );
  INV3 U285 ( .A(n1809), .Q(n1936) );
  NAND26 U286 ( .A(n250), .B(n1112), .Q(n1914) );
  NAND31 U287 ( .A(n1840), .B(n1618), .C(n386), .Q(n936) );
  INV3 U288 ( .A(n611), .Q(n2414) );
  NOR21 U289 ( .A(n1168), .B(n1795), .Q(n1973) );
  NAND23 U290 ( .A(n372), .B(n409), .Q(n611) );
  NOR23 U291 ( .A(n1782), .B(n1781), .Q(n2419) );
  NAND23 U292 ( .A(n2027), .B(n2124), .Q(n2107) );
  INV6 U293 ( .A(n3185), .Q(n406) );
  AOI221 U294 ( .A(n1973), .B(n362), .C(n2180), .D(n1167), .Q(n2053) );
  NOR22 U295 ( .A(n436), .B(u_alu_lt_x_11_B_9_), .Q(n2436) );
  NOR22 U296 ( .A(n1266), .B(n1265), .Q(n232) );
  NOR21 U297 ( .A(n1262), .B(n352), .Q(n1266) );
  NAND23 U298 ( .A(n974), .B(n2429), .Q(n973) );
  INV3 U299 ( .A(n2345), .Q(n2154) );
  NOR21 U300 ( .A(n2209), .B(n1156), .Q(n2218) );
  INV3 U301 ( .A(n403), .Q(n336) );
  INV3 U302 ( .A(n169), .Q(n168) );
  NOR21 U303 ( .A(n969), .B(n1958), .Q(n651) );
  INV3 U304 ( .A(n1012), .Q(n171) );
  INV3 U305 ( .A(n1118), .Q(n428) );
  NAND23 U306 ( .A(n2422), .B(n972), .Q(n1118) );
  NOR22 U307 ( .A(n403), .B(u_alu_lt_x_11_B_14_), .Q(u_alu_lt_x_11_n84) );
  NAND23 U308 ( .A(u_alu_lt_x_11_B_14_), .B(n403), .Q(n2439) );
  NAND22 U309 ( .A(n2307), .B(n528), .Q(n665) );
  NAND22 U310 ( .A(n2463), .B(n139), .Q(n1670) );
  NAND26 U311 ( .A(n1952), .B(n1954), .Q(u_alu_lt_x_11_B_1_) );
  NAND22 U312 ( .A(compare_i_data_rs[17]), .B(n2479), .Q(n2658) );
  NAND23 U313 ( .A(n2518), .B(n2517), .Q(n2659) );
  NOR21 U314 ( .A(n1365), .B(n353), .Q(n1461) );
  INV6 U315 ( .A(n374), .Q(n452) );
  NAND22 U316 ( .A(n441), .B(compare_i_data_rs[21]), .Q(n2845) );
  NAND26 U317 ( .A(n450), .B(u_alu_lt_x_11_B_21_), .Q(u_alu_lt_x_11_n50) );
  NAND22 U318 ( .A(n2778), .B(n362), .Q(n538) );
  BUF6 U319 ( .A(n2926), .Q(n370) );
  INV3 U320 ( .A(u_alu_DP_OP_84J3_125_2615_n50), .Q(n266) );
  INV3 U321 ( .A(n2974), .Q(n586) );
  NOR23 U322 ( .A(n164), .B(n163), .Q(n453) );
  AOI211 U323 ( .A(n3035), .B(n401), .C(n2945), .Q(n2979) );
  NOR22 U324 ( .A(u_alu_DP_OP_84J3_125_2615_n145), .B(
        u_alu_DP_OP_84J3_125_2615_n137), .Q(u_alu_DP_OP_84J3_125_2615_n36) );
  NAND23 U325 ( .A(n2963), .B(n1070), .Q(n3012) );
  NAND22 U326 ( .A(n977), .B(n3042), .Q(n3016) );
  NAND23 U327 ( .A(n928), .B(n3042), .Q(n3047) );
  INV3 U328 ( .A(n3056), .Q(n749) );
  NOR22 U329 ( .A(n650), .B(n749), .Q(n642) );
  NAND22 U330 ( .A(n647), .B(n3175), .Q(n646) );
  NOR22 U331 ( .A(n3129), .B(n3131), .Q(n3091) );
  NAND22 U332 ( .A(n384), .B(n447), .Q(u_alu_lt_x_11_n8) );
  IMUX21 U333 ( .A(n3164), .B(n3163), .S(n145), .Q(n3170) );
  NAND23 U334 ( .A(n882), .B(n881), .Q(n2428) );
  NOR22 U335 ( .A(n1290), .B(n1291), .Q(n2442) );
  INV3 U336 ( .A(n1147), .Q(n1148) );
  INV3 U337 ( .A(n451), .Q(n359) );
  NAND23 U338 ( .A(n398), .B(i_data_rs[19]), .Q(n2559) );
  NAND22 U339 ( .A(n1315), .B(n340), .Q(n339) );
  INV3 U340 ( .A(n770), .Q(n742) );
  NOR23 U341 ( .A(n1310), .B(n663), .Q(n901) );
  INV3 U342 ( .A(n766), .Q(n663) );
  NOR22 U343 ( .A(n1359), .B(n1130), .Q(n828) );
  INV3 U344 ( .A(n1536), .Q(n1938) );
  NAND23 U345 ( .A(n338), .B(i_data_FWmemout[6]), .Q(n1533) );
  NAND22 U346 ( .A(n1134), .B(i_data_FMalures[7]), .Q(n1231) );
  NAND33 U347 ( .A(n581), .B(n1354), .C(n1355), .Q(n583) );
  NAND22 U348 ( .A(n1134), .B(i_data_FMalures[11]), .Q(n543) );
  NOR21 U349 ( .A(n564), .B(n2384), .Q(n1657) );
  INV3 U350 ( .A(u_alu_lt_x_11_B_1_), .Q(n2895) );
  CLKBU12 U351 ( .A(n3184), .Q(n371) );
  NOR22 U352 ( .A(n218), .B(n217), .Q(n216) );
  NAND26 U353 ( .A(n735), .B(n734), .Q(u_alu_lt_x_11_A_5_) );
  NAND22 U354 ( .A(n1815), .B(n1809), .Q(n630) );
  AOI221 U355 ( .A(n1793), .B(n1167), .C(n362), .D(n1990), .Q(n1867) );
  INV6 U356 ( .A(n357), .Q(n358) );
  INV6 U357 ( .A(n887), .Q(n357) );
  INV6 U358 ( .A(i_data_immext[7]), .Q(n1166) );
  AOI211 U359 ( .A(n1857), .B(n2390), .C(n1856), .Q(n1858) );
  NAND24 U360 ( .A(n1478), .B(n1477), .Q(u_alu_lt_x_11_A_10_) );
  INV12 U361 ( .A(n1153), .Q(n422) );
  INV3 U362 ( .A(u_alu_lt_x_11_A_10_), .Q(n440) );
  INV3 U363 ( .A(n1631), .Q(n201) );
  NAND22 U364 ( .A(n973), .B(n417), .Q(n2361) );
  AOI211 U365 ( .A(n2326), .B(n428), .C(n2327), .Q(n2269) );
  NAND22 U366 ( .A(n2328), .B(n423), .Q(n2329) );
  NOR21 U367 ( .A(n2734), .B(n2700), .Q(n2664) );
  INV6 U368 ( .A(n1931), .Q(n372) );
  INV3 U369 ( .A(n2832), .Q(n2859) );
  INV3 U370 ( .A(n2820), .Q(n2729) );
  INV6 U371 ( .A(n3167), .Q(n3121) );
  INV3 U372 ( .A(n928), .Q(n3041) );
  NAND22 U373 ( .A(u_alu_DP_OP_84J3_125_2615_n134), .B(compare_i_data_rs[24]), 
        .Q(u_alu_DP_OP_84J3_125_2615_n50) );
  NAND23 U374 ( .A(n797), .B(n433), .Q(n796) );
  INV3 U375 ( .A(u_alu_DP_OP_84J3_125_2615_n46), .Q(
        u_alu_DP_OP_84J3_125_2615_n45) );
  NAND22 U376 ( .A(n294), .B(n2924), .Q(n2956) );
  NAND22 U377 ( .A(n923), .B(n3008), .Q(n924) );
  NAND31 U378 ( .A(n3016), .B(n1053), .C(n3045), .Q(n1052) );
  NAND24 U379 ( .A(n1635), .B(n1634), .Q(n1638) );
  NAND23 U380 ( .A(n2728), .B(n2727), .Q(n2811) );
  NAND22 U381 ( .A(n1137), .B(i_data_FMmemout[1]), .Q(n259) );
  NOR22 U382 ( .A(n1363), .B(n281), .Q(n1736) );
  INV3 U383 ( .A(n1935), .Q(n732) );
  NOR21 U384 ( .A(n1307), .B(n1158), .Q(n1271) );
  NAND23 U385 ( .A(n1161), .B(i_data_rt[9]), .Q(n2145) );
  NOR22 U386 ( .A(n1230), .B(n482), .Q(n495) );
  NAND23 U387 ( .A(n338), .B(i_data_FWmemout[18]), .Q(n344) );
  NAND23 U388 ( .A(n1161), .B(i_data_rt[19]), .Q(n2553) );
  NAND22 U389 ( .A(n454), .B(i_data_FEalures[19]), .Q(n208) );
  NAND23 U390 ( .A(n338), .B(i_data_FWmemout[21]), .Q(n1488) );
  NAND22 U391 ( .A(n1161), .B(i_data_rt[27]), .Q(n1196) );
  NAND22 U392 ( .A(n1137), .B(i_data_FMmemout[31]), .Q(n1173) );
  INV6 U393 ( .A(n378), .Q(n379) );
  INV12 U394 ( .A(n1164), .Q(n400) );
  INV3 U395 ( .A(n1967), .Q(n304) );
  NOR21 U396 ( .A(n303), .B(n305), .Q(n297) );
  NAND22 U397 ( .A(n1911), .B(n400), .Q(n305) );
  NAND22 U398 ( .A(n1968), .B(n404), .Q(n302) );
  IMUX21 U399 ( .A(n1963), .B(n1962), .S(n1138), .Q(n1968) );
  NOR21 U400 ( .A(n2112), .B(n1156), .Q(n2117) );
  XNR21 U401 ( .A(n2292), .B(n2291), .Q(n2320) );
  NAND22 U402 ( .A(n2698), .B(n571), .Q(n955) );
  INV3 U403 ( .A(n956), .Q(n2515) );
  NAND22 U404 ( .A(n2698), .B(n570), .Q(n956) );
  AOI211 U405 ( .A(n2533), .B(n2907), .C(n2532), .Q(n2536) );
  NAND22 U406 ( .A(n317), .B(n2907), .Q(n2605) );
  INV6 U407 ( .A(n2784), .Q(n2690) );
  NOR22 U408 ( .A(n2758), .B(n952), .Q(n671) );
  INV3 U409 ( .A(n2783), .Q(n149) );
  NAND22 U410 ( .A(n2910), .B(n2909), .Q(n2911) );
  AOI211 U411 ( .A(n378), .B(n2904), .C(n2903), .Q(n2910) );
  NOR22 U412 ( .A(n567), .B(n1076), .Q(n1075) );
  INV3 U413 ( .A(n3141), .Q(n3137) );
  AOI211 U414 ( .A(u_alu_DP_OP_84J3_125_2615_n16), .B(
        u_alu_DP_OP_84J3_125_2615_n108), .C(u_alu_DP_OP_84J3_125_2615_n70), 
        .Q(u_alu_DP_OP_84J3_125_2615_n11) );
  NAND24 U415 ( .A(n2464), .B(n2465), .Q(n191) );
  INV12 U416 ( .A(n269), .Q(n270) );
  NAND26 U417 ( .A(n2451), .B(n1638), .Q(n1627) );
  NOR21 U418 ( .A(n1171), .B(n1168), .Q(n2671) );
  INV3 U419 ( .A(n2726), .Q(n2724) );
  NAND22 U420 ( .A(n988), .B(n2636), .Q(n2621) );
  INV12 U421 ( .A(n363), .Q(n365) );
  INV3 U422 ( .A(n290), .Q(n289) );
  INV3 U423 ( .A(n1339), .Q(n155) );
  NOR23 U424 ( .A(n869), .B(n1347), .Q(n327) );
  INV3 U425 ( .A(n1191), .Q(n222) );
  NAND31 U426 ( .A(n1821), .B(n1820), .C(n1819), .Q(alu_o_data_AluRes[5]) );
  AOI211 U427 ( .A(n1155), .B(n1987), .C(n1986), .Q(n2009) );
  NAND33 U428 ( .A(u_alu_pre_sum_4b[4]), .B(n2919), .C(n659), .Q(n3053) );
  NAND31 U429 ( .A(n659), .B(n2919), .C(u_alu_pre_sum_4b[6]), .Q(n1059) );
  NAND22 U430 ( .A(n517), .B(n139), .Q(n2478) );
  NOR22 U431 ( .A(n2467), .B(n191), .Q(n2475) );
  INV3 U432 ( .A(n1167), .Q(n399) );
  NOR22 U433 ( .A(n1471), .B(n1470), .Q(n2469) );
  NOR21 U434 ( .A(n1637), .B(n1627), .Q(n388) );
  AOI221 U435 ( .A(i_data_FMmemout[26]), .B(n142), .C(i_data_FMalures[26]), 
        .D(n456), .Q(n10) );
  INV3 U436 ( .A(n10), .Q(n1429) );
  OAI222 U437 ( .A(n1387), .B(n353), .C(n1386), .D(n220), .Q(n11) );
  INV3 U438 ( .A(n11), .Q(n1691) );
  AOI211 U439 ( .A(n945), .B(n386), .C(n2928), .Q(n12) );
  NAND20 U440 ( .A(n680), .B(n322), .Q(n13) );
  NAND22 U441 ( .A(n12), .B(n13), .Q(n1652) );
  NAND31 U442 ( .A(n1635), .B(n329), .C(n1634), .Q(n14) );
  NOR22 U443 ( .A(n1636), .B(n14), .Q(n3158) );
  AOI210 U444 ( .A(n1153), .B(n3115), .C(n3116), .Q(n15) );
  IMUX21 U445 ( .A(n3118), .B(n3117), .S(compare_i_data_rs[30]), .Q(n16) );
  OAI212 U446 ( .A(n380), .B(n3123), .C(n3122), .Q(n17) );
  NOR31 U447 ( .A(n15), .B(n16), .C(n17), .Q(n3124) );
  INV3 U448 ( .A(i_data_FWmemout[25]), .Q(n18) );
  OAI212 U449 ( .A(n941), .B(n18), .C(n1180), .Q(n19) );
  INV6 U450 ( .A(n19), .Q(n696) );
  CLKIN0 U451 ( .A(n2112), .Q(n20) );
  INV3 U452 ( .A(n2119), .Q(n21) );
  NOR41 U453 ( .A(n1156), .B(n2326), .C(n20), .D(n21), .Q(n2123) );
  AOI211 U454 ( .A(n365), .B(n1940), .C(n1775), .Q(n626) );
  AOI221 U455 ( .A(n9), .B(i_data_FMalures[0]), .C(i_data_FMmemout[0]), .D(
        n141), .Q(n22) );
  NAND22 U456 ( .A(n22), .B(n468), .Q(n467) );
  OAI222 U457 ( .A(n1307), .B(n351), .C(n1306), .D(n347), .Q(n23) );
  INV3 U458 ( .A(n23), .Q(n1133) );
  OAI212 U459 ( .A(n1171), .B(n2895), .C(n2486), .Q(n24) );
  AOI221 U460 ( .A(n410), .B(n2487), .C(n386), .D(n24), .Q(n2675) );
  OAI212 U461 ( .A(n3167), .B(n1946), .C(n2804), .Q(n25) );
  NAND20 U462 ( .A(n2801), .B(n1153), .Q(n26) );
  AOI211 U463 ( .A(n26), .B(n387), .C(n25), .Q(n2805) );
  AOI210 U464 ( .A(n413), .B(n367), .C(n422), .Q(n27) );
  NAND20 U465 ( .A(n146), .B(n367), .Q(n28) );
  IMUX20 U466 ( .A(n27), .B(n28), .S(n418), .Q(n1747) );
  NOR21 U467 ( .A(n2415), .B(n2416), .Q(n29) );
  NAND31 U468 ( .A(n29), .B(n2417), .C(n611), .Q(n2418) );
  OAI222 U469 ( .A(n1305), .B(n353), .C(n1304), .D(n347), .Q(n30) );
  INV3 U470 ( .A(n30), .Q(n1139) );
  NAND31 U471 ( .A(n1547), .B(n1546), .C(n1548), .Q(n31) );
  NAND20 U472 ( .A(n364), .B(n1549), .Q(n32) );
  NAND22 U473 ( .A(n31), .B(n32), .Q(n1952) );
  OAI311 U474 ( .A(n2561), .B(n2560), .C(n662), .D(n377), .Q(n33) );
  INV3 U475 ( .A(n2574), .Q(n34) );
  NOR22 U476 ( .A(n33), .B(n34), .Q(n2637) );
  AOI210 U477 ( .A(n413), .B(n2982), .C(n422), .Q(n35) );
  NAND20 U478 ( .A(n146), .B(n2982), .Q(n36) );
  IMUX20 U479 ( .A(n35), .B(n36), .S(n406), .Q(n2082) );
  INV3 U480 ( .A(n537), .Q(n37) );
  NAND22 U481 ( .A(n538), .B(n37), .Q(n38) );
  AOI221 U482 ( .A(n1166), .B(n38), .C(n2779), .D(n401), .Q(n2852) );
  IMUX20 U483 ( .A(n413), .B(n376), .S(u_alu_lt_x_11_A_3_), .Q(n39) );
  AOI210 U484 ( .A(n1153), .B(n39), .C(n367), .Q(n1746) );
  NAND20 U485 ( .A(n628), .B(n1775), .Q(n40) );
  OAI210 U486 ( .A(u_alu_lt_x_11_n129), .B(n40), .C(u_alu_lt_x_11_n130), .Q(
        n41) );
  OAI210 U487 ( .A(u_alu_lt_x_11_n115), .B(u_alu_lt_x_11_n118), .C(
        u_alu_lt_x_11_n116), .Q(n42) );
  AOI210 U488 ( .A(u_alu_lt_x_11_n113), .B(n41), .C(n42), .Q(
        u_alu_lt_x_11_n112) );
  AOI212 U489 ( .A(i_data_FMmemout[5]), .B(n141), .C(n1289), .Q(n43) );
  AOI212 U490 ( .A(n1157), .B(i_data_FWmemout[5]), .C(n1287), .Q(n44) );
  NAND22 U491 ( .A(n43), .B(n44), .Q(n1807) );
  IMUX20 U492 ( .A(n425), .B(n1154), .S(n242), .Q(n45) );
  OAI210 U493 ( .A(n422), .B(n45), .C(n372), .Q(n46) );
  OAI210 U494 ( .A(n1872), .B(n2654), .C(n46), .Q(n1843) );
  INV3 U495 ( .A(n1695), .Q(n47) );
  NOR22 U496 ( .A(n1542), .B(n47), .Q(n1036) );
  AOI211 U497 ( .A(n141), .B(i_data_FMmemout[9]), .C(n237), .Q(n49) );
  NAND22 U498 ( .A(n48), .B(n49), .Q(n236) );
  OAI210 U499 ( .A(n1942), .B(n1941), .C(n626), .Q(n50) );
  NOR21 U500 ( .A(n1935), .B(n968), .Q(n51) );
  OAI212 U501 ( .A(n1943), .B(n51), .C(n50), .Q(n1944) );
  CLKIN0 U502 ( .A(i_data_FWmemout[21]), .Q(n52) );
  NOR22 U503 ( .A(n220), .B(n52), .Q(n1455) );
  OAI212 U504 ( .A(n386), .B(n193), .C(n1607), .Q(n53) );
  NAND22 U505 ( .A(n2671), .B(n253), .Q(n54) );
  OAI2112 U506 ( .A(n3162), .B(n2896), .C(n53), .D(n54), .Q(n1754) );
  OAI212 U507 ( .A(n386), .B(n2981), .C(n55), .Q(n2403) );
  NAND22 U508 ( .A(n1135), .B(i_data_FMalures[16]), .Q(n56) );
  OAI212 U509 ( .A(n1159), .B(n1506), .C(n56), .Q(n1507) );
  AOI220 U510 ( .A(n369), .B(n3121), .C(compare_i_data_rs[19]), .D(n806), .Q(
        n57) );
  NAND22 U511 ( .A(n808), .B(n57), .Q(n58) );
  AOI211 U512 ( .A(n2627), .B(n1874), .C(n58), .Q(n2604) );
  NAND34 U513 ( .A(n636), .B(n1445), .C(n637), .Q(compare_i_data_rs[24]) );
  IMUX20 U514 ( .A(n425), .B(n1154), .S(u_alu_lt_x_11_A_5_), .Q(n59) );
  OAI210 U515 ( .A(n422), .B(n59), .C(u_alu_lt_x_11_B_5_), .Q(n60) );
  OAI210 U516 ( .A(n1812), .B(n3074), .C(n60), .Q(n1813) );
  NOR31 U517 ( .A(n1882), .B(n1879), .C(n1880), .Q(n61) );
  AOI311 U518 ( .A(n1881), .B(n1883), .C(n1879), .D(n61), .Q(n1897) );
  IMUX20 U519 ( .A(n2852), .B(n2780), .S(n400), .Q(n2787) );
  NAND33 U520 ( .A(n2363), .B(n2286), .C(n2364), .Q(n2349) );
  AOI2110 U521 ( .A(n383), .B(i_data_rt[3]), .C(n1735), .D(n1736), .Q(n62) );
  CLKIN0 U522 ( .A(n364), .Q(n63) );
  AOI311 U523 ( .A(n1739), .B(n62), .C(n63), .D(n2593), .Q(n64) );
  NAND22 U524 ( .A(u_alu_lt_x_11_A_3_), .B(n64), .Q(n2386) );
  OAI212 U525 ( .A(n1300), .B(n220), .C(n1302), .Q(n65) );
  NOR22 U526 ( .A(n761), .B(n65), .Q(n876) );
  NOR20 U527 ( .A(n3054), .B(compare_i_data_rs[29]), .Q(n66) );
  INV3 U528 ( .A(n66), .Q(u_alu_DP_OP_84J3_125_2615_n109) );
  AOI221 U529 ( .A(i_data_FMalures[16]), .B(n1135), .C(i_data_FEalures[16]), 
        .D(n454), .Q(n67) );
  NAND22 U530 ( .A(n393), .B(i_data_rt[16]), .Q(n68) );
  NAND22 U531 ( .A(n67), .B(n68), .Q(n290) );
  IMUX20 U532 ( .A(n413), .B(n376), .S(n625), .Q(n69) );
  AOI210 U533 ( .A(n1153), .B(n69), .C(n1774), .Q(n1788) );
  XNR21 U534 ( .A(n1862), .B(n1861), .Q(n70) );
  OAI212 U535 ( .A(n1868), .B(n2238), .C(n711), .Q(n71) );
  AOI212 U536 ( .A(n70), .B(n404), .C(n71), .Q(n1900) );
  INV3 U537 ( .A(n2044), .Q(n72) );
  IMUX21 U538 ( .A(n2056), .B(n72), .S(n400), .Q(n2045) );
  IMUX20 U539 ( .A(n2851), .B(n2850), .S(compare_i_data_rs[24]), .Q(n73) );
  AOI210 U540 ( .A(u_alu_lt_x_11_B_8_), .B(n3121), .C(n73), .Q(n74) );
  OAI212 U541 ( .A(n3074), .B(n2852), .C(n74), .Q(n2884) );
  NAND22 U542 ( .A(n456), .B(i_data_FMalures[15]), .Q(n75) );
  INV3 U543 ( .A(n75), .Q(n790) );
  AOI212 U544 ( .A(n2440), .B(u_alu_lt_x_11_n84), .C(n2431), .Q(n2432) );
  INV3 U545 ( .A(n1481), .Q(n76) );
  NAND33 U546 ( .A(n1691), .B(n1385), .C(n76), .Q(n251) );
  OAI212 U547 ( .A(n1261), .B(n220), .C(n1267), .Q(n77) );
  INV3 U548 ( .A(n77), .Q(n233) );
  NOR21 U549 ( .A(n397), .B(n2043), .Q(n78) );
  INV3 U550 ( .A(n2503), .Q(n79) );
  IMUX21 U551 ( .A(n79), .B(n2568), .S(n401), .Q(n2545) );
  NAND20 U552 ( .A(n2624), .B(n2620), .Q(n80) );
  INV3 U553 ( .A(n80), .Q(n2589) );
  CLKIN0 U554 ( .A(u_alu_DP_OP_84J3_125_2615_n5), .Q(n81) );
  OAI212 U555 ( .A(u_alu_DP_OP_84J3_125_2615_n39), .B(
        u_alu_DP_OP_84J3_125_2615_n45), .C(u_alu_DP_OP_84J3_125_2615_n40), .Q(
        n82) );
  IMUX21 U556 ( .A(n81), .B(u_alu_DP_OP_84J3_125_2615_n5), .S(n82), .Q(n567)
         );
  XNR20 U557 ( .A(n145), .B(alu_i_data_B[31]), .Q(u_alu_DP_OP_84J3_125_2615_n1) );
  INV3 U558 ( .A(compare_i_data_rs[21]), .Q(n83) );
  NAND33 U559 ( .A(n2669), .B(n2668), .C(n83), .Q(n2726) );
  NAND22 U560 ( .A(n1134), .B(i_data_FMalures[26]), .Q(n84) );
  OAI212 U561 ( .A(n1159), .B(n1384), .C(n84), .Q(n1199) );
  IMUX20 U562 ( .A(n413), .B(n376), .S(n3192), .Q(n85) );
  AOI210 U563 ( .A(n1153), .B(n85), .C(n2895), .Q(n1666) );
  AOI210 U564 ( .A(n413), .B(n1774), .C(n422), .Q(n86) );
  NAND20 U565 ( .A(n146), .B(n1774), .Q(n87) );
  IMUX20 U566 ( .A(n86), .B(n87), .S(n1775), .Q(n1787) );
  NAND31 U567 ( .A(n421), .B(n953), .C(n404), .Q(n88) );
  INV3 U568 ( .A(n88), .Q(n2447) );
  AOI221 U569 ( .A(n400), .B(n1715), .C(n1164), .D(n1676), .Q(n89) );
  AOI211 U570 ( .A(n1155), .B(n1708), .C(n1707), .Q(n90) );
  OAI212 U571 ( .A(n380), .B(n89), .C(n90), .Q(alu_o_data_AluRes[2]) );
  CLKIN0 U572 ( .A(i_data_FMalures[1]), .Q(n91) );
  NOR21 U573 ( .A(n1111), .B(n91), .Q(n349) );
  INV3 U574 ( .A(u_alu_lt_x_11_n91), .Q(n92) );
  AOI310 U575 ( .A(n408), .B(n446), .C(n1003), .D(n92), .Q(u_alu_lt_x_11_n87)
         );
  INV3 U576 ( .A(n1385), .Q(n93) );
  NOR22 U577 ( .A(n1481), .B(n93), .Q(n1692) );
  NAND22 U578 ( .A(n1242), .B(n1805), .Q(n94) );
  AOI310 U579 ( .A(n2145), .B(n2150), .C(n2149), .D(n2144), .Q(n95) );
  AOI212 U580 ( .A(n227), .B(n226), .C(n95), .Q(n2348) );
  INV3 U581 ( .A(n2725), .Q(n96) );
  NAND33 U582 ( .A(n374), .B(u_alu_lt_x_11_n50), .C(n96), .Q(n2844) );
  NAND30 U583 ( .A(n444), .B(n146), .C(n431), .Q(n97) );
  OAI210 U584 ( .A(n3068), .B(n3167), .C(n97), .Q(n3063) );
  OAI212 U585 ( .A(i_con_Ealuop[3]), .B(n1556), .C(i_con_Ealuop[1]), .Q(n98)
         );
  NOR21 U586 ( .A(n1555), .B(i_con_Ealuop[2]), .Q(n99) );
  OAI212 U587 ( .A(n98), .B(n99), .C(n1148), .Q(n1582) );
  NAND22 U588 ( .A(n1167), .B(n185), .Q(n100) );
  AOI211 U589 ( .A(n1907), .B(n1168), .C(n100), .Q(n101) );
  AOI211 U590 ( .A(n1908), .B(n362), .C(n101), .Q(n2043) );
  OAI212 U591 ( .A(n2384), .B(n2385), .C(n2383), .Q(n102) );
  NAND22 U592 ( .A(n1961), .B(n102), .Q(n170) );
  INV3 U593 ( .A(n2357), .Q(n103) );
  NOR22 U594 ( .A(n2359), .B(n103), .Q(n2304) );
  INV3 U595 ( .A(n2600), .Q(n104) );
  AOI222 U596 ( .A(n362), .B(n104), .C(n2778), .D(n1167), .Q(n2677) );
  OAI222 U597 ( .A(n1323), .B(n220), .C(n1324), .D(n352), .Q(n105) );
  INV3 U598 ( .A(n105), .Q(n831) );
  NAND22 U599 ( .A(n757), .B(n427), .Q(n106) );
  NAND22 U600 ( .A(u_alu_DP_OP_84J3_125_2615_n40), .B(n106), .Q(
        u_alu_DP_OP_84J3_125_2615_n95) );
  IMUX20 U601 ( .A(n425), .B(n1154), .S(u_alu_lt_x_11_A_10_), .Q(n107) );
  OAI210 U602 ( .A(n422), .B(n107), .C(n2027), .Q(n108) );
  OAI212 U603 ( .A(n2035), .B(n2017), .C(n108), .Q(n2025) );
  NAND22 U604 ( .A(n2504), .B(n1163), .Q(n109) );
  OAI212 U605 ( .A(n2545), .B(n1164), .C(n109), .Q(n2509) );
  AOI210 U606 ( .A(n2588), .B(n2621), .C(n412), .Q(n110) );
  XNR20 U607 ( .A(n110), .B(n2589), .Q(n2607) );
  AOI212 U608 ( .A(n2818), .B(n2729), .C(n2811), .Q(n111) );
  NOR21 U609 ( .A(n111), .B(n2757), .Q(n112) );
  AOI2111 U610 ( .A(n111), .B(n2757), .C(n2784), .D(n112), .Q(n2730) );
  XNR21 U611 ( .A(n2792), .B(n2791), .Q(n113) );
  OAI212 U612 ( .A(n380), .B(n2806), .C(n2805), .Q(n114) );
  AOI212 U613 ( .A(n113), .B(n3175), .C(n114), .Q(n2807) );
  CLKIN0 U614 ( .A(u_alu_DP_OP_84J3_125_2615_n50), .Q(n115) );
  NOR21 U615 ( .A(u_alu_DP_OP_84J3_125_2615_n49), .B(n115), .Q(
        u_alu_pre_sum_4a[0]) );
  OAI212 U616 ( .A(n1326), .B(n1158), .C(n1327), .Q(n116) );
  INV3 U617 ( .A(n116), .Q(n2474) );
  NOR21 U618 ( .A(n1541), .B(n1542), .Q(n117) );
  CLKIN0 U619 ( .A(n1804), .Q(n118) );
  NOR31 U620 ( .A(n1786), .B(n1788), .C(n1787), .Q(n119) );
  OAI2112 U621 ( .A(n426), .B(n118), .C(n1789), .D(n119), .Q(
        alu_o_data_AluRes[4]) );
  MUX21 U622 ( .A(n2487), .B(n1972), .S(n410), .Q(n2180) );
  OAI210 U623 ( .A(n452), .B(u_alu_lt_x_11_B_20_), .C(u_alu_lt_x_11_n47), .Q(
        u_alu_lt_x_11_n45) );
  NOR30 U624 ( .A(n379), .B(n400), .C(n458), .Q(n308) );
  AOI210 U625 ( .A(u_alu_lt_x_11_B_1_), .B(n875), .C(n2413), .Q(n120) );
  NOR20 U626 ( .A(n1660), .B(u_alu_lt_x_11_A_0_), .Q(n121) );
  XNR20 U627 ( .A(n120), .B(n121), .Q(n1661) );
  CLKIN0 U628 ( .A(n2833), .Q(n122) );
  IMUX20 U629 ( .A(n122), .B(n2833), .S(n2546), .Q(n459) );
  NAND20 U630 ( .A(alu_i_data_B[31]), .B(n144), .Q(n123) );
  NAND20 U631 ( .A(n1591), .B(n123), .Q(n124) );
  OAI310 U632 ( .A(n445), .B(n1603), .C(n1636), .D(n124), .Q(n602) );
  IMUX20 U633 ( .A(n413), .B(n376), .S(u_alu_lt_x_11_A_12_), .Q(n125) );
  AOI210 U634 ( .A(n1153), .B(n125), .C(n2113), .Q(n2122) );
  OAI210 U635 ( .A(n425), .B(u_alu_lt_x_11_B_15_), .C(n1153), .Q(n126) );
  NOR20 U636 ( .A(u_alu_lt_x_11_B_15_), .B(n2948), .Q(n127) );
  OAI210 U637 ( .A(n424), .B(n2322), .C(u_alu_lt_x_11_B_15_), .Q(n128) );
  IMUX20 U638 ( .A(n126), .B(n127), .S(n2363), .Q(n129) );
  NAND20 U639 ( .A(n128), .B(n129), .Q(n2323) );
  IMUX20 U640 ( .A(u_alu_pre_sum_4a[0]), .B(n927), .S(n943), .Q(n2888) );
  XNR20 U641 ( .A(n757), .B(u_alu_DP_OP_84J3_125_2615_n6), .Q(
        u_alu_pre_sum_4b[2]) );
  NAND40 U642 ( .A(n1110), .B(n1487), .C(n1405), .D(n864), .Q(n130) );
  CLKIN0 U643 ( .A(n130), .Q(n131) );
  NAND20 U644 ( .A(n1488), .B(n131), .Q(n3190) );
  NAND33 U645 ( .A(n651), .B(n1959), .C(n652), .Q(n169) );
  NAND23 U646 ( .A(n652), .B(n630), .Q(n629) );
  NAND33 U647 ( .A(n2604), .B(n2605), .C(n2603), .Q(n2606) );
  NAND26 U648 ( .A(n398), .B(i_data_rs[4]), .Q(n219) );
  AOI211 U649 ( .A(n1135), .B(i_data_FMalures[23]), .C(n1329), .Q(n1408) );
  NAND24 U650 ( .A(n1201), .B(n730), .Q(n729) );
  NOR31 U651 ( .A(n380), .B(n280), .C(n279), .Q(n820) );
  NAND22 U652 ( .A(n1511), .B(n391), .Q(n576) );
  NAND34 U653 ( .A(n2317), .B(n2318), .C(n2316), .Q(n2319) );
  NAND33 U654 ( .A(u_alu_pre_sum_4b[7]), .B(n2919), .C(n659), .Q(n3179) );
  AOI212 U655 ( .A(n2040), .B(n404), .C(n2039), .Q(n2047) );
  NAND24 U656 ( .A(n1134), .B(i_data_FMalures[22]), .Q(n1337) );
  NAND22 U657 ( .A(n2350), .B(n2349), .Q(n2352) );
  NAND23 U658 ( .A(n1210), .B(n1209), .Q(n1211) );
  NAND33 U659 ( .A(n2271), .B(n2269), .C(n2235), .Q(n2236) );
  NAND23 U660 ( .A(n2300), .B(n478), .Q(n2271) );
  INV15 U661 ( .A(n420), .Q(n132) );
  XNR22 U662 ( .A(n3087), .B(n3086), .Q(n3126) );
  NAND23 U663 ( .A(n991), .B(n2832), .Q(n990) );
  NAND23 U664 ( .A(n2477), .B(n591), .Q(n590) );
  NAND23 U665 ( .A(n1136), .B(i_data_FMmemout[17]), .Q(n2472) );
  NOR32 U666 ( .A(n1645), .B(n1644), .C(n1643), .Q(n1646) );
  INV3 U667 ( .A(n2595), .Q(n1740) );
  NAND26 U668 ( .A(n710), .B(n1174), .Q(n1120) );
  INV12 U669 ( .A(n2186), .Q(n1138) );
  NAND23 U670 ( .A(n1934), .B(n1933), .Q(n1959) );
  INV8 U671 ( .A(n1757), .Q(n913) );
  AOI211 U672 ( .A(n1137), .B(i_data_FMmemout[1]), .C(n1544), .Q(n1547) );
  NAND28 U673 ( .A(n204), .B(n2441), .Q(n202) );
  NAND26 U674 ( .A(n1028), .B(n2441), .Q(n2847) );
  NOR22 U675 ( .A(n2425), .B(n2424), .Q(n2426) );
  NAND24 U676 ( .A(n902), .B(n901), .Q(n942) );
  NAND24 U677 ( .A(n2020), .B(n2019), .Q(n2257) );
  INV6 U678 ( .A(n809), .Q(n2673) );
  AOI212 U679 ( .A(n1163), .B(n2570), .C(n2569), .Q(n2571) );
  CLKBU15 U680 ( .A(n594), .Q(n220) );
  NOR24 U681 ( .A(n709), .B(n1097), .Q(n1096) );
  INV15 U682 ( .A(n741), .Q(n1097) );
  CLKBU12 U683 ( .A(n1160), .Q(n454) );
  NAND26 U684 ( .A(n165), .B(n391), .Q(n2063) );
  NAND23 U685 ( .A(n514), .B(n744), .Q(n1117) );
  AOI212 U686 ( .A(n747), .B(n2424), .C(n513), .Q(n514) );
  CLKBU12 U687 ( .A(n594), .Q(n292) );
  NAND24 U688 ( .A(n706), .B(n705), .Q(n898) );
  NOR23 U689 ( .A(i_data_immext[2]), .B(n1564), .Q(n716) );
  NOR23 U690 ( .A(n498), .B(n497), .Q(n545) );
  NAND22 U691 ( .A(n2855), .B(n2854), .Q(n2858) );
  NAND24 U692 ( .A(n3183), .B(n139), .Q(n254) );
  NAND22 U693 ( .A(n1135), .B(i_data_FMalures[29]), .Q(n1189) );
  NAND22 U694 ( .A(n1134), .B(i_data_FMalures[10]), .Q(n1229) );
  NAND22 U695 ( .A(n1135), .B(i_data_FMalures[25]), .Q(n1181) );
  NAND22 U696 ( .A(n1135), .B(i_data_FMalures[31]), .Q(n1175) );
  NAND22 U697 ( .A(n1134), .B(i_data_FMalures[30]), .Q(n1185) );
  NAND22 U698 ( .A(n1134), .B(i_data_FMalures[17]), .Q(n1327) );
  NAND23 U699 ( .A(n2835), .B(n451), .Q(n2836) );
  NAND34 U700 ( .A(n862), .B(n1220), .C(n861), .Q(n133) );
  NAND28 U701 ( .A(n617), .B(n377), .Q(alu_i_data_B[31]) );
  AOI212 U702 ( .A(n1161), .B(i_data_rt[26]), .C(n1199), .Q(n670) );
  OAI212 U703 ( .A(n2333), .B(n3074), .C(n2332), .Q(n2334) );
  NAND26 U704 ( .A(n1098), .B(n725), .Q(n1099) );
  NOR22 U705 ( .A(n3192), .B(u_alu_lt_x_11_B_1_), .Q(n1764) );
  INV6 U706 ( .A(n1061), .Q(n1146) );
  INV6 U707 ( .A(n2828), .Q(n291) );
  NAND26 U708 ( .A(n781), .B(n780), .Q(n895) );
  NAND26 U709 ( .A(n1120), .B(n1097), .Q(n739) );
  INV6 U710 ( .A(i_data_immext[5]), .Q(n1561) );
  NAND23 U711 ( .A(compare_i_data_rt[27]), .B(n139), .Q(n1605) );
  NAND26 U712 ( .A(n1197), .B(n1196), .Q(compare_i_data_rt[27]) );
  AOI212 U713 ( .A(n2690), .B(n2607), .C(n2606), .Q(n2608) );
  INV3 U714 ( .A(n2190), .Q(n2167) );
  NAND33 U715 ( .A(n1492), .B(n1491), .C(n1490), .Q(n1493) );
  NOR23 U716 ( .A(n374), .B(n2725), .Q(n2723) );
  NOR24 U717 ( .A(n893), .B(n895), .Q(n889) );
  NAND28 U718 ( .A(n779), .B(n776), .Q(n893) );
  NOR24 U719 ( .A(n777), .B(n778), .Q(n776) );
  NAND34 U720 ( .A(n1450), .B(n152), .C(n1341), .Q(n1343) );
  INV6 U721 ( .A(u_alu_lt_x_11_A_12_), .Q(n408) );
  INV8 U722 ( .A(n2127), .Q(n448) );
  AOI212 U723 ( .A(n2289), .B(n2199), .C(n799), .Q(n2200) );
  NAND23 U724 ( .A(n2952), .B(n440), .Q(n2156) );
  NAND28 U725 ( .A(n234), .B(n228), .Q(n1310) );
  NOR33 U726 ( .A(n1167), .B(n458), .C(n3101), .Q(n3102) );
  OAI212 U727 ( .A(n2869), .B(n2868), .C(n1168), .Q(n1065) );
  NAND34 U728 ( .A(n258), .B(n1679), .C(n1680), .Q(compare_i_data_rt[1]) );
  NOR22 U729 ( .A(n1501), .B(n364), .Q(n1502) );
  NAND24 U730 ( .A(n1670), .B(n2477), .Q(u_alu_lt_x_11_B_17_) );
  NAND26 U731 ( .A(n221), .B(n377), .Q(n3054) );
  NOR24 U732 ( .A(n506), .B(n505), .Q(n2103) );
  AOI212 U733 ( .A(n383), .B(i_data_rt[10]), .C(n481), .Q(n480) );
  NAND26 U734 ( .A(n2554), .B(n2553), .Q(n1325) );
  NAND24 U735 ( .A(n134), .B(n135), .Q(n137) );
  NAND24 U736 ( .A(n136), .B(n137), .Q(n772) );
  CLKIN6 U737 ( .A(u_alu_lt_x_11_A_0_), .Q(n135) );
  INV8 U738 ( .A(compare_i_data_rt[0]), .Q(n360) );
  INV12 U739 ( .A(n604), .Q(n354) );
  NAND24 U740 ( .A(n604), .B(n411), .Q(n725) );
  NOR22 U741 ( .A(n1162), .B(n1127), .Q(n1126) );
  NOR22 U742 ( .A(n1356), .B(n1159), .Q(n582) );
  NOR33 U743 ( .A(n1483), .B(n1482), .C(n1484), .Q(n1486) );
  OAI222 U744 ( .A(n3036), .B(n400), .C(n3062), .D(n1163), .Q(n3039) );
  NAND24 U745 ( .A(n623), .B(n1198), .Q(n1200) );
  INV3 U746 ( .A(n624), .Q(n623) );
  AOI212 U747 ( .A(n378), .B(n2953), .C(n964), .Q(n963) );
  NAND23 U748 ( .A(n1006), .B(n1275), .Q(n1686) );
  AOI211 U749 ( .A(n2640), .B(n410), .C(n2643), .Q(n2399) );
  NAND28 U750 ( .A(n1215), .B(n1214), .Q(n242) );
  NOR22 U751 ( .A(n1116), .B(n1115), .Q(n835) );
  NOR22 U752 ( .A(n416), .B(n2139), .Q(n252) );
  NOR23 U753 ( .A(n436), .B(n2139), .Q(n2368) );
  NAND24 U754 ( .A(n583), .B(n139), .Q(n633) );
  NOR23 U755 ( .A(n1595), .B(n1574), .Q(n1578) );
  AOI211 U756 ( .A(n3160), .B(n1153), .C(n3162), .Q(n3171) );
  INV12 U757 ( .A(n140), .Q(n142) );
  INV8 U758 ( .A(n1390), .Q(n140) );
  NAND28 U759 ( .A(n432), .B(n1649), .Q(n2518) );
  NOR32 U760 ( .A(n3171), .B(n3170), .C(n3169), .Q(n3172) );
  NOR22 U761 ( .A(n1569), .B(n1576), .Q(n1635) );
  NAND24 U762 ( .A(n1582), .B(n1557), .Q(n1576) );
  NOR24 U763 ( .A(n400), .B(n379), .Q(n850) );
  INV6 U764 ( .A(n2834), .Q(n1162) );
  NAND22 U765 ( .A(i_data_immext[16]), .B(i_con_Ealusrc), .Q(n2834) );
  INV12 U766 ( .A(n1171), .Q(n1170) );
  INV15 U767 ( .A(i_data_immext[10]), .Q(n1171) );
  INV6 U768 ( .A(n144), .Q(n145) );
  NAND22 U769 ( .A(n201), .B(n200), .Q(n375) );
  INV6 U770 ( .A(n375), .Q(n376) );
  BUF2 U771 ( .A(n387), .Q(n253) );
  NOR22 U772 ( .A(u_alu_lt_x_11_B_14_), .B(n336), .Q(n2353) );
  NAND22 U773 ( .A(n393), .B(i_data_rt[5]), .Q(n1243) );
  NAND24 U774 ( .A(n634), .B(n633), .Q(u_alu_lt_x_11_B_9_) );
  INV6 U775 ( .A(n355), .Q(n356) );
  CLKIN4 U776 ( .A(n979), .Q(n355) );
  INV8 U777 ( .A(n1153), .Q(n424) );
  INV3 U778 ( .A(n368), .Q(n367) );
  INV3 U779 ( .A(n2636), .Q(compare_i_data_rs[18]) );
  INV3 U780 ( .A(n378), .Q(n380) );
  INV8 U781 ( .A(n1151), .Q(n378) );
  INV3 U782 ( .A(n329), .Q(n445) );
  BUF6 U783 ( .A(n1637), .Q(n329) );
  NAND26 U784 ( .A(n3009), .B(n414), .Q(n3010) );
  BUF6 U785 ( .A(n3177), .Q(n1145) );
  INV3 U786 ( .A(n410), .Q(n186) );
  INV12 U787 ( .A(n140), .Q(n141) );
  NAND22 U788 ( .A(n1647), .B(n308), .Q(n307) );
  INV3 U789 ( .A(n2896), .Q(n322) );
  NAND26 U790 ( .A(n1013), .B(n1822), .Q(n1931) );
  INV3 U791 ( .A(n2129), .Q(n164) );
  INV6 U792 ( .A(n2165), .Q(n786) );
  INV12 U793 ( .A(n1172), .Q(n363) );
  INV8 U794 ( .A(n389), .Q(n391) );
  INV6 U795 ( .A(u_alu_lt_x_11_B_9_), .Q(n2905) );
  NAND23 U796 ( .A(n1539), .B(n754), .Q(n1543) );
  NAND26 U797 ( .A(n1274), .B(n1273), .Q(compare_i_data_rt[8]) );
  INV6 U798 ( .A(compare_i_data_rt[8]), .Q(n264) );
  INV6 U799 ( .A(n3054), .Q(n431) );
  INV3 U800 ( .A(compare_i_data_rs[31]), .Q(n144) );
  BUF8 U801 ( .A(n1169), .Q(n386) );
  NOR23 U802 ( .A(n1162), .B(n833), .Q(n2477) );
  OAI212 U803 ( .A(n401), .B(n2936), .C(n2899), .Q(n2902) );
  NOR22 U804 ( .A(n2654), .B(n2937), .Q(n2899) );
  INV3 U805 ( .A(n349), .Q(n1303) );
  NAND28 U806 ( .A(n189), .B(n188), .Q(compare_i_data_rs[30]) );
  INV6 U807 ( .A(n1410), .Q(n188) );
  NAND24 U808 ( .A(n1942), .B(n391), .Q(n1756) );
  NOR23 U809 ( .A(n138), .B(i_data_immext[3]), .Q(n2593) );
  INV12 U810 ( .A(n1914), .Q(u_alu_lt_x_11_B_5_) );
  NOR23 U811 ( .A(n1471), .B(n191), .Q(n558) );
  INV3 U812 ( .A(n582), .Q(n581) );
  NOR33 U813 ( .A(n791), .B(n790), .C(n1224), .Q(n789) );
  NAND28 U814 ( .A(n787), .B(n785), .Q(compare_i_data_rt[13]) );
  AOI212 U815 ( .A(n2958), .B(n2516), .C(n2515), .Q(n2551) );
  INV12 U816 ( .A(n203), .Q(n2958) );
  INV6 U817 ( .A(n1358), .Q(n1129) );
  NOR22 U818 ( .A(n1736), .B(n1725), .Q(n1364) );
  NAND33 U819 ( .A(n3011), .B(n3010), .C(compare_i_data_rs[24]), .Q(n3015) );
  INV8 U820 ( .A(compare_i_data_rs[24]), .Q(n433) );
  NOR22 U821 ( .A(n2695), .B(n203), .Q(n2696) );
  NOR23 U822 ( .A(n203), .B(n2666), .Q(n1032) );
  NOR23 U823 ( .A(n203), .B(n2917), .Q(n2918) );
  NOR22 U824 ( .A(n203), .B(n919), .Q(n915) );
  NOR23 U825 ( .A(n203), .B(n3000), .Q(n1079) );
  NOR22 U826 ( .A(n379), .B(n2708), .Q(n2709) );
  INV6 U827 ( .A(n522), .Q(n869) );
  AOI212 U828 ( .A(n2379), .B(n2378), .C(n2377), .Q(n839) );
  OAI222 U829 ( .A(n3146), .B(n386), .C(n3145), .D(n410), .Q(n3151) );
  AOI222 U830 ( .A(n1754), .B(n362), .C(n1608), .D(n1167), .Q(n1675) );
  NAND24 U831 ( .A(n2463), .B(n391), .Q(n591) );
  AOI211 U832 ( .A(n2335), .B(n2336), .C(n2334), .Q(n2337) );
  AOI212 U833 ( .A(n2458), .B(n3175), .C(n2457), .Q(n2459) );
  INV15 U834 ( .A(n2847), .Q(n3175) );
  NOR22 U835 ( .A(n1208), .B(n351), .Q(n1212) );
  INV12 U836 ( .A(n350), .Q(n351) );
  CLKBU15 U837 ( .A(n1545), .Q(n1137) );
  AOI222 U838 ( .A(n362), .B(n2403), .C(n2101), .D(n1167), .Q(n2258) );
  BUF15 U839 ( .A(n392), .Q(n138) );
  BUF15 U840 ( .A(n392), .Q(n139) );
  INV8 U841 ( .A(n389), .Q(n392) );
  OAI212 U842 ( .A(n1150), .B(n1094), .C(n1309), .Q(n880) );
  NOR23 U843 ( .A(n872), .B(n871), .Q(n906) );
  NAND26 U844 ( .A(n446), .B(n1171), .Q(n1790) );
  NOR22 U845 ( .A(n2396), .B(n2395), .Q(n257) );
  AOI211 U846 ( .A(n456), .B(i_data_FMalures[22]), .C(n1449), .Q(n1450) );
  INV3 U847 ( .A(n2835), .Q(n1863) );
  NAND26 U848 ( .A(n821), .B(n377), .Q(n2835) );
  NAND23 U849 ( .A(n495), .B(n480), .Q(compare_i_data_rt[10]) );
  INV6 U850 ( .A(n2635), .Q(n2829) );
  NOR21 U851 ( .A(n364), .B(n2243), .Q(n2244) );
  NAND28 U852 ( .A(n192), .B(compare_i_data_rs[15]), .Q(n2357) );
  AOI212 U853 ( .A(n458), .B(n1992), .C(n1991), .Q(n2023) );
  INV6 U854 ( .A(n2822), .Q(n2771) );
  OAI212 U855 ( .A(n362), .B(n2716), .C(n2522), .Q(n2523) );
  INV6 U856 ( .A(n140), .Q(n143) );
  NAND24 U857 ( .A(n393), .B(i_data_rt[24]), .Q(n522) );
  NAND23 U858 ( .A(n694), .B(n1456), .Q(n690) );
  OAI212 U859 ( .A(n2197), .B(n2188), .C(n2187), .Q(n2195) );
  NAND24 U860 ( .A(n454), .B(i_data_FEalures[13]), .Q(n2188) );
  NOR24 U861 ( .A(n420), .B(n1863), .Q(n2565) );
  AOI222 U862 ( .A(n362), .B(n1905), .C(n1754), .D(n1167), .Q(n1827) );
  NAND23 U863 ( .A(n554), .B(n553), .Q(n681) );
  NAND26 U864 ( .A(n1554), .B(n1568), .Q(n1588) );
  OAI212 U865 ( .A(n1553), .B(n1570), .C(n457), .Q(n1554) );
  NOR23 U866 ( .A(n2124), .B(n2027), .Q(n2109) );
  NAND26 U867 ( .A(n848), .B(n1006), .Q(compare_i_data_rt[0]) );
  NAND24 U868 ( .A(n868), .B(n866), .Q(compare_i_data_rt[4]) );
  OAI210 U869 ( .A(n422), .B(n1965), .C(u_alu_lt_x_11_B_8_), .Q(n1966) );
  NOR24 U870 ( .A(n3178), .B(n1145), .Q(n2919) );
  BUF15 U871 ( .A(n388), .Q(n146) );
  NAND22 U872 ( .A(n2204), .B(n850), .Q(n2205) );
  AOI212 U873 ( .A(n850), .B(n1773), .C(n1772), .Q(n1789) );
  XOR22 U874 ( .A(n149), .B(n147), .Q(n2785) );
  OAI212 U875 ( .A(n2782), .B(n2820), .C(n2781), .Q(n147) );
  AOI212 U876 ( .A(n2811), .B(n2770), .C(n2769), .Q(n2781) );
  NOR24 U877 ( .A(n148), .B(n2660), .Q(n2820) );
  AOI212 U878 ( .A(n2659), .B(n2658), .C(n2657), .Q(n148) );
  NOR24 U879 ( .A(n442), .B(n2763), .Q(n2815) );
  NOR24 U880 ( .A(n879), .B(n880), .Q(n150) );
  NAND26 U881 ( .A(n150), .B(n1133), .Q(n1039) );
  NAND24 U882 ( .A(n264), .B(n150), .Q(n263) );
  NOR24 U883 ( .A(n2362), .B(n151), .Q(n667) );
  OAI212 U884 ( .A(n2169), .B(n151), .C(n2198), .Q(n2170) );
  OAI212 U885 ( .A(n2254), .B(n151), .C(n2302), .Q(n2255) );
  XNR21 U886 ( .A(n2142), .B(n151), .Q(n948) );
  NOR24 U887 ( .A(n951), .B(n949), .Q(n151) );
  XOR22 U888 ( .A(n3187), .B(n1343), .Q(n777) );
  AOI212 U889 ( .A(n343), .B(i_data_rs[22]), .C(n153), .Q(n152) );
  AOI212 U890 ( .A(n382), .B(i_data_rt[22]), .C(n1338), .Q(n154) );
  NOR24 U891 ( .A(n2198), .B(n156), .Q(n2228) );
  NOR20 U892 ( .A(n156), .B(n2229), .Q(n2201) );
  CLKIN6 U893 ( .A(n2227), .Q(n156) );
  NAND24 U894 ( .A(n2445), .B(u_alu_lt_x_11_B_16_), .Q(n2855) );
  NOR24 U895 ( .A(n2444), .B(n157), .Q(n2445) );
  CLKIN6 U896 ( .A(n2443), .Q(n157) );
  NOR24 U897 ( .A(n1474), .B(n496), .Q(n2443) );
  CLKIN15 U898 ( .A(n1150), .Q(n398) );
  NAND28 U899 ( .A(n1100), .B(n1099), .Q(n1150) );
  NAND28 U900 ( .A(n473), .B(n268), .Q(n1100) );
  AOI212 U901 ( .A(n1187), .B(n139), .C(n1162), .Q(n158) );
  CLKIN6 U902 ( .A(n1187), .Q(n160) );
  NAND24 U903 ( .A(n159), .B(n160), .Q(compare_i_data_rt[30]) );
  OAI212 U904 ( .A(n159), .B(n364), .C(n158), .Q(
        u_alu_DP_OP_84J3_125_2615_n140) );
  AOI212 U905 ( .A(n393), .B(i_data_rt[30]), .C(n1186), .Q(n159) );
  NOR24 U906 ( .A(n161), .B(n1672), .Q(n1829) );
  NOR24 U907 ( .A(n1168), .B(n1671), .Q(n161) );
  NOR24 U908 ( .A(n2487), .B(n162), .Q(n1671) );
  CLKIN6 U909 ( .A(n518), .Q(n162) );
  CLKIN6 U910 ( .A(n870), .Q(n163) );
  NAND24 U911 ( .A(n541), .B(n989), .Q(n165) );
  NAND28 U912 ( .A(n167), .B(n166), .Q(n2186) );
  INV6 U913 ( .A(n2393), .Q(n166) );
  NOR23 U914 ( .A(n1763), .B(n654), .Q(n1961) );
  NAND32 U915 ( .A(n1945), .B(n1944), .C(n1959), .Q(n172) );
  NOR24 U916 ( .A(n1937), .B(n173), .Q(n1815) );
  AOI212 U917 ( .A(n1113), .B(n1241), .C(n1172), .Q(n173) );
  NAND22 U918 ( .A(n175), .B(n1171), .Q(n182) );
  OAI212 U919 ( .A(n2952), .B(n1171), .C(n175), .Q(n174) );
  NAND24 U920 ( .A(n2715), .B(n2714), .Q(n3097) );
  NAND24 U921 ( .A(n179), .B(n176), .Q(n183) );
  NOR24 U922 ( .A(n178), .B(n177), .Q(n176) );
  NOR24 U923 ( .A(n184), .B(n2715), .Q(n177) );
  NOR24 U924 ( .A(n184), .B(n2714), .Q(n178) );
  NOR24 U925 ( .A(n2934), .B(n183), .Q(n3029) );
  NOR24 U926 ( .A(n420), .B(n1142), .Q(n2933) );
  CLKIN3 U927 ( .A(n187), .Q(n2640) );
  NAND28 U928 ( .A(n2147), .B(n2146), .Q(u_alu_lt_x_11_B_8_) );
  XOR22 U929 ( .A(compare_i_data_rt[30]), .B(compare_i_data_rs[30]), .Q(n609)
         );
  NOR33 U930 ( .A(n1411), .B(n1412), .C(n190), .Q(n189) );
  NAND28 U931 ( .A(n2439), .B(n2440), .Q(n1119) );
  NAND28 U932 ( .A(u_alu_lt_x_11_B_15_), .B(n2363), .Q(n2440) );
  NAND28 U933 ( .A(n2286), .B(n2364), .Q(u_alu_lt_x_11_B_15_) );
  BUF8 U934 ( .A(u_alu_lt_x_11_B_15_), .Q(n192) );
  OAI212 U935 ( .A(n197), .B(n194), .C(n1041), .Q(n1040) );
  AOI212 U936 ( .A(n3066), .B(n195), .C(n385), .Q(n194) );
  CLKIN6 U937 ( .A(n196), .Q(n195) );
  NOR24 U938 ( .A(n1171), .B(n1914), .Q(n196) );
  OAI222 U939 ( .A(n3068), .B(n3069), .C(n431), .D(n2870), .Q(n197) );
  CLKIN15 U940 ( .A(n1632), .Q(n200) );
  NAND28 U941 ( .A(n202), .B(n423), .Q(n203) );
  NAND28 U942 ( .A(n2428), .B(n2427), .Q(n2441) );
  INV6 U943 ( .A(n2954), .Q(n204) );
  OAI212 U944 ( .A(n2358), .B(n2359), .C(n2357), .Q(n2380) );
  INV6 U945 ( .A(n205), .Q(n2554) );
  AOI222 U946 ( .A(n1135), .B(i_data_FMalures[19]), .C(n1137), .D(
        i_data_FMmemout[19]), .Q(n207) );
  NAND26 U947 ( .A(n335), .B(n209), .Q(n334) );
  AOI2112 U948 ( .A(n343), .B(i_data_rs[14]), .C(n210), .D(n801), .Q(n209) );
  OAI2112 U949 ( .A(n365), .B(n1197), .C(n377), .D(n212), .Q(n2963) );
  NAND28 U950 ( .A(u_alu_lt_x_11_B_20_), .B(n1171), .Q(n3025) );
  NAND28 U951 ( .A(n2618), .B(n2632), .Q(u_alu_lt_x_11_B_20_) );
  NAND28 U952 ( .A(n628), .B(n1170), .Q(n3024) );
  NAND28 U953 ( .A(n913), .B(n1756), .Q(n628) );
  AOI212 U954 ( .A(n2822), .B(n2818), .C(n2811), .Q(n214) );
  NAND43 U955 ( .A(n1204), .B(n219), .C(n216), .D(n215), .Q(n625) );
  NOR24 U956 ( .A(n1202), .B(n347), .Q(n217) );
  NAND24 U957 ( .A(compare_i_data_rt[29]), .B(n391), .Q(n221) );
  NAND24 U958 ( .A(n223), .B(n222), .Q(compare_i_data_rt[29]) );
  AOI212 U959 ( .A(n1161), .B(i_data_rt[29]), .C(n1190), .Q(n223) );
  NAND24 U960 ( .A(n2155), .B(n224), .Q(n2157) );
  AOI212 U961 ( .A(n2348), .B(n2344), .C(n225), .Q(n224) );
  NAND20 U962 ( .A(n2147), .B(n2146), .Q(n226) );
  CLKIN6 U963 ( .A(n407), .Q(n227) );
  NAND26 U964 ( .A(n233), .B(n232), .Q(u_alu_lt_x_11_A_12_) );
  NOR24 U965 ( .A(n231), .B(n229), .Q(n228) );
  NOR24 U966 ( .A(u_alu_lt_x_11_A_12_), .B(n230), .Q(n229) );
  AOI212 U967 ( .A(n233), .B(n232), .C(compare_i_data_rt[12]), .Q(n231) );
  NAND24 U968 ( .A(n1624), .B(n1260), .Q(compare_i_data_rt[12]) );
  NOR23 U969 ( .A(n346), .B(n345), .Q(n1624) );
  OAI221 U970 ( .A(n263), .B(n1132), .C(n235), .D(n264), .Q(n234) );
  NOR24 U971 ( .A(n236), .B(n802), .Q(n803) );
  NOR24 U972 ( .A(n239), .B(n2192), .Q(n2193) );
  CLKIN6 U973 ( .A(n240), .Q(n239) );
  NAND24 U974 ( .A(n2190), .B(n2189), .Q(n241) );
  NAND28 U975 ( .A(n771), .B(n1238), .Q(n887) );
  CLKIN15 U976 ( .A(n242), .Q(n409) );
  NOR24 U977 ( .A(n246), .B(n243), .Q(n975) );
  XNR22 U978 ( .A(compare_i_data_rt[6]), .B(n409), .Q(n243) );
  NAND24 U979 ( .A(n245), .B(n244), .Q(compare_i_data_rt[6]) );
  NOR24 U980 ( .A(n767), .B(n768), .Q(n244) );
  CLKIN6 U981 ( .A(n1535), .Q(n245) );
  XOR22 U982 ( .A(compare_i_data_rt[7]), .B(n887), .Q(n246) );
  NAND24 U983 ( .A(n248), .B(n247), .Q(compare_i_data_rt[7]) );
  NOR24 U984 ( .A(n551), .B(n549), .Q(n247) );
  CLKIN6 U985 ( .A(n1528), .Q(n248) );
  XOR22 U986 ( .A(n251), .B(n3191), .Q(n572) );
  NAND24 U987 ( .A(n752), .B(n1540), .Q(n1542) );
  CLKIN6 U988 ( .A(n2424), .Q(n2438) );
  NAND24 U989 ( .A(n2108), .B(n2107), .Q(n2424) );
  OAI212 U990 ( .A(n2434), .B(n2436), .C(n2438), .Q(n1005) );
  NOR24 U991 ( .A(n1610), .B(n1611), .Q(n2139) );
  NOR22 U992 ( .A(n387), .B(u_alu_lt_x_11_A_23_), .Q(n2812) );
  NAND28 U993 ( .A(n254), .B(n377), .Q(n387) );
  NAND34 U994 ( .A(n1408), .B(n1407), .C(n1406), .Q(n3183) );
  NAND24 U995 ( .A(n856), .B(n255), .Q(n1779) );
  NAND24 U996 ( .A(n855), .B(n256), .Q(n255) );
  NAND24 U997 ( .A(n419), .B(n257), .Q(n256) );
  NAND28 U998 ( .A(n382), .B(i_data_rt[1]), .Q(n1680) );
  INV6 U999 ( .A(n1681), .Q(n258) );
  NAND22 U1000 ( .A(n1135), .B(i_data_FMalures[1]), .Q(n1546) );
  NOR31 U1001 ( .A(n2423), .B(n260), .C(n593), .Q(n592) );
  NAND34 U1002 ( .A(n2439), .B(n2422), .C(n2440), .Q(n260) );
  CLKIN15 U1003 ( .A(n1107), .Q(u_alu_lt_x_11_B_14_) );
  XNR22 U1004 ( .A(n261), .B(compare_i_data_rt[27]), .Q(n706) );
  NAND43 U1005 ( .A(n1426), .B(n1427), .C(n262), .D(n2810), .Q(n261) );
  NOR24 U1006 ( .A(n1381), .B(n1382), .Q(n2810) );
  MUX22 U1007 ( .A(compare_i_data_rt[3]), .B(i_data_immext[3]), .S(n364), .Q(
        n368) );
  CLKIN6 U1008 ( .A(u_alu_lt_x_11_B_21_), .Q(n441) );
  AOI312 U1009 ( .A(i_data_rt[21]), .B(n391), .C(n383), .D(n1162), .Q(n2668)
         );
  NAND24 U1010 ( .A(n265), .B(u_alu_DP_OP_84J3_125_2615_n48), .Q(
        u_alu_DP_OP_84J3_125_2615_n46) );
  NAND24 U1011 ( .A(n756), .B(n266), .Q(n265) );
  CLKIN6 U1012 ( .A(u_alu_lt_x_11_B_16_), .Q(n1649) );
  CLKIN6 U1013 ( .A(n267), .Q(n2868) );
  BUF15 U1014 ( .A(n270), .Q(n268) );
  CLKIN6 U1015 ( .A(i_con_Efamux[1]), .Q(n269) );
  NOR33 U1016 ( .A(i_con_Efamux[0]), .B(n604), .C(n270), .Q(n1390) );
  CLKIN15 U1017 ( .A(i_con_Efamux[2]), .Q(n604) );
  NAND22 U1018 ( .A(u_alu_lt_x_11_B_21_), .B(n1171), .Q(n3066) );
  CLKIN6 U1019 ( .A(n271), .Q(n2672) );
  NAND33 U1020 ( .A(n2407), .B(n274), .C(n272), .Q(n2408) );
  CLKIN6 U1021 ( .A(n273), .Q(n272) );
  NOR23 U1022 ( .A(n2654), .B(n2485), .Q(n273) );
  AOI222 U1023 ( .A(n2525), .B(n397), .C(n2400), .D(n401), .Q(n2485) );
  AOI222 U1024 ( .A(n849), .B(n2504), .C(n2401), .D(n850), .Q(n274) );
  OAI212 U1025 ( .A(n397), .B(n2503), .C(n275), .Q(n2401) );
  AOI212 U1026 ( .A(n2295), .B(n1041), .C(n2294), .Q(n2503) );
  NAND24 U1027 ( .A(n277), .B(n276), .Q(n2504) );
  NAND24 U1028 ( .A(n2542), .B(n401), .Q(n276) );
  CLKIN6 U1029 ( .A(n278), .Q(n277) );
  NOR24 U1030 ( .A(n401), .B(n2406), .Q(n278) );
  AOI222 U1031 ( .A(n1625), .B(n1167), .C(n1652), .D(n362), .Q(n279) );
  NAND24 U1032 ( .A(n397), .B(n1164), .Q(n280) );
  INV6 U1033 ( .A(n526), .Q(n455) );
  NAND28 U1034 ( .A(n769), .B(n1097), .Q(n526) );
  BUF15 U1035 ( .A(n526), .Q(n281) );
  NAND24 U1036 ( .A(n283), .B(n282), .Q(n770) );
  XNR22 U1037 ( .A(n133), .B(n792), .Q(n282) );
  NAND33 U1038 ( .A(n286), .B(n284), .C(n285), .Q(n283) );
  NAND24 U1039 ( .A(n1292), .B(n289), .Q(compare_i_data_rt[16]) );
  INV6 U1040 ( .A(n792), .Q(n2363) );
  NOR22 U1041 ( .A(n2870), .B(n3011), .Q(n1064) );
  NOR23 U1042 ( .A(n1162), .B(n291), .Q(n3011) );
  NAND28 U1043 ( .A(n3186), .B(n138), .Q(n2828) );
  XOR22 U1044 ( .A(n2636), .B(n3182), .Q(n501) );
  NAND24 U1045 ( .A(n548), .B(n1403), .Q(n3182) );
  CLKIN6 U1046 ( .A(n292), .Q(n1157) );
  CLKIN6 U1047 ( .A(n293), .Q(n1438) );
  NAND24 U1048 ( .A(n1157), .B(i_data_FWmemout[25]), .Q(n293) );
  NAND22 U1049 ( .A(n928), .B(n295), .Q(n294) );
  NAND28 U1050 ( .A(n3089), .B(n3088), .Q(n928) );
  NOR24 U1051 ( .A(n1156), .B(n2954), .Q(n2971) );
  NAND31 U1052 ( .A(n2956), .B(n2971), .C(n2955), .Q(n960) );
  NOR23 U1053 ( .A(n1970), .B(n1971), .Q(n300) );
  NAND24 U1054 ( .A(n299), .B(n296), .Q(alu_o_data_AluRes[8]) );
  NOR24 U1055 ( .A(n298), .B(n297), .Q(n296) );
  OAI212 U1056 ( .A(n1969), .B(n1156), .C(n304), .Q(n298) );
  NOR24 U1057 ( .A(n301), .B(n300), .Q(n299) );
  OAI312 U1058 ( .A(n400), .B(n303), .C(n1976), .D(n302), .Q(n301) );
  AOI212 U1059 ( .A(n1165), .B(n1910), .C(n1909), .Q(n1976) );
  NAND22 U1060 ( .A(n306), .B(n1168), .Q(n2020) );
  NOR23 U1061 ( .A(n1170), .B(n405), .Q(n306) );
  NAND24 U1062 ( .A(n310), .B(n309), .Q(n1647) );
  AOI312 U1063 ( .A(n938), .B(n1167), .C(n615), .D(n930), .Q(n309) );
  INV15 U1064 ( .A(n314), .Q(n313) );
  NAND24 U1065 ( .A(n313), .B(n525), .Q(n312) );
  OAI222 U1066 ( .A(n347), .B(n1316), .C(n351), .D(n1317), .Q(n314) );
  NAND24 U1067 ( .A(alu_i_data_B[13]), .B(n1171), .Q(n809) );
  NOR24 U1068 ( .A(n1516), .B(n315), .Q(alu_i_data_B[13]) );
  NOR33 U1069 ( .A(n1515), .B(n316), .C(n786), .Q(n315) );
  OAI212 U1070 ( .A(n2647), .B(n396), .C(n2526), .Q(n317) );
  NAND22 U1071 ( .A(n317), .B(n1874), .Q(n2537) );
  OAI222 U1072 ( .A(n351), .B(n1227), .C(n220), .D(n1226), .Q(n333) );
  CLKIN10 U1073 ( .A(i_con_Efamux[0]), .Q(n411) );
  NOR24 U1074 ( .A(n401), .B(n2875), .Q(n2718) );
  NOR33 U1075 ( .A(n320), .B(n2717), .C(n318), .Q(n2875) );
  OAI212 U1076 ( .A(n2943), .B(n3104), .C(n319), .Q(n318) );
  NOR24 U1077 ( .A(n1066), .B(n1067), .Q(n3104) );
  NOR24 U1078 ( .A(n1167), .B(n2716), .Q(n320) );
  NAND33 U1079 ( .A(n2898), .B(n1043), .C(n321), .Q(n3070) );
  AOI222 U1080 ( .A(u_alu_lt_x_11_B_1_), .B(n322), .C(n3009), .D(n3067), .Q(
        n321) );
  NAND22 U1081 ( .A(n366), .B(n139), .Q(n2131) );
  NAND32 U1082 ( .A(n541), .B(n1246), .C(n989), .Q(n366) );
  NAND26 U1083 ( .A(compare_i_data_rt[8]), .B(n139), .Q(n2147) );
  OAI211 U1084 ( .A(n1172), .B(n323), .C(n1039), .Q(n631) );
  NAND28 U1085 ( .A(n324), .B(n494), .Q(n1111) );
  NOR24 U1086 ( .A(n270), .B(n354), .Q(n324) );
  NAND31 U1087 ( .A(n494), .B(n324), .C(i_data_FMalures[4]), .Q(n798) );
  CLKIN6 U1088 ( .A(n387), .Q(n2763) );
  NAND22 U1089 ( .A(n325), .B(n682), .Q(n553) );
  NOR23 U1090 ( .A(n326), .B(n3186), .Q(n325) );
  NAND28 U1091 ( .A(n328), .B(n327), .Q(n3186) );
  INV6 U1092 ( .A(n636), .Q(n326) );
  NOR23 U1093 ( .A(n1444), .B(n484), .Q(n636) );
  NOR33 U1094 ( .A(n1348), .B(n1054), .C(n1350), .Q(n328) );
  CLKIN6 U1095 ( .A(n1604), .Q(n1628) );
  NAND24 U1096 ( .A(n1597), .B(n1596), .Q(n1604) );
  NAND33 U1097 ( .A(n1597), .B(n1596), .C(n1634), .Q(n1631) );
  BUF8 U1098 ( .A(n1637), .Q(n330) );
  NAND28 U1099 ( .A(n331), .B(n1049), .Q(n1637) );
  NOR24 U1100 ( .A(n1588), .B(n1592), .Q(n331) );
  NAND24 U1101 ( .A(n1637), .B(n200), .Q(n332) );
  CLKIN6 U1102 ( .A(n333), .Q(n335) );
  INV15 U1103 ( .A(n334), .Q(n403) );
  XNR22 U1104 ( .A(n3193), .B(n403), .Q(n773) );
  IMUX21 U1105 ( .A(n425), .B(n1154), .S(n336), .Q(n2274) );
  INV15 U1106 ( .A(n337), .Q(n338) );
  CLKIN6 U1107 ( .A(n455), .Q(n337) );
  NOR24 U1108 ( .A(n341), .B(n339), .Q(n525) );
  NAND22 U1109 ( .A(n143), .B(i_data_FMmemout[18]), .Q(n340) );
  CLKIN6 U1110 ( .A(n342), .Q(n341) );
  NAND24 U1111 ( .A(n343), .B(i_data_rs[18]), .Q(n342) );
  NAND24 U1112 ( .A(n1498), .B(n344), .Q(n1124) );
  NAND24 U1113 ( .A(n596), .B(n1257), .Q(n345) );
  OAI212 U1114 ( .A(n1159), .B(n1262), .C(n1258), .Q(n346) );
  NAND24 U1115 ( .A(n348), .B(i_data_FWmemout[29]), .Q(n608) );
  CLKIN6 U1116 ( .A(n220), .Q(n348) );
  NAND24 U1117 ( .A(n343), .B(i_data_rs[29]), .Q(n1418) );
  NAND23 U1118 ( .A(n463), .B(n2998), .Q(n1084) );
  NOR22 U1119 ( .A(n3023), .B(n2654), .Q(n2990) );
  NOR24 U1120 ( .A(n2197), .B(n2193), .Q(n2194) );
  INV6 U1121 ( .A(n2194), .Q(n1047) );
  NOR22 U1122 ( .A(n1023), .B(n1021), .Q(n3073) );
  BUF8 U1123 ( .A(i_con_Efamux[0]), .Q(n494) );
  NOR23 U1124 ( .A(n1039), .B(n438), .Q(n2425) );
  NOR32 U1125 ( .A(n1735), .B(n1736), .C(n364), .Q(n1738) );
  INV6 U1126 ( .A(n1362), .Q(n1735) );
  NAND34 U1127 ( .A(n3156), .B(n3155), .C(n400), .Q(n3157) );
  NOR22 U1128 ( .A(n904), .B(n900), .Q(n899) );
  INV3 U1129 ( .A(n2189), .Q(n2166) );
  IMUX21 U1130 ( .A(n2305), .B(n2304), .S(n2303), .Q(n2306) );
  OAI212 U1131 ( .A(n2362), .B(n2302), .C(n2358), .Q(n2303) );
  NAND26 U1132 ( .A(n793), .B(n794), .Q(n1757) );
  INV6 U1133 ( .A(n1538), .Q(n794) );
  NAND24 U1134 ( .A(n684), .B(n681), .Q(n1351) );
  INV12 U1135 ( .A(n350), .Q(n353) );
  OAI212 U1136 ( .A(n1280), .B(n1159), .C(n1175), .Q(n1176) );
  NAND24 U1137 ( .A(compare_i_data_rt[31]), .B(n391), .Q(n617) );
  AOI221 U1138 ( .A(n3165), .B(n400), .C(n3120), .D(n1163), .Q(n3123) );
  NAND24 U1139 ( .A(n338), .B(i_data_FWmemout[14]), .Q(n1105) );
  NOR24 U1140 ( .A(n516), .B(n1116), .Q(n515) );
  NOR24 U1141 ( .A(n2677), .B(n401), .Q(n613) );
  NAND26 U1142 ( .A(n990), .B(n2853), .Q(n2860) );
  NAND28 U1143 ( .A(n2830), .B(n2829), .Q(n2856) );
  INV15 U1144 ( .A(n655), .Q(n1161) );
  NOR24 U1145 ( .A(n270), .B(n411), .Q(n585) );
  NOR24 U1146 ( .A(n397), .B(n2176), .Q(n506) );
  NOR24 U1147 ( .A(n394), .B(n2058), .Q(n2059) );
  INV3 U1148 ( .A(n904), .Q(n902) );
  NOR33 U1149 ( .A(n1299), .B(n1298), .C(n1297), .Q(n800) );
  NAND28 U1150 ( .A(n3004), .B(n295), .Q(n3131) );
  NAND24 U1151 ( .A(n796), .B(n3010), .Q(n795) );
  NAND24 U1152 ( .A(n1442), .B(n1441), .Q(n1443) );
  XNR22 U1153 ( .A(u_alu_lt_x_11_A_3_), .B(compare_i_data_rt[3]), .Q(n826) );
  NAND22 U1154 ( .A(n876), .B(n805), .Q(n804) );
  NOR32 U1155 ( .A(n704), .B(n1436), .C(n697), .Q(n699) );
  NAND24 U1156 ( .A(n1435), .B(n1434), .Q(n1436) );
  NOR33 U1157 ( .A(n1213), .B(n1212), .C(n1211), .Q(n1215) );
  NAND33 U1158 ( .A(n696), .B(n1183), .C(n695), .Q(n565) );
  NAND34 U1159 ( .A(n2941), .B(n963), .C(n962), .Q(n961) );
  NOR32 U1160 ( .A(n3074), .B(n2938), .C(n2937), .Q(n2939) );
  NOR22 U1161 ( .A(n1328), .B(n281), .Q(n2471) );
  NOR22 U1162 ( .A(n1261), .B(n281), .Q(n1259) );
  CLKIN4 U1163 ( .A(n1259), .Q(n596) );
  AOI212 U1164 ( .A(n2913), .B(n2912), .C(n2911), .Q(n2920) );
  NOR23 U1165 ( .A(n7), .B(n1114), .Q(n1113) );
  OAI222 U1166 ( .A(n2675), .B(n362), .C(n1041), .D(n2488), .Q(n2590) );
  NOR24 U1167 ( .A(n890), .B(n888), .Q(n1089) );
  NAND33 U1168 ( .A(n2713), .B(n2712), .C(n2711), .Q(alu_o_data_AluRes[21]) );
  AOI212 U1169 ( .A(n2698), .B(n2697), .C(n2696), .Q(n2712) );
  INV12 U1170 ( .A(n1141), .Q(n1142) );
  NAND24 U1171 ( .A(n670), .B(n669), .Q(compare_i_data_rt[26]) );
  INV6 U1172 ( .A(n1200), .Q(n669) );
  AOI212 U1173 ( .A(n2737), .B(n2736), .C(n1163), .Q(n2706) );
  INV8 U1174 ( .A(alu_i_data_B[13]), .Q(n3068) );
  NAND22 U1175 ( .A(n3152), .B(n401), .Q(n3153) );
  NOR22 U1176 ( .A(n1232), .B(n281), .Q(n1529) );
  AOI212 U1177 ( .A(u_alu_lt_x_11_n110), .B(u_alu_lt_x_11_n56), .C(
        u_alu_lt_x_11_n57), .Q(u_alu_lt_x_11_n55) );
  NOR23 U1178 ( .A(u_alu_lt_x_11_n80), .B(u_alu_lt_x_11_n58), .Q(
        u_alu_lt_x_11_n56) );
  NOR24 U1179 ( .A(n704), .B(n701), .Q(n700) );
  INV6 U1180 ( .A(n1048), .Q(n769) );
  NAND34 U1181 ( .A(n720), .B(n1014), .C(n1531), .Q(n1013) );
  NOR23 U1182 ( .A(n916), .B(n3017), .Q(n919) );
  NOR23 U1183 ( .A(n2471), .B(n1500), .Q(n2462) );
  AOI212 U1184 ( .A(n2321), .B(n2240), .C(n2239), .Q(n2285) );
  NAND28 U1185 ( .A(n2157), .B(n430), .Q(n2289) );
  NAND24 U1186 ( .A(n1433), .B(n1432), .Q(n979) );
  NAND33 U1187 ( .A(n2551), .B(n2550), .C(n2549), .Q(alu_o_data_AluRes[18]) );
  NOR21 U1188 ( .A(n979), .B(n1142), .Q(n3003) );
  NOR22 U1189 ( .A(n1380), .B(n351), .Q(n1381) );
  NAND24 U1190 ( .A(n1105), .B(n1106), .Q(n1511) );
  XNR22 U1191 ( .A(n1019), .B(n500), .Q(n499) );
  NAND34 U1192 ( .A(n547), .B(n546), .C(n1425), .Q(n500) );
  NOR23 U1193 ( .A(n406), .B(n471), .Q(n2073) );
  OAI212 U1194 ( .A(n406), .B(n471), .C(n2433), .Q(n2435) );
  OAI212 U1195 ( .A(n1279), .B(n941), .C(n1173), .Q(n1177) );
  NOR24 U1196 ( .A(n364), .B(n941), .Q(n1523) );
  AOI220 U1197 ( .A(n1136), .B(i_data_FMmemout[16]), .C(n338), .D(
        i_data_FWmemout[16]), .Q(n1292) );
  AOI212 U1198 ( .A(n1587), .B(n1586), .C(n1585), .Q(n1601) );
  AOI212 U1199 ( .A(n1161), .B(n1495), .C(n1162), .Q(n2632) );
  OAI212 U1200 ( .A(n2838), .B(n2790), .C(n2754), .Q(n2735) );
  NAND22 U1201 ( .A(n632), .B(n1524), .Q(n1610) );
  NOR22 U1202 ( .A(n436), .B(n2905), .Q(n2030) );
  IMUX20 U1203 ( .A(n425), .B(n1154), .S(n358), .Q(n1892) );
  INV6 U1204 ( .A(n1453), .Q(n694) );
  NAND24 U1205 ( .A(n1452), .B(n1451), .Q(n1453) );
  INV6 U1206 ( .A(n1182), .Q(n695) );
  OAI222 U1207 ( .A(n1771), .B(n3178), .C(n1812), .D(n2654), .Q(n1772) );
  NAND24 U1208 ( .A(i_data_immext[1]), .B(n365), .Q(n1549) );
  NAND24 U1209 ( .A(n343), .B(i_data_rs[24]), .Q(n1445) );
  AOI212 U1210 ( .A(n1897), .B(n1896), .C(n1895), .Q(n1898) );
  NOR22 U1211 ( .A(n1326), .B(n352), .Q(n1470) );
  NAND24 U1212 ( .A(n2432), .B(n423), .Q(n1115) );
  NOR24 U1213 ( .A(n200), .B(n1604), .Q(n1639) );
  NOR23 U1214 ( .A(n1595), .B(n1594), .Q(n1596) );
  OAI212 U1215 ( .A(n2068), .B(n2065), .C(n2344), .Q(n2066) );
  CLKIN4 U1216 ( .A(n1095), .Q(n2371) );
  OAI210 U1217 ( .A(n1170), .B(u_alu_lt_x_11_B_15_), .C(n1902), .Q(n1903) );
  NOR22 U1218 ( .A(n1349), .B(n220), .Q(n1444) );
  OAI212 U1219 ( .A(n2374), .B(n406), .C(n2373), .Q(n621) );
  NAND24 U1220 ( .A(n1756), .B(n913), .Q(n1960) );
  XNR22 U1221 ( .A(n3143), .B(n3142), .Q(n3176) );
  NOR24 U1222 ( .A(n364), .B(n495), .Q(n2127) );
  NAND33 U1223 ( .A(n1900), .B(n1899), .C(n1898), .Q(alu_o_data_AluRes[7]) );
  OAI212 U1224 ( .A(n1379), .B(n941), .C(n1192), .Q(n1195) );
  NAND24 U1225 ( .A(n826), .B(n832), .Q(n838) );
  NAND33 U1226 ( .A(n2512), .B(n2511), .C(n2510), .Q(alu_o_data_AluRes[17]) );
  NOR32 U1227 ( .A(n2499), .B(n2498), .C(n2497), .Q(n2511) );
  AOI212 U1228 ( .A(n2958), .B(n2482), .C(n2481), .Q(n2512) );
  NOR24 U1229 ( .A(n417), .B(n973), .Q(n2229) );
  NAND24 U1230 ( .A(n1421), .B(n1420), .Q(n1422) );
  NAND24 U1231 ( .A(n3134), .B(n921), .Q(n3140) );
  AOI212 U1232 ( .A(n3133), .B(u_alu_lt_x_11_n8), .C(u_alu_lt_x_11_n7), .Q(
        n3134) );
  NAND28 U1233 ( .A(n2172), .B(n377), .Q(n680) );
  NOR22 U1234 ( .A(n1282), .B(n352), .Q(n1283) );
  INV8 U1235 ( .A(n3009), .Q(n405) );
  AOI212 U1236 ( .A(u_alu_DP_OP_84J3_125_2615_n136), .B(n2940), .C(n2939), .Q(
        n2941) );
  NOR22 U1237 ( .A(n1124), .B(n1125), .Q(n971) );
  NAND33 U1238 ( .A(n2048), .B(n2047), .C(n2046), .Q(alu_o_data_AluRes[10]) );
  NOR22 U1239 ( .A(n1758), .B(u_alu_lt_x_11_A_2_), .Q(n2411) );
  IMUX21 U1240 ( .A(n1630), .B(n1629), .S(u_alu_lt_x_11_A_0_), .Q(n1645) );
  NAND24 U1241 ( .A(n1027), .B(n2968), .Q(n2972) );
  NAND24 U1242 ( .A(n877), .B(n2853), .Q(n3089) );
  INV12 U1243 ( .A(i_con_Efbmux[0]), .Q(n710) );
  NOR24 U1244 ( .A(n508), .B(n507), .Q(n851) );
  INV3 U1245 ( .A(n523), .Q(n497) );
  NOR32 U1246 ( .A(n1588), .B(n1598), .C(n1601), .Q(n1589) );
  NAND23 U1247 ( .A(n418), .B(n1741), .Q(n1101) );
  NAND28 U1248 ( .A(n2063), .B(n453), .Q(n471) );
  NAND24 U1249 ( .A(n343), .B(i_data_rs[17]), .Q(n1469) );
  AOI212 U1250 ( .A(n2766), .B(u_alu_lt_x_11_n44), .C(u_alu_lt_x_11_n43), .Q(
        n2788) );
  NOR24 U1251 ( .A(n2634), .B(n2633), .Q(n2734) );
  AOI212 U1252 ( .A(n2731), .B(n1155), .C(n2730), .Q(n2762) );
  NOR22 U1253 ( .A(n1170), .B(n1946), .Q(n2308) );
  NOR23 U1254 ( .A(n1233), .B(n1159), .Q(n490) );
  NAND28 U1255 ( .A(n2828), .B(n377), .Q(u_alu_DP_OP_84J3_125_2615_n134) );
  NOR22 U1256 ( .A(n1170), .B(n2849), .Q(n2500) );
  INV12 U1257 ( .A(u_alu_DP_OP_84J3_125_2615_n134), .Q(n2849) );
  NOR22 U1258 ( .A(n2057), .B(n397), .Q(n1991) );
  OAI212 U1259 ( .A(n1142), .B(n356), .C(n3012), .Q(n3013) );
  NOR24 U1260 ( .A(n417), .B(u_alu_lt_x_11_B_13_), .Q(u_alu_lt_x_11_n90) );
  NOR23 U1261 ( .A(n408), .B(n446), .Q(u_alu_lt_x_11_n94) );
  INV6 U1262 ( .A(n2073), .Q(u_alu_lt_x_11_n100) );
  NOR22 U1263 ( .A(n875), .B(u_alu_lt_x_11_B_1_), .Q(n2413) );
  NAND24 U1264 ( .A(n387), .B(n442), .Q(u_alu_lt_x_11_n40) );
  NAND28 U1265 ( .A(n421), .B(n1077), .Q(n2827) );
  INV6 U1266 ( .A(n658), .Q(n2959) );
  CLKBU12 U1267 ( .A(n399), .Q(n362) );
  NAND24 U1268 ( .A(n2300), .B(n475), .Q(n2077) );
  NOR22 U1269 ( .A(n1207), .B(n220), .Q(n1213) );
  NAND22 U1270 ( .A(n3165), .B(n850), .Q(n3166) );
  OAI212 U1271 ( .A(n2882), .B(n203), .C(n2881), .Q(n2883) );
  INV3 U1272 ( .A(n2559), .Q(n2561) );
  NOR31 U1273 ( .A(n895), .B(n896), .C(n838), .Q(n1091) );
  INV3 U1274 ( .A(n2527), .Q(n2533) );
  NAND33 U1275 ( .A(n2461), .B(n2460), .C(n2459), .Q(alu_o_data_AluRes[16]) );
  AOI212 U1276 ( .A(n2958), .B(n2448), .C(n2447), .Q(n2460) );
  AOI212 U1277 ( .A(n3027), .B(n3026), .C(n410), .Q(n3107) );
  AOI211 U1278 ( .A(n1170), .B(u_alu_lt_x_11_B_14_), .C(n3105), .Q(n3106) );
  NOR23 U1279 ( .A(n2869), .B(n2868), .Q(n2397) );
  NOR22 U1280 ( .A(n2425), .B(n2202), .Q(n1996) );
  CLKBU12 U1281 ( .A(i_con_Ealusrc), .Q(n1172) );
  INV15 U1282 ( .A(n363), .Q(n364) );
  INV6 U1283 ( .A(n1469), .Q(n2467) );
  AOI212 U1284 ( .A(n2715), .B(n2714), .C(n2932), .Q(n2717) );
  NAND24 U1285 ( .A(n2410), .B(n2409), .Q(n2421) );
  NAND33 U1286 ( .A(n1917), .B(n611), .C(n1919), .Q(n2410) );
  INV3 U1287 ( .A(n1283), .Q(n468) );
  INV6 U1288 ( .A(n1439), .Q(n704) );
  CLKIN4 U1289 ( .A(n1827), .Q(n1832) );
  NOR24 U1290 ( .A(n1278), .B(n723), .Q(n848) );
  OAI212 U1291 ( .A(n3074), .B(n2974), .C(n2996), .Q(n465) );
  NOR24 U1292 ( .A(n588), .B(n587), .Q(n2974) );
  NAND24 U1293 ( .A(n1052), .B(n1051), .Q(n3017) );
  NAND33 U1294 ( .A(n1560), .B(i_data_immext[1]), .C(n1583), .Q(n1571) );
  OAI212 U1295 ( .A(n410), .B(n1622), .C(n1621), .Q(n1625) );
  XOR22 U1296 ( .A(n3185), .B(n366), .Q(n871) );
  NAND26 U1297 ( .A(n1179), .B(n1178), .Q(compare_i_data_rt[31]) );
  NOR23 U1298 ( .A(n1177), .B(n1176), .Q(n1179) );
  AOI2112 U1299 ( .A(n2631), .B(n378), .C(n1030), .D(n2655), .Q(n1029) );
  OAI212 U1300 ( .A(n400), .B(n2617), .C(n2616), .Q(n2631) );
  OAI212 U1301 ( .A(n2654), .B(n2653), .C(n2652), .Q(n2655) );
  AOI212 U1302 ( .A(n849), .B(n2401), .C(n2301), .Q(n2318) );
  NOR24 U1303 ( .A(n2329), .B(n2335), .Q(n2301) );
  AOI212 U1304 ( .A(n3025), .B(n3024), .C(n410), .Q(n2927) );
  OAI212 U1305 ( .A(n1504), .B(n941), .C(n1503), .Q(n1508) );
  INV6 U1306 ( .A(n1550), .Q(n1552) );
  NAND33 U1307 ( .A(n382), .B(i_data_rt[1]), .C(n391), .Q(n1550) );
  XOR22 U1308 ( .A(n483), .B(compare_i_data_rt[10]), .Q(n872) );
  NOR22 U1309 ( .A(n1379), .B(n220), .Q(n1382) );
  NOR23 U1310 ( .A(n1168), .B(n2397), .Q(n2643) );
  NAND22 U1311 ( .A(n1050), .B(n3132), .Q(n3090) );
  NAND26 U1312 ( .A(n1044), .B(n943), .Q(n1061) );
  INV6 U1313 ( .A(n3177), .Q(n943) );
  NOR22 U1314 ( .A(n2436), .B(n2011), .Q(n2074) );
  NOR22 U1315 ( .A(n1922), .B(n1921), .Q(n2412) );
  NOR23 U1316 ( .A(n1687), .B(n1686), .Q(n2395) );
  NOR22 U1317 ( .A(n2223), .B(n2222), .Q(n2224) );
  OAI212 U1318 ( .A(n362), .B(n2600), .C(n2312), .Q(n2489) );
  AOI212 U1319 ( .A(n3035), .B(n397), .C(n3034), .Q(n3062) );
  NAND28 U1320 ( .A(n3130), .B(u_alu_lt_x_11_n8), .Q(n3135) );
  NAND26 U1321 ( .A(n1044), .B(n404), .Q(n2784) );
  NAND23 U1322 ( .A(n1639), .B(n1638), .Q(n470) );
  NOR23 U1323 ( .A(n1638), .B(n330), .Q(n2450) );
  AOI221 U1324 ( .A(n1167), .B(n3151), .C(n3150), .D(n362), .Q(n3154) );
  NAND24 U1325 ( .A(n1147), .B(i_con_Ealuop[1]), .Q(n1585) );
  CLKIN4 U1326 ( .A(i_con_Ealuop[0]), .Q(n1147) );
  NAND33 U1327 ( .A(n2920), .B(n660), .C(n656), .Q(alu_o_data_AluRes[25]) );
  NAND33 U1328 ( .A(n2226), .B(n2225), .C(n2224), .Q(n3194) );
  AOI211 U1329 ( .A(n2307), .B(n2185), .C(n2184), .Q(n2226) );
  OAI212 U1330 ( .A(n2723), .B(n2820), .C(n2691), .Q(n2670) );
  NAND33 U1331 ( .A(n696), .B(n695), .C(n1183), .Q(compare_i_data_rt[25]) );
  NOR33 U1332 ( .A(n2556), .B(n2557), .C(n2558), .Q(n2635) );
  NAND33 U1333 ( .A(n2285), .B(n2284), .C(n2283), .Q(n3195) );
  AOI212 U1334 ( .A(n2307), .B(n2263), .C(n2262), .Q(n2284) );
  NOR23 U1335 ( .A(n1195), .B(n1194), .Q(n1197) );
  OAI212 U1336 ( .A(i_data_immext[2]), .B(i_data_immext[0]), .C(n1561), .Q(
        n1562) );
  NOR22 U1337 ( .A(n1221), .B(n220), .Q(n1224) );
  NOR22 U1338 ( .A(n1294), .B(n220), .Q(n1299) );
  AOI212 U1339 ( .A(i_data_FMmemout[23]), .B(n1136), .C(n1330), .Q(n1407) );
  NOR23 U1340 ( .A(n2436), .B(n2434), .Q(n746) );
  AOI222 U1341 ( .A(n2541), .B(n362), .C(n2257), .D(n1167), .Q(n2406) );
  AOI222 U1342 ( .A(n1563), .B(n1562), .C(n717), .D(n716), .Q(n715) );
  OAI212 U1343 ( .A(n351), .B(n1301), .C(n1303), .Q(n761) );
  OAI212 U1344 ( .A(n1508), .B(n1507), .C(n391), .Q(n825) );
  INV15 U1345 ( .A(n952), .Q(n2698) );
  NAND28 U1346 ( .A(n421), .B(n404), .Q(n952) );
  NAND24 U1347 ( .A(n685), .B(n689), .Q(n686) );
  NOR24 U1348 ( .A(n863), .B(n687), .Q(n685) );
  AOI212 U1349 ( .A(n2988), .B(n2987), .C(n397), .Q(n2989) );
  NOR24 U1350 ( .A(n3103), .B(n3102), .Q(n3156) );
  NOR22 U1351 ( .A(n465), .B(n464), .Q(n463) );
  OAI212 U1352 ( .A(n1305), .B(n1159), .C(n1229), .Q(n482) );
  OAI212 U1353 ( .A(n364), .B(n1624), .C(n1623), .Q(n2360) );
  NAND33 U1354 ( .A(n411), .B(n604), .C(n270), .Q(n1388) );
  NOR24 U1355 ( .A(n896), .B(n894), .Q(n891) );
  OAI212 U1356 ( .A(n2363), .B(n2358), .C(n2357), .Q(n2342) );
  NAND33 U1357 ( .A(n2339), .B(n2338), .C(n2337), .Q(n3196) );
  NAND33 U1358 ( .A(n2687), .B(n2686), .C(n2685), .Q(n2688) );
  NAND33 U1359 ( .A(n2684), .B(n1155), .C(n400), .Q(n2685) );
  NOR22 U1360 ( .A(n138), .B(n385), .Q(n1522) );
  NAND33 U1361 ( .A(n383), .B(n139), .C(i_data_rt[11]), .Q(n870) );
  NOR22 U1362 ( .A(n139), .B(i_data_immext[0]), .Q(n2396) );
  INV3 U1363 ( .A(n2198), .Q(n799) );
  NOR24 U1364 ( .A(n394), .B(n2862), .Q(n532) );
  NOR24 U1365 ( .A(n394), .B(n2488), .Q(n2179) );
  INV8 U1366 ( .A(n1167), .Q(n394) );
  NOR23 U1367 ( .A(n2094), .B(n1791), .Q(n1792) );
  NAND22 U1368 ( .A(compare_i_data_rt[10]), .B(n391), .Q(n2138) );
  INV6 U1369 ( .A(n1070), .Q(u_alu_DP_OP_84J3_125_2615_n145) );
  OAI212 U1370 ( .A(n3100), .B(n3099), .C(n3098), .Q(n3103) );
  NAND33 U1371 ( .A(n1038), .B(n753), .C(n1036), .Q(n1035) );
  INV6 U1372 ( .A(u_alu_DP_OP_83J3_124_3384_n154), .Q(n432) );
  NAND24 U1373 ( .A(u_alu_lt_x_11_B_14_), .B(n1171), .Q(n1617) );
  INV6 U1374 ( .A(n367), .Q(n369) );
  NAND26 U1375 ( .A(n1117), .B(n515), .Q(n2954) );
  NAND33 U1376 ( .A(n2216), .B(n2215), .C(n2214), .Q(n2223) );
  NOR23 U1377 ( .A(n3075), .B(n3074), .Q(n645) );
  NOR22 U1378 ( .A(n416), .B(n2345), .Q(n2346) );
  NOR23 U1379 ( .A(n2153), .B(n631), .Q(n2345) );
  NAND24 U1380 ( .A(n1136), .B(i_data_FMmemout[13]), .Q(n2190) );
  NAND24 U1381 ( .A(n1035), .B(n1037), .Q(n1758) );
  NAND22 U1382 ( .A(n2590), .B(n401), .Q(n616) );
  NAND24 U1383 ( .A(n676), .B(n3082), .Q(n3129) );
  INV8 U1384 ( .A(n3080), .Q(n3082) );
  NAND33 U1385 ( .A(n1033), .B(n1029), .C(n1031), .Q(alu_o_data_AluRes[20]) );
  AOI312 U1386 ( .A(n2626), .B(n404), .C(n421), .D(n1032), .Q(n1031) );
  XNR22 U1387 ( .A(n1335), .B(n3183), .Q(n778) );
  NAND23 U1388 ( .A(n2878), .B(n2877), .Q(n2879) );
  NAND33 U1389 ( .A(n2908), .B(n1155), .C(n1163), .Q(n2878) );
  AOI222 U1390 ( .A(n2094), .B(n386), .C(n2093), .D(n410), .Q(n2398) );
  NOR22 U1391 ( .A(n2414), .B(n1878), .Q(n1882) );
  NOR24 U1392 ( .A(n666), .B(n665), .Q(n664) );
  NOR32 U1393 ( .A(n2026), .B(n2025), .C(n2024), .Q(n2048) );
  NAND24 U1394 ( .A(n1931), .B(n409), .Q(n2390) );
  NAND24 U1395 ( .A(n2475), .B(n2469), .Q(compare_i_data_rs[17]) );
  NOR24 U1396 ( .A(n394), .B(n1829), .Q(n1830) );
  AOI210 U1397 ( .A(n859), .B(n1153), .C(n407), .Q(n858) );
  CLKIN4 U1398 ( .A(n1039), .Q(n407) );
  NAND23 U1399 ( .A(n1135), .B(i_data_FMalures[13]), .Q(n2189) );
  NOR24 U1400 ( .A(n474), .B(n2081), .Q(n2086) );
  NOR24 U1401 ( .A(n477), .B(n2077), .Q(n474) );
  NOR22 U1402 ( .A(n419), .B(n1660), .Q(n1690) );
  INV15 U1403 ( .A(u_alu_lt_x_11_B_0_), .Q(n1660) );
  OAI212 U1404 ( .A(n362), .B(n2740), .C(n2739), .Q(n2864) );
  NAND23 U1405 ( .A(n852), .B(n2419), .Q(n1824) );
  NAND23 U1406 ( .A(n1241), .B(n1240), .Q(n1935) );
  NOR24 U1407 ( .A(n1103), .B(n1239), .Q(n1241) );
  OAI212 U1408 ( .A(n1322), .B(n941), .C(n1321), .Q(n1482) );
  NOR22 U1409 ( .A(n1119), .B(n748), .Q(n1116) );
  INV6 U1410 ( .A(n788), .Q(n2415) );
  NAND22 U1411 ( .A(n1960), .B(n1775), .Q(n788) );
  AOI212 U1412 ( .A(n2719), .B(n401), .C(n2718), .Q(n2780) );
  NAND33 U1413 ( .A(n1600), .B(n1599), .C(i_con_Ealuop[1]), .Q(n1602) );
  OAI222 U1414 ( .A(n2929), .B(n458), .C(n589), .D(n3101), .Q(n588) );
  NOR23 U1415 ( .A(n2368), .B(n2029), .Q(n2065) );
  INV3 U1416 ( .A(n2141), .Q(n2029) );
  XNR22 U1417 ( .A(n783), .B(n1367), .Q(n462) );
  INV6 U1418 ( .A(n2625), .Q(n412) );
  NAND24 U1419 ( .A(u_alu_lt_x_11_B_18_), .B(compare_i_data_rs[18]), .Q(n2625)
         );
  IMUX21 U1420 ( .A(n1834), .B(n1833), .S(n409), .Q(n1835) );
  AOI212 U1421 ( .A(n603), .B(n1591), .C(n820), .Q(n600) );
  AOI212 U1422 ( .A(n1919), .B(n1920), .C(n1069), .Q(n2409) );
  XOR22 U1423 ( .A(compare_i_data_rs[31]), .B(compare_i_data_rt[31]), .Q(n782)
         );
  OAI212 U1424 ( .A(n1380), .B(n1159), .C(n1193), .Q(n1194) );
  AOI212 U1425 ( .A(u_alu_DP_OP_84J3_125_2615_n46), .B(
        u_alu_DP_OP_84J3_125_2615_n91), .C(u_alu_DP_OP_84J3_125_2615_n92), .Q(
        u_alu_DP_OP_84J3_125_2615_n33) );
  NAND22 U1426 ( .A(n807), .B(n1153), .Q(n806) );
  NAND28 U1427 ( .A(n828), .B(n827), .Q(u_alu_lt_x_11_A_3_) );
  NOR33 U1428 ( .A(n1360), .B(n1129), .C(n743), .Q(n827) );
  NOR24 U1429 ( .A(n722), .B(n721), .Q(n720) );
  NAND33 U1430 ( .A(n1532), .B(n1206), .C(n1533), .Q(n721) );
  NOR23 U1431 ( .A(n1956), .B(n1955), .Q(n653) );
  OAI222 U1432 ( .A(n1785), .B(n1156), .C(n1784), .D(n3074), .Q(n1786) );
  NAND24 U1433 ( .A(n892), .B(n891), .Q(n890) );
  NOR22 U1434 ( .A(n838), .B(n897), .Q(n892) );
  NAND24 U1435 ( .A(n452), .B(u_alu_lt_x_11_B_20_), .Q(n2837) );
  INV15 U1436 ( .A(n1172), .Q(n395) );
  NOR22 U1437 ( .A(n364), .B(n2145), .Q(n635) );
  IMUX21 U1438 ( .A(n2803), .B(n2802), .S(u_alu_lt_x_11_A_23_), .Q(n2804) );
  NAND24 U1439 ( .A(n1046), .B(n1047), .Q(n2227) );
  NOR22 U1440 ( .A(n2195), .B(compare_i_data_rs[13]), .Q(n1046) );
  AOI212 U1441 ( .A(n458), .B(n2489), .C(n2314), .Q(n2456) );
  NOR24 U1442 ( .A(n1937), .B(u_alu_lt_x_11_A_5_), .Q(n1933) );
  IMUX21 U1443 ( .A(n1799), .B(n1798), .S(u_alu_lt_x_11_A_5_), .Q(n1800) );
  NAND24 U1444 ( .A(n668), .B(n2834), .Q(n1141) );
  INV6 U1445 ( .A(n1277), .Q(n1006) );
  NAND24 U1446 ( .A(n1465), .B(n1466), .Q(n662) );
  NOR23 U1447 ( .A(n1807), .B(n1808), .Q(n1809) );
  OAI212 U1448 ( .A(n2932), .B(n3104), .C(n2931), .Q(n2934) );
  NOR23 U1449 ( .A(n610), .B(n609), .Q(n780) );
  NOR32 U1450 ( .A(n1455), .B(n1454), .C(n1453), .Q(n1457) );
  AOI212 U1451 ( .A(n2690), .B(n2539), .C(n2538), .Q(n2550) );
  NAND33 U1452 ( .A(n2536), .B(n2537), .C(n2535), .Q(n2538) );
  NAND22 U1453 ( .A(n922), .B(n3044), .Q(n921) );
  NAND26 U1454 ( .A(n1761), .B(n1762), .Q(n2387) );
  AOI212 U1455 ( .A(n1760), .B(n418), .C(n439), .Q(n1761) );
  IMUX21 U1456 ( .A(n413), .B(n376), .S(compare_i_data_rs[29]), .Q(n3060) );
  AOI211 U1457 ( .A(n3064), .B(compare_i_data_rs[29]), .C(n3063), .Q(n3065) );
  INV6 U1458 ( .A(compare_i_data_rs[29]), .Q(n444) );
  NAND26 U1459 ( .A(n1419), .B(n1418), .Q(compare_i_data_rs[29]) );
  AOI212 U1460 ( .A(n757), .B(u_alu_DP_OP_84J3_125_2615_n91), .C(
        u_alu_DP_OP_84J3_125_2615_n92), .Q(u_alu_DP_OP_84J3_125_2615_n90) );
  NAND24 U1461 ( .A(n758), .B(u_alu_DP_OP_84J3_125_2615_n48), .Q(n757) );
  OAI212 U1462 ( .A(u_alu_DP_OP_84J3_125_2615_n40), .B(
        u_alu_DP_OP_84J3_125_2615_n36), .C(u_alu_DP_OP_84J3_125_2615_n37), .Q(
        u_alu_DP_OP_84J3_125_2615_n92) );
  NOR22 U1463 ( .A(n1150), .B(n1131), .Q(n743) );
  NAND22 U1464 ( .A(n2554), .B(n492), .Q(n2555) );
  OAI212 U1465 ( .A(n422), .B(n2900), .C(n3009), .Q(n2901) );
  NOR32 U1466 ( .A(n1417), .B(n1416), .C(n638), .Q(n1419) );
  NOR22 U1467 ( .A(n444), .B(n3054), .Q(u_alu_lt_x_11_n15) );
  OAI222 U1468 ( .A(n3062), .B(n400), .C(n1164), .D(n1025), .Q(n1024) );
  AOI222 U1469 ( .A(n1041), .B(n1990), .C(n1989), .D(n362), .Q(n2057) );
  NAND24 U1470 ( .A(compare_i_data_rt[26]), .B(n391), .Q(n668) );
  NAND23 U1471 ( .A(n1142), .B(n356), .Q(n3008) );
  NAND33 U1472 ( .A(n2762), .B(n2761), .C(n2760), .Q(alu_o_data_AluRes[22]) );
  AOI212 U1473 ( .A(n2958), .B(n2759), .C(n671), .Q(n2760) );
  AOI212 U1474 ( .A(n2913), .B(n2752), .C(n2751), .Q(n2761) );
  NOR32 U1475 ( .A(n2348), .B(n2347), .C(n2346), .Q(n2355) );
  NOR32 U1476 ( .A(n2304), .B(n2303), .C(n667), .Q(n666) );
  NOR23 U1477 ( .A(n1163), .B(n2617), .Q(n2569) );
  AOI222 U1478 ( .A(n2703), .B(n1165), .C(n2568), .D(n397), .Q(n2617) );
  INV12 U1479 ( .A(alu_i_data_B[31]), .Q(n3162) );
  OAI212 U1480 ( .A(u_alu_lt_x_11_B_18_), .B(n425), .C(n1153), .Q(n2529) );
  AOI212 U1481 ( .A(n3093), .B(n3175), .C(n1058), .Q(n1056) );
  NOR24 U1482 ( .A(n3007), .B(n3008), .Q(n982) );
  NAND23 U1483 ( .A(n2108), .B(n2109), .Q(n2110) );
  NOR23 U1484 ( .A(n1577), .B(n1576), .Q(n1593) );
  NOR24 U1485 ( .A(n1957), .B(n653), .Q(n2385) );
  NAND33 U1486 ( .A(n1951), .B(n1950), .C(u_alu_lt_x_11_A_0_), .Q(n1957) );
  NOR22 U1487 ( .A(n2414), .B(n1876), .Q(n1881) );
  NOR22 U1488 ( .A(n544), .B(n1493), .Q(n783) );
  NOR33 U1489 ( .A(n898), .B(n572), .C(n1391), .Q(n524) );
  AOI211 U1490 ( .A(n2326), .B(n2117), .C(n2116), .Q(n2118) );
  NAND23 U1491 ( .A(n1005), .B(n747), .Q(n2326) );
  NOR24 U1492 ( .A(n1310), .B(n770), .Q(n903) );
  NAND22 U1493 ( .A(n1754), .B(n811), .Q(n810) );
  NOR22 U1494 ( .A(n1328), .B(n220), .Q(n1471) );
  NOR24 U1495 ( .A(n1726), .B(n1725), .Q(n1739) );
  NOR23 U1496 ( .A(n1726), .B(n760), .Q(n759) );
  NOR22 U1497 ( .A(n1361), .B(n1158), .Q(n1726) );
  NAND33 U1498 ( .A(n2971), .B(n2972), .C(n2970), .Q(n2973) );
  NOR32 U1499 ( .A(n2885), .B(n2884), .C(n2883), .Q(n2886) );
  AOI2112 U1500 ( .A(n2865), .B(n400), .C(n2800), .D(n2799), .Q(n2806) );
  OAI212 U1501 ( .A(n400), .B(n2798), .C(n2797), .Q(n2799) );
  NOR33 U1502 ( .A(n2343), .B(n2342), .C(n2341), .Q(n1007) );
  NOR22 U1503 ( .A(n2358), .B(n3168), .Q(n2343) );
  NOR33 U1504 ( .A(n2359), .B(n2353), .C(n2340), .Q(n2341) );
  NOR22 U1505 ( .A(n401), .B(n3029), .Q(n587) );
  NOR22 U1506 ( .A(n3003), .B(n3007), .Q(n3004) );
  NOR21 U1507 ( .A(n1682), .B(n1681), .Q(n1683) );
  NAND31 U1508 ( .A(n1680), .B(n1679), .C(n139), .Q(n1682) );
  OAI2112 U1509 ( .A(n2353), .B(n2340), .C(n2290), .D(n2358), .Q(n2291) );
  AOI212 U1510 ( .A(n2707), .B(n1163), .C(n2706), .Q(n2708) );
  OAI222 U1511 ( .A(n2741), .B(n1166), .C(n401), .D(n2615), .Q(n2707) );
  NOR22 U1512 ( .A(n1422), .B(n1423), .Q(n547) );
  NOR24 U1513 ( .A(compare_i_data_rs[29]), .B(n431), .Q(n3080) );
  NOR32 U1514 ( .A(n2282), .B(n2281), .C(n2280), .Q(n2283) );
  NAND33 U1515 ( .A(n2279), .B(n2278), .C(n2277), .Q(n2280) );
  AOI212 U1516 ( .A(n2524), .B(n362), .C(n2523), .Q(n2647) );
  NAND24 U1517 ( .A(n889), .B(n524), .Q(n888) );
  NAND28 U1518 ( .A(n678), .B(n677), .Q(compare_i_data_rs[28]) );
  NOR24 U1519 ( .A(n458), .B(n2102), .Q(n508) );
  OAI222 U1520 ( .A(n2258), .B(n1166), .C(n2102), .D(n401), .Q(n2204) );
  AOI222 U1521 ( .A(n362), .B(n2257), .C(n2021), .D(n1167), .Q(n2102) );
  INV3 U1522 ( .A(n1829), .Q(n1673) );
  NOR22 U1523 ( .A(n242), .B(n372), .Q(n1932) );
  NOR21 U1524 ( .A(n409), .B(n372), .Q(u_alu_lt_x_11_n125) );
  NAND23 U1525 ( .A(u_alu_lt_x_11_B_5_), .B(n1809), .Q(n2417) );
  NAND33 U1526 ( .A(n2962), .B(n2961), .C(n2960), .Q(alu_o_data_AluRes[26]) );
  AOI2112 U1527 ( .A(n2957), .B(n2958), .C(n959), .D(n961), .Q(n2962) );
  NAND33 U1528 ( .A(n3159), .B(n1155), .C(n3157), .Q(n3173) );
  OAI2112 U1529 ( .A(n1165), .B(n3154), .C(n3153), .D(n1163), .Q(n3159) );
  NOR32 U1530 ( .A(n1541), .B(n1542), .C(n1543), .Q(n1619) );
  INV3 U1531 ( .A(n1543), .Q(n1038) );
  NOR23 U1532 ( .A(n462), .B(n782), .Q(n781) );
  NOR24 U1533 ( .A(n534), .B(n532), .Q(n2944) );
  NAND28 U1534 ( .A(n1486), .B(n1485), .Q(n1019) );
  AOI212 U1535 ( .A(n2326), .B(n2422), .C(u_alu_lt_x_11_n94), .Q(n2217) );
  NAND33 U1536 ( .A(n2469), .B(n2465), .C(n2464), .Q(n2466) );
  NAND33 U1537 ( .A(n2315), .B(n1155), .C(n1164), .Q(n2316) );
  NAND24 U1538 ( .A(n1161), .B(i_data_rt[0]), .Q(n574) );
  XNR22 U1539 ( .A(compare_i_data_rt[1]), .B(n3192), .Q(n874) );
  AOI212 U1540 ( .A(n383), .B(n1510), .C(n1162), .Q(n2394) );
  AOI312 U1541 ( .A(n2386), .B(n2387), .C(n2388), .D(n845), .Q(n844) );
  XNR22 U1542 ( .A(n606), .B(compare_i_data_rt[29]), .Q(n610) );
  AOI212 U1543 ( .A(n2958), .B(n2774), .C(n2773), .Q(n2809) );
  INV3 U1544 ( .A(n608), .Q(n1417) );
  NAND24 U1545 ( .A(n847), .B(n846), .Q(n845) );
  OAI212 U1546 ( .A(n1369), .B(n1158), .C(n1189), .Q(n1190) );
  NAND23 U1547 ( .A(n398), .B(i_data_rs[1]), .Q(n1953) );
  NOR22 U1548 ( .A(n364), .B(n1679), .Q(n1551) );
  NAND33 U1549 ( .A(n621), .B(n2375), .C(n2376), .Q(n2377) );
  AOI222 U1550 ( .A(n2252), .B(n2251), .C(n417), .D(n2250), .Q(n2376) );
  OAI210 U1551 ( .A(n3108), .B(n3107), .C(n1167), .Q(n3028) );
  NOR32 U1552 ( .A(n458), .B(n3108), .C(n3107), .Q(n3109) );
  AOI212 U1553 ( .A(n2734), .B(u_alu_lt_x_11_n50), .C(n2733), .Q(n2754) );
  NOR24 U1554 ( .A(n362), .B(n2986), .Q(n537) );
  NOR24 U1555 ( .A(n539), .B(n2777), .Q(n2986) );
  AOI212 U1556 ( .A(n458), .B(n2864), .C(n2863), .Q(n2893) );
  NOR22 U1557 ( .A(n2944), .B(n458), .Q(n2863) );
  NAND33 U1558 ( .A(n2289), .B(n2288), .C(n2287), .Q(n2290) );
  AOI212 U1559 ( .A(n2089), .B(n404), .C(n2088), .Q(n2090) );
  NAND33 U1560 ( .A(n2087), .B(n2086), .C(n2085), .Q(n2088) );
  OAI312 U1561 ( .A(n2956), .B(n2955), .C(n1149), .D(n960), .Q(n959) );
  NAND22 U1562 ( .A(n1065), .B(n1063), .Q(n2925) );
  NOR22 U1563 ( .A(n1511), .B(n1512), .Q(n2243) );
  AOI212 U1564 ( .A(n3071), .B(n397), .C(n2989), .Q(n3023) );
  NAND24 U1565 ( .A(n1020), .B(n2985), .Q(n3071) );
  NOR23 U1566 ( .A(n2843), .B(n2838), .Q(n2853) );
  NAND24 U1567 ( .A(n2837), .B(u_alu_lt_x_11_n50), .Q(n2838) );
  NOR22 U1568 ( .A(n2013), .B(n1140), .Q(n1477) );
  NOR23 U1569 ( .A(u_alu_DP_OP_84J3_125_2615_n36), .B(
        u_alu_DP_OP_84J3_125_2615_n39), .Q(u_alu_DP_OP_84J3_125_2615_n91) );
  NOR22 U1570 ( .A(n356), .B(u_alu_DP_OP_84J3_125_2615_n136), .Q(
        u_alu_DP_OP_84J3_125_2615_n39) );
  NAND42 U1571 ( .A(n1488), .B(n1487), .C(n1110), .D(n864), .Q(n1489) );
  CLKIN4 U1572 ( .A(n2432), .Q(n516) );
  NOR23 U1573 ( .A(n2467), .B(n2466), .Q(n2468) );
  AOI212 U1574 ( .A(n928), .B(n3057), .C(n3056), .Q(n3058) );
  NAND26 U1575 ( .A(n1019), .B(n139), .Q(n2172) );
  OAI2112 U1576 ( .A(n1019), .B(n1162), .C(n678), .D(n672), .Q(n676) );
  NAND24 U1577 ( .A(n405), .B(compare_i_data_rs[25]), .Q(n3014) );
  INV12 U1578 ( .A(compare_i_data_rs[25]), .Q(n414) );
  OAI210 U1579 ( .A(n422), .B(n2995), .C(u_alu_DP_OP_84J3_125_2615_n137), .Q(
        n2996) );
  INV8 U1580 ( .A(u_alu_DP_OP_84J3_125_2615_n137), .Q(n434) );
  NAND24 U1581 ( .A(n1605), .B(n377), .Q(u_alu_DP_OP_84J3_125_2615_n137) );
  NOR24 U1582 ( .A(n1165), .B(n2022), .Q(n507) );
  AOI222 U1583 ( .A(n1167), .B(n1905), .C(n2101), .D(n362), .Q(n2022) );
  NAND24 U1584 ( .A(i_data_immext[4]), .B(n364), .Q(n1940) );
  NOR22 U1585 ( .A(n942), .B(n1088), .Q(n1087) );
  NAND33 U1586 ( .A(n975), .B(n742), .C(n976), .Q(n1088) );
  NAND24 U1587 ( .A(n503), .B(n502), .Q(n896) );
  XNR22 U1588 ( .A(n556), .B(n3180), .Q(n502) );
  NAND28 U1589 ( .A(n762), .B(n519), .Q(u_alu_lt_x_11_A_23_) );
  INV6 U1590 ( .A(n520), .Q(n519) );
  OAI212 U1591 ( .A(n2385), .B(n2384), .C(n2383), .Q(n2388) );
  NOR22 U1592 ( .A(n359), .B(n2835), .Q(n2722) );
  INV8 U1593 ( .A(n1343), .Q(n451) );
  NAND24 U1594 ( .A(n143), .B(i_data_FMmemout[17]), .Q(n2465) );
  MUX26 U1595 ( .A(compare_i_data_rt[0]), .B(i_data_immext[0]), .S(n364), .Q(
        u_alu_lt_x_11_B_0_) );
  INV6 U1596 ( .A(compare_i_data_rs[17]), .Q(n415) );
  OAI212 U1597 ( .A(n662), .B(n830), .C(n1325), .Q(n829) );
  AOI212 U1598 ( .A(n1325), .B(n2592), .C(n2591), .Q(n2597) );
  OAI312 U1599 ( .A(n662), .B(n1325), .C(n830), .D(n829), .Q(n832) );
  NAND24 U1600 ( .A(n766), .B(n975), .Q(n900) );
  XNR22 U1601 ( .A(compare_i_data_rs[13]), .B(compare_i_data_rt[13]), .Q(n766)
         );
  INV8 U1602 ( .A(compare_i_data_rs[21]), .Q(n450) );
  AOI212 U1603 ( .A(n1523), .B(i_data_FWmemout[9]), .C(n1522), .Q(n1524) );
  NAND24 U1604 ( .A(n1008), .B(n1007), .Q(n1010) );
  AOI212 U1605 ( .A(n700), .B(n565), .C(n698), .Q(n705) );
  AOI212 U1606 ( .A(n1245), .B(i_data_FEalures[11]), .C(n542), .Q(n541) );
  NAND24 U1607 ( .A(n543), .B(n595), .Q(n542) );
  AOI212 U1608 ( .A(n2321), .B(n2320), .C(n2319), .Q(n2339) );
  NOR22 U1609 ( .A(n2944), .B(n401), .Q(n2945) );
  INV8 U1610 ( .A(n795), .Q(n295) );
  OAI212 U1611 ( .A(u_alu_DP_OP_84J3_125_2615_n17), .B(
        u_alu_DP_OP_84J3_125_2615_n90), .C(u_alu_DP_OP_84J3_125_2615_n18), .Q(
        u_alu_DP_OP_84J3_125_2615_n73) );
  NOR24 U1612 ( .A(n2425), .B(n2423), .Q(n2111) );
  INV6 U1613 ( .A(u_alu_lt_x_11_n109), .Q(n2423) );
  NAND22 U1614 ( .A(n1946), .B(n357), .Q(n1947) );
  NOR24 U1615 ( .A(n1202), .B(n281), .Q(n1536) );
  NAND33 U1616 ( .A(n521), .B(n1447), .C(n1446), .Q(n1334) );
  NOR24 U1617 ( .A(n590), .B(n415), .Q(n823) );
  NAND24 U1618 ( .A(n981), .B(n2468), .Q(n2854) );
  OAI212 U1619 ( .A(n1162), .B(n139), .C(n831), .Q(n2558) );
  INV6 U1620 ( .A(n545), .Q(n496) );
  NOR24 U1621 ( .A(n1694), .B(n1693), .Q(n1780) );
  INV6 U1622 ( .A(n2416), .Q(n1919) );
  INV6 U1623 ( .A(compare_i_data_rs[20]), .Q(n373) );
  INV12 U1624 ( .A(n373), .Q(n374) );
  INV6 U1625 ( .A(n466), .Q(n1592) );
  AOI212 U1626 ( .A(n1832), .B(n458), .C(n1831), .Q(n1868) );
  NOR22 U1627 ( .A(n1222), .B(n352), .Q(n791) );
  NAND22 U1628 ( .A(n591), .B(n2477), .Q(n981) );
  NAND22 U1629 ( .A(n2478), .B(n2477), .Q(n2479) );
  AOI212 U1630 ( .A(n2765), .B(n2837), .C(n2734), .Q(n2694) );
  NOR24 U1631 ( .A(n397), .B(n2313), .Q(n2314) );
  AOI212 U1632 ( .A(n2180), .B(n362), .C(n2179), .Q(n2313) );
  NAND33 U1633 ( .A(n1925), .B(n611), .C(n2417), .Q(n1926) );
  NAND24 U1634 ( .A(n408), .B(n446), .Q(n2422) );
  CLKBU15 U1635 ( .A(n2360), .Q(n446) );
  OAI212 U1636 ( .A(n3168), .B(n3167), .C(n3166), .Q(n3169) );
  NOR24 U1637 ( .A(n1530), .B(n1875), .Q(alu_i_data_B[7]) );
  INV6 U1638 ( .A(n1045), .Q(n1875) );
  OAI311 U1639 ( .A(n362), .B(n370), .C(n2925), .D(n2873), .Q(n2874) );
  AOI311 U1640 ( .A(n362), .B(n2872), .C(n2871), .D(n1165), .Q(n2873) );
  AOI212 U1641 ( .A(n928), .B(n3141), .C(n3140), .Q(n3142) );
  NAND28 U1642 ( .A(n2574), .B(n377), .Q(u_alu_lt_x_11_B_19_) );
  NAND24 U1643 ( .A(n1325), .B(n391), .Q(n2574) );
  NAND24 U1644 ( .A(n906), .B(n905), .Q(n904) );
  NOR23 U1645 ( .A(n773), .B(n772), .Q(n905) );
  NAND22 U1646 ( .A(n682), .B(n636), .Q(n552) );
  NAND24 U1647 ( .A(n2028), .B(n2371), .Q(n2141) );
  INV6 U1648 ( .A(n1627), .Q(n1060) );
  OAI212 U1649 ( .A(n2127), .B(n2126), .C(n2125), .Q(n2128) );
  INV6 U1650 ( .A(n2126), .Q(n449) );
  NAND33 U1651 ( .A(n1521), .B(n1520), .C(n2132), .Q(n2126) );
  NOR32 U1652 ( .A(n1780), .B(n371), .C(n1143), .Q(n1781) );
  NOR24 U1653 ( .A(n1101), .B(n1740), .Q(n1143) );
  NOR22 U1654 ( .A(n1280), .B(n351), .Q(n1375) );
  NOR24 U1655 ( .A(n2229), .B(n2228), .Q(n2340) );
  NOR24 U1656 ( .A(n2637), .B(n878), .Q(n2832) );
  AOI212 U1657 ( .A(n1924), .B(n357), .C(n2415), .Q(n1925) );
  INV6 U1658 ( .A(n583), .Q(n2150) );
  NOR32 U1659 ( .A(n1462), .B(n1461), .C(n1460), .Q(n1464) );
  INV3 U1660 ( .A(n3132), .Q(n3133) );
  AOI212 U1661 ( .A(n3083), .B(n3082), .C(u_alu_lt_x_11_n15), .Q(n3132) );
  NOR23 U1662 ( .A(n1448), .B(n1334), .Q(n1335) );
  NOR24 U1663 ( .A(n579), .B(n575), .Q(n1107) );
  NOR32 U1664 ( .A(n2121), .B(n2122), .C(n2123), .Q(n2162) );
  NOR42 U1665 ( .A(n1156), .B(n2038), .C(n2037), .D(n2036), .Q(n2039) );
  NOR22 U1666 ( .A(n1371), .B(n351), .Q(n1411) );
  AOI222 U1667 ( .A(n2178), .B(n1168), .C(u_alu_lt_x_11_B_13_), .D(n3067), .Q(
        n2488) );
  NAND33 U1668 ( .A(n2462), .B(n2474), .C(n555), .Q(n3180) );
  NOR24 U1669 ( .A(n619), .B(n2362), .Q(n2375) );
  OAI212 U1670 ( .A(n2875), .B(n397), .C(n2874), .Q(n2908) );
  OAI212 U1671 ( .A(n2856), .B(n2833), .C(n2832), .Q(n877) );
  INV3 U1672 ( .A(n2367), .Q(n950) );
  AOI212 U1673 ( .A(n406), .B(n2374), .C(n2128), .Q(n2367) );
  IMUX20 U1674 ( .A(n2276), .B(n2275), .S(n403), .Q(n2277) );
  BUF15 U1675 ( .A(n2834), .Q(n377) );
  OAI210 U1676 ( .A(n2763), .B(u_alu_lt_x_11_A_23_), .C(n2842), .Q(n2792) );
  INV6 U1677 ( .A(u_alu_lt_x_11_A_23_), .Q(n442) );
  OAI212 U1678 ( .A(n1765), .B(n2384), .C(n2383), .Q(n1766) );
  AOI212 U1679 ( .A(n458), .B(n3031), .C(n3030), .Q(n3075) );
  NAND24 U1680 ( .A(n1587), .B(n1567), .Q(n1574) );
  AOI212 U1681 ( .A(n2021), .B(n362), .C(n1830), .Q(n1906) );
  AOI212 U1682 ( .A(n2975), .B(n362), .C(n2794), .Q(n2891) );
  NOR23 U1683 ( .A(n2943), .B(n2793), .Q(n2794) );
  NAND33 U1684 ( .A(n2810), .B(n1426), .C(n1427), .Q(n1122) );
  NAND24 U1685 ( .A(n977), .B(n3057), .Q(n751) );
  NOR23 U1686 ( .A(n3055), .B(n3131), .Q(n3057) );
  NAND24 U1687 ( .A(n3158), .B(n1163), .Q(n2654) );
  NAND28 U1688 ( .A(n1639), .B(n2450), .Q(n3178) );
  INV15 U1689 ( .A(n381), .Q(n382) );
  NAND22 U1690 ( .A(n2839), .B(n1171), .Q(n1068) );
  NOR22 U1691 ( .A(n1171), .B(n1931), .Q(n1066) );
  NAND43 U1692 ( .A(n903), .B(n1092), .C(n1093), .D(n899), .Q(n1399) );
  NAND28 U1693 ( .A(n605), .B(n1285), .Q(u_alu_lt_x_11_A_0_) );
  NOR23 U1694 ( .A(n3178), .B(n1138), .Q(n2307) );
  BUF15 U1695 ( .A(u_alu_DP_OP_84J3_125_2615_n140), .Q(n384) );
  AOI211 U1696 ( .A(n413), .B(n3116), .C(n422), .Q(n3117) );
  OAI210 U1697 ( .A(n422), .B(n1703), .C(n371), .Q(n1704) );
  NOR22 U1698 ( .A(n1279), .B(n347), .Q(n1376) );
  NOR22 U1699 ( .A(n1248), .B(n220), .Q(n1254) );
  NOR23 U1700 ( .A(n1363), .B(n347), .Q(n1360) );
  NOR22 U1701 ( .A(n1333), .B(n352), .Q(n763) );
  NAND24 U1702 ( .A(n1590), .B(n1589), .Q(n1626) );
  OAI212 U1703 ( .A(n1585), .B(n1578), .C(n1593), .Q(n1590) );
  INV8 U1704 ( .A(n655), .Q(n393) );
  NAND33 U1705 ( .A(n2476), .B(n2478), .C(n2475), .Q(n2517) );
  NOR24 U1706 ( .A(n370), .B(n2925), .Q(n3101) );
  NOR24 U1707 ( .A(n691), .B(n690), .Q(n689) );
  NAND24 U1708 ( .A(n693), .B(n692), .Q(n691) );
  NOR32 U1709 ( .A(n1272), .B(n1271), .C(n1270), .Q(n1274) );
  NOR24 U1710 ( .A(n1551), .B(n1552), .Q(n1954) );
  NAND42 U1711 ( .A(n2133), .B(n1476), .C(n2134), .D(n1139), .Q(n483) );
  NAND26 U1712 ( .A(n1010), .B(n1009), .Q(n1011) );
  NOR22 U1713 ( .A(n2167), .B(n2166), .Q(n2168) );
  NOR32 U1714 ( .A(n1438), .B(n8), .C(n1436), .Q(n1440) );
  INV12 U1715 ( .A(n803), .Q(n416) );
  NAND33 U1716 ( .A(n558), .B(n1469), .C(n557), .Q(n556) );
  INV15 U1717 ( .A(n2665), .Q(n1156) );
  NOR24 U1718 ( .A(n470), .B(n329), .Q(n2665) );
  NAND34 U1719 ( .A(n1225), .B(n789), .C(n1223), .Q(n792) );
  INV6 U1720 ( .A(n2593), .Q(n1741) );
  AOI212 U1721 ( .A(n2639), .B(n2638), .C(n2859), .Q(n2790) );
  INV6 U1722 ( .A(n1626), .Q(n2451) );
  INV15 U1723 ( .A(n1156), .Q(n423) );
  NOR22 U1724 ( .A(n2268), .B(n1156), .Q(n2272) );
  NAND28 U1725 ( .A(n985), .B(n984), .Q(n3044) );
  NAND26 U1726 ( .A(n986), .B(n987), .Q(n984) );
  NOR22 U1727 ( .A(n983), .B(n982), .Q(n985) );
  NOR22 U1728 ( .A(n1332), .B(n220), .Q(n764) );
  NOR24 U1729 ( .A(n2421), .B(n1927), .Q(n2202) );
  NAND33 U1730 ( .A(n2300), .B(n2299), .C(n2325), .Q(n2335) );
  INV15 U1731 ( .A(i_data_immext[8]), .Q(n1167) );
  INV3 U1732 ( .A(n2442), .Q(n2444) );
  NAND34 U1733 ( .A(n862), .B(n1220), .C(n861), .Q(n3197) );
  INV6 U1734 ( .A(n1219), .Q(n861) );
  XOR22 U1735 ( .A(n1775), .B(compare_i_data_rt[4]), .Q(n907) );
  INV12 U1736 ( .A(n625), .Q(n1775) );
  AOI211 U1737 ( .A(n458), .B(n2866), .C(n2865), .Q(n2867) );
  NOR22 U1738 ( .A(n397), .B(n2891), .Q(n2865) );
  NAND24 U1739 ( .A(n489), .B(n487), .Q(n1045) );
  INV12 U1740 ( .A(n3068), .Q(u_alu_lt_x_11_B_13_) );
  NOR24 U1741 ( .A(n1697), .B(n1696), .Q(n2381) );
  NOR24 U1742 ( .A(n467), .B(n1284), .Q(n605) );
  AOI312 U1743 ( .A(n524), .B(n1090), .C(n1091), .D(n1086), .Q(n1085) );
  INV15 U1744 ( .A(n988), .Q(u_alu_lt_x_11_B_18_) );
  NAND26 U1745 ( .A(n511), .B(n510), .Q(n988) );
  NOR23 U1746 ( .A(n763), .B(n764), .Q(n521) );
  NOR24 U1747 ( .A(n980), .B(n1429), .Q(n1433) );
  NOR23 U1748 ( .A(n1430), .B(n1431), .Q(n1432) );
  BUF6 U1749 ( .A(n1169), .Q(n385) );
  CLKIN4 U1750 ( .A(i_data_immext[9]), .Q(n1169) );
  NAND28 U1751 ( .A(n1256), .B(n1255), .Q(compare_i_data_rs[13]) );
  NOR32 U1752 ( .A(n1254), .B(n1253), .C(n1252), .Q(n1256) );
  NAND28 U1753 ( .A(n448), .B(n449), .Q(n2027) );
  OAI2112 U1754 ( .A(n2373), .B(n2141), .C(n430), .D(n950), .Q(n949) );
  NOR22 U1755 ( .A(n2496), .B(n2784), .Q(n2497) );
  AOI312 U1756 ( .A(n1649), .B(n824), .C(n2854), .D(n823), .Q(n2833) );
  NOR23 U1757 ( .A(u_alu_lt_x_11_n94), .B(n2233), .Q(n2112) );
  AOI212 U1758 ( .A(n2430), .B(u_alu_lt_x_11_n94), .C(u_alu_lt_x_11_n90), .Q(
        n748) );
  NOR24 U1759 ( .A(n420), .B(n1815), .Q(n2178) );
  AOI210 U1760 ( .A(n413), .B(n1914), .C(n422), .Q(n1798) );
  INV6 U1761 ( .A(n376), .Q(n1154) );
  AOI212 U1762 ( .A(n378), .B(n2880), .C(n2879), .Q(n2881) );
  OAI222 U1763 ( .A(n2893), .B(n1163), .C(n2867), .D(n400), .Q(n2880) );
  NAND28 U1764 ( .A(n1401), .B(n1400), .Q(o_con_ifbranch) );
  AOI212 U1765 ( .A(n1399), .B(n1398), .C(n1397), .Q(n1400) );
  CLKIN4 U1766 ( .A(n2124), .Q(n2125) );
  NAND33 U1767 ( .A(n2191), .B(n1514), .C(n2190), .Q(n1515) );
  OAI210 U1768 ( .A(n2928), .B(n2927), .C(n1167), .Q(n2645) );
  INV3 U1769 ( .A(n2928), .Q(n2872) );
  NOR22 U1770 ( .A(n386), .B(n1790), .Q(n2928) );
  INV12 U1771 ( .A(n146), .Q(n2948) );
  NOR22 U1772 ( .A(u_alu_lt_x_11_A_3_), .B(n1759), .Q(n2382) );
  NOR23 U1773 ( .A(n875), .B(n2895), .Q(n2384) );
  INV15 U1774 ( .A(n395), .Q(n389) );
  INV6 U1775 ( .A(n389), .Q(n390) );
  NAND24 U1776 ( .A(n559), .B(n1628), .Q(n1151) );
  NAND28 U1777 ( .A(n1062), .B(n1011), .Q(n1044) );
  AOI220 U1778 ( .A(n3067), .B(u_alu_lt_x_11_B_8_), .C(n2868), .D(n410), .Q(
        n1650) );
  NOR24 U1779 ( .A(n406), .B(n2374), .Q(n2369) );
  OAI210 U1780 ( .A(n1924), .B(n425), .C(n1153), .Q(n1891) );
  OAI210 U1781 ( .A(n2027), .B(n425), .C(n1153), .Q(n2015) );
  OAI210 U1782 ( .A(n371), .B(n425), .C(n1153), .Q(n1702) );
  AOI210 U1783 ( .A(n1633), .B(n1153), .C(n1660), .Q(n1644) );
  AOI210 U1784 ( .A(n2080), .B(n1153), .C(n2982), .Q(n2081) );
  AOI210 U1785 ( .A(n1998), .B(n1153), .C(n2905), .Q(n1999) );
  AOI210 U1786 ( .A(n3037), .B(n1153), .C(n435), .Q(n3038) );
  AOI210 U1787 ( .A(n2744), .B(n1153), .C(n1863), .Q(n2745) );
  OAI210 U1788 ( .A(u_alu_lt_x_11_B_13_), .B(n425), .C(n1153), .Q(n2213) );
  INV12 U1789 ( .A(compare_i_data_rs[13]), .Q(n417) );
  INV8 U1790 ( .A(n416), .Q(n436) );
  INV15 U1791 ( .A(n413), .Q(n425) );
  INV15 U1792 ( .A(n1152), .Q(n413) );
  NAND28 U1793 ( .A(n739), .B(n1123), .Q(n655) );
  AOI211 U1794 ( .A(n1641), .B(n423), .C(n1640), .Q(n1642) );
  AOI212 U1795 ( .A(n2420), .B(n2419), .C(n1926), .Q(n1927) );
  CLKIN3 U1796 ( .A(n1081), .Q(n1080) );
  NOR21 U1797 ( .A(n642), .B(n641), .Q(n640) );
  NOR31 U1798 ( .A(n2970), .B(n2972), .C(n1149), .Q(n2999) );
  OAI211 U1799 ( .A(n1164), .B(n2023), .C(n1994), .Q(n2007) );
  OAI212 U1800 ( .A(n2654), .B(n3075), .C(n3040), .Q(n3051) );
  OAI221 U1801 ( .A(n2100), .B(n1164), .C(n400), .D(n2221), .Q(n2106) );
  XNR21 U1802 ( .A(n2846), .B(n3041), .Q(n2848) );
  NAND21 U1803 ( .A(n2720), .B(n400), .Q(n2721) );
  NAND21 U1804 ( .A(n1851), .B(n404), .Q(n1852) );
  OAI212 U1805 ( .A(n1885), .B(n1887), .C(n1884), .Q(n1886) );
  IMUX20 U1806 ( .A(n2115), .B(n2114), .S(n408), .Q(n2116) );
  IMUX21 U1807 ( .A(n2747), .B(n2746), .S(n451), .Q(n2748) );
  NAND21 U1808 ( .A(n2525), .B(n401), .Q(n2526) );
  INV2 U1809 ( .A(n2779), .Q(n2678) );
  OAI212 U1810 ( .A(n2075), .B(n2074), .C(n2433), .Q(n2084) );
  CLKIN3 U1811 ( .A(n2393), .Q(n1009) );
  INV3 U1812 ( .A(n530), .Q(n529) );
  NAND21 U1813 ( .A(n2976), .B(n458), .Q(n2977) );
  NAND21 U1814 ( .A(n2501), .B(n362), .Q(n2174) );
  OAI211 U1815 ( .A(u_alu_lt_x_11_n84), .B(u_alu_lt_x_11_n87), .C(
        u_alu_lt_x_11_n85), .Q(u_alu_lt_x_11_n83) );
  INV3 U1816 ( .A(n2448), .Q(n2458) );
  NAND22 U1817 ( .A(n1929), .B(n2371), .Q(n1962) );
  CLKIN3 U1818 ( .A(n535), .Q(n534) );
  OAI222 U1819 ( .A(n1620), .B(n933), .C(n939), .D(n931), .Q(n930) );
  INV2 U1820 ( .A(n2304), .Q(n2292) );
  NAND21 U1821 ( .A(n2050), .B(n1167), .Q(n2051) );
  INV2 U1822 ( .A(n1864), .Q(n935) );
  INV3 U1823 ( .A(n2446), .Q(n953) );
  NAND22 U1824 ( .A(n378), .B(n817), .Q(n816) );
  INV3 U1825 ( .A(n2612), .Q(n1904) );
  INV2 U1826 ( .A(n2031), .Q(n1929) );
  NAND21 U1827 ( .A(n2361), .B(n2365), .Q(n2171) );
  CLKIN3 U1828 ( .A(n2714), .Q(n1709) );
  INV2 U1829 ( .A(n2417), .Q(n1823) );
  INV2 U1830 ( .A(u_alu_lt_x_11_n26), .Q(u_alu_lt_x_11_n24) );
  INV2 U1831 ( .A(n2942), .Q(n2738) );
  INV3 U1832 ( .A(u_alu_DP_OP_84J3_125_2615_n22), .Q(
        u_alu_DP_OP_84J3_125_2615_n77) );
  INV2 U1833 ( .A(n1068), .Q(n1067) );
  INV2 U1834 ( .A(n1764), .Q(n1689) );
  INV2 U1835 ( .A(n680), .Q(n435) );
  INV2 U1836 ( .A(n2837), .Q(n2700) );
  NAND22 U1837 ( .A(n552), .B(n3186), .Q(n554) );
  INV3 U1838 ( .A(n1759), .Q(n1760) );
  INV1 U1839 ( .A(n409), .Q(n775) );
  NAND21 U1840 ( .A(n1523), .B(i_data_FWmemout[10]), .Q(n1520) );
  INV3 U1841 ( .A(n1126), .Q(n1125) );
  INV3 U1842 ( .A(n1445), .Q(n683) );
  INV3 U1843 ( .A(n1721), .Q(n1722) );
  INV3 U1844 ( .A(n1638), .Q(n1603) );
  INV2 U1845 ( .A(n1691), .Q(n1694) );
  NAND22 U1846 ( .A(n1161), .B(i_data_rt[31]), .Q(n1178) );
  NAND22 U1847 ( .A(n393), .B(n1502), .Q(n834) );
  CLKIN3 U1848 ( .A(n1588), .Q(n1600) );
  CLKIN3 U1849 ( .A(n1240), .Q(n1114) );
  NAND22 U1850 ( .A(n456), .B(i_data_FMalures[12]), .Q(n1264) );
  NAND22 U1851 ( .A(n456), .B(i_data_FMalures[2]), .Q(n1479) );
  NAND21 U1852 ( .A(n9), .B(i_data_FMalures[7]), .Q(n460) );
  NAND22 U1853 ( .A(n9), .B(i_data_FMalures[18]), .Q(n1315) );
  NAND22 U1854 ( .A(n141), .B(i_data_FMmemout[6]), .Q(n1209) );
  INV2 U1855 ( .A(n2671), .Q(n3069) );
  INV2 U1856 ( .A(n1575), .Q(n1577) );
  INV1 U1857 ( .A(n3096), .Q(n3100) );
  NAND22 U1858 ( .A(n141), .B(i_data_FMmemout[12]), .Q(n1263) );
  NAND22 U1859 ( .A(n142), .B(i_data_FMmemout[4]), .Q(n1204) );
  INV6 U1860 ( .A(n401), .Q(n397) );
  NAND21 U1861 ( .A(i_con_Ealuop[4]), .B(n1148), .Q(n1575) );
  NOR21 U1862 ( .A(i_con_bop[2]), .B(n1311), .Q(n976) );
  CLKIN6 U1863 ( .A(n1166), .Q(n1165) );
  INV2 U1864 ( .A(i_data_FMalures[14]), .Q(n784) );
  NAND21 U1865 ( .A(n1901), .B(n849), .Q(n711) );
  INV3 U1866 ( .A(n2271), .Q(n2273) );
  NOR22 U1867 ( .A(n650), .B(n751), .Q(n641) );
  NAND31 U1868 ( .A(n751), .B(n749), .C(n650), .Q(n639) );
  OAI211 U1869 ( .A(n426), .B(n2261), .C(n2260), .Q(n2262) );
  OAI211 U1870 ( .A(n2074), .B(n2017), .C(n2016), .Q(n2026) );
  NAND22 U1871 ( .A(n2299), .B(n428), .Q(n479) );
  NAND21 U1872 ( .A(n2707), .B(n400), .Q(n2616) );
  AOI210 U1873 ( .A(n3121), .B(n628), .C(n2651), .Q(n2652) );
  INV2 U1874 ( .A(n2329), .Q(n2330) );
  OAI211 U1875 ( .A(n2790), .B(n2789), .C(n2788), .Q(n2791) );
  OAI211 U1876 ( .A(n2700), .B(n2790), .C(n2699), .Q(n2701) );
  CLKIN3 U1877 ( .A(n2175), .Q(n1989) );
  OAI221 U1878 ( .A(n1871), .B(n1166), .C(n1974), .D(n401), .Q(n1911) );
  NAND31 U1879 ( .A(n3097), .B(n1168), .C(n3096), .Q(n3098) );
  INV3 U1880 ( .A(n2740), .Q(n2540) );
  INV3 U1881 ( .A(n2833), .Q(n2639) );
  NAND21 U1882 ( .A(n146), .B(n434), .Q(n2993) );
  NAND21 U1883 ( .A(n3033), .B(n362), .Q(n535) );
  OAI211 U1884 ( .A(n386), .B(n1753), .C(n1606), .Q(n1608) );
  NAND21 U1885 ( .A(n146), .B(n3116), .Q(n3118) );
  CLKIN3 U1886 ( .A(u_alu_lt_x_11_n126), .Q(u_alu_lt_x_11_n124) );
  NAND21 U1887 ( .A(n146), .B(n2490), .Q(n2491) );
  NAND21 U1888 ( .A(n146), .B(n435), .Q(n3020) );
  CLKIN1 U1889 ( .A(n2813), .Q(n2769) );
  INV2 U1890 ( .A(n2845), .Q(n2733) );
  NAND22 U1891 ( .A(n1809), .B(u_alu_lt_x_11_B_5_), .Q(n910) );
  INV2 U1892 ( .A(n3147), .Q(n3149) );
  CLKIN3 U1893 ( .A(n929), .Q(n1972) );
  CLKIN2 U1894 ( .A(u_alu_lt_x_11_n54), .Q(u_alu_lt_x_11_n52) );
  CLKIN3 U1895 ( .A(n2981), .Q(n533) );
  INV3 U1896 ( .A(n1592), .Q(n1597) );
  INV2 U1897 ( .A(n1534), .Q(n722) );
  NAND21 U1898 ( .A(n383), .B(i_data_rt[18]), .Q(n1403) );
  INV3 U1899 ( .A(n1525), .Q(n551) );
  NAND21 U1900 ( .A(n1136), .B(i_data_FMmemout[16]), .Q(n1503) );
  NAND22 U1901 ( .A(n1136), .B(i_data_FMmemout[12]), .Q(n1257) );
  INV2 U1902 ( .A(n1454), .Q(n693) );
  INV3 U1903 ( .A(n1472), .Q(n498) );
  NAND22 U1904 ( .A(n1136), .B(i_data_FMmemout[25]), .Q(n1180) );
  NAND22 U1905 ( .A(n1136), .B(i_data_FMmemout[8]), .Q(n1269) );
  NAND22 U1906 ( .A(n9), .B(i_data_FMalures[16]), .Q(n1472) );
  NAND22 U1907 ( .A(n1135), .B(i_data_FMalures[15]), .Q(n1217) );
  NAND22 U1908 ( .A(n456), .B(i_data_FMalures[27]), .Q(n1426) );
  INV1 U1909 ( .A(n2641), .Q(n2095) );
  NAND21 U1910 ( .A(n1805), .B(n364), .Q(n1112) );
  INV2 U1911 ( .A(n3067), .Q(n2870) );
  INV3 U1912 ( .A(n361), .Q(n1041) );
  NAND21 U1913 ( .A(n1695), .B(n365), .Q(n1037) );
  INV6 U1914 ( .A(n385), .Q(n410) );
  INV2 U1915 ( .A(i_con_bop[2]), .Q(n1313) );
  OAI211 U1916 ( .A(n379), .B(n1669), .C(n1668), .Q(alu_o_data_AluRes[1]) );
  OAI221 U1917 ( .A(n2238), .B(n2023), .C(n851), .D(n426), .Q(n2024) );
  OAI211 U1918 ( .A(n2221), .B(n3074), .C(n2220), .Q(n2222) );
  NAND22 U1919 ( .A(n2902), .B(n2901), .Q(n2903) );
  OAI211 U1920 ( .A(n2210), .B(n2206), .C(n2205), .Q(n2207) );
  NOR31 U1921 ( .A(n2202), .B(n2203), .C(n2233), .Q(n2210) );
  NAND22 U1922 ( .A(n1983), .B(n404), .Q(n1984) );
  INV2 U1923 ( .A(n1867), .Q(n713) );
  NOR21 U1924 ( .A(n2176), .B(n401), .Q(n2177) );
  AOI221 U1925 ( .A(n362), .B(n1793), .C(n1652), .D(n1167), .Q(n1714) );
  IMUX20 U1926 ( .A(n2682), .B(n2681), .S(n450), .Q(n2683) );
  INV2 U1927 ( .A(n2765), .Q(n2767) );
  NAND31 U1928 ( .A(n2796), .B(n1163), .C(n458), .Q(n2797) );
  INV2 U1929 ( .A(n3092), .Q(n3087) );
  OAI210 U1930 ( .A(n2928), .B(n2927), .C(n362), .Q(n2929) );
  INV2 U1931 ( .A(n2028), .Q(n1977) );
  NOR21 U1932 ( .A(n2298), .B(n1118), .Q(n2325) );
  INV1 U1933 ( .A(n2381), .Q(n1729) );
  INV2 U1934 ( .A(n2156), .Q(n2068) );
  CLKIN2 U1935 ( .A(u_alu_lt_x_11_n43), .Q(n2732) );
  INV2 U1936 ( .A(u_alu_DP_OP_84J3_125_2615_n39), .Q(n427) );
  NAND22 U1937 ( .A(n3033), .B(n1167), .Q(n3119) );
  NAND21 U1938 ( .A(n1742), .B(n1778), .Q(n1688) );
  NOR21 U1939 ( .A(u_alu_lt_x_11_n15), .B(n3080), .Q(n3059) );
  NOR21 U1940 ( .A(u_alu_lt_x_11_n7), .B(n3079), .Q(n3092) );
  INV3 U1941 ( .A(n540), .Q(n539) );
  INV1 U1942 ( .A(n2362), .Q(n2246) );
  INV3 U1943 ( .A(u_alu_lt_x_11_B_19_), .Q(n1752) );
  INV2 U1944 ( .A(n2411), .Q(n1778) );
  INV2 U1945 ( .A(n823), .Q(n2857) );
  NAND22 U1946 ( .A(n3144), .B(n386), .Q(n540) );
  INV1 U1947 ( .A(u_alu_DP_OP_84J3_125_2615_n36), .Q(
        u_alu_DP_OP_84J3_125_2615_n111) );
  INV1 U1948 ( .A(n2376), .Q(n2254) );
  NAND22 U1949 ( .A(n3181), .B(n416), .Q(n504) );
  INV1 U1950 ( .A(n2734), .Q(n2699) );
  NAND22 U1951 ( .A(n3009), .B(n1170), .Q(n518) );
  INV3 U1952 ( .A(n1758), .Q(n1762) );
  INV2 U1953 ( .A(n1639), .Q(n1636) );
  INV1 U1954 ( .A(n1143), .Q(n1777) );
  INV2 U1955 ( .A(n371), .Q(n2531) );
  INV2 U1956 ( .A(n2470), .Q(n2476) );
  INV1 U1957 ( .A(n676), .Q(n3055) );
  INV2 U1958 ( .A(n1610), .Q(n634) );
  INV2 U1959 ( .A(compare_i_data_rs[30]), .Q(n447) );
  NAND41 U1960 ( .A(i_con_bop[0]), .B(i_con_bop[2]), .C(n1394), .D(n145), .Q(
        n1395) );
  NOR21 U1961 ( .A(n1208), .B(n1159), .Q(n1015) );
  NAND21 U1962 ( .A(n393), .B(i_data_rt[11]), .Q(n1246) );
  INV1 U1963 ( .A(n831), .Q(n2560) );
  INV2 U1964 ( .A(n1443), .Q(n637) );
  INV6 U1965 ( .A(n655), .Q(n402) );
  INV3 U1966 ( .A(n1228), .Q(n1230) );
  INV8 U1967 ( .A(n455), .Q(n941) );
  NAND22 U1968 ( .A(n1136), .B(i_data_FMmemout[2]), .Q(n754) );
  NAND22 U1969 ( .A(n1136), .B(i_data_FMmemout[10]), .Q(n1228) );
  INV2 U1970 ( .A(n1446), .Q(n765) );
  INV3 U1971 ( .A(n1357), .Q(n1130) );
  NAND22 U1972 ( .A(n9), .B(i_data_FMalures[3]), .Q(n1358) );
  NAND22 U1973 ( .A(n1134), .B(i_data_FMalures[12]), .Q(n1258) );
  NAND22 U1974 ( .A(n456), .B(i_data_FMalures[19]), .Q(n1465) );
  NAND22 U1975 ( .A(n1135), .B(i_data_FMalures[18]), .Q(n1318) );
  NAND22 U1976 ( .A(n1135), .B(i_data_FMalures[2]), .Q(n752) );
  INV3 U1977 ( .A(n1308), .Q(n879) );
  NAND22 U1978 ( .A(n1134), .B(i_data_FMalures[24]), .Q(n1345) );
  NAND22 U1979 ( .A(n1135), .B(i_data_FMalures[4]), .Q(n730) );
  NAND22 U1980 ( .A(n141), .B(i_data_FMmemout[3]), .Q(n1357) );
  NAND22 U1981 ( .A(n141), .B(i_data_FMmemout[19]), .Q(n1466) );
  NAND22 U1982 ( .A(n141), .B(i_data_FMmemout[8]), .Q(n1308) );
  NAND22 U1983 ( .A(n142), .B(i_data_FMmemout[1]), .Q(n1302) );
  INV2 U1984 ( .A(n386), .Q(n615) );
  INV3 U1985 ( .A(n1171), .Q(n420) );
  INV6 U1986 ( .A(n1165), .Q(n458) );
  INV1 U1987 ( .A(i_data_immext[13]), .Q(n2164) );
  CLKIN6 U1988 ( .A(i_data_immext[6]), .Q(n1163) );
  XNR21 U1989 ( .A(n3092), .B(n920), .Q(n3093) );
  NOR21 U1990 ( .A(n3178), .B(n2186), .Q(n2321) );
  AOI210 U1991 ( .A(n3121), .B(u_alu_lt_x_11_B_0_), .C(n2454), .Q(n2455) );
  OAI210 U1992 ( .A(n424), .B(n2402), .C(u_alu_lt_x_11_B_16_), .Q(n2407) );
  AOI221 U1993 ( .A(n2099), .B(n401), .C(n397), .D(n2266), .Q(n2221) );
  OAI210 U1994 ( .A(n414), .B(n738), .C(n736), .Q(n2906) );
  IMUX20 U1995 ( .A(n425), .B(n1154), .S(n374), .Q(n2628) );
  IMUX20 U1996 ( .A(n425), .B(n1154), .S(compare_i_data_rs[13]), .Q(n2211) );
  IMUX20 U1997 ( .A(n425), .B(n1154), .S(compare_i_data_rs[17]), .Q(n2483) );
  NOR21 U1998 ( .A(n2436), .B(n2423), .Q(n1997) );
  IMUX20 U1999 ( .A(n425), .B(n1154), .S(compare_i_data_rs[18]), .Q(n2534) );
  NAND21 U2000 ( .A(n2358), .B(n2246), .Q(n2256) );
  NOR21 U2001 ( .A(n2415), .B(n1823), .Q(n1879) );
  INV2 U2002 ( .A(n1064), .Q(n1063) );
  CLKIN3 U2003 ( .A(n1797), .Q(n1717) );
  INV1 U2004 ( .A(n1920), .Q(n562) );
  INV3 U2005 ( .A(n3006), .Q(n983) );
  INV2 U2006 ( .A(n3011), .Q(n797) );
  AOI211 U2007 ( .A(n3148), .B(n410), .C(n362), .Q(n2983) );
  INV1 U2008 ( .A(u_alu_lt_x_11_n84), .Q(n2234) );
  NAND21 U2009 ( .A(n146), .B(n1660), .Q(n1630) );
  NAND21 U2010 ( .A(n2417), .B(n1915), .Q(n1811) );
  INV2 U2011 ( .A(n850), .Q(n2238) );
  AOI211 U2012 ( .A(n3162), .B(n1170), .C(n410), .Q(n1902) );
  INV6 U2013 ( .A(n3178), .Q(n404) );
  INV2 U2014 ( .A(n860), .Q(n1840) );
  INV2 U2015 ( .A(n2422), .Q(n2233) );
  NOR21 U2016 ( .A(n2813), .B(n2812), .Q(n2814) );
  OAI212 U2017 ( .A(n416), .B(n3181), .C(n504), .Q(n503) );
  NOR21 U2018 ( .A(u_alu_lt_x_11_A_12_), .B(n446), .Q(n2169) );
  NOR21 U2019 ( .A(n420), .B(n1931), .Q(n860) );
  CLKIN2 U2020 ( .A(u_alu_lt_x_11_n50), .Q(u_alu_lt_x_11_n48) );
  NAND21 U2021 ( .A(n732), .B(n1244), .Q(n3188) );
  INV1 U2022 ( .A(u_alu_DP_OP_84J3_125_2615_n145), .Q(u_alu_lt_x_11_n171) );
  NAND21 U2023 ( .A(n2477), .B(n2469), .Q(n2470) );
  INV3 U2024 ( .A(n865), .Q(n688) );
  NAND22 U2025 ( .A(n1464), .B(n1463), .Q(n1367) );
  NAND22 U2026 ( .A(n1487), .B(n1488), .Q(n865) );
  INV2 U2027 ( .A(n1455), .Q(n692) );
  INV2 U2028 ( .A(n1593), .Q(n1594) );
  NAND22 U2029 ( .A(n1136), .B(i_data_FMmemout[3]), .Q(n1719) );
  INV3 U2030 ( .A(n1288), .Q(n1289) );
  NAND22 U2031 ( .A(n1136), .B(i_data_FMmemout[26]), .Q(n1198) );
  NAND22 U2032 ( .A(n456), .B(i_data_FMalures[5]), .Q(n1288) );
  NAND21 U2033 ( .A(n456), .B(i_data_FMalures[13]), .Q(n1251) );
  NAND22 U2034 ( .A(n1135), .B(i_data_FMalures[6]), .Q(n1206) );
  NAND22 U2035 ( .A(n1135), .B(i_data_FMalures[14]), .Q(n1108) );
  NAND21 U2036 ( .A(n9), .B(i_data_FMalures[8]), .Q(n1309) );
  NAND22 U2037 ( .A(n1135), .B(i_data_FMalures[20]), .Q(n1490) );
  NAND21 U2038 ( .A(n456), .B(i_data_FMalures[6]), .Q(n1210) );
  NAND22 U2039 ( .A(n141), .B(i_data_FMmemout[15]), .Q(n1223) );
  INV2 U2040 ( .A(n1570), .Q(n527) );
  INV2 U2041 ( .A(n1568), .Q(n1569) );
  NAND21 U2042 ( .A(n141), .B(i_data_FMmemout[11]), .Q(n1296) );
  NAND21 U2043 ( .A(n143), .B(i_data_FMmemout[7]), .Q(n1234) );
  INV3 U2044 ( .A(n397), .Q(n396) );
  INV2 U2045 ( .A(n1163), .Q(n509) );
  NOR21 U2046 ( .A(n599), .B(n598), .Q(n597) );
  NOR21 U2047 ( .A(n379), .B(n2060), .Q(n2061) );
  AOI221 U2048 ( .A(n1163), .B(n1654), .C(n1676), .D(n400), .Q(n1669) );
  INV2 U2049 ( .A(n3091), .Q(n3085) );
  MUX22 U2050 ( .A(n851), .B(n2103), .S(n509), .Q(n2060) );
  NAND21 U2051 ( .A(n2946), .B(n1163), .Q(n2947) );
  CLKIN3 U2052 ( .A(n885), .Q(n884) );
  OAI211 U2053 ( .A(n3074), .B(n2485), .C(n2484), .Q(n2499) );
  AOI211 U2054 ( .A(n413), .B(n435), .C(n422), .Q(n3019) );
  AOI211 U2055 ( .A(n413), .B(n434), .C(n422), .Q(n2992) );
  INV2 U2056 ( .A(n2074), .Q(n2038) );
  OAI210 U2057 ( .A(n424), .B(n2211), .C(u_alu_lt_x_11_B_13_), .Q(n2215) );
  AOI221 U2058 ( .A(n2266), .B(n401), .C(n458), .D(n2400), .Q(n2333) );
  OAI210 U2059 ( .A(n424), .B(n2483), .C(u_alu_lt_x_11_B_17_), .Q(n2484) );
  OAI221 U2060 ( .A(n1678), .B(n1163), .C(n1718), .D(n400), .Q(n1708) );
  OAI210 U2061 ( .A(n424), .B(n2628), .C(u_alu_lt_x_11_B_20_), .Q(n2629) );
  OAI210 U2062 ( .A(n424), .B(n2534), .C(u_alu_lt_x_11_B_18_), .Q(n2535) );
  OAI222 U2063 ( .A(n1871), .B(n1165), .C(n1797), .D(n458), .Q(n1836) );
  IMUX20 U2064 ( .A(n425), .B(n1154), .S(compare_i_data_rs[19]), .Q(n2602) );
  OAI220 U2065 ( .A(n410), .B(n1612), .C(n1671), .D(n386), .Q(n1614) );
  CLKIN2 U2066 ( .A(n940), .Q(n938) );
  BUF6 U2067 ( .A(n3158), .Q(n1155) );
  NAND21 U2068 ( .A(n146), .B(n2648), .Q(n2649) );
  INV1 U2069 ( .A(n2439), .Q(n2298) );
  INV3 U2070 ( .A(n1293), .Q(n1093) );
  NAND31 U2071 ( .A(n2738), .B(n362), .C(n386), .Q(n2739) );
  NAND21 U2072 ( .A(n2297), .B(n2440), .Q(n2328) );
  INV3 U2073 ( .A(n2369), .Q(n430) );
  INV2 U2074 ( .A(n628), .Q(n1774) );
  NAND21 U2075 ( .A(n3188), .B(n392), .Q(n1934) );
  INV2 U2076 ( .A(n2363), .Q(compare_i_data_rs[15]) );
  NAND22 U2077 ( .A(n144), .B(n1312), .Q(n1392) );
  NOR21 U2078 ( .A(n1632), .B(n1603), .Q(n559) );
  INV2 U2079 ( .A(n493), .Q(n492) );
  NAND22 U2080 ( .A(n343), .B(i_data_rs[31]), .Q(n1377) );
  NAND21 U2081 ( .A(n1161), .B(i_data_rt[17]), .Q(n555) );
  NAND22 U2082 ( .A(n1136), .B(i_data_FMmemout[5]), .Q(n1104) );
  NAND22 U2083 ( .A(n456), .B(i_data_FMalures[31]), .Q(n1372) );
  NAND22 U2084 ( .A(n142), .B(i_data_FMmemout[23]), .Q(n1447) );
  NAND22 U2085 ( .A(n143), .B(i_data_FMmemout[31]), .Q(n1373) );
  INV6 U2086 ( .A(n385), .Q(n1168) );
  OAI211 U2087 ( .A(n3074), .B(n2456), .C(n2455), .Q(n2457) );
  OAI211 U2088 ( .A(n2654), .B(n2527), .C(n2494), .Q(n2498) );
  INV2 U2089 ( .A(n3044), .Q(n1053) );
  NAND22 U2090 ( .A(n3044), .B(n676), .Q(n750) );
  AOI210 U2091 ( .A(n3121), .B(n372), .C(n2745), .Q(n2749) );
  CLKIN3 U2092 ( .A(n1712), .Q(n1713) );
  AOI210 U2093 ( .A(n3121), .B(u_alu_lt_x_11_B_5_), .C(n2683), .Q(n2686) );
  OAI210 U2094 ( .A(n424), .B(n2274), .C(u_alu_lt_x_11_B_14_), .Q(n2278) );
  OAI210 U2095 ( .A(n424), .B(n2602), .C(u_alu_lt_x_11_B_19_), .Q(n2603) );
  NAND22 U2096 ( .A(n936), .B(n934), .Q(n1712) );
  NOR21 U2097 ( .A(n458), .B(n3119), .Q(n3034) );
  AOI211 U2098 ( .A(u_alu_lt_x_11_n42), .B(u_alu_lt_x_11_n35), .C(
        u_alu_lt_x_11_n36), .Q(n469) );
  NAND21 U2099 ( .A(n2287), .B(n2358), .Q(n2232) );
  INV3 U2100 ( .A(n849), .Q(n426) );
  NOR22 U2101 ( .A(n2815), .B(n2814), .Q(n2816) );
  INV2 U2102 ( .A(n2353), .Q(n2287) );
  CLKIN3 U2103 ( .A(n2722), .Q(n2770) );
  INV2 U2104 ( .A(alu_i_data_B[7]), .Q(n429) );
  NAND21 U2105 ( .A(n2598), .B(n615), .Q(n614) );
  INV3 U2106 ( .A(n2027), .Q(n2952) );
  CLKIN3 U2107 ( .A(u_alu_lt_x_11_n49), .Q(u_alu_lt_x_11_n47) );
  NAND31 U2108 ( .A(n732), .B(u_alu_lt_x_11_A_5_), .C(n1244), .Q(n731) );
  INV2 U2109 ( .A(n1392), .Q(n1393) );
  INV1 U2110 ( .A(n2618), .Q(n2633) );
  AOI211 U2111 ( .A(n2595), .B(n1741), .C(n418), .Q(n1782) );
  NAND31 U2112 ( .A(n145), .B(i_con_bop[1]), .C(n1313), .Q(n1314) );
  INV2 U2113 ( .A(n490), .Q(n485) );
  INV2 U2114 ( .A(n1473), .Q(n1474) );
  NAND22 U2115 ( .A(n1243), .B(n1242), .Q(n967) );
  NAND22 U2116 ( .A(n1463), .B(n1464), .Q(compare_i_data_rs[20]) );
  NAND22 U2117 ( .A(n864), .B(n1110), .Q(n863) );
  INV1 U2118 ( .A(n2471), .Q(n2473) );
  NAND22 U2119 ( .A(n1572), .B(n457), .Q(n1634) );
  NOR21 U2120 ( .A(n1344), .B(n352), .Q(n1454) );
  INV2 U2121 ( .A(n1576), .Q(n1559) );
  NOR21 U2122 ( .A(n1573), .B(n1585), .Q(n1595) );
  INV3 U2123 ( .A(n1585), .Q(n457) );
  INV3 U2124 ( .A(n270), .Q(n1098) );
  INV2 U2125 ( .A(i_data_rt[12]), .Q(n1517) );
  AOI211 U2126 ( .A(n2690), .B(n2446), .C(n2408), .Q(n2461) );
  OAI2111 U2127 ( .A(n379), .B(n1751), .C(n1750), .D(n1749), .Q(
        alu_o_data_AluRes[3]) );
  AOI211 U2128 ( .A(n1155), .B(n2062), .C(n2061), .Q(n2091) );
  AOI211 U2129 ( .A(n2007), .B(n378), .C(n2006), .Q(n2008) );
  OAI211 U2130 ( .A(n1868), .B(n426), .C(n1837), .Q(n1838) );
  AOI221 U2131 ( .A(n1773), .B(n400), .C(n1164), .D(n1715), .Q(n1751) );
  AOI221 U2132 ( .A(n1674), .B(n1167), .C(n1673), .D(n362), .Q(n1755) );
  AOI210 U2133 ( .A(n3121), .B(u_alu_lt_x_11_B_1_), .C(n2493), .Q(n2494) );
  OAI210 U2134 ( .A(u_alu_lt_x_11_B_9_), .B(n425), .C(n1153), .Q(n2002) );
  NOR21 U2135 ( .A(n894), .B(n893), .Q(n1090) );
  OAI222 U2136 ( .A(n362), .B(n2399), .C(n1041), .D(n2398), .Q(n2525) );
  INV3 U2137 ( .A(n2391), .Q(n847) );
  AOI220 U2138 ( .A(n1700), .B(n423), .C(n1699), .D(n404), .Q(n1706) );
  NAND21 U2139 ( .A(n2976), .B(n401), .Q(n2890) );
  NAND22 U2140 ( .A(n2390), .B(n2389), .Q(n2391) );
  NAND21 U2141 ( .A(n1608), .B(n813), .Q(n812) );
  NAND22 U2142 ( .A(n755), .B(n756), .Q(n758) );
  INV3 U2143 ( .A(n2109), .Q(n2433) );
  NAND22 U2144 ( .A(n733), .B(n731), .Q(n1293) );
  INV2 U2145 ( .A(n2178), .Q(n1795) );
  INV2 U2146 ( .A(n1689), .Q(n564) );
  INV1 U2147 ( .A(n2723), .Q(n2619) );
  INV2 U2148 ( .A(n446), .Q(n2113) );
  NAND22 U2149 ( .A(n1392), .B(n1314), .Q(n1398) );
  INV2 U2150 ( .A(n2196), .Q(n974) );
  NOR21 U2151 ( .A(n2249), .B(n2248), .Q(n2196) );
  INV3 U2152 ( .A(n1808), .Q(n734) );
  INV3 U2153 ( .A(n7), .Q(n1244) );
  INV3 U2154 ( .A(u_alu_lt_x_11_A_0_), .Q(n419) );
  INV3 U2155 ( .A(n1806), .Q(n1808) );
  INV3 U2156 ( .A(n1404), .Q(n544) );
  INV1 U2157 ( .A(n1133), .Q(n1132) );
  NAND22 U2158 ( .A(n1574), .B(n457), .Q(n466) );
  INV3 U2159 ( .A(n1071), .Q(n1049) );
  NAND22 U2160 ( .A(n1148), .B(i_con_Ealuop[5]), .Q(n1568) );
  NAND21 U2161 ( .A(i_data_immext[12]), .B(n365), .Q(n1518) );
  AOI211 U2162 ( .A(n1394), .B(n1313), .C(i_con_bop[0]), .Q(n1312) );
  NOR21 U2163 ( .A(n400), .B(n1901), .Q(n1971) );
  AOI211 U2164 ( .A(n1814), .B(n423), .C(n1813), .Q(n1820) );
  NAND21 U2165 ( .A(n1044), .B(u_alu_pre_sum_4a[0]), .Q(n927) );
  OAI211 U2166 ( .A(n1164), .B(n2056), .C(n2055), .Q(n2062) );
  INV2 U2167 ( .A(n2289), .Q(n2230) );
  AOI210 U2168 ( .A(n413), .B(n2113), .C(n422), .Q(n2115) );
  INV3 U2169 ( .A(n1824), .Q(n1876) );
  OAI211 U2170 ( .A(n422), .B(n1892), .C(n1924), .Q(n1893) );
  IMUX21 U2171 ( .A(n1982), .B(n1981), .S(n1138), .Q(n1983) );
  INV3 U2172 ( .A(n2203), .Q(n2299) );
  OAI222 U2173 ( .A(n2053), .B(n1165), .C(n1974), .D(n458), .Q(n2044) );
  AOI210 U2174 ( .A(n2679), .B(n1153), .C(n441), .Q(n2680) );
  AOI210 U2175 ( .A(n3060), .B(n1153), .C(n431), .Q(n3072) );
  NAND20 U2176 ( .A(n2935), .B(n1153), .Q(n2940) );
  INV2 U2177 ( .A(n2589), .Q(n2579) );
  INV2 U2178 ( .A(n2986), .Q(n1026) );
  INV2 U2179 ( .A(n2117), .Q(n2120) );
  NOR21 U2180 ( .A(n2392), .B(n1845), .Q(n1855) );
  AOI221 U2181 ( .A(n1717), .B(n397), .C(n1716), .D(n401), .Q(n1784) );
  IMUX20 U2182 ( .A(n413), .B(n376), .S(u_alu_lt_x_11_A_0_), .Q(n1633) );
  INV3 U2183 ( .A(n1877), .Q(n1878) );
  INV1 U2184 ( .A(n2927), .Q(n2871) );
  NAND21 U2185 ( .A(n652), .B(n1949), .Q(n1862) );
  NAND22 U2186 ( .A(n2389), .B(n1847), .Q(n1767) );
  INV2 U2187 ( .A(n3081), .Q(n3083) );
  INV1 U2188 ( .A(n2431), .Q(n2297) );
  NOR21 U2189 ( .A(n420), .B(n1758), .Q(n2041) );
  INV2 U2190 ( .A(u_alu_lt_x_11_B_15_), .Q(n3168) );
  NOR21 U2191 ( .A(n2363), .B(u_alu_lt_x_11_B_15_), .Q(n2431) );
  NOR20 U2192 ( .A(n1775), .B(n1757), .Q(n912) );
  INV1 U2193 ( .A(compare_i_data_rs[28]), .Q(u_alu_lt_x_11_n172) );
  XOR21 U2194 ( .A(compare_i_data_rt[26]), .B(n979), .Q(n1391) );
  INV2 U2195 ( .A(n2145), .Q(n1353) );
  NAND22 U2196 ( .A(n383), .B(i_data_rt[21]), .Q(n1405) );
  NAND22 U2197 ( .A(n1161), .B(i_data_rt[3]), .Q(n1737) );
  NOR21 U2198 ( .A(n1317), .B(n1158), .Q(n1497) );
  INV2 U2199 ( .A(n1930), .Q(n1530) );
  NOR21 U2200 ( .A(n1369), .B(n353), .Q(n1416) );
  NAND22 U2201 ( .A(i_data_immext[15]), .B(n365), .Q(n2364) );
  INV3 U2202 ( .A(i_data_FEalures[29]), .Q(n1369) );
  AOI221 U2203 ( .A(n3175), .B(n2656), .C(n2690), .D(n2667), .Q(n1033) );
  AOI211 U2204 ( .A(n2710), .B(n3175), .C(n2709), .Q(n2711) );
  NAND28 U2205 ( .A(n1077), .B(n404), .Q(n1076) );
  AOI211 U2206 ( .A(n423), .B(n1839), .C(n1838), .Q(n1854) );
  AOI311 U2207 ( .A(n1889), .B(n1888), .C(n1887), .D(n1886), .Q(n1896) );
  OAI211 U2208 ( .A(n400), .B(n2780), .C(n2721), .Q(n2731) );
  NOR21 U2209 ( .A(n2270), .B(n2269), .Q(n2281) );
  NAND22 U2210 ( .A(n3071), .B(n401), .Q(n3094) );
  AOI211 U2211 ( .A(n2324), .B(n850), .C(n2323), .Q(n2338) );
  INV2 U2212 ( .A(n3135), .Q(n922) );
  NAND22 U2213 ( .A(n2719), .B(n458), .Q(n2646) );
  OAI222 U2214 ( .A(n2678), .B(n1165), .C(n397), .D(n2677), .Q(n2720) );
  NOR21 U2215 ( .A(n3002), .B(n2914), .Q(n2861) );
  AOI211 U2216 ( .A(n1848), .B(n1855), .C(n1857), .Q(n1849) );
  INV3 U2217 ( .A(n1848), .Q(n1859) );
  INV2 U2218 ( .A(n1855), .Q(n1860) );
  NOR21 U2219 ( .A(n2580), .B(n2582), .Q(n2546) );
  NAND22 U2220 ( .A(n428), .B(n512), .Q(n513) );
  INV3 U2221 ( .A(n2753), .Q(n2756) );
  INV10 U2222 ( .A(n2823), .Q(n2824) );
  INV2 U2223 ( .A(n2856), .Q(n993) );
  INV3 U2224 ( .A(n2654), .Q(n1874) );
  INV2 U2225 ( .A(n2351), .Q(n2288) );
  INV2 U2226 ( .A(n2368), .Q(n2140) );
  NOR21 U2227 ( .A(u_alu_lt_x_11_B_1_), .B(n2948), .Q(n1658) );
  INV2 U2228 ( .A(n947), .Q(n2093) );
  CLKIN3 U2229 ( .A(n822), .Q(n3105) );
  INV3 U2230 ( .A(n1742), .Q(n1743) );
  NOR21 U2231 ( .A(n1143), .B(n2411), .Q(n1923) );
  NAND20 U2232 ( .A(n3162), .B(n145), .Q(n908) );
  NAND22 U2233 ( .A(n2531), .B(u_alu_lt_x_11_A_2_), .Q(n1742) );
  INV2 U2234 ( .A(n1946), .Q(n1924) );
  NOR20 U2235 ( .A(n414), .B(n3009), .Q(u_alu_lt_x_11_n31) );
  INV2 U2236 ( .A(n2012), .Q(n1478) );
  INV2 U2237 ( .A(n635), .Q(n632) );
  NOR21 U2238 ( .A(n2143), .B(n1353), .Q(n1402) );
  INV1 U2239 ( .A(n2191), .Q(n2192) );
  NAND22 U2240 ( .A(n2165), .B(n2191), .Q(n2249) );
  NOR21 U2241 ( .A(n1203), .B(n1158), .Q(n727) );
  NAND22 U2242 ( .A(n398), .B(i_data_rs[5]), .Q(n1806) );
  NAND22 U2243 ( .A(n338), .B(i_data_FWmemout[5]), .Q(n1242) );
  INV3 U2244 ( .A(n1529), .Q(n550) );
  NOR21 U2245 ( .A(n1352), .B(n281), .Q(n2143) );
  INV3 U2246 ( .A(n1719), .Q(n1725) );
  INV3 U2247 ( .A(n1275), .Q(n1278) );
  NOR21 U2248 ( .A(n1506), .B(n353), .Q(n1290) );
  NOR21 U2249 ( .A(n1346), .B(n351), .Q(n484) );
  INV3 U2250 ( .A(i_data_FEalures[28]), .Q(n1319) );
  INV2 U2251 ( .A(i_data_FEalures[2]), .Q(n1387) );
  INV3 U2252 ( .A(i_data_FEalures[30]), .Q(n1371) );
  INV3 U2253 ( .A(i_data_FEalures[27]), .Q(n1380) );
  INV2 U2254 ( .A(i_data_FEalures[13]), .Q(n1249) );
  INV3 U2255 ( .A(i_data_FEalures[16]), .Q(n1506) );
  IMUX21 U2256 ( .A(i_addr_rt[2]), .B(i_data_immext[13]), .S(i_con_Eregdst), 
        .Q(n3200) );
  INV2 U2257 ( .A(i_data_FWmemout[14]), .Q(n1226) );
  INV3 U2258 ( .A(i_data_immext[3]), .Q(n1583) );
  INV2 U2259 ( .A(i_data_FEalures[11]), .Q(n1295) );
  INV2 U2260 ( .A(i_data_FEalures[1]), .Q(n1301) );
  AOI211 U2261 ( .A(n2698), .B(n2587), .C(n2586), .Q(n2609) );
  AOI211 U2262 ( .A(n2690), .B(n2689), .C(n2688), .Q(n2713) );
  INV3 U2263 ( .A(n1149), .Q(n2913) );
  NAND24 U2264 ( .A(n1061), .B(n661), .Q(n658) );
  NOR21 U2265 ( .A(n2507), .B(n2847), .Q(n2508) );
  NOR21 U2266 ( .A(n459), .B(n2847), .Q(n2547) );
  INV3 U2267 ( .A(n1844), .Q(n1802) );
  INV2 U2268 ( .A(n1881), .Q(n1888) );
  NAND22 U2269 ( .A(n2210), .B(n2218), .Q(n2216) );
  INV3 U2270 ( .A(n2092), .Q(n2100) );
  NAND21 U2271 ( .A(n2946), .B(n400), .Q(n2892) );
  NAND28 U2272 ( .A(n2860), .B(n3088), .Q(n977) );
  OAI211 U2273 ( .A(n2531), .B(n3167), .C(n2530), .Q(n2532) );
  INV2 U2274 ( .A(n2217), .Q(n2219) );
  NAND22 U2275 ( .A(n2044), .B(n1163), .Q(n1975) );
  OAI222 U2276 ( .A(n1165), .B(n2054), .C(n2053), .D(n397), .Q(n2092) );
  NAND22 U2277 ( .A(n3152), .B(n458), .Q(n3095) );
  OAI211 U2278 ( .A(n1167), .B(n3101), .C(n3028), .Q(n3031) );
  AOI211 U2279 ( .A(n413), .B(n1660), .C(n422), .Q(n1629) );
  NAND21 U2280 ( .A(n3046), .B(n3044), .Q(n1051) );
  INV3 U2281 ( .A(n924), .Q(n2968) );
  IMUX21 U2282 ( .A(n2492), .B(n2491), .S(n415), .Q(n2493) );
  INV2 U2283 ( .A(n2083), .Q(n477) );
  NAND22 U2284 ( .A(n2542), .B(n458), .Q(n2543) );
  INV2 U2285 ( .A(n2866), .Q(n2795) );
  NAND22 U2286 ( .A(n2111), .B(n2438), .Q(n2203) );
  NAND22 U2287 ( .A(n412), .B(n2620), .Q(n978) );
  NOR20 U2288 ( .A(n2376), .B(n2304), .Q(n2305) );
  NOR21 U2289 ( .A(n2373), .B(n2140), .Q(n951) );
  NAND22 U2290 ( .A(n2403), .B(n1167), .Q(n2404) );
  INV3 U2291 ( .A(n2754), .Q(n2766) );
  INV3 U2292 ( .A(n755), .Q(u_alu_DP_OP_84J3_125_2615_n49) );
  INV1 U2293 ( .A(n2370), .Q(n1979) );
  NAND21 U2294 ( .A(n146), .B(n1914), .Q(n1799) );
  NOR21 U2295 ( .A(n2635), .B(n2637), .Q(n2584) );
  NAND21 U2296 ( .A(n146), .B(n1649), .Q(n2452) );
  NOR21 U2297 ( .A(n1171), .B(n2849), .Q(n1648) );
  AOI2110 U2298 ( .A(n419), .B(n1660), .C(n1690), .D(n3178), .Q(n1640) );
  INV3 U2299 ( .A(u_alu_DP_OP_84J3_125_2615_n30), .Q(
        u_alu_DP_OP_84J3_125_2615_n81) );
  INV3 U2300 ( .A(u_alu_DP_OP_84J3_125_2615_n31), .Q(
        u_alu_DP_OP_84J3_125_2615_n86) );
  INV3 U2301 ( .A(n1918), .Q(n1069) );
  INV3 U2302 ( .A(n3010), .Q(n3001) );
  NAND22 U2303 ( .A(n384), .B(n1171), .Q(n822) );
  NOR20 U2304 ( .A(u_alu_lt_x_11_n159), .B(u_alu_lt_x_11_B_15_), .Q(
        u_alu_lt_x_11_n78) );
  NOR21 U2305 ( .A(u_alu_lt_x_11_B_17_), .B(n415), .Q(u_alu_lt_x_11_n72) );
  INV2 U2306 ( .A(n2413), .Q(n856) );
  INV1 U2307 ( .A(u_alu_lt_x_11_B_17_), .Q(n2490) );
  NAND22 U2308 ( .A(n2575), .B(n2574), .Q(n2620) );
  INV3 U2309 ( .A(n972), .Q(n593) );
  INV3 U2310 ( .A(n633), .Q(n1611) );
  NAND22 U2311 ( .A(n1402), .B(n2150), .Q(n3181) );
  OAI211 U2312 ( .A(n1937), .B(n139), .C(n1936), .Q(n1943) );
  INV2 U2313 ( .A(n1684), .Q(n805) );
  AOI211 U2314 ( .A(n383), .B(n1519), .C(n2247), .Q(n1623) );
  INV3 U2315 ( .A(n531), .Q(n980) );
  INV3 U2316 ( .A(n560), .Q(n802) );
  NAND21 U2317 ( .A(n2553), .B(n377), .Q(n493) );
  NAND22 U2318 ( .A(n382), .B(i_data_rt[20]), .Q(n1404) );
  NAND22 U2319 ( .A(n398), .B(i_data_rs[10]), .Q(n1476) );
  NOR21 U2320 ( .A(n1304), .B(n941), .Q(n481) );
  NOR21 U2321 ( .A(n1383), .B(n281), .Q(n624) );
  INV3 U2322 ( .A(n2472), .Q(n1500) );
  INV2 U2323 ( .A(n1424), .Q(n546) );
  NOR21 U2324 ( .A(n1232), .B(n347), .Q(n1237) );
  NOR21 U2325 ( .A(n1366), .B(n347), .Q(n1462) );
  NOR21 U2326 ( .A(n1322), .B(n220), .Q(n1424) );
  INV2 U2327 ( .A(n1470), .Q(n557) );
  INV3 U2328 ( .A(n2134), .Q(n2013) );
  NAND21 U2329 ( .A(n456), .B(i_data_FMalures[30]), .Q(n472) );
  NAND21 U2330 ( .A(n142), .B(i_data_FMmemout[25]), .Q(n1434) );
  INV2 U2331 ( .A(n1549), .Q(n1544) );
  NAND31 U2332 ( .A(n1584), .B(n1583), .C(n561), .Q(n1586) );
  NAND22 U2333 ( .A(n719), .B(i_data_immext[1]), .Q(n718) );
  INV3 U2334 ( .A(n1561), .Q(n561) );
  INV3 U2335 ( .A(i_data_FEalures[22]), .Q(n1342) );
  INV2 U2336 ( .A(i_data_FWmemout[29]), .Q(n1368) );
  INV2 U2337 ( .A(i_data_rt[16]), .Q(n1509) );
  INV2 U2338 ( .A(i_data_rt[17]), .Q(n1501) );
  INV2 U2339 ( .A(i_data_rs[3]), .Q(n1131) );
  NOR22 U2340 ( .A(n1084), .B(n1083), .Q(n1082) );
  NAND31 U2341 ( .A(n2610), .B(n2609), .C(n2608), .Q(alu_o_data_AluRes[19]) );
  NAND33 U2342 ( .A(n659), .B(n404), .C(n943), .Q(n3077) );
  NAND22 U2343 ( .A(n996), .B(n995), .Q(n994) );
  NOR23 U2344 ( .A(n568), .B(n658), .Q(n657) );
  NOR22 U2345 ( .A(n380), .B(n2104), .Q(n2105) );
  NOR22 U2346 ( .A(n883), .B(n884), .Q(n2104) );
  NOR22 U2347 ( .A(n3178), .B(n3128), .Q(n661) );
  AOI211 U2348 ( .A(n2991), .B(n378), .C(n2990), .Q(n2998) );
  NAND22 U2349 ( .A(n2300), .B(n2299), .Q(n2119) );
  NAND22 U2350 ( .A(n2300), .B(n2111), .Q(n2035) );
  INV3 U2351 ( .A(n1034), .Q(n1028) );
  NOR22 U2352 ( .A(n400), .B(n2103), .Q(n883) );
  INV3 U2353 ( .A(n2684), .Q(n2653) );
  NAND22 U2354 ( .A(n667), .B(n529), .Q(n528) );
  NAND22 U2355 ( .A(n2570), .B(n400), .Q(n2544) );
  NAND31 U2356 ( .A(n2217), .B(n423), .C(n2209), .Q(n2206) );
  INV3 U2357 ( .A(n479), .Q(n478) );
  OAI211 U2358 ( .A(n2876), .B(n422), .C(u_alu_DP_OP_84J3_125_2615_n134), .Q(
        n2877) );
  IMUX21 U2359 ( .A(n1702), .B(n1701), .S(n439), .Q(n1705) );
  IMUX21 U2360 ( .A(n2002), .B(n2001), .S(n436), .Q(n2003) );
  NOR24 U2361 ( .A(n2821), .B(n2820), .Q(n944) );
  IMUX21 U2362 ( .A(n2453), .B(n2452), .S(n432), .Q(n2454) );
  OAI222 U2363 ( .A(n2258), .B(n1165), .C(n2406), .D(n397), .Q(n2324) );
  INV3 U2364 ( .A(n476), .Q(n475) );
  NAND21 U2365 ( .A(n1661), .B(n423), .Q(n1662) );
  NOR21 U2366 ( .A(n2932), .B(n2793), .Q(n2564) );
  IMUX21 U2367 ( .A(n425), .B(n1154), .S(u_alu_lt_x_11_A_2_), .Q(n1703) );
  IMUX21 U2368 ( .A(n425), .B(n1154), .S(compare_i_data_rs[15]), .Q(n2322) );
  IMUX21 U2369 ( .A(n425), .B(n1154), .S(u_alu_DP_OP_83J3_124_3384_n154), .Q(
        n2402) );
  NAND21 U2370 ( .A(n2111), .B(n2107), .Q(n476) );
  IMUX21 U2371 ( .A(n425), .B(n1154), .S(u_alu_DP_OP_84J3_125_2615_n145), .Q(
        n2995) );
  INV3 U2372 ( .A(n2437), .Q(n747) );
  IMUX20 U2373 ( .A(n425), .B(n1154), .S(compare_i_data_rs[24]), .Q(n2876) );
  INV2 U2374 ( .A(n2495), .Q(n2480) );
  INV3 U2375 ( .A(n1351), .Q(n779) );
  INV2 U2376 ( .A(n1727), .Q(n1730) );
  NOR21 U2377 ( .A(n2513), .B(n2623), .Q(n2495) );
  INV2 U2378 ( .A(u_alu_lt_x_11_n30), .Q(u_alu_lt_x_11_n28) );
  OAI211 U2379 ( .A(n386), .B(n2049), .C(n2309), .Q(n2050) );
  NAND22 U2380 ( .A(n2849), .B(n433), .Q(n755) );
  NOR21 U2381 ( .A(u_alu_lt_x_11_B_14_), .B(n2948), .Q(n2275) );
  NAND21 U2382 ( .A(n429), .B(n358), .Q(u_alu_lt_x_11_n119) );
  NAND22 U2383 ( .A(n2704), .B(n410), .Q(n2173) );
  INV2 U2384 ( .A(n911), .Q(n1913) );
  INV3 U2385 ( .A(n2387), .Q(n654) );
  NOR21 U2386 ( .A(n371), .B(n2948), .Q(n1701) );
  NAND22 U2387 ( .A(n2841), .B(n2842), .Q(n926) );
  INV3 U2388 ( .A(n3027), .Q(n2704) );
  INV2 U2389 ( .A(n2350), .Q(n2064) );
  NAND22 U2390 ( .A(n2775), .B(n1018), .Q(n2777) );
  NAND22 U2391 ( .A(n2621), .B(n2620), .Q(n2657) );
  INV2 U2392 ( .A(n1960), .Q(n1776) );
  NOR31 U2393 ( .A(n819), .B(n1167), .C(n380), .Q(n811) );
  NAND22 U2394 ( .A(u_alu_lt_x_11_B_5_), .B(u_alu_lt_x_11_A_5_), .Q(n1846) );
  NOR21 U2395 ( .A(n2776), .B(n3162), .Q(n2613) );
  NOR21 U2396 ( .A(n3069), .B(n438), .Q(n2926) );
  NAND20 U2397 ( .A(u_alu_lt_x_11_B_15_), .B(u_alu_lt_x_11_n159), .Q(
        u_alu_lt_x_11_n79) );
  INV3 U2398 ( .A(n774), .Q(n1920) );
  NAND22 U2399 ( .A(n622), .B(n2372), .Q(n2373) );
  AOI220 U2400 ( .A(alu_i_data_B[31]), .B(n1171), .C(u_alu_lt_x_11_B_15_), .D(
        n1170), .Q(n3145) );
  NAND31 U2401 ( .A(n387), .B(n386), .C(n1171), .Q(n2775) );
  NAND22 U2402 ( .A(n3009), .B(compare_i_data_rs[25]), .Q(
        u_alu_DP_OP_84J3_125_2615_n48) );
  NAND21 U2403 ( .A(n446), .B(n1170), .Q(n3026) );
  INV3 U2404 ( .A(u_alu_lt_x_11_A_2_), .Q(n439) );
  INV2 U2405 ( .A(n471), .Q(n2982) );
  INV2 U2406 ( .A(n2395), .Q(n1951) );
  INV2 U2407 ( .A(n1692), .Q(n1693) );
  NAND22 U2408 ( .A(n2443), .B(n2442), .Q(u_alu_DP_OP_83J3_124_3384_n154) );
  NOR21 U2409 ( .A(n1162), .B(compare_i_data_rs[19]), .Q(n2575) );
  NAND22 U2410 ( .A(compare_i_data_rt[25]), .B(n139), .Q(n1609) );
  NAND24 U2411 ( .A(n3187), .B(n391), .Q(n821) );
  NAND22 U2412 ( .A(n577), .B(n576), .Q(n575) );
  INV3 U2413 ( .A(n704), .Q(n563) );
  NAND22 U2414 ( .A(n485), .B(n1231), .Q(n1528) );
  INV1 U2415 ( .A(n1952), .Q(n1956) );
  INV3 U2416 ( .A(n1247), .Q(n787) );
  INV3 U2417 ( .A(n1015), .Q(n1014) );
  INV2 U2418 ( .A(n702), .Q(n697) );
  NAND22 U2419 ( .A(n1527), .B(n550), .Q(n549) );
  NAND22 U2420 ( .A(n1527), .B(n1525), .Q(n488) );
  NAND22 U2421 ( .A(n383), .B(i_data_rt[8]), .Q(n1273) );
  NAND22 U2422 ( .A(n550), .B(n1231), .Q(n486) );
  NAND22 U2423 ( .A(n1737), .B(n1362), .Q(n760) );
  NAND31 U2424 ( .A(n1685), .B(n574), .C(n138), .Q(n1687) );
  NAND22 U2425 ( .A(n398), .B(i_data_rs[21]), .Q(n1456) );
  NAND22 U2426 ( .A(n343), .B(i_data_rs[16]), .Q(n1473) );
  NAND22 U2427 ( .A(n343), .B(i_data_rs[9]), .Q(n560) );
  NAND22 U2428 ( .A(n521), .B(n1447), .Q(n520) );
  NAND22 U2429 ( .A(n1108), .B(n1109), .Q(n1512) );
  NAND22 U2430 ( .A(n338), .B(i_data_FWmemout[0]), .Q(n1685) );
  NAND22 U2431 ( .A(n398), .B(i_data_rs[26]), .Q(n531) );
  INV3 U2432 ( .A(n1139), .Q(n1140) );
  NOR21 U2433 ( .A(n1319), .B(n1158), .Q(n1484) );
  INV2 U2434 ( .A(n1436), .Q(n703) );
  NOR21 U2435 ( .A(n1349), .B(n281), .Q(n1350) );
  NOR21 U2436 ( .A(n1383), .B(n220), .Q(n1431) );
  INV1 U2437 ( .A(n1123), .Q(n1245) );
  NAND21 U2438 ( .A(n9), .B(i_data_FMalures[11]), .Q(n461) );
  NOR21 U2439 ( .A(n1233), .B(n353), .Q(n1236) );
  NAND22 U2440 ( .A(n1571), .B(n527), .Q(n1572) );
  NAND21 U2441 ( .A(n2641), .B(n1172), .Q(n2151) );
  INV2 U2442 ( .A(n932), .Q(n931) );
  NAND21 U2443 ( .A(n456), .B(i_data_FMalures[29]), .Q(n1414) );
  NOR21 U2444 ( .A(n1361), .B(n352), .Q(n1359) );
  NOR21 U2445 ( .A(n1342), .B(n353), .Q(n1449) );
  NAND21 U2446 ( .A(n456), .B(i_data_FMalures[20]), .Q(n1458) );
  NAND21 U2447 ( .A(n9), .B(i_data_FMalures[28]), .Q(n1420) );
  NAND21 U2448 ( .A(n456), .B(i_data_FMalures[21]), .Q(n1451) );
  NAND21 U2449 ( .A(n9), .B(i_data_FMalures[24]), .Q(n1441) );
  NOR21 U2450 ( .A(n1319), .B(n352), .Q(n1423) );
  NAND21 U2451 ( .A(n143), .B(i_data_FMmemout[30]), .Q(n1409) );
  NAND22 U2452 ( .A(n364), .B(n1514), .Q(n1513) );
  NAND21 U2453 ( .A(n142), .B(i_data_FMmemout[16]), .Q(n523) );
  NAND21 U2454 ( .A(n143), .B(i_data_FMmemout[21]), .Q(n1452) );
  NAND22 U2455 ( .A(n1041), .B(n385), .Q(n2943) );
  INV2 U2456 ( .A(i_data_rs[8]), .Q(n1094) );
  INV3 U2457 ( .A(i_data_FEalures[23]), .Q(n1333) );
  INV3 U2458 ( .A(i_data_FEalures[9]), .Q(n1356) );
  INV3 U2459 ( .A(i_data_FEalures[18]), .Q(n1317) );
  INV2 U2460 ( .A(i_data_FEalures[20]), .Q(n1365) );
  INV3 U2461 ( .A(i_data_FEalures[10]), .Q(n1305) );
  INV3 U2462 ( .A(i_data_FWmemout[10]), .Q(n1304) );
  NAND22 U2463 ( .A(n2091), .B(n2090), .Q(alu_o_data_AluRes[11]) );
  NAND33 U2464 ( .A(u_alu_pre_sum_4b[2]), .B(n2919), .C(n659), .Q(n2961) );
  NAND33 U2465 ( .A(n646), .B(n3073), .C(n644), .Q(n643) );
  AOI212 U2466 ( .A(n2509), .B(n378), .C(n2508), .Q(n2510) );
  NAND22 U2467 ( .A(n601), .B(n597), .Q(alu_o_data_AluRes[0]) );
  AOI211 U2468 ( .A(n3175), .B(n2573), .C(n2572), .Q(n2610) );
  AOI212 U2469 ( .A(n2548), .B(n378), .C(n2547), .Q(n2549) );
  NAND22 U2470 ( .A(n640), .B(n639), .Q(n649) );
  BUF15 U2471 ( .A(n2827), .Q(n659) );
  NAND31 U2472 ( .A(n1854), .B(n1853), .C(n1852), .Q(alu_o_data_AluRes[6]) );
  NAND22 U2473 ( .A(n2997), .B(n2973), .Q(n464) );
  NOR22 U2474 ( .A(n2785), .B(n2784), .Q(n2786) );
  INV8 U2475 ( .A(n3128), .Q(n1077) );
  NAND22 U2476 ( .A(n2306), .B(n664), .Q(n2317) );
  OAI211 U2477 ( .A(n2723), .B(n2771), .C(n2691), .Q(n2692) );
  AOI211 U2478 ( .A(n850), .B(n1844), .C(n1843), .Q(n1853) );
  OAI211 U2479 ( .A(n2979), .B(n1163), .C(n2947), .Q(n2953) );
  AOI212 U2480 ( .A(n928), .B(n3091), .C(n3090), .Q(n920) );
  NAND31 U2481 ( .A(n3155), .B(n3156), .C(n1163), .Q(n3113) );
  XOR21 U2482 ( .A(u_alu_DP_OP_84J3_125_2615_n1), .B(
        u_alu_DP_OP_84J3_125_2615_n68), .Q(u_alu_pre_sum_4b[7]) );
  OAI211 U2483 ( .A(n400), .B(n2893), .C(n2892), .Q(n2904) );
  AOI211 U2484 ( .A(n2908), .B(n2907), .C(n2906), .Q(n2909) );
  OAI211 U2485 ( .A(n1164), .B(n1976), .C(n1975), .Q(n1987) );
  OAI311 U2486 ( .A(n1958), .B(n1860), .C(n1859), .D(n1858), .Q(n1861) );
  OAI211 U2487 ( .A(n2979), .B(n400), .C(n2978), .Q(n2991) );
  IMUX21 U2488 ( .A(n3020), .B(n3019), .S(compare_i_data_rs[28]), .Q(n3021) );
  NAND22 U2489 ( .A(n3065), .B(n1022), .Q(n1021) );
  NAND22 U2490 ( .A(n750), .B(n3081), .Q(n3056) );
  INV2 U2491 ( .A(n2272), .Q(n2270) );
  IMUX21 U2492 ( .A(n2213), .B(n2212), .S(n417), .Q(n2214) );
  NAND22 U2493 ( .A(n1865), .B(n1167), .Q(n1866) );
  OAI211 U2494 ( .A(n401), .B(n2313), .C(n2182), .Q(n2259) );
  INV2 U2495 ( .A(n2324), .Q(n2261) );
  IMUX21 U2496 ( .A(n1659), .B(n1658), .S(n875), .Q(n1663) );
  INV2 U2497 ( .A(n3032), .Q(n3036) );
  OAI211 U2498 ( .A(n401), .B(n2891), .C(n2890), .Q(n2946) );
  AOI211 U2499 ( .A(n378), .B(n1024), .C(n3072), .Q(n1022) );
  NOR21 U2500 ( .A(n401), .B(n2936), .Q(n2938) );
  NAND22 U2501 ( .A(n616), .B(n612), .Q(n2627) );
  IMUX21 U2502 ( .A(n1891), .B(n1890), .S(n357), .Q(n1894) );
  XNR21 U2503 ( .A(n1783), .B(n1824), .Q(n1785) );
  AOI221 U2504 ( .A(n1734), .B(n1155), .C(n1733), .D(n404), .Q(n1750) );
  IMUX20 U2505 ( .A(n2529), .B(n2528), .S(n2636), .Q(n2530) );
  NOR31 U2506 ( .A(n401), .B(n1163), .C(n2795), .Q(n2800) );
  OAI221 U2507 ( .A(n1678), .B(n400), .C(n1656), .D(n1164), .Q(n1667) );
  INV2 U2508 ( .A(n1997), .Q(n1995) );
  INV3 U2509 ( .A(n613), .Q(n612) );
  OAI211 U2510 ( .A(n2654), .B(n1656), .C(n1642), .Q(n1643) );
  OAI221 U2511 ( .A(n1784), .B(n400), .C(n1718), .D(n1163), .Q(n1734) );
  NAND21 U2512 ( .A(n2181), .B(n401), .Q(n2182) );
  OAI221 U2513 ( .A(n1615), .B(n401), .C(n1675), .D(n1166), .Q(n1654) );
  NAND22 U2514 ( .A(n746), .B(n745), .Q(n744) );
  NOR21 U2515 ( .A(u_alu_lt_x_11_n115), .B(u_alu_lt_x_11_n117), .Q(
        u_alu_lt_x_11_n113) );
  OAI211 U2516 ( .A(n2582), .B(n2662), .C(n2581), .Q(n2583) );
  AOI211 U2517 ( .A(n2565), .B(n2611), .C(n2564), .Q(n2566) );
  NOR31 U2518 ( .A(n2010), .B(n1156), .C(n1997), .Q(n2000) );
  NAND22 U2519 ( .A(n1042), .B(n1040), .Q(n3152) );
  NAND22 U2520 ( .A(n1779), .B(n853), .Q(n852) );
  AOI211 U2521 ( .A(n2639), .B(n2562), .C(n2580), .Q(n2563) );
  NAND22 U2522 ( .A(n538), .B(n396), .Q(n536) );
  INV2 U2523 ( .A(n2965), .Q(n2924) );
  NAND21 U2524 ( .A(n3070), .B(n394), .Q(n1042) );
  OAI211 U2525 ( .A(n2577), .B(n2576), .C(n2625), .Q(n2578) );
  OAI211 U2526 ( .A(n2068), .B(n2067), .C(n2344), .Q(n2069) );
  AOI211 U2527 ( .A(u_alu_lt_x_11_n119), .B(u_alu_lt_x_11_n124), .C(
        u_alu_lt_x_11_n120), .Q(u_alu_lt_x_11_n118) );
  INV2 U2528 ( .A(n3120), .Q(n1025) );
  NAND22 U2529 ( .A(n3070), .B(n1167), .Q(n2987) );
  NAND22 U2530 ( .A(u_alu_lt_x_11_n100), .B(u_alu_lt_x_11_n104), .Q(
        u_alu_lt_x_11_n98) );
  NOR21 U2531 ( .A(n401), .B(n3119), .Q(n3165) );
  NOR21 U2532 ( .A(n2381), .B(n1728), .Q(n1698) );
  NAND22 U2533 ( .A(n2894), .B(n394), .Q(n2988) );
  NOR21 U2534 ( .A(n401), .B(n3061), .Q(n3120) );
  NOR21 U2535 ( .A(n2641), .B(n187), .Q(n2642) );
  NAND21 U2536 ( .A(n146), .B(n2113), .Q(n2114) );
  INV2 U2537 ( .A(u_alu_lt_x_11_n125), .Q(u_alu_lt_x_11_n123) );
  INV2 U2538 ( .A(n1908), .Q(n1769) );
  NAND21 U2539 ( .A(n146), .B(n3162), .Q(n3164) );
  INV2 U2540 ( .A(u_alu_lt_x_11_n76), .Q(u_alu_lt_x_11_n74) );
  AOI221 U2541 ( .A(n2613), .B(n1167), .C(n2612), .D(n2611), .Q(n2614) );
  INV2 U2542 ( .A(u_alu_lt_x_11_n107), .Q(u_alu_lt_x_11_n105) );
  INV2 U2543 ( .A(n2365), .Q(n2253) );
  INV2 U2544 ( .A(u_alu_lt_x_11_n106), .Q(u_alu_lt_x_11_n104) );
  NOR21 U2545 ( .A(n2027), .B(n2948), .Q(n2014) );
  NOR21 U2546 ( .A(u_alu_lt_x_11_B_9_), .B(n2948), .Q(n2001) );
  INV2 U2547 ( .A(u_alu_lt_x_11_n122), .Q(u_alu_lt_x_11_n120) );
  NAND21 U2548 ( .A(n409), .B(n372), .Q(u_alu_lt_x_11_n126) );
  INV1 U2549 ( .A(n2580), .Q(n2581) );
  INV1 U2550 ( .A(n2621), .Q(n2577) );
  INV2 U2551 ( .A(n908), .Q(n603) );
  NOR21 U2552 ( .A(u_alu_lt_x_11_B_13_), .B(n2948), .Q(n2212) );
  INV2 U2553 ( .A(u_alu_lt_x_11_n29), .Q(u_alu_lt_x_11_n27) );
  INV2 U2554 ( .A(u_alu_lt_x_11_n73), .Q(u_alu_lt_x_11_n71) );
  INV2 U2555 ( .A(u_alu_lt_x_11_n77), .Q(u_alu_lt_x_11_n75) );
  OAI210 U2556 ( .A(n410), .B(n3149), .C(n3148), .Q(n3150) );
  INV1 U2557 ( .A(n2425), .Q(n1912) );
  INV2 U2558 ( .A(n966), .Q(n965) );
  NAND22 U2559 ( .A(n909), .B(n403), .Q(n618) );
  INV2 U2560 ( .A(u_alu_lt_x_11_n94), .Q(u_alu_lt_x_11_n92) );
  INV2 U2561 ( .A(n1398), .Q(n1086) );
  INV2 U2562 ( .A(n2445), .Q(n824) );
  INV2 U2563 ( .A(n1796), .Q(n1655) );
  NOR21 U2564 ( .A(n1143), .B(n1782), .Q(n1745) );
  NAND22 U2565 ( .A(n533), .B(n186), .Q(n2862) );
  INV2 U2566 ( .A(n2486), .Q(n2018) );
  NOR21 U2567 ( .A(u_alu_lt_x_11_B_16_), .B(n2445), .Q(n2831) );
  NAND22 U2568 ( .A(n1780), .B(n1695), .Q(n1697) );
  NAND22 U2569 ( .A(n1931), .B(n775), .Q(n774) );
  INV3 U2570 ( .A(n2980), .Q(n2599) );
  AOI210 U2571 ( .A(n1170), .B(u_alu_lt_x_11_B_17_), .C(n1972), .Q(n1612) );
  INV1 U2572 ( .A(n2107), .Q(n2075) );
  AOI221 U2573 ( .A(n369), .B(n3067), .C(n2671), .D(u_alu_lt_x_11_B_19_), .Q(
        n1606) );
  INV3 U2574 ( .A(n1790), .Q(n2094) );
  NOR22 U2575 ( .A(n2722), .B(n2812), .Q(n2819) );
  INV2 U2576 ( .A(u_alu_lt_x_11_n103), .Q(u_alu_lt_x_11_n101) );
  INV2 U2577 ( .A(n680), .Q(n3005) );
  INV1 U2578 ( .A(compare_i_data_rs[15]), .Q(u_alu_lt_x_11_n159) );
  NOR21 U2579 ( .A(n409), .B(n1931), .Q(n1856) );
  NAND22 U2580 ( .A(n2597), .B(n2596), .Q(n2980) );
  NAND22 U2581 ( .A(n680), .B(compare_i_data_rs[28]), .Q(
        u_alu_DP_OP_84J3_125_2615_n31) );
  INV2 U2582 ( .A(n384), .Q(n3116) );
  INV1 U2583 ( .A(u_alu_lt_x_11_B_20_), .Q(n2648) );
  NAND21 U2584 ( .A(n875), .B(n1954), .Q(n1955) );
  NAND21 U2585 ( .A(compare_i_data_rt[12]), .B(n139), .Q(n2251) );
  NAND21 U2586 ( .A(u_alu_lt_x_11_B_20_), .B(n1170), .Q(n946) );
  NAND22 U2587 ( .A(n2632), .B(n2618), .Q(n2725) );
  INV2 U2588 ( .A(compare_i_data_rs[19]), .Q(n443) );
  NAND22 U2589 ( .A(n1499), .B(n971), .Q(n511) );
  NAND21 U2590 ( .A(n374), .B(n2632), .Q(n2634) );
  INV3 U2591 ( .A(n679), .Q(n678) );
  NOR21 U2592 ( .A(n2247), .B(u_alu_lt_x_11_A_12_), .Q(n2252) );
  NAND21 U2593 ( .A(n1244), .B(n1805), .Q(n968) );
  NAND22 U2594 ( .A(n831), .B(n2559), .Q(n830) );
  NAND22 U2595 ( .A(n1476), .B(n2133), .Q(n2012) );
  NAND31 U2596 ( .A(n2474), .B(n2473), .C(n2472), .Q(n517) );
  OAI211 U2597 ( .A(i_data_immext[1]), .B(n391), .C(n1953), .Q(n1684) );
  INV3 U2598 ( .A(n488), .Q(n487) );
  INV1 U2599 ( .A(n1476), .Q(n2135) );
  OAI211 U2600 ( .A(n2249), .B(n2248), .C(n2429), .Q(n2250) );
  NAND41 U2601 ( .A(n1492), .B(n1491), .C(n1490), .D(n1404), .Q(n3189) );
  NAND22 U2602 ( .A(n398), .B(i_data_rs[2]), .Q(n1385) );
  NAND22 U2603 ( .A(n343), .B(i_data_rs[12]), .Q(n1267) );
  NAND22 U2604 ( .A(n1685), .B(n574), .Q(n723) );
  NAND21 U2605 ( .A(n1536), .B(n138), .Q(n1537) );
  NAND22 U2606 ( .A(n1161), .B(i_data_rt[7]), .Q(n1527) );
  NAND22 U2607 ( .A(n1161), .B(i_data_rt[6]), .Q(n1534) );
  NAND21 U2608 ( .A(n1719), .B(n391), .Q(n1720) );
  NAND22 U2609 ( .A(n1459), .B(n1458), .Q(n1460) );
  NOR21 U2610 ( .A(n1332), .B(n281), .Q(n1330) );
  NAND22 U2611 ( .A(n1136), .B(i_data_FMmemout[6]), .Q(n1531) );
  NAND22 U2612 ( .A(n1136), .B(i_data_FMmemout[7]), .Q(n1525) );
  NOR21 U2613 ( .A(n1286), .B(n353), .Q(n1287) );
  NAND22 U2614 ( .A(n1136), .B(i_data_FMmemout[21]), .Q(n1487) );
  INV2 U2615 ( .A(n2932), .Q(n2097) );
  NAND21 U2616 ( .A(n142), .B(i_data_FMmemout[2]), .Q(n1480) );
  NAND21 U2617 ( .A(n141), .B(i_data_FMmemout[28]), .Q(n1421) );
  NAND21 U2618 ( .A(n142), .B(i_data_FMmemout[24]), .Q(n1442) );
  NAND21 U2619 ( .A(n142), .B(i_data_FMmemout[22]), .Q(n1341) );
  NAND22 U2620 ( .A(n1134), .B(i_data_FMalures[3]), .Q(n1362) );
  NAND21 U2621 ( .A(n142), .B(i_data_FMmemout[29]), .Q(n1415) );
  NAND21 U2622 ( .A(n142), .B(i_data_FMmemout[20]), .Q(n1459) );
  NAND21 U2623 ( .A(n377), .B(n364), .Q(n674) );
  BUF15 U2624 ( .A(n1505), .Q(n1135) );
  NAND21 U2625 ( .A(n400), .B(n401), .Q(n819) );
  NAND22 U2626 ( .A(n410), .B(n361), .Q(n2641) );
  INV2 U2627 ( .A(n1526), .Q(n491) );
  INV2 U2628 ( .A(n2396), .Q(n1950) );
  INV2 U2629 ( .A(i_data_FWmemout[1]), .Q(n1300) );
  INV3 U2630 ( .A(i_data_FWmemout[30]), .Q(n1370) );
  INV2 U2631 ( .A(i_con_bop[1]), .Q(n1394) );
  INV2 U2632 ( .A(i_data_FEalures[14]), .Q(n1227) );
  INV2 U2633 ( .A(i_data_FWmemout[6]), .Q(n1207) );
  INV2 U2634 ( .A(i_data_FWmemout[20]), .Q(n1366) );
  INV2 U2635 ( .A(i_data_FWmemout[11]), .Q(n1294) );
  INV2 U2636 ( .A(i_data_FEalures[19]), .Q(n1324) );
  INV2 U2637 ( .A(i_data_FWmemout[19]), .Q(n1323) );
  INV2 U2638 ( .A(i_data_FWmemout[0]), .Q(n1281) );
  INV3 U2639 ( .A(i_data_FEalures[3]), .Q(n1361) );
  INV3 U2640 ( .A(i_data_FEalures[4]), .Q(n1203) );
  INV2 U2641 ( .A(i_data_FWmemout[13]), .Q(n1248) );
  INV2 U2642 ( .A(i_con_Ealuop[3]), .Q(n1579) );
  INV3 U2643 ( .A(i_data_FEalures[26]), .Q(n1384) );
  INV2 U2644 ( .A(i_con_Ealuop[2]), .Q(n1580) );
  INV2 U2645 ( .A(i_data_FEalures[21]), .Q(n1344) );
  INV2 U2646 ( .A(i_data_FWmemout[18]), .Q(n1316) );
  INV1 U2647 ( .A(i_con_bop[0]), .Q(n1311) );
  INV2 U2648 ( .A(i_data_FWmemout[2]), .Q(n1386) );
  XOR22 U2649 ( .A(n2783), .B(n2772), .Q(n569) );
  INV3 U2650 ( .A(i_data_FWmemout[27]), .Q(n1379) );
  NAND22 U2651 ( .A(n1234), .B(n460), .Q(n1235) );
  NAND23 U2652 ( .A(n1137), .B(i_data_FMmemout[27]), .Q(n1192) );
  OAI212 U2653 ( .A(n469), .B(u_alu_lt_x_11_n11), .C(u_alu_lt_x_11_n12), .Q(
        u_alu_lt_x_11_n10) );
  NAND22 U2654 ( .A(n143), .B(i_data_FMmemout[10]), .Q(n2134) );
  AOI222 U2655 ( .A(n2565), .B(n410), .C(n386), .D(n1864), .Q(n2058) );
  NOR31 U2656 ( .A(n2396), .B(n2395), .C(u_alu_lt_x_11_A_0_), .Q(n1921) );
  CLKIN6 U2657 ( .A(i_con_Efbmux[1]), .Q(n740) );
  AOI222 U2658 ( .A(i_data_FMmemout[20]), .B(n1137), .C(n338), .D(
        i_data_FWmemout[20]), .Q(n1492) );
  CLKIN6 U2659 ( .A(i_con_Efbmux[2]), .Q(n708) );
  INV12 U2660 ( .A(n740), .Q(n741) );
  NAND31 U2661 ( .A(n383), .B(i_data_rt[3]), .C(n391), .Q(n1721) );
  NAND24 U2662 ( .A(n2811), .B(n2819), .Q(n2817) );
  NAND28 U2663 ( .A(n2817), .B(n2816), .Q(n2823) );
  NOR21 U2664 ( .A(u_alu_lt_x_11_B_21_), .B(n450), .Q(u_alu_lt_x_11_n49) );
  NOR31 U2665 ( .A(n2136), .B(n1140), .C(n2135), .Q(n2137) );
  AOI211 U2666 ( .A(n3121), .B(n446), .C(n3021), .Q(n3022) );
  NOR21 U2667 ( .A(n407), .B(u_alu_lt_x_11_B_8_), .Q(u_alu_lt_x_11_n115) );
  NAND22 U2668 ( .A(n1135), .B(i_data_FMalures[27]), .Q(n1193) );
  AOI222 U2669 ( .A(n362), .B(n1865), .C(n1713), .D(n1167), .Q(n1794) );
  AOI2112 U2670 ( .A(n1080), .B(n2919), .C(n1079), .D(n2999), .Q(n1078) );
  XNR22 U2671 ( .A(n2916), .B(n2915), .Q(n2917) );
  NOR21 U2672 ( .A(n386), .B(n3104), .Q(n3112) );
  INV3 U2673 ( .A(n645), .Q(n644) );
  AOI212 U2674 ( .A(n850), .B(n1804), .C(n1803), .Q(n1821) );
  AOI212 U2675 ( .A(n2787), .B(n1155), .C(n2786), .Q(n2808) );
  NOR23 U2676 ( .A(n2918), .B(n657), .Q(n656) );
  NAND33 U2677 ( .A(n2809), .B(n2808), .C(n2807), .Q(alu_o_data_AluRes[23]) );
  NAND24 U2678 ( .A(n1137), .B(i_data_FMmemout[28]), .Q(n1321) );
  NOR21 U2679 ( .A(n1111), .B(n784), .Q(n801) );
  NOR20 U2680 ( .A(n442), .B(n387), .Q(u_alu_lt_x_11_n39) );
  NAND20 U2681 ( .A(u_alu_lt_x_11_B_1_), .B(n875), .Q(u_alu_lt_x_11_n142) );
  NAND20 U2682 ( .A(n369), .B(n418), .Q(u_alu_lt_x_11_n137) );
  NAND20 U2683 ( .A(u_alu_lt_x_11_B_5_), .B(n437), .Q(u_alu_lt_x_11_n130) );
  NAND20 U2684 ( .A(u_alu_lt_x_11_B_8_), .B(n407), .Q(u_alu_lt_x_11_n116) );
  NOR20 U2685 ( .A(n436), .B(u_alu_lt_x_11_B_9_), .Q(u_alu_lt_x_11_n108) );
  NAND20 U2686 ( .A(alu_i_data_B[31]), .B(n144), .Q(u_alu_lt_x_11_n6) );
  NOR21 U2687 ( .A(n144), .B(alu_i_data_B[31]), .Q(u_alu_lt_x_11_n5) );
  INV3 U2688 ( .A(u_alu_lt_x_11_n72), .Q(u_alu_lt_x_11_n70) );
  NAND20 U2689 ( .A(n371), .B(n439), .Q(u_alu_lt_x_11_n139) );
  NAND20 U2690 ( .A(n415), .B(u_alu_lt_x_11_B_17_), .Q(u_alu_lt_x_11_n73) );
  NAND22 U2691 ( .A(u_alu_DP_OP_84J3_125_2615_n145), .B(n434), .Q(n566) );
  NOR20 U2692 ( .A(n437), .B(u_alu_lt_x_11_B_5_), .Q(u_alu_lt_x_11_n129) );
  NOR20 U2693 ( .A(n439), .B(n371), .Q(u_alu_lt_x_11_n138) );
  XNR22 U2694 ( .A(n3059), .B(n3058), .Q(n647) );
  NAND22 U2695 ( .A(n1137), .B(i_data_FMmemout[30]), .Q(n1184) );
  INV3 U2696 ( .A(i_data_FWmemout[4]), .Q(n1202) );
  NOR24 U2697 ( .A(n2823), .B(n944), .Q(n3177) );
  AOI212 U2698 ( .A(u_alu_pre_sum_4a[4]), .B(n3078), .C(n915), .Q(n914) );
  NAND22 U2699 ( .A(n709), .B(i_con_Efbmux[0]), .Q(n1048) );
  CLKBU15 U2700 ( .A(n1545), .Q(n1136) );
  NAND34 U2701 ( .A(n1174), .B(n741), .C(n710), .Q(n1123) );
  CLKBU15 U2702 ( .A(n1505), .Q(n1134) );
  OAI212 U2703 ( .A(n1342), .B(n1159), .C(n1337), .Q(n1338) );
  INV15 U2704 ( .A(n724), .Q(n1160) );
  NAND26 U2705 ( .A(n1096), .B(n710), .Q(n724) );
  INV15 U2706 ( .A(n1160), .Q(n1159) );
  AOI211 U2707 ( .A(n413), .B(n3162), .C(n422), .Q(n3163) );
  OAI212 U2708 ( .A(n2413), .B(n2412), .C(n1923), .Q(n2420) );
  NAND28 U2709 ( .A(n2825), .B(n2824), .Q(n3128) );
  XNR22 U2710 ( .A(n2970), .B(n2967), .Q(n3000) );
  AOI212 U2711 ( .A(n977), .B(n2966), .C(n924), .Q(n2967) );
  NOR32 U2712 ( .A(n3052), .B(n3051), .C(n3050), .Q(n918) );
  NOR32 U2713 ( .A(n3049), .B(n3048), .C(n1149), .Q(n3050) );
  OAI212 U2714 ( .A(n1167), .B(n2058), .C(n1866), .Q(n1992) );
  AOI212 U2715 ( .A(n1155), .B(n2106), .C(n2105), .Q(n2163) );
  IMUX21 U2716 ( .A(n2993), .B(n2992), .S(u_alu_DP_OP_84J3_125_2615_n145), .Q(
        n2994) );
  AOI212 U2717 ( .A(n997), .B(n2958), .C(n994), .Q(n1000) );
  NOR32 U2718 ( .A(n3045), .B(n3044), .C(n3043), .Q(n3049) );
  NAND33 U2719 ( .A(n914), .B(n3053), .C(n918), .Q(alu_o_data_AluRes[28]) );
  AOI212 U2720 ( .A(n977), .B(n796), .C(n2914), .Q(n2915) );
  NOR33 U2721 ( .A(n709), .B(n741), .C(n710), .Q(n1505) );
  AOI212 U2722 ( .A(n362), .B(n2295), .C(n2059), .Q(n2176) );
  NAND33 U2723 ( .A(n1000), .B(n998), .C(n3179), .Q(alu_o_data_AluRes[31]) );
  NOR22 U2724 ( .A(n1168), .B(n1170), .Q(n3067) );
  AOI212 U2725 ( .A(n1165), .B(n2296), .C(n2177), .Q(n2237) );
  NOR33 U2726 ( .A(n1174), .B(i_con_Efbmux[0]), .C(n741), .Q(n1545) );
  INV12 U2727 ( .A(n709), .Q(n1174) );
  AOI2112 U2728 ( .A(n2959), .B(u_alu_pre_sum_4a[5]), .C(n648), .D(n643), .Q(
        n3076) );
  AOI212 U2729 ( .A(n2844), .B(n2845), .C(n2843), .Q(n925) );
  NAND24 U2730 ( .A(n1137), .B(i_data_FMmemout[14]), .Q(n1106) );
  NAND22 U2731 ( .A(n821), .B(n2834), .Q(n2839) );
  NOR24 U2732 ( .A(n926), .B(n925), .Q(n3088) );
  NAND33 U2733 ( .A(n2162), .B(n2163), .C(n2161), .Q(alu_o_data_AluRes[12]) );
  NAND42 U2734 ( .A(n1057), .B(n1056), .C(n3127), .D(n1059), .Q(
        alu_o_data_AluRes[30]) );
  NOR32 U2735 ( .A(n3128), .B(n3178), .C(n1146), .Q(n3078) );
  INV3 U2736 ( .A(i_con_Malupc8), .Q(n3203) );
  NOR21 U2737 ( .A(n2382), .B(n1763), .Q(n1732) );
  NOR31 U2738 ( .A(n445), .B(n1638), .C(n1626), .Q(n1591) );
  IMUX21 U2739 ( .A(n2015), .B(n2014), .S(n440), .Q(n2016) );
  NOR21 U2740 ( .A(n1920), .B(n2414), .Q(n1826) );
  NAND22 U2741 ( .A(n630), .B(n1846), .Q(n1817) );
  NAND22 U2742 ( .A(n1885), .B(n562), .Q(n1880) );
  AOI210 U2743 ( .A(n1946), .B(n386), .C(n1170), .Q(n1607) );
  OAI210 U2744 ( .A(n410), .B(n3106), .C(n458), .Q(n3111) );
  IMUX21 U2745 ( .A(n2650), .B(n2649), .S(n452), .Q(n2651) );
  AOI221 U2746 ( .A(n1870), .B(n362), .C(n1869), .D(n1167), .Q(n1974) );
  NAND22 U2747 ( .A(n2621), .B(n2625), .Q(n2519) );
  NAND22 U2748 ( .A(n2659), .B(n2658), .Q(n2588) );
  NAND22 U2749 ( .A(u_alu_lt_x_11_B_18_), .B(n2636), .Q(n2562) );
  NAND22 U2750 ( .A(n2845), .B(u_alu_lt_x_11_n50), .Q(n2702) );
  NAND22 U2751 ( .A(u_alu_lt_x_11_B_20_), .B(n374), .Q(n2691) );
  NAND22 U2752 ( .A(n2726), .B(n2727), .Q(n2693) );
  NOR31 U2753 ( .A(n2353), .B(n2352), .C(n2351), .Q(n2354) );
  INV3 U2754 ( .A(n2449), .Q(n2427) );
  INV3 U2755 ( .A(n897), .Q(n1092) );
  NAND22 U2756 ( .A(u_alu_lt_x_11_n100), .B(n2108), .Q(n2078) );
  INV3 U2757 ( .A(i_data_FWmemout[9]), .Q(n1352) );
  INV3 U2758 ( .A(i_data_FWmemout[22]), .Q(n1340) );
  INV3 U2759 ( .A(i_data_FWmemout[16]), .Q(n1504) );
  INV3 U2760 ( .A(i_data_FEalures[24]), .Q(n1346) );
  INV3 U2761 ( .A(i_data_rt[20]), .Q(n1494) );
  INV3 U2762 ( .A(i_data_FWmemout[28]), .Q(n1322) );
  AOI211 U2763 ( .A(n1170), .B(n3054), .C(n2673), .Q(n1828) );
  INV3 U2764 ( .A(i_data_FWmemout[17]), .Q(n1328) );
  INV3 U2765 ( .A(i_data_FEalures[17]), .Q(n1326) );
  INV3 U2766 ( .A(i_data_FEalures[31]), .Q(n1280) );
  AOI211 U2767 ( .A(n2963), .B(n1170), .C(n2598), .Q(n1753) );
  INV3 U2768 ( .A(i_data_FEalures[5]), .Q(n1286) );
  NAND22 U2769 ( .A(i_data_immext[11]), .B(n364), .Q(n2129) );
  INV3 U2770 ( .A(i_data_FWmemout[7]), .Q(n1232) );
  INV3 U2771 ( .A(i_data_FEalures[0]), .Q(n1282) );
  NOR21 U2772 ( .A(n1168), .B(n947), .Q(n1908) );
  NAND31 U2773 ( .A(n1123), .B(n739), .C(i_data_rt[2]), .Q(n753) );
  INV12 U2774 ( .A(n708), .Q(n709) );
  NAND41 U2775 ( .A(n1148), .B(i_con_Ealuop[2]), .C(i_con_Ealuop[3]), .D(n1556), .Q(n1557) );
  INV3 U2776 ( .A(i_data_FWmemout[26]), .Q(n1383) );
  INV3 U2777 ( .A(i_data_FWmemout[24]), .Q(n1349) );
  INV3 U2778 ( .A(i_data_FEalures[12]), .Q(n1262) );
  INV3 U2779 ( .A(i_data_FWmemout[31]), .Q(n1279) );
  INV3 U2780 ( .A(i_data_FWmemout[3]), .Q(n1363) );
  INV3 U2781 ( .A(i_data_FEalures[7]), .Q(n1233) );
  INV3 U2782 ( .A(i_data_FEalures[8]), .Q(n1307) );
  INV3 U2783 ( .A(i_data_FWmemout[8]), .Q(n1306) );
  INV3 U2784 ( .A(i_data_FEalures[6]), .Q(n1208) );
  INV3 U2785 ( .A(i_data_FEalures[15]), .Q(n1222) );
  NAND22 U2786 ( .A(n1160), .B(i_data_FEalures[1]), .Q(n1548) );
  NAND31 U2787 ( .A(n1099), .B(n1100), .C(i_data_rs[23]), .Q(n1331) );
  NOR21 U2788 ( .A(n3074), .B(n1872), .Q(n1873) );
  NAND22 U2789 ( .A(n2565), .B(n186), .Q(n2293) );
  NAND31 U2790 ( .A(n2150), .B(n2149), .C(n2148), .Q(n2152) );
  NOR21 U2791 ( .A(n365), .B(n2143), .Q(n2149) );
  NAND22 U2792 ( .A(n9), .B(i_data_FMalures[17]), .Q(n2464) );
  NAND22 U2793 ( .A(n1480), .B(n1479), .Q(n1481) );
  NAND22 U2794 ( .A(n1160), .B(i_data_FEalures[14]), .Q(n1109) );
  NAND22 U2795 ( .A(n1137), .B(i_data_FMmemout[29]), .Q(n1188) );
  NAND22 U2796 ( .A(n338), .B(i_data_FWmemout[11]), .Q(n989) );
  NAND22 U2797 ( .A(n1135), .B(i_data_FMalures[8]), .Q(n1268) );
  NAND22 U2798 ( .A(n1160), .B(i_data_FEalures[2]), .Q(n1540) );
  OAI2111 U2799 ( .A(n1165), .B(n2741), .C(n2798), .D(n400), .Q(n2742) );
  OAI212 U2800 ( .A(n426), .B(n2237), .C(n2183), .Q(n2184) );
  NAND31 U2801 ( .A(n2259), .B(n1155), .C(n1164), .Q(n2183) );
  IMUX21 U2802 ( .A(n2034), .B(n2033), .S(n1138), .Q(n2040) );
  NAND31 U2803 ( .A(u_alu_lt_x_11_B_9_), .B(n1170), .C(n386), .Q(n2898) );
  NAND20 U2804 ( .A(n146), .B(n441), .Q(n2681) );
  NAND22 U2805 ( .A(n1466), .B(n1465), .Q(n1467) );
  NAND41 U2806 ( .A(i_data_FMalures[23]), .B(n1098), .C(n604), .D(n494), .Q(
        n1446) );
  NOR31 U2807 ( .A(n1156), .B(n2078), .C(n2084), .Q(n2076) );
  NOR31 U2808 ( .A(n1736), .B(n1720), .C(n1735), .Q(n1724) );
  NAND31 U2809 ( .A(n1939), .B(n1938), .C(n1940), .Q(n1941) );
  NAND22 U2810 ( .A(n454), .B(i_data_FEalures[20]), .Q(n1491) );
  NAND22 U2811 ( .A(n1135), .B(i_data_FMalures[28]), .Q(n1320) );
  NAND22 U2812 ( .A(n1137), .B(i_data_FMmemout[9]), .Q(n1354) );
  NAND22 U2813 ( .A(n1137), .B(i_data_FMmemout[0]), .Q(n1276) );
  NAND31 U2814 ( .A(n393), .B(i_data_rt[10]), .C(n138), .Q(n1521) );
  NAND31 U2815 ( .A(n2259), .B(n1155), .C(n400), .Q(n2260) );
  NAND31 U2816 ( .A(n2737), .B(n2736), .C(n1163), .Q(n2743) );
  NAND31 U2817 ( .A(n3095), .B(n3094), .C(n400), .Q(n3114) );
  NAND22 U2818 ( .A(u_alu_lt_x_11_B_22_), .B(n1170), .Q(n1618) );
  NAND22 U2819 ( .A(n3176), .B(n3175), .Q(n996) );
  OAI212 U2820 ( .A(n400), .B(n2545), .C(n2544), .Q(n2548) );
  OAI212 U2821 ( .A(n3061), .B(n397), .C(n2977), .Q(n3032) );
  NAND22 U2822 ( .A(n2975), .B(n1167), .Q(n3061) );
  IMUX21 U2823 ( .A(n948), .B(n2159), .S(n1138), .Q(n2160) );
  NAND22 U2824 ( .A(n2703), .B(n458), .Q(n2737) );
  NOR21 U2825 ( .A(n1168), .B(n1617), .Q(n2264) );
  AOI211 U2826 ( .A(n2720), .B(n1874), .C(n2680), .Q(n2687) );
  NAND22 U2827 ( .A(n2864), .B(n401), .Q(n2798) );
  OAI2111 U2828 ( .A(i_con_Ealusrc), .B(compare_i_data_rt[13]), .C(n417), .D(
        n2429), .Q(n2430) );
  IMUX21 U2829 ( .A(n2072), .B(n2071), .S(n1138), .Q(n2089) );
  NAND22 U2830 ( .A(n9), .B(i_data_FMalures[10]), .Q(n2133) );
  NAND22 U2831 ( .A(n384), .B(n1170), .Q(n1616) );
  AOI311 U2832 ( .A(n391), .B(n382), .C(i_data_rt[14]), .D(n578), .Q(n577) );
  NAND22 U2833 ( .A(i_data_immext[14]), .B(n365), .Q(n2241) );
  OAI222 U2834 ( .A(n2793), .B(n386), .C(n1168), .D(n2714), .Q(n2295) );
  NOR21 U2835 ( .A(n1128), .B(n655), .Q(n1127) );
  NAND22 U2836 ( .A(n1136), .B(i_data_FMmemout[18]), .Q(n1498) );
  NAND22 U2837 ( .A(n1135), .B(i_data_FMalures[21]), .Q(n864) );
  OAI212 U2838 ( .A(n1389), .B(n1159), .C(n1181), .Q(n1182) );
  OAI212 U2839 ( .A(n1222), .B(n1159), .C(n1217), .Q(n1218) );
  NOR21 U2840 ( .A(n1333), .B(n1158), .Q(n1329) );
  NAND22 U2841 ( .A(n1135), .B(i_data_FMalures[9]), .Q(n1355) );
  NAND31 U2842 ( .A(n383), .B(n139), .C(i_data_rt[4]), .Q(n793) );
  OAI222 U2843 ( .A(n1794), .B(n1166), .C(n1714), .D(n1165), .Q(n1773) );
  AOI310 U2844 ( .A(n414), .B(n146), .C(n405), .D(n737), .Q(n736) );
  NAND31 U2845 ( .A(n2743), .B(n2742), .C(n378), .Q(n2750) );
  NOR31 U2846 ( .A(n1156), .B(n2328), .C(n2331), .Q(n2336) );
  AOI211 U2847 ( .A(n2327), .B(n2439), .C(u_alu_lt_x_11_n84), .Q(n1002) );
  AOI221 U2848 ( .A(n1770), .B(n397), .C(n1677), .D(n401), .Q(n1718) );
  OAI212 U2849 ( .A(n426), .B(n1802), .C(n1801), .Q(n1803) );
  AOI211 U2850 ( .A(n1836), .B(n1874), .C(n1800), .Q(n1801) );
  OAI222 U2851 ( .A(n1165), .B(n1794), .C(n1867), .D(n458), .Q(n1844) );
  OAI212 U2852 ( .A(n3074), .B(n3023), .C(n3022), .Q(n3052) );
  AOI210 U2853 ( .A(n413), .B(n2648), .C(n424), .Q(n2650) );
  NAND22 U2854 ( .A(n1993), .B(n1163), .Q(n1994) );
  AOI210 U2855 ( .A(n413), .B(n2490), .C(n424), .Q(n2492) );
  AOI211 U2856 ( .A(u_alu_pre_sum_4a[0]), .B(n3128), .C(n3178), .Q(n2826) );
  OAI212 U2857 ( .A(n2615), .B(n397), .C(n2543), .Q(n2570) );
  OAI212 U2858 ( .A(n362), .B(n2175), .C(n2174), .Q(n2296) );
  OAI212 U2859 ( .A(n410), .B(n3025), .C(n2173), .Q(n2501) );
  NAND31 U2860 ( .A(n2344), .B(n2154), .C(n436), .Q(n2155) );
  NAND22 U2861 ( .A(n2866), .B(n401), .Q(n2736) );
  OAI212 U2862 ( .A(n362), .B(n2567), .C(n2566), .Q(n2703) );
  OAI222 U2863 ( .A(n2942), .B(n386), .C(n3066), .D(n410), .Q(n2541) );
  OAI212 U2864 ( .A(n397), .B(n2647), .C(n2646), .Q(n2684) );
  AOI210 U2865 ( .A(n413), .B(n441), .C(n424), .Q(n2682) );
  OAI212 U2866 ( .A(n1167), .B(n2862), .C(n2614), .Q(n2796) );
  NAND22 U2867 ( .A(n3054), .B(n1171), .Q(n2942) );
  OAI222 U2868 ( .A(n362), .B(n2705), .C(n2889), .D(n1167), .Q(n2866) );
  OAI212 U2869 ( .A(n1914), .B(n3069), .C(n2674), .Q(n2894) );
  OAI212 U2870 ( .A(n410), .B(n2599), .C(n614), .Q(n2778) );
  OAI212 U2871 ( .A(u_alu_lt_x_11_A_12_), .B(n446), .C(n2227), .Q(n2351) );
  NAND31 U2872 ( .A(n2286), .B(n2364), .C(n2363), .Q(n620) );
  NAND22 U2873 ( .A(n2763), .B(u_alu_lt_x_11_A_23_), .Q(n2842) );
  OAI212 U2874 ( .A(n1935), .B(n7), .C(n437), .Q(n733) );
  OAI212 U2875 ( .A(n1172), .B(n1619), .C(n1695), .Q(n3184) );
  NAND22 U2876 ( .A(n343), .B(i_data_rs[0]), .Q(n1285) );
  NOR21 U2877 ( .A(n1281), .B(n220), .Q(n1284) );
  NAND22 U2878 ( .A(n2905), .B(n436), .Q(n2028) );
  NAND22 U2879 ( .A(n1137), .B(i_data_FMmemout[22]), .Q(n1336) );
  NOR21 U2880 ( .A(n1497), .B(n1496), .Q(n1499) );
  NOR21 U2881 ( .A(n1171), .B(n3005), .Q(n1791) );
  OAI222 U2882 ( .A(n1828), .B(n1168), .C(n3066), .D(n386), .Q(n2021) );
  OAI212 U2883 ( .A(n1221), .B(n941), .C(n1216), .Q(n1219) );
  NAND22 U2884 ( .A(n2092), .B(n1163), .Q(n2055) );
  OAI212 U2885 ( .A(n2052), .B(n1167), .C(n2051), .Q(n2181) );
  NAND22 U2886 ( .A(n3203), .B(n3200), .Q(o_addr_Erd[2]) );
  AOI2111 U2887 ( .A(n1748), .B(n423), .C(n1747), .D(n1746), .Q(n1749) );
  AOI211 U2888 ( .A(n1779), .B(n1778), .C(n1743), .Q(n1744) );
  AOI211 U2889 ( .A(n1730), .B(n1729), .C(n1728), .Q(n1731) );
  NOR21 U2890 ( .A(n1913), .B(n2415), .Q(n1783) );
  NAND22 U2891 ( .A(n814), .B(n1646), .Q(n598) );
  NOR21 U2892 ( .A(n818), .B(n815), .Q(n814) );
  NOR21 U2893 ( .A(n816), .B(n1615), .Q(n815) );
  NAND22 U2894 ( .A(n812), .B(n810), .Q(n818) );
  NAND22 U2895 ( .A(n307), .B(n600), .Q(n599) );
  NAND22 U2896 ( .A(u_alu_N306), .B(n602), .Q(n601) );
  NAND31 U2897 ( .A(n2827), .B(n2919), .C(u_alu_pre_sum_4b[1]), .Q(n660) );
  NAND22 U2898 ( .A(n1102), .B(n2921), .Q(n1144) );
  NAND22 U2899 ( .A(n928), .B(n796), .Q(n1102) );
  NAND22 U2900 ( .A(n3010), .B(n3014), .Q(n2916) );
  NAND22 U2901 ( .A(n1966), .B(n857), .Q(n1967) );
  AOI211 U2902 ( .A(n1964), .B(n407), .C(n858), .Q(n857) );
  NAND22 U2903 ( .A(n1912), .B(n2010), .Q(n1928) );
  OAI212 U2904 ( .A(n1164), .B(n1993), .C(n378), .Q(n1970) );
  NAND22 U2905 ( .A(n2273), .B(n2272), .Q(n2279) );
  INV3 U2906 ( .A(n2267), .Q(n2268) );
  OAI212 U2907 ( .A(n2238), .B(n2237), .C(n2236), .Q(n2239) );
  NAND22 U2908 ( .A(n2234), .B(n2439), .Q(n2267) );
  OAI212 U2909 ( .A(n2351), .B(n2230), .C(n2340), .Q(n2231) );
  AOI211 U2910 ( .A(n2765), .B(n2764), .C(n2766), .Q(n2755) );
  NAND31 U2911 ( .A(n2750), .B(n2749), .C(n2748), .Q(n2751) );
  NAND22 U2912 ( .A(n2732), .B(n2836), .Q(n2753) );
  NAND22 U2913 ( .A(n2770), .B(n2813), .Q(n2757) );
  NAND22 U2914 ( .A(n2219), .B(n2218), .Q(n2220) );
  NOR21 U2915 ( .A(u_alu_lt_x_11_n90), .B(n593), .Q(n2209) );
  NAND22 U2916 ( .A(u_alu_pre_sum_4a[2]), .B(n2959), .Q(n2960) );
  NAND22 U2917 ( .A(n1874), .B(n586), .Q(n962) );
  NAND22 U2918 ( .A(n2988), .B(n2987), .Q(n2936) );
  NAND22 U2919 ( .A(n2951), .B(n965), .Q(n964) );
  IMUX20 U2920 ( .A(n2950), .B(n2949), .S(n356), .Q(n2951) );
  AOI211 U2921 ( .A(n977), .B(n295), .C(n2965), .Q(n2922) );
  INV3 U2922 ( .A(n2955), .Q(n2923) );
  NAND22 U2923 ( .A(n2964), .B(n3008), .Q(n2955) );
  NAND22 U2924 ( .A(n2331), .B(n2330), .Q(n2332) );
  NAND22 U2925 ( .A(n1004), .B(n1002), .Q(n2331) );
  OAI212 U2926 ( .A(n593), .B(u_alu_lt_x_11_n92), .C(n1003), .Q(n2327) );
  NAND22 U2927 ( .A(n2326), .B(n2325), .Q(n1004) );
  AOI211 U2928 ( .A(n799), .B(n2361), .C(n2253), .Q(n2302) );
  NAND22 U2929 ( .A(n2045), .B(n1155), .Q(n2046) );
  INV3 U2930 ( .A(n2035), .Q(n2036) );
  NAND22 U2931 ( .A(n2156), .B(n2344), .Q(n2032) );
  NAND22 U2932 ( .A(n2037), .B(n423), .Q(n2017) );
  NAND22 U2933 ( .A(n2433), .B(n2107), .Q(n2037) );
  NAND31 U2934 ( .A(n1706), .B(n1705), .C(n1704), .Q(n1707) );
  NOR21 U2935 ( .A(n439), .B(n2531), .Q(n1728) );
  OAI222 U2936 ( .A(n1755), .B(n1166), .C(n1675), .D(n401), .Q(n1715) );
  NAND22 U2937 ( .A(u_alu_pre_sum_4a[6]), .B(n3078), .Q(n3127) );
  NAND22 U2938 ( .A(n3125), .B(n3124), .Q(n1058) );
  OAI212 U2939 ( .A(n3138), .B(n3085), .C(n3084), .Q(n3086) );
  INV3 U2940 ( .A(n3090), .Q(n3084) );
  NAND22 U2941 ( .A(n3044), .B(n3130), .Q(n1050) );
  INV3 U2942 ( .A(u_alu_lt_x_11_n8), .Q(n3079) );
  NOR21 U2943 ( .A(n1856), .B(n1958), .Q(n1850) );
  AOI211 U2944 ( .A(n1824), .B(n1879), .C(n1877), .Q(n1825) );
  AOI2111 U2945 ( .A(n1667), .B(n1155), .C(n1666), .D(n1665), .Q(n1668) );
  OAI2111 U2946 ( .A(n3178), .B(n1664), .C(n1663), .D(n1662), .Q(n1665) );
  NAND22 U2947 ( .A(n1677), .B(n458), .Q(n1656) );
  NOR21 U2948 ( .A(n394), .B(n1768), .Q(n1677) );
  NAND22 U2949 ( .A(n1716), .B(n458), .Q(n1678) );
  NOR21 U2950 ( .A(n394), .B(n1655), .Q(n1716) );
  OAI222 U2951 ( .A(n1653), .B(n1165), .C(n1714), .D(n397), .Q(n1676) );
  NAND22 U2952 ( .A(n947), .B(n946), .Q(n945) );
  INV3 U2953 ( .A(n1647), .Q(n1653) );
  NOR21 U2954 ( .A(n386), .B(n394), .Q(n932) );
  AOI221 U2955 ( .A(n1167), .B(n1614), .C(n1674), .D(n362), .Q(n1615) );
  NAND22 U2956 ( .A(n1818), .B(n404), .Q(n1819) );
  OAI212 U2957 ( .A(n1845), .B(n1859), .C(n1847), .Q(n1816) );
  AOI221 U2958 ( .A(n1770), .B(n401), .C(n1842), .D(n458), .Q(n1812) );
  NOR21 U2959 ( .A(n394), .B(n1841), .Q(n1770) );
  OAI212 U2960 ( .A(n2415), .B(n1876), .C(n911), .Q(n1810) );
  NAND22 U2961 ( .A(n1870), .B(n1167), .Q(n1797) );
  NAND22 U2962 ( .A(n935), .B(n410), .Q(n934) );
  OAI222 U2963 ( .A(n1755), .B(n1165), .C(n1827), .D(n458), .Q(n1804) );
  OAI222 U2964 ( .A(n1828), .B(n386), .C(n410), .D(n1613), .Q(n1674) );
  AOI211 U2965 ( .A(n1170), .B(u_alu_lt_x_11_B_21_), .C(n2178), .Q(n1613) );
  NAND22 U2966 ( .A(n1894), .B(n1893), .Q(n1895) );
  NOR21 U2967 ( .A(n1924), .B(n2948), .Q(n1890) );
  INV3 U2968 ( .A(n1882), .Q(n1887) );
  INV3 U2969 ( .A(n1880), .Q(n1889) );
  OAI212 U2970 ( .A(n911), .B(n1823), .C(n1915), .Q(n1877) );
  NAND22 U2971 ( .A(n912), .B(n1756), .Q(n911) );
  INV3 U2972 ( .A(n854), .Q(n853) );
  NAND22 U2973 ( .A(n1777), .B(n1778), .Q(n854) );
  INV3 U2974 ( .A(n1885), .Q(n1883) );
  NAND22 U2975 ( .A(n1919), .B(n1918), .Q(n1885) );
  AOI211 U2976 ( .A(n1874), .B(n1911), .C(n1873), .Q(n1899) );
  AOI221 U2977 ( .A(n1166), .B(n1910), .C(n1842), .D(n401), .Q(n1872) );
  OAI222 U2978 ( .A(n1769), .B(n362), .C(n1768), .D(n1041), .Q(n1842) );
  NAND22 U2979 ( .A(n2096), .B(n386), .Q(n1768) );
  AOI221 U2980 ( .A(n1973), .B(n1167), .C(n1796), .D(n362), .Q(n1871) );
  NOR21 U2981 ( .A(n1168), .B(n929), .Q(n1796) );
  NAND22 U2982 ( .A(n714), .B(n712), .Q(n1901) );
  NAND22 U2983 ( .A(n713), .B(n397), .Q(n712) );
  NAND22 U2984 ( .A(n1650), .B(n1651), .Q(n1793) );
  NAND22 U2985 ( .A(n1648), .B(n386), .Q(n1651) );
  NAND22 U2986 ( .A(n1992), .B(n396), .Q(n714) );
  OAI212 U2987 ( .A(n1847), .B(n2392), .C(n1846), .Q(n1857) );
  NAND22 U2988 ( .A(n625), .B(n628), .Q(n1847) );
  NAND22 U2989 ( .A(n1961), .B(n1766), .Q(n1848) );
  NOR31 U2990 ( .A(n419), .B(n1764), .C(n1660), .Q(n1765) );
  INV3 U2991 ( .A(n2389), .Q(n1845) );
  NAND22 U2992 ( .A(n999), .B(u_alu_pre_sum_4a[7]), .Q(n998) );
  INV3 U2993 ( .A(u_alu_DP_OP_84J3_125_2615_n15), .Q(
        u_alu_DP_OP_84J3_125_2615_n70) );
  INV3 U2994 ( .A(u_alu_DP_OP_84J3_125_2615_n14), .Q(
        u_alu_DP_OP_84J3_125_2615_n108) );
  INV3 U2995 ( .A(n1001), .Q(n999) );
  NAND22 U2996 ( .A(n1061), .B(n1073), .Q(n1001) );
  INV3 U2997 ( .A(n1076), .Q(n1073) );
  INV3 U2998 ( .A(n3174), .Q(n995) );
  NAND22 U2999 ( .A(n3172), .B(n3173), .Q(n3174) );
  OAI212 U3000 ( .A(n3112), .B(n3111), .C(n3110), .Q(n3155) );
  XOR21 U3001 ( .A(n3143), .B(n3139), .Q(n997) );
  OAI212 U3002 ( .A(n3138), .B(n3137), .C(n3136), .Q(n3139) );
  INV3 U3003 ( .A(n3140), .Q(n3136) );
  INV3 U3004 ( .A(n3047), .Q(n3043) );
  INV3 U3005 ( .A(n3046), .Q(n3045) );
  INV3 U3006 ( .A(n917), .Q(n916) );
  NAND22 U3007 ( .A(n3018), .B(n3046), .Q(n917) );
  NAND22 U3008 ( .A(n676), .B(n3081), .Q(n3046) );
  INV3 U3009 ( .A(n3016), .Q(n3018) );
  INV3 U3010 ( .A(n3131), .Q(n3042) );
  NAND22 U3011 ( .A(n2629), .B(n2630), .Q(n1030) );
  NAND22 U3012 ( .A(n2627), .B(n2907), .Q(n2630) );
  NAND22 U3013 ( .A(n2619), .B(n2691), .Q(n2661) );
  NAND22 U3014 ( .A(n2009), .B(n2008), .Q(alu_o_data_AluRes[9]) );
  NAND31 U3015 ( .A(n2005), .B(n2004), .C(n2003), .Q(n2006) );
  NOR21 U3016 ( .A(n2000), .B(n1999), .Q(n2004) );
  NAND31 U3017 ( .A(n1996), .B(n423), .C(n1995), .Q(n2005) );
  OAI222 U3018 ( .A(n2022), .B(n397), .C(n1906), .D(n401), .Q(n1993) );
  NOR21 U3019 ( .A(n186), .B(n2486), .Q(n1672) );
  OAI212 U3020 ( .A(n1168), .B(n1711), .C(n1710), .Q(n1865) );
  NAND22 U3021 ( .A(n1709), .B(n1168), .Q(n1710) );
  INV3 U3022 ( .A(n937), .Q(n1711) );
  NAND22 U3023 ( .A(u_alu_DP_OP_84J3_125_2615_n136), .B(n1170), .Q(n940) );
  OAI212 U3024 ( .A(n1996), .B(n1985), .C(n1984), .Q(n1986) );
  NOR21 U3025 ( .A(n1979), .B(n2030), .Q(n1980) );
  NOR21 U3026 ( .A(n2368), .B(n1977), .Q(n1978) );
  NAND31 U3027 ( .A(n1997), .B(n423), .C(n2010), .Q(n1985) );
  INV3 U3028 ( .A(n2052), .Q(n1869) );
  NOR21 U3029 ( .A(n1168), .B(n2049), .Q(n1870) );
  NOR21 U3030 ( .A(n401), .B(n2043), .Q(n1909) );
  OAI222 U3031 ( .A(n1841), .B(n1167), .C(n2042), .D(n362), .Q(n1910) );
  NAND22 U3032 ( .A(n2041), .B(n386), .Q(n1841) );
  INV3 U3033 ( .A(n3074), .Q(n2907) );
  XOR21 U3034 ( .A(n2519), .B(n2576), .Q(n570) );
  INV3 U3035 ( .A(n955), .Q(n2481) );
  XOR21 U3036 ( .A(n2514), .B(n2480), .Q(n571) );
  NAND22 U3037 ( .A(n2857), .B(n2854), .Q(n2505) );
  NAND22 U3038 ( .A(n1082), .B(n1078), .Q(alu_o_data_AluRes[27]) );
  NAND22 U3039 ( .A(n2827), .B(u_alu_pre_sum_4b[3]), .Q(n1081) );
  INV3 U3040 ( .A(n1074), .Q(n1083) );
  NAND22 U3041 ( .A(n1061), .B(n1075), .Q(n1074) );
  NAND22 U3042 ( .A(n3006), .B(n3012), .Q(n2970) );
  NAND22 U3043 ( .A(n2965), .B(n2964), .Q(n923) );
  OAI212 U3044 ( .A(n3001), .B(n2921), .C(n3014), .Q(n2965) );
  INV3 U3045 ( .A(n2969), .Q(n2966) );
  NAND22 U3046 ( .A(n295), .B(n2964), .Q(n2969) );
  INV3 U3047 ( .A(n3003), .Q(n2964) );
  AOI211 U3048 ( .A(n3121), .B(n471), .C(n2994), .Q(n2997) );
  OAI212 U3049 ( .A(n2888), .B(n2887), .C(n2886), .Q(alu_o_data_AluRes[24]) );
  INV3 U3050 ( .A(n2861), .Q(n2846) );
  INV3 U3051 ( .A(n2921), .Q(n2914) );
  NAND22 U3052 ( .A(n2849), .B(compare_i_data_rs[24]), .Q(n2921) );
  INV3 U3053 ( .A(n796), .Q(n3002) );
  OAI212 U3054 ( .A(u_alu_pre_sum_4a[0]), .B(n2827), .C(n2826), .Q(n2887) );
  OAI212 U3055 ( .A(n3077), .B(n573), .C(n3076), .Q(alu_o_data_AluRes[29]) );
  NOR21 U3056 ( .A(n2943), .B(n2942), .Q(n3035) );
  AOI211 U3057 ( .A(n3094), .B(n3095), .C(n2654), .Q(n1023) );
  NAND22 U3058 ( .A(n410), .B(n1170), .Q(n2896) );
  OAI212 U3059 ( .A(n2984), .B(n3147), .C(n2983), .Q(n2985) );
  INV3 U3060 ( .A(n3148), .Q(n2984) );
  NAND22 U3061 ( .A(n2980), .B(n410), .Q(n3148) );
  NAND22 U3062 ( .A(n1026), .B(n394), .Q(n1020) );
  NAND22 U3063 ( .A(u_alu_lt_x_11_n40), .B(n2840), .Q(n2841) );
  NOR21 U3064 ( .A(n451), .B(n2839), .Q(n2840) );
  NAND22 U3065 ( .A(n993), .B(n992), .Q(n991) );
  NAND22 U3066 ( .A(n2858), .B(n2857), .Q(n992) );
  INV3 U3067 ( .A(n673), .Q(n672) );
  NAND22 U3068 ( .A(n677), .B(n674), .Q(n673) );
  INV3 U3069 ( .A(n3013), .Q(n987) );
  NAND22 U3070 ( .A(n434), .B(u_alu_DP_OP_84J3_125_2615_n145), .Q(n3006) );
  INV3 U3071 ( .A(n3059), .Q(n650) );
  INV3 U3072 ( .A(u_alu_DP_OP_84J3_125_2615_n33), .Q(
        u_alu_DP_OP_84J3_125_2615_n32) );
  INV3 U3073 ( .A(n1422), .Q(n677) );
  NAND22 U3074 ( .A(n1425), .B(n675), .Q(n679) );
  NOR21 U3075 ( .A(n1424), .B(n1423), .Q(n675) );
  INV3 U3076 ( .A(u_alu_DP_OP_84J3_125_2615_n90), .Q(
        u_alu_DP_OP_84J3_125_2615_n89) );
  NAND22 U3077 ( .A(n2601), .B(n443), .Q(n808) );
  INV3 U3078 ( .A(n2562), .Q(n2582) );
  NOR21 U3079 ( .A(n2623), .B(n2622), .Q(n2576) );
  NOR21 U3080 ( .A(n2571), .B(n380), .Q(n2572) );
  OAI212 U3081 ( .A(n2705), .B(n1167), .C(n2502), .Q(n2568) );
  NAND22 U3082 ( .A(n2501), .B(n1167), .Q(n2502) );
  AOI211 U3083 ( .A(n2311), .B(n369), .C(n2310), .Q(n2312) );
  NAND22 U3084 ( .A(n2506), .B(n2855), .Q(n2448) );
  INV3 U3085 ( .A(n2831), .Q(n2506) );
  OAI212 U3086 ( .A(n1041), .B(n2405), .C(n2404), .Q(n2542) );
  AOI211 U3087 ( .A(n2612), .B(n386), .C(n2613), .Q(n2405) );
  OAI222 U3088 ( .A(n362), .B(n2520), .C(n1041), .D(n2265), .Q(n2400) );
  AOI211 U3089 ( .A(n2293), .B(n2567), .C(n1041), .Q(n2294) );
  NAND22 U3090 ( .A(n2518), .B(n2514), .Q(n2446) );
  NAND22 U3091 ( .A(n2160), .B(n404), .Q(n2161) );
  INV3 U3092 ( .A(n2142), .Q(n2158) );
  NAND22 U3093 ( .A(n2199), .B(n2198), .Q(n2142) );
  INV3 U3094 ( .A(n2169), .Q(n2199) );
  OAI212 U3095 ( .A(n2120), .B(n2119), .C(n2118), .Q(n2121) );
  OAI212 U3096 ( .A(n362), .B(n2398), .C(n2098), .Q(n2266) );
  AOI221 U3097 ( .A(n2640), .B(n2097), .C(n2096), .D(n2095), .Q(n2098) );
  INV3 U3098 ( .A(n1907), .Q(n2096) );
  NAND22 U3099 ( .A(n3105), .B(n1168), .Q(n2567) );
  AOI221 U3100 ( .A(n2541), .B(n1167), .C(n2540), .D(n362), .Q(n2615) );
  INV3 U3101 ( .A(n2796), .Q(n2741) );
  INV3 U3102 ( .A(n2943), .Q(n2611) );
  NAND22 U3103 ( .A(n2704), .B(n186), .Q(n2889) );
  NAND22 U3104 ( .A(n2500), .B(n186), .Q(n2705) );
  NAND22 U3105 ( .A(n1117), .B(n835), .Q(n1034) );
  INV3 U3106 ( .A(n2663), .Q(n2638) );
  NAND22 U3107 ( .A(n386), .B(n362), .Q(n2932) );
  NAND22 U3108 ( .A(n2644), .B(n2645), .Q(n2719) );
  AOI211 U3109 ( .A(n2643), .B(n362), .C(n2642), .Q(n2644) );
  OAI222 U3110 ( .A(n2676), .B(n362), .C(n2675), .D(n1167), .Q(n2779) );
  INV3 U3111 ( .A(n2894), .Q(n2676) );
  INV3 U3112 ( .A(n954), .Q(n2773) );
  NAND22 U3113 ( .A(n2698), .B(n569), .Q(n954) );
  OAI212 U3114 ( .A(n2782), .B(n2771), .C(n2781), .Q(n2772) );
  NAND22 U3115 ( .A(n2835), .B(n359), .Q(n2813) );
  NAND22 U3116 ( .A(u_alu_lt_x_11_B_21_), .B(compare_i_data_rs[21]), .Q(n2727)
         );
  NAND31 U3117 ( .A(n2726), .B(n2725), .C(n374), .Q(n2728) );
  NAND22 U3118 ( .A(u_alu_lt_x_11_B_19_), .B(compare_i_data_rs[19]), .Q(n2624)
         );
  INV3 U3119 ( .A(n1467), .Q(n1468) );
  OAI212 U3120 ( .A(n2356), .B(n2355), .C(n2354), .Q(n1008) );
  INV3 U3121 ( .A(n2429), .Q(n2197) );
  NAND22 U3122 ( .A(n2152), .B(n2151), .Q(n2153) );
  NOR21 U3123 ( .A(u_alu_lt_x_11_A_10_), .B(n2027), .Q(n2347) );
  NAND22 U3124 ( .A(n2344), .B(n430), .Q(n2356) );
  OAI222 U3125 ( .A(n844), .B(n2393), .C(n840), .D(n839), .Q(n1062) );
  NAND22 U3126 ( .A(n2138), .B(n2137), .Q(n2372) );
  NAND22 U3127 ( .A(n2130), .B(n2131), .Q(n622) );
  NAND22 U3128 ( .A(n2371), .B(n2370), .Q(n2378) );
  NOR31 U3129 ( .A(n2367), .B(n2369), .C(n2368), .Q(n2379) );
  INV3 U3130 ( .A(n2380), .Q(n841) );
  NAND22 U3131 ( .A(n843), .B(n2375), .Q(n842) );
  NOR21 U3132 ( .A(n2245), .B(n2244), .Q(n909) );
  INV3 U3133 ( .A(n620), .Q(n619) );
  NAND22 U3134 ( .A(n2366), .B(n2365), .Q(n843) );
  NAND22 U3135 ( .A(u_alu_lt_x_11_B_13_), .B(compare_i_data_rs[13]), .Q(n2365)
         );
  NAND22 U3136 ( .A(n799), .B(n2361), .Q(n2366) );
  INV3 U3137 ( .A(n629), .Q(n846) );
  NAND22 U3138 ( .A(n1776), .B(n1775), .Q(n2389) );
  OAI212 U3139 ( .A(n2789), .B(n2767), .C(n2788), .Q(n2768) );
  OAI212 U3140 ( .A(n2663), .B(n2662), .C(n2832), .Q(n2765) );
  NAND22 U3141 ( .A(n2829), .B(n2830), .Q(n2663) );
  NAND22 U3142 ( .A(n2764), .B(n2836), .Q(n2789) );
  NAND22 U3143 ( .A(n592), .B(n2426), .Q(n2449) );
  NAND22 U3144 ( .A(n2420), .B(n2419), .Q(n957) );
  INV3 U3145 ( .A(n2418), .Q(n958) );
  NAND22 U3146 ( .A(n417), .B(alu_i_data_B[13]), .Q(n972) );
  INV3 U3147 ( .A(n2435), .Q(n745) );
  NAND22 U3148 ( .A(n2110), .B(u_alu_lt_x_11_n100), .Q(n2437) );
  NAND22 U3149 ( .A(n1396), .B(n1395), .Q(n1397) );
  NAND31 U3150 ( .A(n1393), .B(i_con_bop[1]), .C(i_con_bop[2]), .Q(n1396) );
  AOI312 U3151 ( .A(n1093), .B(n1089), .C(n1087), .D(n1085), .Q(n1401) );
  INV3 U3152 ( .A(n1533), .Q(n767) );
  NAND22 U3153 ( .A(n1534), .B(n1531), .Q(n768) );
  NAND22 U3154 ( .A(n1014), .B(n1206), .Q(n1535) );
  NAND22 U3155 ( .A(n343), .B(i_data_rs[15]), .Q(n1225) );
  NAND22 U3156 ( .A(n2188), .B(n2191), .Q(n1247) );
  NAND22 U3157 ( .A(n398), .B(i_data_rs[13]), .Q(n1255) );
  NAND22 U3158 ( .A(n1251), .B(n1250), .Q(n1252) );
  NOR21 U3159 ( .A(n1249), .B(n353), .Q(n1253) );
  NAND22 U3160 ( .A(n1264), .B(n1263), .Q(n1265) );
  NAND22 U3161 ( .A(n383), .B(i_data_rt[12]), .Q(n1260) );
  NAND22 U3162 ( .A(n702), .B(n703), .Q(n701) );
  NOR21 U3163 ( .A(n1384), .B(n353), .Q(n1430) );
  INV3 U3164 ( .A(n1331), .Q(n1448) );
  OAI212 U3165 ( .A(n685), .B(n689), .C(n686), .Q(n684) );
  NAND22 U3166 ( .A(n688), .B(n1405), .Q(n687) );
  NAND22 U3167 ( .A(n1415), .B(n1414), .Q(n638) );
  NAND22 U3168 ( .A(n1373), .B(n1372), .Q(n1374) );
  NAND22 U3169 ( .A(n343), .B(i_data_rs[20]), .Q(n1463) );
  NAND22 U3170 ( .A(n398), .B(i_data_rs[28]), .Q(n1425) );
  NAND22 U3171 ( .A(n1939), .B(n1938), .Q(n867) );
  AOI211 U3172 ( .A(n2084), .B(n2083), .C(n2082), .Q(n2085) );
  NOR21 U3173 ( .A(n2079), .B(n1156), .Q(n2083) );
  INV3 U3174 ( .A(n2078), .Q(n2079) );
  NAND22 U3175 ( .A(n2077), .B(n2076), .Q(n2087) );
  INV3 U3176 ( .A(n2374), .Q(n1121) );
  NAND22 U3177 ( .A(n1946), .B(n358), .Q(n1918) );
  NAND31 U3178 ( .A(n771), .B(n1238), .C(n1930), .Q(n886) );
  NAND22 U3179 ( .A(n1916), .B(n1915), .Q(n1917) );
  NAND22 U3180 ( .A(n1914), .B(n1936), .Q(n1915) );
  NAND22 U3181 ( .A(n910), .B(n627), .Q(n1916) );
  NOR21 U3182 ( .A(n1960), .B(n625), .Q(n969) );
  NAND22 U3183 ( .A(n357), .B(n429), .Q(n652) );
  NOR21 U3184 ( .A(n1172), .B(n1619), .Q(n1696) );
  OAI212 U3185 ( .A(n2593), .B(n1724), .C(n1723), .Q(n1759) );
  INV3 U3186 ( .A(n2386), .Q(n1763) );
  NAND22 U3187 ( .A(n1948), .B(n1949), .Q(n1012) );
  NAND22 U3188 ( .A(alu_i_data_B[7]), .B(n358), .Q(n1949) );
  NAND31 U3189 ( .A(n1947), .B(n372), .C(n242), .Q(n1948) );
  NOR21 U3190 ( .A(n1203), .B(n352), .Q(n1205) );
  NAND22 U3191 ( .A(n382), .B(i_data_rt[4]), .Q(n1939) );
  INV3 U3192 ( .A(n1807), .Q(n735) );
  AOI211 U3193 ( .A(n357), .B(n1946), .C(n1932), .Q(n1945) );
  NAND22 U3194 ( .A(n343), .B(i_data_rs[6]), .Q(n1214) );
  AOI211 U3195 ( .A(n2031), .B(n2370), .C(n2030), .Q(n2067) );
  NAND22 U3196 ( .A(n2027), .B(u_alu_lt_x_11_A_10_), .Q(n2344) );
  NOR21 U3197 ( .A(n2369), .B(n2064), .Q(n2070) );
  NAND22 U3198 ( .A(n2374), .B(n406), .Q(n2350) );
  NAND22 U3199 ( .A(n398), .B(i_data_rs[11]), .Q(n1475) );
  OAI212 U3200 ( .A(n1371), .B(n1159), .C(n1185), .Q(n1186) );
  OAI212 U3201 ( .A(n1370), .B(n941), .C(n1184), .Q(n1187) );
  INV3 U3202 ( .A(n2241), .Q(n578) );
  INV3 U3203 ( .A(n580), .Q(n579) );
  NAND22 U3204 ( .A(n1512), .B(n139), .Q(n580) );
  OAI212 U3205 ( .A(n1340), .B(n941), .C(n1336), .Q(n1339) );
  INV3 U3206 ( .A(n1125), .Q(n970) );
  INV3 U3207 ( .A(n1318), .Q(n1496) );
  NOR21 U3208 ( .A(n1509), .B(n365), .Q(n1510) );
  INV3 U3209 ( .A(n1055), .Q(n1054) );
  OAI222 U3210 ( .A(n1792), .B(n1168), .C(n3025), .D(n386), .Q(n1990) );
  NOR21 U3211 ( .A(n1494), .B(n365), .Q(n1495) );
  INV3 U3212 ( .A(n1320), .Q(n1483) );
  INV3 U3213 ( .A(n1518), .Q(n2247) );
  NOR21 U3214 ( .A(n1517), .B(n365), .Q(n1519) );
  INV3 U3215 ( .A(i_data_FWmemout[12]), .Q(n1261) );
  INV3 U3216 ( .A(n1513), .Q(n1516) );
  NAND22 U3217 ( .A(i_data_immext[13]), .B(n364), .Q(n1514) );
  OAI212 U3218 ( .A(n1368), .B(n941), .C(n1188), .Q(n1191) );
  NAND22 U3219 ( .A(n2018), .B(n186), .Q(n2019) );
  NAND22 U3220 ( .A(u_alu_lt_x_11_B_17_), .B(n1171), .Q(n2486) );
  INV3 U3221 ( .A(n834), .Q(n833) );
  INV3 U3222 ( .A(i_data_FEalures[25]), .Q(n1389) );
  NAND22 U3223 ( .A(n393), .B(i_data_rt[25]), .Q(n1183) );
  OAI212 U3224 ( .A(n386), .B(n1904), .C(n1903), .Q(n2101) );
  INV3 U3225 ( .A(i_data_FWmemout[15]), .Q(n1221) );
  NAND22 U3226 ( .A(n382), .B(i_data_rt[15]), .Q(n1220) );
  INV3 U3227 ( .A(n1218), .Q(n862) );
  NAND22 U3228 ( .A(n393), .B(i_data_rt[23]), .Q(n1406) );
  INV3 U3229 ( .A(i_data_FWmemout[23]), .Q(n1332) );
  OAI222 U3230 ( .A(n1753), .B(n1168), .C(n1752), .D(n2776), .Q(n1905) );
  INV3 U3231 ( .A(n2897), .Q(n2776) );
  NOR21 U3232 ( .A(n386), .B(n1170), .Q(n2897) );
  NAND22 U3233 ( .A(u_alu_lt_x_11_B_1_), .B(n1171), .Q(n929) );
  INV3 U3234 ( .A(n1104), .Q(n1103) );
  INV3 U3235 ( .A(n1805), .Q(n1937) );
  NAND22 U3236 ( .A(n561), .B(n364), .Q(n1805) );
  INV3 U3237 ( .A(n2181), .Q(n2054) );
  NAND22 U3238 ( .A(n368), .B(n1171), .Q(n2049) );
  NAND22 U3239 ( .A(n2308), .B(n186), .Q(n2052) );
  NAND22 U3240 ( .A(n1526), .B(n364), .Q(n1930) );
  NAND22 U3241 ( .A(n365), .B(n394), .Q(n2146) );
  NAND22 U3242 ( .A(n1268), .B(n1269), .Q(n1270) );
  NOR21 U3243 ( .A(n1306), .B(n281), .Q(n1272) );
  NAND22 U3244 ( .A(u_alu_lt_x_11_B_0_), .B(n1171), .Q(n1907) );
  OAI212 U3245 ( .A(n1282), .B(n1159), .C(n1276), .Q(n1277) );
  NAND22 U3246 ( .A(n1135), .B(i_data_FMalures[0]), .Q(n1275) );
  NAND22 U3247 ( .A(n628), .B(n1171), .Q(n947) );
  INV3 U3248 ( .A(n727), .Q(n726) );
  INV3 U3249 ( .A(n729), .Q(n728) );
  NAND22 U3250 ( .A(n1537), .B(n1940), .Q(n1538) );
  OAI222 U3251 ( .A(n2265), .B(n362), .C(n2042), .D(n1167), .Q(n2099) );
  NAND22 U3252 ( .A(n860), .B(n386), .Q(n2042) );
  NAND22 U3253 ( .A(n1532), .B(n365), .Q(n1822) );
  NAND22 U3254 ( .A(n400), .B(n364), .Q(n1532) );
  AOI221 U3255 ( .A(n2521), .B(n386), .C(n2041), .D(n1168), .Q(n2265) );
  NAND22 U3256 ( .A(i_data_immext[2]), .B(n365), .Q(n1695) );
  INV3 U3257 ( .A(n753), .Q(n1541) );
  NAND22 U3258 ( .A(n338), .B(i_data_FWmemout[2]), .Q(n1539) );
  NAND22 U3259 ( .A(n1170), .B(n365), .Q(n2132) );
  INV3 U3260 ( .A(n1598), .Q(n1599) );
  NAND22 U3261 ( .A(n1582), .B(n1581), .Q(n1598) );
  NAND31 U3262 ( .A(n1580), .B(n1579), .C(n1148), .Q(n1581) );
  NAND22 U3263 ( .A(n1559), .B(n1072), .Q(n1071) );
  AOI311 U3264 ( .A(n1148), .B(n1580), .C(i_con_Ealuop[3]), .D(n1558), .Q(
        n1072) );
  INV3 U3265 ( .A(i_data_immext[2]), .Q(n1584) );
  INV3 U3266 ( .A(i_con_Ealuop[4]), .Q(n1556) );
  NAND22 U3267 ( .A(n1566), .B(n1565), .Q(n1567) );
  NAND22 U3268 ( .A(n1564), .B(n1573), .Q(n1566) );
  NAND22 U3269 ( .A(i_data_immext[2]), .B(i_data_immext[1]), .Q(n1573) );
  OAI212 U3270 ( .A(i_data_immext[4]), .B(n1571), .C(n715), .Q(n1587) );
  INV3 U3271 ( .A(n718), .Q(n717) );
  NAND22 U3272 ( .A(n1561), .B(i_data_immext[2]), .Q(n1560) );
  NOR21 U3273 ( .A(i_data_immext[1]), .B(i_data_immext[5]), .Q(n1553) );
  NAND22 U3274 ( .A(n383), .B(i_data_rt[14]), .Q(n2242) );
  XNR21 U3275 ( .A(n1745), .B(n1744), .Q(n1748) );
  XNR21 U3276 ( .A(n1732), .B(n1731), .Q(n1733) );
  XNR21 U3277 ( .A(n1767), .B(n1859), .Q(n1771) );
  XNR21 U3278 ( .A(u_alu_lt_x_11_A_0_), .B(n1660), .Q(n1641) );
  NOR20 U3279 ( .A(n401), .B(n1164), .Q(n817) );
  NOR30 U3280 ( .A(n819), .B(n394), .C(n379), .Q(n813) );
  OAI210 U3281 ( .A(n2640), .B(n1648), .C(n1168), .Q(n1621) );
  AOI220 U3282 ( .A(n1170), .B(u_alu_lt_x_11_B_16_), .C(u_alu_lt_x_11_B_0_), 
        .D(n1171), .Q(n1622) );
  NOR20 U3283 ( .A(n2905), .B(n3167), .Q(n737) );
  AOI210 U3284 ( .A(n413), .B(n405), .C(n424), .Q(n738) );
  IMUX20 U3285 ( .A(n425), .B(n1154), .S(compare_i_data_rs[25]), .Q(n2900) );
  NAND20 U3286 ( .A(n413), .B(n438), .Q(n859) );
  NOR20 U3287 ( .A(u_alu_lt_x_11_B_8_), .B(n2948), .Q(n1964) );
  IMUX20 U3288 ( .A(n425), .B(n1154), .S(n1039), .Q(n1965) );
  OAI210 U3289 ( .A(u_alu_lt_x_11_B_14_), .B(n425), .C(n1153), .Q(n2276) );
  XNR21 U3290 ( .A(n2256), .B(n2255), .Q(n2263) );
  NOR20 U3291 ( .A(n2267), .B(n1156), .Q(n2235) );
  XNR21 U3292 ( .A(n2232), .B(n2231), .Q(n2240) );
  XNR21 U3293 ( .A(n2756), .B(n2755), .Q(n2759) );
  NOR20 U3294 ( .A(n2835), .B(n2948), .Q(n2746) );
  OAI210 U3295 ( .A(n2835), .B(n425), .C(n1153), .Q(n2747) );
  IMUX20 U3296 ( .A(n413), .B(n376), .S(n359), .Q(n2744) );
  XNR21 U3297 ( .A(n2753), .B(n2735), .Q(n2752) );
  XNR21 U3298 ( .A(n2201), .B(n2200), .Q(n2208) );
  XNR21 U3299 ( .A(n2171), .B(n2170), .Q(n2185) );
  IMUX20 U3300 ( .A(n413), .B(n376), .S(n356), .Q(n2935) );
  OAI210 U3301 ( .A(u_alu_DP_OP_84J3_125_2615_n136), .B(n425), .C(n1153), .Q(
        n2949) );
  NOR20 U3302 ( .A(u_alu_DP_OP_84J3_125_2615_n136), .B(n2948), .Q(n2950) );
  XNR21 U3303 ( .A(n2923), .B(n2922), .Q(n2957) );
  XNR21 U3304 ( .A(n2032), .B(n2067), .Q(n2033) );
  XNR21 U3305 ( .A(n2032), .B(n2065), .Q(n2034) );
  XNR21 U3306 ( .A(n1727), .B(n1698), .Q(n1699) );
  XNR21 U3307 ( .A(n1779), .B(n1688), .Q(n1700) );
  NAND20 U3308 ( .A(n3121), .B(u_alu_lt_x_11_B_14_), .Q(n3122) );
  IMUX20 U3309 ( .A(n413), .B(n376), .S(compare_i_data_rs[30]), .Q(n3115) );
  XNR21 U3310 ( .A(n1850), .B(n1849), .Q(n1851) );
  NAND20 U3311 ( .A(n146), .B(n1931), .Q(n1833) );
  AOI210 U3312 ( .A(n413), .B(n1931), .C(n422), .Q(n1834) );
  XNR21 U3313 ( .A(n1826), .B(n1825), .Q(n1839) );
  OAI210 U3314 ( .A(u_alu_lt_x_11_B_1_), .B(n425), .C(n1153), .Q(n1659) );
  XNR21 U3315 ( .A(n1690), .B(n1657), .Q(n1664) );
  NAND20 U3316 ( .A(n386), .B(n1167), .Q(n933) );
  AOI210 U3317 ( .A(n1170), .B(u_alu_lt_x_11_B_18_), .C(n2041), .Q(n1620) );
  XNR21 U3318 ( .A(n1817), .B(n1816), .Q(n1818) );
  XNR21 U3319 ( .A(n1811), .B(n1810), .Q(n1814) );
  IMUX20 U3320 ( .A(n413), .B(n376), .S(n145), .Q(n3160) );
  NOR20 U3321 ( .A(n401), .B(n1167), .Q(n3096) );
  IMUX20 U3322 ( .A(n413), .B(n376), .S(compare_i_data_rs[28]), .Q(n3037) );
  XNR21 U3323 ( .A(n2664), .B(n2765), .Q(n2666) );
  XNR21 U3324 ( .A(n2661), .B(n2822), .Q(n2626) );
  XNR21 U3325 ( .A(n2661), .B(n2729), .Q(n2667) );
  XNR21 U3326 ( .A(n2664), .B(n2790), .Q(n2656) );
  IMUX20 U3327 ( .A(n413), .B(n376), .S(n416), .Q(n1998) );
  XNR21 U3328 ( .A(n2031), .B(n1980), .Q(n1981) );
  XNR21 U3329 ( .A(n2371), .B(n1978), .Q(n1982) );
  NOR20 U3330 ( .A(u_alu_lt_x_11_B_18_), .B(n2948), .Q(n2528) );
  XNR21 U3331 ( .A(n2519), .B(n2588), .Q(n2539) );
  XNR21 U3332 ( .A(n2546), .B(n2662), .Q(n2516) );
  XNR21 U3333 ( .A(n2506), .B(n2505), .Q(n2507) );
  XNR21 U3334 ( .A(n2518), .B(n2495), .Q(n2496) );
  XNR21 U3335 ( .A(n2855), .B(n2505), .Q(n2482) );
  NAND20 U3336 ( .A(n1165), .B(n1167), .Q(n589) );
  XNR21 U3337 ( .A(n2861), .B(n977), .Q(n2882) );
  AOI210 U3338 ( .A(n413), .B(n2849), .C(n424), .Q(n2850) );
  NAND20 U3339 ( .A(n146), .B(n2849), .Q(n2851) );
  OAI210 U3340 ( .A(n3054), .B(n425), .C(n1153), .Q(n3064) );
  NAND20 U3341 ( .A(n413), .B(n1752), .Q(n807) );
  NOR20 U3342 ( .A(u_alu_lt_x_11_B_19_), .B(n2948), .Q(n2601) );
  XNR21 U3343 ( .A(n2584), .B(n2583), .Q(n2585) );
  XNR21 U3344 ( .A(n2579), .B(n2578), .Q(n2587) );
  XNR21 U3345 ( .A(n2584), .B(n2563), .Q(n2573) );
  AOI210 U3346 ( .A(n413), .B(n1649), .C(n424), .Q(n2453) );
  NOR30 U3347 ( .A(n420), .B(n186), .C(n1167), .Q(n2311) );
  XNR21 U3348 ( .A(n2158), .B(n2289), .Q(n2159) );
  XNR21 U3349 ( .A(n2702), .B(n2701), .Q(n2710) );
  XNR21 U3350 ( .A(n2702), .B(n2694), .Q(n2695) );
  XNR21 U3351 ( .A(n2693), .B(n2692), .Q(n2697) );
  IMUX20 U3352 ( .A(n413), .B(n376), .S(compare_i_data_rs[21]), .Q(n2679) );
  XNR21 U3353 ( .A(n2693), .B(n2670), .Q(n2689) );
  OAI210 U3354 ( .A(n387), .B(n425), .C(n1153), .Q(n2802) );
  NOR20 U3355 ( .A(n387), .B(n2948), .Q(n2803) );
  IMUX20 U3356 ( .A(n413), .B(n376), .S(u_alu_lt_x_11_A_23_), .Q(n2801) );
  NOR20 U3357 ( .A(n377), .B(n1170), .Q(n2591) );
  NOR20 U3358 ( .A(n364), .B(n1170), .Q(n2592) );
  OAI2110 U3359 ( .A(n1017), .B(n3197), .C(n2897), .D(n1016), .Q(n1018) );
  NAND20 U3360 ( .A(n2364), .B(n364), .Q(n1016) );
  INV0 U3361 ( .A(n2364), .Q(n1017) );
  NAND30 U3362 ( .A(n383), .B(i_data_rt[13]), .C(n391), .Q(n2187) );
  NAND20 U3363 ( .A(n383), .B(i_data_rt[9]), .Q(n2148) );
  NOR20 U3364 ( .A(n139), .B(n410), .Q(n2144) );
  NAND30 U3365 ( .A(n2134), .B(n2133), .C(n2132), .Q(n2136) );
  OAI210 U3366 ( .A(n365), .B(n2242), .C(n2241), .Q(n2245) );
  XNR21 U3367 ( .A(n2792), .B(n2768), .Q(n2774) );
  INV3 U3368 ( .A(n867), .Q(n866) );
  INV3 U3369 ( .A(n1942), .Q(n868) );
  IMUX20 U3370 ( .A(n413), .B(n376), .S(n3185), .Q(n2080) );
  XNR21 U3371 ( .A(n2070), .B(n2069), .Q(n2071) );
  XNR21 U3372 ( .A(n2070), .B(n2066), .Q(n2072) );
  NAND22 U3373 ( .A(n383), .B(i_data_rt[28]), .Q(n1485) );
  NAND22 U3374 ( .A(n1135), .B(i_data_FMalures[5]), .Q(n1240) );
  NOR40 U3375 ( .A(i_data_immext[1]), .B(n1584), .C(n1565), .D(n1585), .Q(
        n1558) );
  XNR21 U3376 ( .A(u_alu_DP_OP_84J3_125_2615_n50), .B(
        u_alu_DP_OP_84J3_125_2615_n7), .Q(n568) );
  XNR21 U3377 ( .A(u_alu_DP_OP_84J3_125_2615_n3), .B(
        u_alu_DP_OP_84J3_125_2615_n80), .Q(n573) );
  AOI210 U3378 ( .A(n1171), .B(n253), .C(n3144), .Q(n3146) );
  AOI210 U3379 ( .A(n1883), .B(n1920), .C(n1156), .Q(n1884) );
  NAND22 U3380 ( .A(n3203), .B(n3202), .Q(o_addr_Erd[4]) );
  XNR21 U3381 ( .A(n407), .B(u_alu_lt_x_11_B_8_), .Q(n1963) );
  XNR21 U3382 ( .A(n145), .B(alu_i_data_B[31]), .Q(n3143) );
  XNR21 U3383 ( .A(n1928), .B(n2202), .Q(n1969) );
  NAND22 U3384 ( .A(n3203), .B(n3198), .Q(o_addr_Erd[0]) );
  NAND22 U3385 ( .A(n3203), .B(n3201), .Q(o_addr_Erd[3]) );
  NAND22 U3386 ( .A(n3203), .B(n3199), .Q(o_addr_Erd[1]) );
  XNR21 U3387 ( .A(n2916), .B(n1144), .Q(n2912) );
  IMUX20 U3388 ( .A(i_addr_rt[0]), .B(i_data_immext[11]), .S(i_con_Eregdst), 
        .Q(n3198) );
  IMUX20 U3389 ( .A(i_addr_rt[1]), .B(i_data_immext[12]), .S(i_con_Eregdst), 
        .Q(n3199) );
  IMUX20 U3390 ( .A(i_addr_rt[3]), .B(i_data_immext[14]), .S(i_con_Eregdst), 
        .Q(n3201) );
  IMUX20 U3391 ( .A(i_addr_rt[4]), .B(i_data_immext[15]), .S(i_con_Eregdst), 
        .Q(n3202) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_con_RegWr, i_addr_Rd, 
        i_data_Rd, o_data_Rs, o_data_Rt, i_addr_Rt_4_, i_addr_Rt_3_, 
        i_addr_Rt_2_, i_addr_Rt_1_, i_addr_Rt_0_ );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr, i_addr_Rt_4_, i_addr_Rt_3_, i_addr_Rt_2_,
         i_addr_Rt_1_, i_addr_Rt_0_;
  wire   n5, n6, n9, n11, n13, n15, n16, n17, n18, n20, n21, n22, n23, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n1, n2, n3, n4, n7, n8, n10, n12, n14, n19, n24,
         n33, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823;
  wire   [1023:0] regs;

  DFEC1 regs_reg_31__31_ ( .D(n262), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1023]) );
  DFEC1 regs_reg_31__30_ ( .D(n260), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(n258), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(n256), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(n254), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(n252), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(n250), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(n248), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(n246), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(n244), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(n242), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(n240), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(n238), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(n236), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(n234), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(n232), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(n230), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(n228), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(n226), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(n224), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(n222), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(n220), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(n218), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(n216), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(n214), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(n212), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(n210), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(n208), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(n206), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(n204), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(n202), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(n200), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[992]) );
  DFEC1 regs_reg_30__31_ ( .D(n262), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(n260), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(n258), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(n256), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(n254), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(n252), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(n250), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(n248), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(n246), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(n244), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(n242), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(n240), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(n238), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(n236), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(n234), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(n232), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(n230), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(n228), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(n226), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(n224), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(n222), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(n220), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(n218), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(n216), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(n214), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(n212), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(n210), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(n208), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(n206), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(n204), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(n202), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(n200), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[960]) );
  DFEC1 regs_reg_29__31_ ( .D(n262), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[959]), .QN(n191) );
  DFEC1 regs_reg_29__30_ ( .D(n260), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[958]), .QN(n188) );
  DFEC1 regs_reg_29__29_ ( .D(n258), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[957]), .QN(n185) );
  DFEC1 regs_reg_29__28_ ( .D(n256), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[956]), .QN(n182) );
  DFEC1 regs_reg_29__27_ ( .D(n254), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[955]), .QN(n179) );
  DFEC1 regs_reg_29__26_ ( .D(n252), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[954]), .QN(n176) );
  DFEC1 regs_reg_29__25_ ( .D(n250), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[953]), .QN(n173) );
  DFEC1 regs_reg_29__24_ ( .D(n248), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[952]), .QN(n170) );
  DFEC1 regs_reg_29__23_ ( .D(n246), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[951]), .QN(n167) );
  DFEC1 regs_reg_29__22_ ( .D(n244), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[950]), .QN(n164) );
  DFEC1 regs_reg_29__21_ ( .D(n242), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[949]), .QN(n110) );
  DFEC1 regs_reg_29__20_ ( .D(n240), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[948]), .QN(n108) );
  DFEC1 regs_reg_29__19_ ( .D(n238), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[947]), .QN(n106) );
  DFEC1 regs_reg_29__18_ ( .D(n236), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[946]), .QN(n104) );
  DFEC1 regs_reg_29__17_ ( .D(n234), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[945]), .QN(n102) );
  DFEC1 regs_reg_29__16_ ( .D(n232), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[944]), .QN(n100) );
  DFEC1 regs_reg_29__15_ ( .D(n230), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[943]), .QN(n98) );
  DFEC1 regs_reg_29__14_ ( .D(n228), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[942]), .QN(n96) );
  DFEC1 regs_reg_29__13_ ( .D(n226), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[941]), .QN(n94) );
  DFEC1 regs_reg_29__12_ ( .D(n224), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[940]), .QN(n92) );
  DFEC1 regs_reg_29__11_ ( .D(n222), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[939]), .QN(n90) );
  DFEC1 regs_reg_29__10_ ( .D(n220), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[938]), .QN(n88) );
  DFEC1 regs_reg_29__9_ ( .D(n218), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[937]), .QN(n86) );
  DFEC1 regs_reg_29__8_ ( .D(n216), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[936]), .QN(n84) );
  DFEC1 regs_reg_29__7_ ( .D(n214), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[935]), .QN(n82) );
  DFEC1 regs_reg_29__6_ ( .D(n212), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[934]), .QN(n80) );
  DFEC1 regs_reg_29__5_ ( .D(n210), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[933]), .QN(n78) );
  DFEC1 regs_reg_29__4_ ( .D(n208), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[932]), .QN(n76) );
  DFEC1 regs_reg_29__3_ ( .D(n206), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[931]), .QN(n74) );
  DFEC1 regs_reg_29__2_ ( .D(n204), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[930]), .QN(n72) );
  DFEC1 regs_reg_29__1_ ( .D(n202), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[929]), .QN(n67) );
  DFEC1 regs_reg_29__0_ ( .D(n200), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[928]), .QN(n121) );
  DFEC1 regs_reg_28__31_ ( .D(n262), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(n260), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(n258), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(n256), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(n254), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(n252), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(n250), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(n248), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(n246), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(n244), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(n242), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(n240), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(n238), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(n236), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(n234), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(n232), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(n230), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(n228), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(n226), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(n224), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(n222), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(n220), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(n218), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(n216), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(n214), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(n212), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(n210), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(n208), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(n206), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(n204), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(n202), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(n200), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(n262), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(n260), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(n258), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(n256), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(n254), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(n252), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(n250), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(n248), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(n246), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(n244), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(n242), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(n240), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(n238), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(n236), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(n234), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(n232), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(n230), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(n228), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(n226), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(n224), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(n222), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(n220), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(n218), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(n216), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(n214), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(n212), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(n210), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(n208), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(n206), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(n204), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(n202), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(n200), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[864]) );
  DFEC1 regs_reg_26__31_ ( .D(n262), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(n260), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(n258), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(n256), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(n254), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(n252), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(n250), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(n248), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(n246), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(n244), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(n242), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(n240), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(n238), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(n236), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(n234), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(n232), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(n230), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(n228), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(n226), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(n224), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(n222), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(n220), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(n218), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(n216), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(n214), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(n212), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(n210), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(n208), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(n206), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(n204), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(n202), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(n200), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[832]) );
  DFEC1 regs_reg_25__31_ ( .D(n262), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(n260), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(n258), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(n256), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(n254), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(n252), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(n250), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(n248), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(n246), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(n244), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(n242), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(n240), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(n238), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(n236), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(n234), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(n232), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(n230), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(n228), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(n226), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(n224), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(n222), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(n220), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(n218), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(n216), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(n214), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(n212), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(n210), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(n208), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(n206), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(n204), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(n202), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(n200), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[800]) );
  DFEC1 regs_reg_24__31_ ( .D(n262), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(n260), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(n258), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(n256), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(n254), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(n252), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(n250), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(n248), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(n246), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(n244), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(n242), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(n240), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(n238), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(n236), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(n234), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(n232), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(n230), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(n228), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(n226), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(n224), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(n222), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(n220), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(n218), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(n216), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(n214), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(n212), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(n210), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(n208), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(n206), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(n204), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(n202), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(n200), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(n263), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(n261), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(n259), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(n257), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(n255), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(n253), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(n251), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(n249), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(n247), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(n245), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(n243), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(n241), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(n239), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(n237), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(n235), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(n233), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(n231), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(n229), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(n227), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(n225), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(n223), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(n221), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(n219), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(n217), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(n215), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(n213), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(n211), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(n209), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(n207), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(n205), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(n203), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(n201), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[736]) );
  DFEC1 regs_reg_22__31_ ( .D(n262), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(n260), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(n258), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(n256), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(n254), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(n252), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(n250), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(n248), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(n246), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(n244), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(n242), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(n240), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(n238), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(n236), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(n234), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(n232), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(n230), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(n228), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(n226), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(n224), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(n222), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(n220), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(n218), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(n216), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(n214), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(n212), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(n210), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(n208), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(n206), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(n204), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(n202), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(n200), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[704]) );
  DFEC1 regs_reg_21__31_ ( .D(n263), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[703]), .QN(n193) );
  DFEC1 regs_reg_21__30_ ( .D(n261), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[702]), .QN(n190) );
  DFEC1 regs_reg_21__29_ ( .D(n259), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[701]), .QN(n187) );
  DFEC1 regs_reg_21__28_ ( .D(n257), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[700]), .QN(n184) );
  DFEC1 regs_reg_21__27_ ( .D(n255), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[699]), .QN(n181) );
  DFEC1 regs_reg_21__26_ ( .D(n253), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[698]), .QN(n178) );
  DFEC1 regs_reg_21__25_ ( .D(n251), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[697]), .QN(n175) );
  DFEC1 regs_reg_21__24_ ( .D(n249), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[696]), .QN(n172) );
  DFEC1 regs_reg_21__23_ ( .D(n247), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[695]), .QN(n169) );
  DFEC1 regs_reg_21__22_ ( .D(n245), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[694]), .QN(n166) );
  DFEC1 regs_reg_21__21_ ( .D(n243), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[693]), .QN(n163) );
  DFEC1 regs_reg_21__20_ ( .D(n241), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[692]), .QN(n161) );
  DFEC1 regs_reg_21__19_ ( .D(n239), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[691]), .QN(n159) );
  DFEC1 regs_reg_21__18_ ( .D(n237), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[690]), .QN(n157) );
  DFEC1 regs_reg_21__17_ ( .D(n235), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[689]), .QN(n155) );
  DFEC1 regs_reg_21__16_ ( .D(n233), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[688]), .QN(n153) );
  DFEC1 regs_reg_21__15_ ( .D(n231), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[687]), .QN(n151) );
  DFEC1 regs_reg_21__14_ ( .D(n229), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[686]), .QN(n149) );
  DFEC1 regs_reg_21__13_ ( .D(n227), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[685]), .QN(n147) );
  DFEC1 regs_reg_21__12_ ( .D(n225), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[684]), .QN(n145) );
  DFEC1 regs_reg_21__11_ ( .D(n223), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[683]), .QN(n143) );
  DFEC1 regs_reg_21__10_ ( .D(n221), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[682]), .QN(n141) );
  DFEC1 regs_reg_21__9_ ( .D(n219), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[681]), .QN(n139) );
  DFEC1 regs_reg_21__8_ ( .D(n217), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[680]), .QN(n137) );
  DFEC1 regs_reg_21__7_ ( .D(n215), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[679]), .QN(n135) );
  DFEC1 regs_reg_21__6_ ( .D(n213), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[678]), .QN(n133) );
  DFEC1 regs_reg_21__5_ ( .D(n211), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[677]), .QN(n131) );
  DFEC1 regs_reg_21__4_ ( .D(n209), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[676]), .QN(n129) );
  DFEC1 regs_reg_21__3_ ( .D(n207), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[675]), .QN(n127) );
  DFEC1 regs_reg_21__2_ ( .D(n205), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[674]), .QN(n125) );
  DFEC1 regs_reg_21__1_ ( .D(n203), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[673]), .QN(n69) );
  DFEC1 regs_reg_21__0_ ( .D(n201), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[672]), .QN(n194) );
  DFEC1 regs_reg_20__31_ ( .D(n263), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(n261), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(n259), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(n257), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(n255), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(n253), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(n251), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(n249), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(n247), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(n245), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(n243), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(n241), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(n239), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(n237), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(n235), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(n233), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(n231), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(n229), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(n227), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(n225), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(n223), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(n221), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(n219), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(n217), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(n215), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(n213), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(n211), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(n209), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(n207), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(n205), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(n203), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(n201), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(n262), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(n260), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(n258), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(n256), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(n254), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(n252), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(n250), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(n248), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(n246), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(n244), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(n242), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(n240), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(n238), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(n236), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(n234), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(n232), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(n230), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(n228), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(n226), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(n224), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(n222), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(n220), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(n218), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(n216), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(n214), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(n212), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(n210), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(n208), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(n206), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(n204), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(n202), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(n200), .E(n63), .C(i_clk), .RN(i_rst_n), .Q(
        regs[608]) );
  DFEC1 regs_reg_18__31_ ( .D(n262), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(n260), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(n258), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(n256), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(n254), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(n252), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(n250), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(n248), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(n246), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(n244), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(n242), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(n240), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(n238), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(n236), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(n234), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(n232), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(n230), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(n228), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(n226), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(n224), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(n222), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(n220), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(n218), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(n216), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(n214), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(n212), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(n210), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(n208), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(n206), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(n204), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(n202), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(n200), .E(n64), .C(i_clk), .RN(i_rst_n), .Q(
        regs[576]) );
  DFEC1 regs_reg_17__31_ ( .D(n263), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(n261), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(n259), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(n257), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(n255), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(n253), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(n251), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(n249), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(n247), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(n245), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(n243), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(n241), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(n239), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(n237), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(n235), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(n233), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(n231), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(n229), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(n227), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(n225), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(n223), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(n221), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(n219), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(n217), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(n215), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(n213), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(n211), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(n209), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(n207), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(n205), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(n203), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(n201), .E(n61), .C(i_clk), .RN(i_rst_n), .Q(
        regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(n262), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(n260), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(n258), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(n256), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(n254), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(n252), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(n250), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(n248), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(n246), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(n244), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(n242), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(n240), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(n238), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(n236), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(n234), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(n232), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(n230), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(n228), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(n226), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(n224), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(n222), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(n220), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(n218), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(n216), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(n214), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(n212), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(n210), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(n208), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(n206), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(n204), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(n202), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(n200), .E(n62), .C(i_clk), .RN(i_rst_n), .Q(
        regs[512]) );
  DFEC1 regs_reg_15__31_ ( .D(i_data_Rd[31]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(i_data_Rd[30]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(i_data_Rd[29]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(i_data_Rd[28]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(i_data_Rd[27]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(i_data_Rd[26]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(i_data_Rd[25]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(i_data_Rd[24]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(i_data_Rd[23]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(i_data_Rd[22]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(i_data_Rd[21]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(i_data_Rd[20]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(i_data_Rd[19]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(i_data_Rd[18]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(i_data_Rd[17]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(i_data_Rd[16]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(i_data_Rd[15]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(i_data_Rd[13]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(i_data_Rd[12]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(i_data_Rd[11]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(i_data_Rd[9]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(i_data_Rd[8]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(i_data_Rd[7]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(i_data_Rd[6]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(i_data_Rd[5]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(i_data_Rd[4]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(i_data_Rd[3]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(i_data_Rd[2]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(i_data_Rd[1]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(i_data_Rd[0]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[480]) );
  DFEC1 regs_reg_14__31_ ( .D(i_data_Rd[31]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(i_data_Rd[30]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(i_data_Rd[29]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(i_data_Rd[28]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(i_data_Rd[27]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(i_data_Rd[26]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(i_data_Rd[25]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(i_data_Rd[24]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(i_data_Rd[23]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(i_data_Rd[22]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(i_data_Rd[21]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(i_data_Rd[20]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(i_data_Rd[19]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(i_data_Rd[18]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(i_data_Rd[17]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(i_data_Rd[16]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(i_data_Rd[15]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(i_data_Rd[13]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(i_data_Rd[12]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(i_data_Rd[11]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(i_data_Rd[9]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(i_data_Rd[8]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(i_data_Rd[7]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(i_data_Rd[6]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(i_data_Rd[5]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(i_data_Rd[4]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(i_data_Rd[3]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(i_data_Rd[2]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(i_data_Rd[1]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(i_data_Rd[0]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[448]) );
  DFEC1 regs_reg_13__31_ ( .D(i_data_Rd[31]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[447]), .QN(n120) );
  DFEC1 regs_reg_13__30_ ( .D(i_data_Rd[30]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[446]), .QN(n119) );
  DFEC1 regs_reg_13__29_ ( .D(i_data_Rd[29]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[445]), .QN(n118) );
  DFEC1 regs_reg_13__28_ ( .D(i_data_Rd[28]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[444]), .QN(n117) );
  DFEC1 regs_reg_13__27_ ( .D(i_data_Rd[27]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[443]), .QN(n116) );
  DFEC1 regs_reg_13__26_ ( .D(i_data_Rd[26]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[442]), .QN(n115) );
  DFEC1 regs_reg_13__25_ ( .D(i_data_Rd[25]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[441]), .QN(n114) );
  DFEC1 regs_reg_13__24_ ( .D(i_data_Rd[24]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[440]), .QN(n113) );
  DFEC1 regs_reg_13__23_ ( .D(i_data_Rd[23]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[439]), .QN(n112) );
  DFEC1 regs_reg_13__22_ ( .D(i_data_Rd[22]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[438]), .QN(n111) );
  DFEC1 regs_reg_13__21_ ( .D(i_data_Rd[21]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[437]), .QN(n109) );
  DFEC1 regs_reg_13__20_ ( .D(i_data_Rd[20]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[436]), .QN(n107) );
  DFEC1 regs_reg_13__19_ ( .D(i_data_Rd[19]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[435]), .QN(n105) );
  DFEC1 regs_reg_13__18_ ( .D(i_data_Rd[18]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[434]), .QN(n103) );
  DFEC1 regs_reg_13__17_ ( .D(i_data_Rd[17]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[433]), .QN(n101) );
  DFEC1 regs_reg_13__16_ ( .D(i_data_Rd[16]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[432]), .QN(n99) );
  DFEC1 regs_reg_13__15_ ( .D(i_data_Rd[15]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[431]), .QN(n97) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[430]), .QN(n95) );
  DFEC1 regs_reg_13__13_ ( .D(i_data_Rd[13]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[429]), .QN(n93) );
  DFEC1 regs_reg_13__12_ ( .D(i_data_Rd[12]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[428]), .QN(n91) );
  DFEC1 regs_reg_13__11_ ( .D(i_data_Rd[11]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[427]), .QN(n89) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[426]), .QN(n87) );
  DFEC1 regs_reg_13__9_ ( .D(i_data_Rd[9]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[425]), .QN(n85) );
  DFEC1 regs_reg_13__8_ ( .D(i_data_Rd[8]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[424]), .QN(n83) );
  DFEC1 regs_reg_13__7_ ( .D(i_data_Rd[7]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[423]), .QN(n81) );
  DFEC1 regs_reg_13__6_ ( .D(i_data_Rd[6]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[422]), .QN(n79) );
  DFEC1 regs_reg_13__5_ ( .D(i_data_Rd[5]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[421]), .QN(n77) );
  DFEC1 regs_reg_13__4_ ( .D(i_data_Rd[4]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[420]), .QN(n75) );
  DFEC1 regs_reg_13__3_ ( .D(i_data_Rd[3]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[419]), .QN(n73) );
  DFEC1 regs_reg_13__2_ ( .D(i_data_Rd[2]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[418]), .QN(n71) );
  DFEC1 regs_reg_13__1_ ( .D(i_data_Rd[1]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[417]), .QN(n68) );
  DFEC1 regs_reg_13__0_ ( .D(i_data_Rd[0]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[416]), .QN(n122) );
  DFEC1 regs_reg_12__31_ ( .D(i_data_Rd[31]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(i_data_Rd[30]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(i_data_Rd[29]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(i_data_Rd[28]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(i_data_Rd[27]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(i_data_Rd[26]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(i_data_Rd[25]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(i_data_Rd[24]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(i_data_Rd[23]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(i_data_Rd[22]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(i_data_Rd[21]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(i_data_Rd[20]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(i_data_Rd[19]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(i_data_Rd[18]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(i_data_Rd[17]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(i_data_Rd[16]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(i_data_Rd[15]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(i_data_Rd[13]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(i_data_Rd[12]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(i_data_Rd[11]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(i_data_Rd[9]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(i_data_Rd[8]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(i_data_Rd[7]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(i_data_Rd[6]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(i_data_Rd[5]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(i_data_Rd[4]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(i_data_Rd[3]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(i_data_Rd[2]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(i_data_Rd[1]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(i_data_Rd[0]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[384]) );
  DFEC1 regs_reg_11__31_ ( .D(i_data_Rd[31]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(i_data_Rd[30]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(i_data_Rd[29]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(i_data_Rd[28]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(i_data_Rd[27]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(i_data_Rd[26]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(i_data_Rd[25]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(i_data_Rd[24]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(i_data_Rd[23]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(i_data_Rd[22]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(i_data_Rd[21]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(i_data_Rd[20]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(i_data_Rd[19]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(i_data_Rd[18]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(i_data_Rd[17]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(i_data_Rd[16]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(i_data_Rd[15]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(i_data_Rd[13]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(i_data_Rd[12]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(i_data_Rd[11]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(i_data_Rd[10]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(i_data_Rd[9]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(i_data_Rd[8]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(i_data_Rd[7]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(i_data_Rd[6]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(i_data_Rd[5]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(i_data_Rd[4]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(i_data_Rd[3]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(i_data_Rd[2]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(i_data_Rd[1]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(i_data_Rd[0]), .E(n58), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[352]) );
  DFEC1 regs_reg_10__31_ ( .D(i_data_Rd[31]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(i_data_Rd[30]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(i_data_Rd[29]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(i_data_Rd[28]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(i_data_Rd[27]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(i_data_Rd[26]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(i_data_Rd[25]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(i_data_Rd[24]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(i_data_Rd[23]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(i_data_Rd[22]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(i_data_Rd[21]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(i_data_Rd[20]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(i_data_Rd[19]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(i_data_Rd[18]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(i_data_Rd[17]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(i_data_Rd[16]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(i_data_Rd[15]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(i_data_Rd[13]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(i_data_Rd[12]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(i_data_Rd[11]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(i_data_Rd[9]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(i_data_Rd[8]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(i_data_Rd[7]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(i_data_Rd[6]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(i_data_Rd[5]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(i_data_Rd[4]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(i_data_Rd[3]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(i_data_Rd[2]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(i_data_Rd[1]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(i_data_Rd[0]), .E(n56), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[320]) );
  DFEC1 regs_reg_9__31_ ( .D(n263), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(n261), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(n259), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(n257), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(n255), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(n253), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(n251), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(n249), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(n247), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(n245), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(n243), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(n241), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(n239), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(n237), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(n235), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(n233), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(n231), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(n229), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(n227), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(n225), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(n223), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(n221), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(n219), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(n217), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(n215), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(n213), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(n211), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(n209), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(n207), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(n205), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(n203), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(n201), .E(n53), .C(i_clk), .RN(i_rst_n), .Q(
        regs[288]) );
  DFEC1 regs_reg_8__31_ ( .D(n262), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(n260), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(n258), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(n256), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(n254), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(n252), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(n250), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(n248), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(n246), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(n244), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(n242), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(n240), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(n238), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(n236), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(n234), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(n232), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(n230), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(n228), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(n226), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(n224), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(n222), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(n220), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(n218), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(n216), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(n214), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(n212), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(n210), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(n208), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(n206), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(n204), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(n202), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(n200), .E(n57), .C(i_clk), .RN(i_rst_n), .Q(
        regs[256]) );
  DFEC1 regs_reg_7__31_ ( .D(n263), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(n261), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(n259), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(n257), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(n255), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(n253), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(n251), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(n249), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(n247), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(n245), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(n243), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(n241), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(n239), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(n237), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(n235), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(n233), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(n231), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(n229), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(n227), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(n225), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(n223), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(n221), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(n219), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(n217), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(n215), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(n213), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(n211), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(n209), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(n207), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(n205), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(n203), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(n201), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[224]) );
  DFEC1 regs_reg_6__31_ ( .D(n263), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(n261), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(n259), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(n257), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(n255), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(n253), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(n251), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(n249), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(n247), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(n245), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(n243), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(n241), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(n239), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(n237), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(n235), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(n233), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(n231), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(n229), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(n227), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(n225), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(n223), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(n221), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(n219), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(n217), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(n215), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(n213), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(n211), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(n209), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(n207), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(n205), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(n203), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(n201), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[192]) );
  DFEC1 regs_reg_5__31_ ( .D(n263), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[191]), .QN(n192) );
  DFEC1 regs_reg_5__30_ ( .D(n261), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[190]), .QN(n189) );
  DFEC1 regs_reg_5__29_ ( .D(n259), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[189]), .QN(n186) );
  DFEC1 regs_reg_5__28_ ( .D(n257), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[188]), .QN(n183) );
  DFEC1 regs_reg_5__27_ ( .D(n255), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[187]), .QN(n180) );
  DFEC1 regs_reg_5__26_ ( .D(n253), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[186]), .QN(n177) );
  DFEC1 regs_reg_5__25_ ( .D(n251), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[185]), .QN(n174) );
  DFEC1 regs_reg_5__24_ ( .D(n249), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[184]), .QN(n171) );
  DFEC1 regs_reg_5__23_ ( .D(n247), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[183]), .QN(n168) );
  DFEC1 regs_reg_5__22_ ( .D(n245), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[182]), .QN(n165) );
  DFEC1 regs_reg_5__21_ ( .D(n243), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[181]), .QN(n162) );
  DFEC1 regs_reg_5__20_ ( .D(n241), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[180]), .QN(n160) );
  DFEC1 regs_reg_5__19_ ( .D(n239), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[179]), .QN(n158) );
  DFEC1 regs_reg_5__18_ ( .D(n237), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[178]), .QN(n156) );
  DFEC1 regs_reg_5__17_ ( .D(n235), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[177]), .QN(n154) );
  DFEC1 regs_reg_5__16_ ( .D(n233), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[176]), .QN(n152) );
  DFEC1 regs_reg_5__15_ ( .D(n231), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[175]), .QN(n150) );
  DFEC1 regs_reg_5__14_ ( .D(n229), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[174]), .QN(n148) );
  DFEC1 regs_reg_5__13_ ( .D(n227), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[173]), .QN(n146) );
  DFEC1 regs_reg_5__12_ ( .D(n225), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[172]), .QN(n144) );
  DFEC1 regs_reg_5__11_ ( .D(n223), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[171]), .QN(n142) );
  DFEC1 regs_reg_5__10_ ( .D(n221), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[170]), .QN(n140) );
  DFEC1 regs_reg_5__9_ ( .D(n219), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[169]), .QN(n138) );
  DFEC1 regs_reg_5__8_ ( .D(n217), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[168]), .QN(n136) );
  DFEC1 regs_reg_5__7_ ( .D(n215), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[167]), .QN(n134) );
  DFEC1 regs_reg_5__6_ ( .D(n213), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[166]), .QN(n132) );
  DFEC1 regs_reg_5__5_ ( .D(n211), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[165]), .QN(n130) );
  DFEC1 regs_reg_5__4_ ( .D(n209), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[164]), .QN(n128) );
  DFEC1 regs_reg_5__3_ ( .D(n207), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[163]), .QN(n126) );
  DFEC1 regs_reg_5__2_ ( .D(n205), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[162]), .QN(n124) );
  DFEC1 regs_reg_5__1_ ( .D(n203), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[161]), .QN(n70) );
  DFEC1 regs_reg_5__0_ ( .D(n201), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[160]), .QN(n123) );
  DFEC1 regs_reg_4__31_ ( .D(n263), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(n261), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(n259), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(n257), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(n255), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(n253), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(n251), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(n249), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(n247), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(n245), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(n243), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(n241), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(n239), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(n237), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(n235), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(n233), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(n231), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(n229), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(n227), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(n225), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(n223), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(n221), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(n219), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(n217), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(n215), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(n213), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(n211), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(n209), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(n207), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(n205), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(n203), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(n201), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[128]) );
  DFEC1 regs_reg_3__31_ ( .D(n263), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(n261), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(n259), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(n257), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(n255), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(n253), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(n251), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(n249), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(n247), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(n245), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(n243), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(n241), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(n239), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(n237), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(n235), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(n233), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(n231), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(n229), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(n227), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(n225), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(n223), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(n221), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(n219), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(n217), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(n215), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(n213), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(n211), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(n209), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(n207), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(n205), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(n203), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(n201), .E(n60), .C(i_clk), .RN(i_rst_n), .Q(
        regs[96]) );
  DFEC1 regs_reg_2__31_ ( .D(n263), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(n261), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(n259), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(n257), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(n255), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(n253), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(n251), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(n249), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(n247), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(n245), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(n243), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(n241), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(n239), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(n237), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(n235), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(n233), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(n231), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(n229), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(n227), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(n225), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(n223), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(n221), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(n219), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(n217), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(n215), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(n213), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(n211), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(n209), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(n207), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(n205), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(n203), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(n201), .E(n55), .C(i_clk), .RN(i_rst_n), .Q(
        regs[64]) );
  DFEC1 regs_reg_1__31_ ( .D(n263), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(n261), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(n259), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(n257), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(n255), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(n253), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(n251), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(n249), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(n247), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(n245), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(n243), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(n241), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(n239), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(n237), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(n235), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(n233), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(n231), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(n229), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(n227), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(n225), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(n223), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(n221), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(n219), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(n217), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(n215), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(n213), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(n211), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(n209), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(n207), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(n205), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(n203), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(n201), .E(n54), .C(i_clk), .RN(i_rst_n), .Q(
        regs[32]) );
  DFEC1 regs_reg_0__31_ ( .D(n263), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(n261), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(n259), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(n257), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(n255), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(n253), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(n251), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(n249), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(n247), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(n245), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(n243), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(n241), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(n239), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(n237), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(n235), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(n233), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(n231), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(n229), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(n227), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(n225), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(n223), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(n221), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(n219), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(n217), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(n215), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(n213), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(n211), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(n209), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(n207), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(n205), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(n203), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(n201), .E(n59), .C(i_clk), .RN(i_rst_n), .Q(
        regs[0]) );
  BUF8 U2 ( .A(n51), .Q(n1) );
  NOR24 U3 ( .A(n2), .B(n1798), .Q(n51) );
  CLKIN6 U4 ( .A(i_addr_Rs[2]), .Q(n2) );
  NOR41 U5 ( .A(n760), .B(n759), .C(n758), .D(n757), .Q(n761) );
  CLKBU12 U6 ( .A(n1061), .Q(n49) );
  CLKBU15 U7 ( .A(n1784), .Q(n48) );
  NOR41 U8 ( .A(n197), .B(n1817), .C(n1818), .D(n1819), .Q(n17) );
  BUF8 U9 ( .A(n15), .Q(n61) );
  BUF8 U10 ( .A(n16), .Q(n64) );
  BUF8 U11 ( .A(n13), .Q(n62) );
  INV3 U12 ( .A(n1075), .Q(n1039) );
  CLKBU12 U13 ( .A(n1057), .Q(n19) );
  CLKBU12 U14 ( .A(n1785), .Q(n8) );
  CLKBU12 U15 ( .A(n1787), .Q(n12) );
  BUF8 U16 ( .A(n1780), .Q(n10) );
  INV3 U17 ( .A(n1073), .Q(n1051) );
  NAND22 U18 ( .A(i_addr_Rs[3]), .B(i_addr_Rs[4]), .Q(n1045) );
  INV3 U19 ( .A(n1074), .Q(n1064) );
  NOR22 U20 ( .A(n1084), .B(n1091), .Q(n1775) );
  NOR22 U21 ( .A(i_addr_Rt_3_), .B(i_addr_Rt_4_), .Q(n1793) );
  BUF2 U22 ( .A(i_addr_Rd[1]), .Q(n196) );
  NAND31 U23 ( .A(i_con_RegWr), .B(i_addr_Rd[4]), .C(n1815), .Q(n1819) );
  BUF2 U24 ( .A(i_addr_Rd[0]), .Q(n195) );
  BUF2 U25 ( .A(n32), .Q(n59) );
  BUF2 U26 ( .A(n34), .Q(n54) );
  BUF2 U27 ( .A(n35), .Q(n55) );
  BUF2 U28 ( .A(n36), .Q(n60) );
  NOR22 U29 ( .A(n1816), .B(n1813), .Q(n37) );
  NOR22 U30 ( .A(n1813), .B(n1822), .Q(n38) );
  NOR22 U31 ( .A(n1813), .B(n1821), .Q(n39) );
  NOR22 U32 ( .A(n1820), .B(n1813), .Q(n40) );
  BUF2 U33 ( .A(n41), .Q(n57) );
  BUF2 U34 ( .A(n42), .Q(n53) );
  BUF2 U35 ( .A(n43), .Q(n56) );
  BUF2 U36 ( .A(n44), .Q(n58) );
  NOR22 U37 ( .A(n1823), .B(n1816), .Q(n5) );
  BUF2 U38 ( .A(n17), .Q(n63) );
  NOR22 U39 ( .A(n1816), .B(n1819), .Q(n18) );
  BUF2 U40 ( .A(i_data_Rd[0]), .Q(n201) );
  BUF2 U41 ( .A(i_data_Rd[1]), .Q(n203) );
  BUF2 U42 ( .A(i_data_Rd[2]), .Q(n205) );
  BUF2 U43 ( .A(i_data_Rd[3]), .Q(n207) );
  BUF2 U44 ( .A(i_data_Rd[4]), .Q(n209) );
  BUF2 U45 ( .A(i_data_Rd[5]), .Q(n211) );
  BUF2 U46 ( .A(i_data_Rd[6]), .Q(n213) );
  BUF2 U47 ( .A(i_data_Rd[7]), .Q(n215) );
  BUF2 U48 ( .A(i_data_Rd[8]), .Q(n217) );
  BUF2 U49 ( .A(i_data_Rd[9]), .Q(n219) );
  BUF2 U50 ( .A(i_data_Rd[10]), .Q(n221) );
  BUF2 U51 ( .A(i_data_Rd[11]), .Q(n223) );
  BUF2 U52 ( .A(i_data_Rd[12]), .Q(n225) );
  BUF2 U53 ( .A(i_data_Rd[13]), .Q(n227) );
  BUF2 U54 ( .A(i_data_Rd[14]), .Q(n229) );
  BUF2 U55 ( .A(i_data_Rd[15]), .Q(n231) );
  BUF2 U56 ( .A(i_data_Rd[16]), .Q(n233) );
  BUF2 U57 ( .A(i_data_Rd[17]), .Q(n235) );
  BUF2 U58 ( .A(i_data_Rd[18]), .Q(n237) );
  BUF2 U59 ( .A(i_data_Rd[19]), .Q(n239) );
  BUF2 U60 ( .A(i_data_Rd[20]), .Q(n241) );
  BUF2 U61 ( .A(i_data_Rd[21]), .Q(n243) );
  BUF2 U62 ( .A(i_data_Rd[22]), .Q(n245) );
  BUF2 U63 ( .A(i_data_Rd[23]), .Q(n247) );
  BUF2 U64 ( .A(i_data_Rd[24]), .Q(n249) );
  BUF2 U65 ( .A(i_data_Rd[25]), .Q(n251) );
  BUF2 U66 ( .A(i_data_Rd[26]), .Q(n253) );
  BUF2 U67 ( .A(i_data_Rd[27]), .Q(n255) );
  BUF2 U68 ( .A(i_data_Rd[28]), .Q(n257) );
  BUF2 U69 ( .A(i_data_Rd[29]), .Q(n259) );
  BUF2 U70 ( .A(i_data_Rd[30]), .Q(n261) );
  BUF2 U71 ( .A(i_data_Rd[31]), .Q(n263) );
  NOR22 U72 ( .A(n1816), .B(n1814), .Q(n28) );
  NOR22 U73 ( .A(n1822), .B(n1814), .Q(n29) );
  NOR22 U74 ( .A(n1821), .B(n1814), .Q(n30) );
  BUF2 U75 ( .A(i_data_Rd[0]), .Q(n200) );
  BUF2 U76 ( .A(i_data_Rd[1]), .Q(n202) );
  BUF2 U77 ( .A(i_data_Rd[2]), .Q(n204) );
  BUF2 U78 ( .A(i_data_Rd[3]), .Q(n206) );
  BUF2 U79 ( .A(i_data_Rd[4]), .Q(n208) );
  BUF2 U80 ( .A(i_data_Rd[5]), .Q(n210) );
  BUF2 U81 ( .A(i_data_Rd[6]), .Q(n212) );
  BUF2 U82 ( .A(i_data_Rd[7]), .Q(n214) );
  BUF2 U83 ( .A(i_data_Rd[8]), .Q(n216) );
  BUF2 U84 ( .A(i_data_Rd[9]), .Q(n218) );
  BUF2 U85 ( .A(i_data_Rd[10]), .Q(n220) );
  BUF2 U86 ( .A(i_data_Rd[11]), .Q(n222) );
  BUF2 U87 ( .A(i_data_Rd[12]), .Q(n224) );
  BUF2 U88 ( .A(i_data_Rd[13]), .Q(n226) );
  BUF2 U89 ( .A(i_data_Rd[14]), .Q(n228) );
  BUF2 U90 ( .A(i_data_Rd[15]), .Q(n230) );
  BUF2 U91 ( .A(i_data_Rd[16]), .Q(n232) );
  BUF2 U92 ( .A(i_data_Rd[17]), .Q(n234) );
  BUF2 U93 ( .A(i_data_Rd[18]), .Q(n236) );
  BUF2 U94 ( .A(i_data_Rd[19]), .Q(n238) );
  BUF2 U95 ( .A(i_data_Rd[20]), .Q(n240) );
  BUF2 U96 ( .A(i_data_Rd[21]), .Q(n242) );
  BUF2 U97 ( .A(i_data_Rd[22]), .Q(n244) );
  BUF2 U98 ( .A(i_data_Rd[23]), .Q(n246) );
  BUF2 U99 ( .A(i_data_Rd[24]), .Q(n248) );
  BUF2 U100 ( .A(i_data_Rd[25]), .Q(n250) );
  BUF2 U101 ( .A(i_data_Rd[26]), .Q(n252) );
  BUF2 U102 ( .A(i_data_Rd[27]), .Q(n254) );
  BUF2 U103 ( .A(i_data_Rd[28]), .Q(n256) );
  BUF2 U104 ( .A(i_data_Rd[29]), .Q(n258) );
  BUF2 U105 ( .A(i_data_Rd[30]), .Q(n260) );
  NOR22 U106 ( .A(n1820), .B(n1814), .Q(n31) );
  BUF2 U107 ( .A(i_data_Rd[31]), .Q(n262) );
  NOR32 U108 ( .A(i_addr_Rt_1_), .B(i_addr_Rt_2_), .C(n1078), .Q(n1784) );
  NOR22 U109 ( .A(n1822), .B(n1819), .Q(n20) );
  NOR22 U110 ( .A(n1821), .B(n1819), .Q(n21) );
  NOR22 U111 ( .A(n1820), .B(n1819), .Q(n22) );
  NOR42 U112 ( .A(n195), .B(n196), .C(n197), .D(n1814), .Q(n23) );
  NOR42 U113 ( .A(n197), .B(n196), .C(n1818), .D(n1814), .Q(n25) );
  NOR42 U114 ( .A(n195), .B(n197), .C(n1817), .D(n1814), .Q(n26) );
  NOR42 U115 ( .A(n197), .B(n1817), .C(n1818), .D(n1814), .Q(n27) );
  BUF8 U116 ( .A(n1061), .Q(n65) );
  NAND24 U117 ( .A(i_addr_Rs[1]), .B(i_addr_Rs[0]), .Q(n1798) );
  NOR33 U118 ( .A(n269), .B(i_addr_Rs[0]), .C(n268), .Q(n1056) );
  CLKBU12 U119 ( .A(n1063), .Q(n3) );
  CLKBU12 U120 ( .A(n1063), .Q(n4) );
  CLKIN3 U121 ( .A(n386), .Q(o_data_Rs[4]) );
  CLKIN3 U122 ( .A(n911), .Q(o_data_Rs[25]) );
  CLKIN3 U123 ( .A(n836), .Q(o_data_Rs[22]) );
  CLKIN3 U124 ( .A(n361), .Q(o_data_Rs[3]) );
  CLKIN3 U125 ( .A(n461), .Q(o_data_Rs[7]) );
  CLKIN3 U126 ( .A(n1011), .Q(o_data_Rs[29]) );
  CLKIN3 U127 ( .A(n336), .Q(o_data_Rs[2]) );
  CLKIN3 U128 ( .A(n661), .Q(o_data_Rs[15]) );
  CLKIN3 U129 ( .A(n1036), .Q(o_data_Rs[30]) );
  CLKIN3 U130 ( .A(n636), .Q(o_data_Rs[14]) );
  CLKIN3 U131 ( .A(n861), .Q(o_data_Rs[23]) );
  CLKIN3 U132 ( .A(n486), .Q(o_data_Rs[8]) );
  CLKIN3 U133 ( .A(n586), .Q(o_data_Rs[12]) );
  CLKIN3 U134 ( .A(n611), .Q(o_data_Rs[13]) );
  CLKIN3 U135 ( .A(n436), .Q(o_data_Rs[6]) );
  CLKIN3 U136 ( .A(n786), .Q(o_data_Rs[20]) );
  CLKIN3 U137 ( .A(n1072), .Q(o_data_Rs[31]) );
  CLKIN3 U138 ( .A(n711), .Q(o_data_Rs[17]) );
  CLKIN3 U139 ( .A(n511), .Q(o_data_Rs[9]) );
  CLKIN3 U140 ( .A(n886), .Q(o_data_Rs[24]) );
  CLKIN3 U141 ( .A(n936), .Q(o_data_Rs[26]) );
  CLKIN3 U142 ( .A(n536), .Q(o_data_Rs[10]) );
  CLKIN3 U143 ( .A(n686), .Q(o_data_Rs[16]) );
  CLKIN3 U144 ( .A(n411), .Q(o_data_Rs[5]) );
  CLKIN3 U145 ( .A(n811), .Q(o_data_Rs[21]) );
  CLKIN3 U146 ( .A(n561), .Q(o_data_Rs[11]) );
  CLKIN3 U147 ( .A(n761), .Q(o_data_Rs[19]) );
  OAI212 U148 ( .A(n100), .B(n49), .C(n667), .Q(n668) );
  OAI212 U149 ( .A(n99), .B(n49), .C(n662), .Q(n663) );
  OAI212 U150 ( .A(n152), .B(n49), .C(n672), .Q(n673) );
  BUF15 U151 ( .A(n1055), .Q(n7) );
  BUF12 U152 ( .A(n1058), .Q(n47) );
  BUF8 U153 ( .A(n1782), .Q(n50) );
  BUF12 U154 ( .A(n1783), .Q(n46) );
  NAND31 U155 ( .A(n197), .B(n1818), .C(n1817), .Q(n1816) );
  NOR32 U156 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .C(n1076), .Q(n1782) );
  BUF15 U157 ( .A(n1781), .Q(n14) );
  BUF15 U158 ( .A(n1786), .Q(n24) );
  BUF15 U159 ( .A(n1056), .Q(n33) );
  BUF15 U160 ( .A(n1059), .Q(n45) );
  CLKIN3 U161 ( .A(n736), .Q(o_data_Rs[18]) );
  AOI211 U162 ( .A(n3), .B(regs[577]), .C(n303), .Q(n306) );
  BUF6 U163 ( .A(n51), .Q(n199) );
  BUF6 U164 ( .A(n1782), .Q(n52) );
  NOR31 U165 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_2_), .C(n1079), .Q(n1787) );
  NAND31 U166 ( .A(n196), .B(n197), .C(n1818), .Q(n1821) );
  NAND31 U167 ( .A(n195), .B(n197), .C(n1817), .Q(n1822) );
  NAND31 U168 ( .A(n195), .B(n196), .C(n197), .Q(n1820) );
  NOR23 U169 ( .A(i_addr_Rt_3_), .B(n1091), .Q(n1795) );
  INV3 U170 ( .A(n195), .Q(n1818) );
  INV3 U171 ( .A(n196), .Q(n1817) );
  BUF6 U172 ( .A(i_addr_Rd[2]), .Q(n197) );
  NOR21 U173 ( .A(i_addr_Rs[4]), .B(i_addr_Rs[3]), .Q(n1073) );
  INV2 U174 ( .A(i_addr_Rs[3]), .Q(n275) );
  INV2 U175 ( .A(i_addr_Rs[4]), .Q(n281) );
  AOI211 U176 ( .A(n3), .B(regs[593]), .C(n703), .Q(n704) );
  AOI211 U177 ( .A(n4), .B(regs[579]), .C(n353), .Q(n354) );
  NOR40 U178 ( .A(n197), .B(n1818), .C(n1823), .D(n1817), .Q(n44) );
  NOR22 U179 ( .A(n1823), .B(n1820), .Q(n11) );
  NOR22 U180 ( .A(n1823), .B(n1821), .Q(n9) );
  NOR22 U181 ( .A(n1823), .B(n1822), .Q(n6) );
  NOR40 U182 ( .A(n195), .B(n197), .C(n1823), .D(n1817), .Q(n43) );
  NAND22 U183 ( .A(n1812), .B(n1815), .Q(n1813) );
  NOR31 U184 ( .A(i_addr_Rt_0_), .B(n1079), .C(n1076), .Q(n1783) );
  NOR31 U185 ( .A(i_addr_Rt_1_), .B(n1078), .C(n1076), .Q(n1780) );
  NOR21 U186 ( .A(n1077), .B(n1076), .Q(n1781) );
  NAND22 U187 ( .A(n1812), .B(i_addr_Rd[3]), .Q(n1823) );
  INV2 U188 ( .A(n1045), .Q(n198) );
  NOR21 U189 ( .A(n281), .B(i_addr_Rs[3]), .Q(n1074) );
  NOR21 U190 ( .A(i_addr_Rd[4]), .B(n1811), .Q(n1812) );
  NOR21 U191 ( .A(n275), .B(i_addr_Rs[4]), .Q(n1075) );
  NOR22 U192 ( .A(i_addr_Rt_4_), .B(n1084), .Q(n1773) );
  INV2 U193 ( .A(n961), .Q(o_data_Rs[27]) );
  INV2 U194 ( .A(n986), .Q(o_data_Rs[28]) );
  NOR40 U195 ( .A(n860), .B(n859), .C(n858), .D(n857), .Q(n861) );
  NOR40 U196 ( .A(n935), .B(n934), .C(n933), .D(n932), .Q(n936) );
  NOR40 U197 ( .A(n1071), .B(n1070), .C(n1069), .D(n1068), .Q(n1072) );
  NOR40 U198 ( .A(n910), .B(n909), .C(n908), .D(n907), .Q(n911) );
  NOR40 U199 ( .A(n835), .B(n834), .C(n833), .D(n832), .Q(n836) );
  NOR40 U200 ( .A(n960), .B(n959), .C(n958), .D(n957), .Q(n961) );
  NOR40 U201 ( .A(n885), .B(n884), .C(n883), .D(n882), .Q(n886) );
  NOR40 U202 ( .A(n635), .B(n634), .C(n633), .D(n632), .Q(n636) );
  NOR40 U203 ( .A(n810), .B(n809), .C(n808), .D(n807), .Q(n811) );
  NOR40 U204 ( .A(n360), .B(n359), .C(n358), .D(n357), .Q(n361) );
  NOR40 U205 ( .A(n785), .B(n784), .C(n783), .D(n782), .Q(n786) );
  NOR40 U206 ( .A(n735), .B(n734), .C(n733), .D(n732), .Q(n736) );
  NOR40 U207 ( .A(n385), .B(n384), .C(n383), .D(n382), .Q(n386) );
  NOR40 U208 ( .A(n660), .B(n659), .C(n658), .D(n657), .Q(n661) );
  NOR40 U209 ( .A(n685), .B(n684), .C(n683), .D(n682), .Q(n686) );
  NOR40 U210 ( .A(n710), .B(n709), .C(n708), .D(n707), .Q(n711) );
  NOR40 U211 ( .A(n1010), .B(n1009), .C(n1008), .D(n1007), .Q(n1011) );
  NOR40 U212 ( .A(n585), .B(n584), .C(n583), .D(n582), .Q(n586) );
  NOR40 U213 ( .A(n1035), .B(n1034), .C(n1033), .D(n1032), .Q(n1036) );
  NOR40 U214 ( .A(n535), .B(n534), .C(n533), .D(n532), .Q(n536) );
  NOR40 U215 ( .A(n985), .B(n984), .C(n983), .D(n982), .Q(n986) );
  NOR40 U216 ( .A(n335), .B(n334), .C(n333), .D(n332), .Q(n336) );
  NOR40 U217 ( .A(n610), .B(n609), .C(n608), .D(n607), .Q(n611) );
  NOR40 U218 ( .A(n485), .B(n484), .C(n483), .D(n482), .Q(n486) );
  NOR40 U219 ( .A(n410), .B(n409), .C(n408), .D(n407), .Q(n411) );
  NOR40 U220 ( .A(n560), .B(n559), .C(n558), .D(n557), .Q(n561) );
  NOR40 U221 ( .A(n510), .B(n509), .C(n508), .D(n507), .Q(n511) );
  NOR40 U222 ( .A(n460), .B(n459), .C(n458), .D(n457), .Q(n461) );
  AOI210 U223 ( .A(n4), .B(regs[65]), .C(n308), .Q(n311) );
  AOI210 U224 ( .A(n3), .B(regs[833]), .C(n293), .Q(n296) );
  OAI211 U225 ( .A(n113), .B(n49), .C(n862), .Q(n863) );
  OAI211 U226 ( .A(n93), .B(n49), .C(n587), .Q(n588) );
  OAI211 U227 ( .A(n191), .B(n49), .C(n1043), .Q(n1044) );
  NOR40 U228 ( .A(n197), .B(n1817), .C(n1818), .D(n1813), .Q(n36) );
  NOR40 U229 ( .A(n196), .B(n197), .C(n1818), .D(n1823), .Q(n42) );
  NOR40 U230 ( .A(n196), .B(n195), .C(n197), .D(n1823), .Q(n41) );
  NOR40 U231 ( .A(n195), .B(n197), .C(n1817), .D(n1813), .Q(n35) );
  NOR40 U232 ( .A(n195), .B(n196), .C(n197), .D(n1813), .Q(n32) );
  NOR40 U233 ( .A(n197), .B(n196), .C(n1818), .D(n1813), .Q(n34) );
  NOR22 U234 ( .A(i_addr_Rt_2_), .B(n1077), .Q(n1785) );
  NOR40 U235 ( .A(n195), .B(n196), .C(n197), .D(n1819), .Q(n13) );
  NOR40 U236 ( .A(n197), .B(n196), .C(n1818), .D(n1819), .Q(n15) );
  NOR40 U237 ( .A(n195), .B(n197), .C(n1817), .D(n1819), .Q(n16) );
  NOR40 U238 ( .A(n435), .B(n434), .C(n433), .D(n432), .Q(n436) );
  OAI211 U239 ( .A(n103), .B(n49), .C(n712), .Q(n713) );
  OAI211 U240 ( .A(n98), .B(n49), .C(n642), .Q(n643) );
  OAI211 U241 ( .A(n132), .B(n49), .C(n422), .Q(n423) );
  OAI211 U242 ( .A(n74), .B(n49), .C(n342), .Q(n343) );
  OAI211 U243 ( .A(n150), .B(n49), .C(n647), .Q(n648) );
  OAI211 U244 ( .A(n97), .B(n49), .C(n637), .Q(n638) );
  NOR21 U245 ( .A(i_addr_Rs[0]), .B(n271), .Q(n1055) );
  INV2 U246 ( .A(n270), .Q(n271) );
  NOR21 U247 ( .A(i_addr_Rs[0]), .B(n267), .Q(n1057) );
  NOR21 U248 ( .A(n266), .B(n267), .Q(n1058) );
  NOR21 U249 ( .A(n268), .B(i_addr_Rs[1]), .Q(n270) );
  NOR31 U250 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .C(i_addr_Rt_2_), .Q(n1786)
         );
  INV3 U251 ( .A(i_addr_Rs[2]), .Q(n268) );
  INV3 U252 ( .A(i_addr_Rs[1]), .Q(n269) );
  AOI221 U253 ( .A(n45), .B(regs[371]), .C(n199), .D(regs[499]), .Q(n737) );
  AOI221 U254 ( .A(n45), .B(regs[372]), .C(n199), .D(regs[500]), .Q(n762) );
  AOI221 U255 ( .A(n45), .B(regs[374]), .C(n199), .D(regs[502]), .Q(n812) );
  AOI221 U256 ( .A(n45), .B(regs[112]), .C(n1), .D(regs[240]), .Q(n672) );
  AOI221 U257 ( .A(n45), .B(regs[882]), .C(n199), .D(regs[1010]), .Q(n717) );
  AOI221 U258 ( .A(n45), .B(regs[623]), .C(n1), .D(regs[751]), .Q(n652) );
  AOI221 U259 ( .A(n45), .B(regs[624]), .C(n1), .D(regs[752]), .Q(n677) );
  AOI221 U260 ( .A(n45), .B(regs[884]), .C(n199), .D(regs[1012]), .Q(n767) );
  AOI221 U261 ( .A(n45), .B(regs[626]), .C(n199), .D(regs[754]), .Q(n727) );
  AOI221 U262 ( .A(n45), .B(regs[116]), .C(n199), .D(regs[244]), .Q(n772) );
  AOI221 U263 ( .A(n45), .B(regs[609]), .C(n1), .D(regs[737]), .Q(n302) );
  AOI221 U264 ( .A(n45), .B(regs[880]), .C(n1), .D(regs[1008]), .Q(n667) );
  AOI221 U265 ( .A(n45), .B(regs[881]), .C(n1), .D(regs[1009]), .Q(n692) );
  AOI221 U266 ( .A(n45), .B(regs[113]), .C(n1), .D(regs[241]), .Q(n697) );
  AOI221 U267 ( .A(n45), .B(regs[117]), .C(n199), .D(regs[245]), .Q(n797) );
  AOI221 U268 ( .A(n45), .B(regs[368]), .C(n1), .D(regs[496]), .Q(n662) );
  AOI221 U269 ( .A(n45), .B(regs[625]), .C(n1), .D(regs[753]), .Q(n702) );
  AOI221 U270 ( .A(n45), .B(regs[621]), .C(n1), .D(regs[749]), .Q(n602) );
  AOI221 U271 ( .A(n45), .B(regs[115]), .C(n199), .D(regs[243]), .Q(n747) );
  AOI221 U272 ( .A(n45), .B(regs[369]), .C(n1), .D(regs[497]), .Q(n687) );
  INV3 U273 ( .A(i_addr_Rt_2_), .Q(n1076) );
  NOR31 U274 ( .A(n269), .B(i_addr_Rs[0]), .C(i_addr_Rs[2]), .Q(n1063) );
  INV2 U275 ( .A(i_addr_Rs[0]), .Q(n266) );
  AOI221 U276 ( .A(n46), .B(regs[462]), .C(n1782), .D(regs[398]), .Q(n1396) );
  AOI221 U277 ( .A(n46), .B(regs[205]), .C(n1782), .D(regs[141]), .Q(n1384) );
  AOI221 U278 ( .A(n46), .B(regs[461]), .C(n1782), .D(regs[397]), .Q(n1374) );
  INV3 U279 ( .A(i_addr_Rt_1_), .Q(n1079) );
  NAND22 U280 ( .A(n268), .B(n269), .Q(n267) );
  NOR21 U281 ( .A(n1798), .B(i_addr_Rs[2]), .Q(n1059) );
  INV3 U282 ( .A(i_addr_Rt_0_), .Q(n1078) );
  INV3 U283 ( .A(i_addr_Rt_4_), .Q(n1091) );
  INV3 U284 ( .A(i_addr_Rt_3_), .Q(n1084) );
  AOI221 U285 ( .A(n46), .B(regs[730]), .C(n1782), .D(regs[666]), .Q(n1666) );
  AOI221 U286 ( .A(n46), .B(regs[218]), .C(n1782), .D(regs[154]), .Q(n1670) );
  AOI221 U287 ( .A(n46), .B(regs[988]), .C(n1782), .D(regs[924]), .Q(n1700) );
  AOI221 U288 ( .A(n46), .B(regs[474]), .C(n1782), .D(regs[410]), .Q(n1660) );
  AOI220 U289 ( .A(n46), .B(regs[475]), .C(n1782), .D(regs[411]), .Q(n1682) );
  NAND22 U290 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .Q(n1077) );
  AOI221 U291 ( .A(n8), .B(regs[622]), .C(n48), .D(regs[558]), .Q(n1401) );
  AOI221 U292 ( .A(n8), .B(regs[110]), .C(n48), .D(regs[46]), .Q(n1405) );
  AOI221 U293 ( .A(n8), .B(regs[619]), .C(n48), .D(regs[555]), .Q(n1335) );
  AOI220 U294 ( .A(n46), .B(regs[473]), .C(n1782), .D(regs[409]), .Q(n1638) );
  AOI221 U295 ( .A(n8), .B(regs[618]), .C(n48), .D(regs[554]), .Q(n1313) );
  AOI221 U296 ( .A(n46), .B(regs[987]), .C(n1782), .D(regs[923]), .Q(n1678) );
  AOI220 U297 ( .A(n46), .B(regs[217]), .C(n1782), .D(regs[153]), .Q(n1648) );
  AOI220 U298 ( .A(n46), .B(regs[472]), .C(n1782), .D(regs[408]), .Q(n1616) );
  AOI220 U299 ( .A(n46), .B(regs[976]), .C(n1782), .D(regs[912]), .Q(n1436) );
  AOI221 U300 ( .A(n8), .B(regs[367]), .C(n48), .D(regs[303]), .Q(n1417) );
  AOI221 U301 ( .A(n8), .B(regs[879]), .C(n48), .D(regs[815]), .Q(n1413) );
  AOI221 U302 ( .A(n46), .B(regs[719]), .C(n1782), .D(regs[655]), .Q(n1424) );
  AOI221 U303 ( .A(n8), .B(regs[113]), .C(n48), .D(regs[49]), .Q(n1471) );
  AOI221 U304 ( .A(n8), .B(regs[623]), .C(n48), .D(regs[559]), .Q(n1423) );
  AOI221 U305 ( .A(n8), .B(regs[368]), .C(n48), .D(regs[304]), .Q(n1439) );
  AOI221 U306 ( .A(n8), .B(regs[880]), .C(n48), .D(regs[816]), .Q(n1435) );
  AOI221 U307 ( .A(n46), .B(regs[223]), .C(n1782), .D(regs[159]), .Q(n1790) );
  AOI221 U308 ( .A(n8), .B(regs[127]), .C(n48), .D(regs[63]), .Q(n1789) );
  AOI221 U309 ( .A(n8), .B(regs[111]), .C(n48), .D(regs[47]), .Q(n1427) );
  AOI221 U310 ( .A(n33), .B(regs[726]), .C(n7), .D(regs[662]), .Q(n831) );
  AOI221 U311 ( .A(n47), .B(regs[572]), .C(n19), .D(regs[540]), .Q(n980) );
  AOI221 U312 ( .A(n47), .B(regs[299]), .C(n19), .D(regs[267]), .Q(n540) );
  AOI221 U313 ( .A(n47), .B(regs[317]), .C(n19), .D(regs[285]), .Q(n990) );
  AOI221 U314 ( .A(n47), .B(regs[557]), .C(n19), .D(regs[525]), .Q(n605) );
  AOI220 U315 ( .A(n46), .B(regs[718]), .C(n1782), .D(regs[654]), .Q(n1402) );
  AOI221 U316 ( .A(n47), .B(regs[828]), .C(n19), .D(regs[796]), .Q(n970) );
  AOI221 U317 ( .A(n47), .B(regs[316]), .C(n19), .D(regs[284]), .Q(n965) );
  AOI221 U318 ( .A(n47), .B(regs[827]), .C(n19), .D(regs[795]), .Q(n945) );
  AOI220 U319 ( .A(n46), .B(regs[463]), .C(n1782), .D(regs[399]), .Q(n1418) );
  AOI221 U320 ( .A(n47), .B(regs[38]), .C(n19), .D(regs[6]), .Q(n425) );
  AOI220 U321 ( .A(n46), .B(regs[207]), .C(n1782), .D(regs[143]), .Q(n1428) );
  AOI220 U322 ( .A(n46), .B(regs[975]), .C(n1782), .D(regs[911]), .Q(n1414) );
  AOI221 U323 ( .A(n47), .B(regs[571]), .C(n19), .D(regs[539]), .Q(n955) );
  AOI221 U324 ( .A(n47), .B(regs[298]), .C(n19), .D(regs[266]), .Q(n515) );
  AOI221 U325 ( .A(n47), .B(regs[302]), .C(n19), .D(regs[270]), .Q(n615) );
  AOI221 U326 ( .A(n47), .B(regs[814]), .C(n19), .D(regs[782]), .Q(n620) );
  AOI221 U327 ( .A(n47), .B(regs[824]), .C(n19), .D(regs[792]), .Q(n870) );
  AOI221 U328 ( .A(n47), .B(regs[56]), .C(n19), .D(regs[24]), .Q(n875) );
  AOI220 U329 ( .A(n46), .B(regs[206]), .C(n1782), .D(regs[142]), .Q(n1406) );
  AOI221 U330 ( .A(n47), .B(regs[548]), .C(n19), .D(regs[516]), .Q(n380) );
  AOI221 U331 ( .A(n47), .B(regs[558]), .C(n19), .D(regs[526]), .Q(n630) );
  AOI221 U332 ( .A(n47), .B(regs[805]), .C(n19), .D(regs[773]), .Q(n395) );
  OAI211 U333 ( .A(n87), .B(n65), .C(n512), .Q(n513) );
  OAI211 U334 ( .A(n143), .B(n65), .C(n552), .Q(n553) );
  OAI211 U335 ( .A(n142), .B(n65), .C(n547), .Q(n548) );
  OAI211 U336 ( .A(n114), .B(n65), .C(n887), .Q(n888) );
  OAI211 U337 ( .A(n73), .B(n65), .C(n337), .Q(n338) );
  OAI211 U338 ( .A(n90), .B(n65), .C(n542), .Q(n543) );
  OAI211 U339 ( .A(n125), .B(n65), .C(n327), .Q(n328) );
  OAI211 U340 ( .A(n172), .B(n65), .C(n877), .Q(n878) );
  OAI211 U341 ( .A(n89), .B(n65), .C(n537), .Q(n538) );
  OAI211 U342 ( .A(n145), .B(n65), .C(n577), .Q(n578) );
  OAI211 U343 ( .A(n144), .B(n65), .C(n572), .Q(n573) );
  OAI211 U344 ( .A(n166), .B(n65), .C(n827), .Q(n828) );
  OAI211 U345 ( .A(n92), .B(n65), .C(n567), .Q(n568) );
  OAI211 U346 ( .A(n124), .B(n65), .C(n322), .Q(n323) );
  OAI211 U347 ( .A(n164), .B(n65), .C(n817), .Q(n818) );
  OAI211 U348 ( .A(n91), .B(n65), .C(n562), .Q(n563) );
  OAI211 U349 ( .A(n69), .B(n65), .C(n302), .Q(n303) );
  OAI211 U350 ( .A(n71), .B(n65), .C(n312), .Q(n313) );
  OAI211 U351 ( .A(n68), .B(n65), .C(n297), .Q(n298) );
  OAI211 U352 ( .A(n70), .B(n65), .C(n307), .Q(n308) );
  OAI211 U353 ( .A(n170), .B(n65), .C(n867), .Q(n868) );
  OAI211 U354 ( .A(n121), .B(n65), .C(n264), .Q(n265) );
  OAI211 U355 ( .A(n139), .B(n65), .C(n502), .Q(n503) );
  OAI211 U356 ( .A(n122), .B(n65), .C(n276), .Q(n277) );
  OAI211 U357 ( .A(n141), .B(n65), .C(n527), .Q(n528) );
  OAI211 U358 ( .A(n111), .B(n65), .C(n812), .Q(n813) );
  OAI211 U359 ( .A(n174), .B(n65), .C(n897), .Q(n898) );
  OAI211 U360 ( .A(n194), .B(n65), .C(n282), .Q(n283) );
  OAI211 U361 ( .A(n123), .B(n65), .C(n287), .Q(n288) );
  OAI211 U362 ( .A(n140), .B(n65), .C(n522), .Q(n523) );
  OAI211 U363 ( .A(n67), .B(n65), .C(n292), .Q(n293) );
  OAI211 U364 ( .A(n72), .B(n65), .C(n317), .Q(n318) );
  OAI211 U365 ( .A(n165), .B(n65), .C(n822), .Q(n823) );
  OAI211 U366 ( .A(n88), .B(n65), .C(n517), .Q(n518) );
  OAI211 U367 ( .A(n185), .B(n65), .C(n992), .Q(n993) );
  OAI211 U368 ( .A(n162), .B(n65), .C(n797), .Q(n798) );
  OAI211 U369 ( .A(n169), .B(n65), .C(n852), .Q(n853) );
  OAI211 U370 ( .A(n186), .B(n65), .C(n997), .Q(n998) );
  OAI211 U371 ( .A(n153), .B(n65), .C(n677), .Q(n678) );
  OAI211 U372 ( .A(n154), .B(n65), .C(n697), .Q(n698) );
  AOI221 U373 ( .A(n46), .B(regs[197]), .C(n52), .D(regs[133]), .Q(n1208) );
  OAI211 U374 ( .A(n95), .B(n65), .C(n612), .Q(n613) );
  OAI211 U375 ( .A(n104), .B(n65), .C(n717), .Q(n718) );
  OAI211 U376 ( .A(n168), .B(n65), .C(n847), .Q(n848) );
  OAI211 U377 ( .A(n159), .B(n65), .C(n752), .Q(n753) );
  OAI211 U378 ( .A(n158), .B(n65), .C(n747), .Q(n748) );
  OAI211 U379 ( .A(n105), .B(n65), .C(n737), .Q(n738) );
  OAI211 U380 ( .A(n161), .B(n65), .C(n777), .Q(n778) );
  OAI211 U381 ( .A(n107), .B(n65), .C(n762), .Q(n763) );
  OAI211 U382 ( .A(n167), .B(n65), .C(n842), .Q(n843) );
  OAI211 U383 ( .A(n112), .B(n65), .C(n837), .Q(n838) );
  OAI211 U384 ( .A(n118), .B(n65), .C(n987), .Q(n988) );
  OAI211 U385 ( .A(n146), .B(n65), .C(n597), .Q(n598) );
  OAI211 U386 ( .A(n96), .B(n65), .C(n617), .Q(n618) );
  OAI211 U387 ( .A(n177), .B(n65), .C(n922), .Q(n923) );
  OAI211 U388 ( .A(n182), .B(n65), .C(n967), .Q(n968) );
  OAI211 U389 ( .A(n149), .B(n65), .C(n627), .Q(n628) );
  OAI211 U390 ( .A(n110), .B(n65), .C(n792), .Q(n793) );
  AOI221 U391 ( .A(n8), .B(regs[352]), .C(n48), .D(regs[288]), .Q(n1086) );
  AOI221 U392 ( .A(n8), .B(regs[878]), .C(n1784), .D(regs[814]), .Q(n1391) );
  AOI221 U393 ( .A(n8), .B(regs[866]), .C(n48), .D(regs[802]), .Q(n1127) );
  AOI221 U394 ( .A(n8), .B(regs[620]), .C(n48), .D(regs[556]), .Q(n1357) );
  AOI221 U395 ( .A(n8), .B(regs[112]), .C(n48), .D(regs[48]), .Q(n1449) );
  AOI221 U396 ( .A(n8), .B(regs[108]), .C(n48), .D(regs[44]), .Q(n1361) );
  AOI221 U397 ( .A(n8), .B(regs[624]), .C(n48), .D(regs[560]), .Q(n1445) );
  AOI221 U398 ( .A(n8), .B(regs[881]), .C(n48), .D(regs[817]), .Q(n1457) );
  AOI221 U399 ( .A(n8), .B(regs[874]), .C(n48), .D(regs[810]), .Q(n1303) );
  AOI221 U400 ( .A(n8), .B(regs[365]), .C(n48), .D(regs[301]), .Q(n1373) );
  AOI221 U401 ( .A(n8), .B(regs[873]), .C(n48), .D(regs[809]), .Q(n1281) );
  AOI221 U402 ( .A(n8), .B(regs[877]), .C(n1784), .D(regs[813]), .Q(n1369) );
  AOI221 U403 ( .A(n8), .B(regs[354]), .C(n48), .D(regs[290]), .Q(n1131) );
  AOI221 U404 ( .A(n8), .B(regs[109]), .C(n48), .D(regs[45]), .Q(n1383) );
  AOI221 U405 ( .A(n8), .B(regs[366]), .C(n48), .D(regs[302]), .Q(n1395) );
  AOI221 U406 ( .A(n8), .B(regs[625]), .C(n48), .D(regs[561]), .Q(n1467) );
  AOI221 U407 ( .A(n8), .B(regs[882]), .C(n48), .D(regs[818]), .Q(n1479) );
  AOI221 U408 ( .A(n8), .B(regs[621]), .C(n48), .D(regs[557]), .Q(n1379) );
  AOI221 U409 ( .A(n8), .B(regs[369]), .C(n48), .D(regs[305]), .Q(n1461) );
  AOI221 U410 ( .A(n8), .B(regs[353]), .C(n48), .D(regs[289]), .Q(n1109) );
  AOI221 U411 ( .A(n8), .B(regs[370]), .C(n48), .D(regs[306]), .Q(n1483) );
  AOI221 U412 ( .A(n8), .B(regs[616]), .C(n48), .D(regs[552]), .Q(n1269) );
  AOI221 U413 ( .A(n8), .B(regs[871]), .C(n48), .D(regs[807]), .Q(n1237) );
  AOI221 U414 ( .A(n8), .B(regs[617]), .C(n48), .D(regs[553]), .Q(n1291) );
  AOI221 U415 ( .A(n47), .B(regs[40]), .C(n19), .D(regs[8]), .Q(n475) );
  AOI221 U416 ( .A(n47), .B(regs[62]), .C(n19), .D(regs[30]), .Q(n1025) );
  AOI221 U417 ( .A(n47), .B(regs[294]), .C(n19), .D(regs[262]), .Q(n415) );
  AOI221 U418 ( .A(n47), .B(regs[806]), .C(n19), .D(regs[774]), .Q(n420) );
  AOI221 U419 ( .A(n47), .B(regs[63]), .C(n19), .D(regs[31]), .Q(n1053) );
  AOI221 U420 ( .A(n47), .B(regs[831]), .C(n19), .D(regs[799]), .Q(n1047) );
  AOI221 U421 ( .A(n47), .B(regs[550]), .C(n19), .D(regs[518]), .Q(n430) );
  AOI221 U422 ( .A(n47), .B(regs[319]), .C(n19), .D(regs[287]), .Q(n1041) );
  AOI221 U423 ( .A(n47), .B(regs[37]), .C(n19), .D(regs[5]), .Q(n400) );
  AOI221 U424 ( .A(n47), .B(regs[549]), .C(n19), .D(regs[517]), .Q(n405) );
  AOI221 U425 ( .A(n47), .B(regs[36]), .C(n19), .D(regs[4]), .Q(n375) );
  AOI221 U426 ( .A(n47), .B(regs[803]), .C(n19), .D(regs[771]), .Q(n345) );
  AOI221 U427 ( .A(n47), .B(regs[801]), .C(n19), .D(regs[769]), .Q(n295) );
  AOI221 U428 ( .A(n47), .B(regs[289]), .C(n19), .D(regs[257]), .Q(n300) );
  AOI221 U429 ( .A(n47), .B(regs[545]), .C(n19), .D(regs[513]), .Q(n305) );
  AOI221 U430 ( .A(n47), .B(regs[33]), .C(n19), .D(regs[1]), .Q(n310) );
  AOI221 U431 ( .A(n47), .B(regs[800]), .C(n19), .D(regs[768]), .Q(n273) );
  AOI221 U432 ( .A(n47), .B(regs[288]), .C(n19), .D(regs[256]), .Q(n279) );
  AOI221 U433 ( .A(n47), .B(regs[544]), .C(n19), .D(regs[512]), .Q(n285) );
  AOI221 U434 ( .A(n47), .B(regs[32]), .C(n19), .D(regs[0]), .Q(n290) );
  AOI221 U435 ( .A(n47), .B(regs[567]), .C(n19), .D(regs[535]), .Q(n855) );
  AOI221 U436 ( .A(n47), .B(regs[310]), .C(n19), .D(regs[278]), .Q(n815) );
  AOI221 U437 ( .A(n47), .B(regs[822]), .C(n19), .D(regs[790]), .Q(n820) );
  AOI221 U438 ( .A(n47), .B(regs[54]), .C(n19), .D(regs[22]), .Q(n825) );
  AOI221 U439 ( .A(n47), .B(regs[566]), .C(n19), .D(regs[534]), .Q(n830) );
  AOI221 U440 ( .A(n47), .B(regs[309]), .C(n19), .D(regs[277]), .Q(n790) );
  AOI221 U441 ( .A(n47), .B(regs[821]), .C(n19), .D(regs[789]), .Q(n795) );
  AOI221 U442 ( .A(n47), .B(regs[53]), .C(n19), .D(regs[21]), .Q(n800) );
  AOI221 U443 ( .A(n47), .B(regs[565]), .C(n19), .D(regs[533]), .Q(n805) );
  AOI221 U444 ( .A(n47), .B(regs[49]), .C(n19), .D(regs[17]), .Q(n700) );
  AOI221 U445 ( .A(n47), .B(regs[561]), .C(n19), .D(regs[529]), .Q(n705) );
  AOI221 U446 ( .A(n47), .B(regs[304]), .C(n19), .D(regs[272]), .Q(n665) );
  AOI221 U447 ( .A(n47), .B(regs[816]), .C(n19), .D(regs[784]), .Q(n670) );
  AOI221 U448 ( .A(n47), .B(regs[48]), .C(n19), .D(regs[16]), .Q(n675) );
  AOI221 U449 ( .A(n47), .B(regs[560]), .C(n19), .D(regs[528]), .Q(n680) );
  AOI221 U450 ( .A(n47), .B(regs[303]), .C(n19), .D(regs[271]), .Q(n640) );
  AOI221 U451 ( .A(n47), .B(regs[815]), .C(n19), .D(regs[783]), .Q(n645) );
  AOI221 U452 ( .A(n47), .B(regs[47]), .C(n19), .D(regs[15]), .Q(n650) );
  AOI221 U453 ( .A(n47), .B(regs[559]), .C(n19), .D(regs[527]), .Q(n655) );
  INV3 U454 ( .A(i_addr_Rd[3]), .Q(n1815) );
  AOI221 U455 ( .A(n14), .B(regs[231]), .C(n10), .D(regs[167]), .Q(n1253) );
  AOI221 U456 ( .A(n46), .B(regs[198]), .C(n52), .D(regs[134]), .Q(n1230) );
  AOI221 U457 ( .A(n14), .B(regs[230]), .C(n10), .D(regs[166]), .Q(n1231) );
  AOI221 U458 ( .A(n46), .B(regs[194]), .C(n52), .D(regs[130]), .Q(n1142) );
  AOI221 U459 ( .A(n46), .B(regs[715]), .C(n50), .D(regs[651]), .Q(n1336) );
  AOI221 U460 ( .A(n46), .B(regs[210]), .C(n50), .D(regs[146]), .Q(n1494) );
  AOI221 U461 ( .A(n14), .B(regs[496]), .C(n10), .D(regs[432]), .Q(n1441) );
  AOI221 U462 ( .A(n14), .B(regs[1000]), .C(n10), .D(regs[936]), .Q(n1261) );
  AOI221 U463 ( .A(n46), .B(regs[199]), .C(n52), .D(regs[135]), .Q(n1252) );
  AOI221 U464 ( .A(n46), .B(regs[211]), .C(n50), .D(regs[147]), .Q(n1516) );
  AOI221 U465 ( .A(n14), .B(regs[488]), .C(n10), .D(regs[424]), .Q(n1265) );
  AOI221 U466 ( .A(n14), .B(regs[487]), .C(n10), .D(regs[423]), .Q(n1243) );
  AOI221 U467 ( .A(n46), .B(regs[201]), .C(n50), .D(regs[137]), .Q(n1296) );
  AOI221 U468 ( .A(n14), .B(regs[497]), .C(n10), .D(regs[433]), .Q(n1463) );
  AOI221 U469 ( .A(n14), .B(regs[1010]), .C(n10), .D(regs[946]), .Q(n1481) );
  AOI221 U470 ( .A(n14), .B(regs[742]), .C(n10), .D(regs[678]), .Q(n1227) );
  AOI221 U471 ( .A(n14), .B(regs[237]), .C(n10), .D(regs[173]), .Q(n1385) );
  AOI221 U472 ( .A(n46), .B(regs[710]), .C(n52), .D(regs[646]), .Q(n1226) );
  AOI221 U473 ( .A(n14), .B(regs[743]), .C(n10), .D(regs[679]), .Q(n1249) );
  AOI221 U474 ( .A(n14), .B(regs[505]), .C(n10), .D(regs[441]), .Q(n1639) );
  AOI221 U475 ( .A(n46), .B(regs[203]), .C(n50), .D(regs[139]), .Q(n1340) );
  AOI221 U476 ( .A(n14), .B(regs[1020]), .C(n10), .D(regs[956]), .Q(n1701) );
  AOI221 U477 ( .A(n14), .B(regs[236]), .C(n10), .D(regs[172]), .Q(n1363) );
  AOI221 U478 ( .A(n14), .B(regs[763]), .C(n10), .D(regs[699]), .Q(n1689) );
  AOI221 U479 ( .A(n14), .B(regs[494]), .C(n10), .D(regs[430]), .Q(n1397) );
  AOI221 U480 ( .A(n14), .B(regs[506]), .C(n10), .D(regs[442]), .Q(n1661) );
  AOI221 U481 ( .A(n14), .B(regs[226]), .C(n10), .D(regs[162]), .Q(n1143) );
  AOI221 U482 ( .A(n14), .B(regs[493]), .C(n10), .D(regs[429]), .Q(n1375) );
  AOI221 U483 ( .A(n46), .B(regs[714]), .C(n50), .D(regs[650]), .Q(n1314) );
  AOI221 U484 ( .A(n14), .B(regs[999]), .C(n10), .D(regs[935]), .Q(n1239) );
  AOI221 U485 ( .A(n46), .B(regs[202]), .C(n50), .D(regs[138]), .Q(n1318) );
  AOI221 U486 ( .A(n8), .B(regs[124]), .C(n48), .D(regs[60]), .Q(n1713) );
  OAI211 U487 ( .A(n176), .B(n49), .C(n917), .Q(n918) );
  OAI211 U488 ( .A(n119), .B(n49), .C(n1012), .Q(n1013) );
  AOI221 U489 ( .A(n12), .B(regs[597]), .C(n24), .D(regs[533]), .Q(n1554) );
  AOI221 U490 ( .A(n8), .B(regs[611]), .C(n48), .D(regs[547]), .Q(n1159) );
  AOI221 U491 ( .A(n8), .B(regs[355]), .C(n48), .D(regs[291]), .Q(n1153) );
  OAI211 U492 ( .A(n188), .B(n49), .C(n1017), .Q(n1018) );
  AOI221 U493 ( .A(n8), .B(regs[99]), .C(n1784), .D(regs[35]), .Q(n1163) );
  AOI221 U494 ( .A(n12), .B(regs[341]), .C(n24), .D(regs[277]), .Q(n1548) );
  AOI221 U495 ( .A(n12), .B(regs[853]), .C(n24), .D(regs[789]), .Q(n1544) );
  AOI221 U496 ( .A(n8), .B(regs[891]), .C(n1784), .D(regs[827]), .Q(n1677) );
  AOI221 U497 ( .A(n46), .B(regs[479]), .C(n50), .D(regs[415]), .Q(n1770) );
  OAI211 U498 ( .A(n106), .B(n49), .C(n742), .Q(n743) );
  OAI211 U499 ( .A(n127), .B(n49), .C(n352), .Q(n353) );
  AOI221 U500 ( .A(n8), .B(regs[875]), .C(n1784), .D(regs[811]), .Q(n1325) );
  AOI221 U501 ( .A(n8), .B(regs[125]), .C(n1784), .D(regs[61]), .Q(n1735) );
  AOI221 U502 ( .A(n12), .B(regs[84]), .C(n24), .D(regs[20]), .Q(n1536) );
  OAI211 U503 ( .A(n129), .B(n49), .C(n377), .Q(n378) );
  AOI221 U504 ( .A(n46), .B(regs[221]), .C(n50), .D(regs[157]), .Q(n1736) );
  OAI211 U505 ( .A(n160), .B(n49), .C(n772), .Q(n773) );
  AOI221 U506 ( .A(n8), .B(regs[357]), .C(n48), .D(regs[293]), .Q(n1197) );
  AOI221 U507 ( .A(n8), .B(regs[637]), .C(n48), .D(regs[573]), .Q(n1731) );
  AOI221 U508 ( .A(n46), .B(regs[733]), .C(n50), .D(regs[669]), .Q(n1732) );
  AOI221 U509 ( .A(n8), .B(regs[892]), .C(n1784), .D(regs[828]), .Q(n1699) );
  AOI221 U510 ( .A(n8), .B(regs[381]), .C(n48), .D(regs[317]), .Q(n1725) );
  OAI211 U511 ( .A(n126), .B(n49), .C(n347), .Q(n348) );
  AOI221 U512 ( .A(n12), .B(regs[596]), .C(n24), .D(regs[532]), .Q(n1532) );
  AOI221 U513 ( .A(n46), .B(regs[477]), .C(n50), .D(regs[413]), .Q(n1726) );
  AOI221 U514 ( .A(n8), .B(regs[893]), .C(n1784), .D(regs[829]), .Q(n1721) );
  AOI221 U515 ( .A(n46), .B(regs[989]), .C(n50), .D(regs[925]), .Q(n1722) );
  OAI211 U516 ( .A(n108), .B(n49), .C(n767), .Q(n768) );
  AOI221 U517 ( .A(n8), .B(regs[868]), .C(n1784), .D(regs[804]), .Q(n1171) );
  AOI221 U518 ( .A(n12), .B(regs[340]), .C(n24), .D(regs[276]), .Q(n1526) );
  AOI221 U519 ( .A(n46), .B(regs[476]), .C(n50), .D(regs[412]), .Q(n1704) );
  AOI221 U520 ( .A(n8), .B(regs[380]), .C(n48), .D(regs[316]), .Q(n1703) );
  AOI221 U521 ( .A(n8), .B(regs[356]), .C(n48), .D(regs[292]), .Q(n1175) );
  AOI221 U522 ( .A(n12), .B(regs[324]), .C(n24), .D(regs[260]), .Q(n1174) );
  AOI221 U523 ( .A(n46), .B(regs[204]), .C(n52), .D(regs[140]), .Q(n1362) );
  OAI211 U524 ( .A(n190), .B(n49), .C(n1027), .Q(n1028) );
  AOI221 U525 ( .A(n46), .B(regs[732]), .C(n50), .D(regs[668]), .Q(n1710) );
  AOI221 U526 ( .A(n8), .B(regs[100]), .C(n48), .D(regs[36]), .Q(n1185) );
  AOI221 U527 ( .A(n8), .B(regs[636]), .C(n48), .D(regs[572]), .Q(n1709) );
  AOI221 U528 ( .A(n46), .B(regs[974]), .C(n52), .D(regs[910]), .Q(n1392) );
  AOI221 U529 ( .A(n12), .B(regs[85]), .C(n24), .D(regs[21]), .Q(n1558) );
  AOI221 U530 ( .A(n46), .B(regs[478]), .C(n50), .D(regs[414]), .Q(n1748) );
  AOI221 U531 ( .A(n8), .B(regs[867]), .C(n48), .D(regs[803]), .Q(n1149) );
  AOI221 U532 ( .A(n8), .B(regs[894]), .C(n48), .D(regs[830]), .Q(n1743) );
  OAI211 U533 ( .A(n189), .B(n49), .C(n1022), .Q(n1023) );
  AOI221 U534 ( .A(n46), .B(regs[990]), .C(n50), .D(regs[926]), .Q(n1744) );
  AOI221 U535 ( .A(n46), .B(regs[208]), .C(n52), .D(regs[144]), .Q(n1450) );
  AOI221 U536 ( .A(n46), .B(regs[220]), .C(n50), .D(regs[156]), .Q(n1714) );
  AOI221 U537 ( .A(n8), .B(regs[876]), .C(n48), .D(regs[812]), .Q(n1347) );
  OAI211 U538 ( .A(n193), .B(n49), .C(n1060), .Q(n1062) );
  AOI221 U539 ( .A(n8), .B(regs[634]), .C(n48), .D(regs[570]), .Q(n1665) );
  OAI211 U540 ( .A(n101), .B(n49), .C(n687), .Q(n688) );
  AOI221 U541 ( .A(n12), .B(regs[855]), .C(n24), .D(regs[791]), .Q(n1588) );
  OAI211 U542 ( .A(n102), .B(n49), .C(n692), .Q(n693) );
  AOI221 U543 ( .A(n8), .B(regs[122]), .C(n1784), .D(regs[58]), .Q(n1669) );
  OAI211 U544 ( .A(n155), .B(n49), .C(n702), .Q(n703) );
  AOI221 U545 ( .A(regs[704]), .B(n46), .C(regs[640]), .D(n50), .Q(n1094) );
  AOI221 U546 ( .A(n46), .B(regs[985]), .C(n50), .D(regs[921]), .Q(n1634) );
  AOI221 U547 ( .A(n8), .B(regs[889]), .C(n48), .D(regs[825]), .Q(n1633) );
  OAI211 U548 ( .A(n109), .B(n49), .C(n787), .Q(n788) );
  OAI211 U549 ( .A(n192), .B(n49), .C(n1049), .Q(n1050) );
  AOI221 U550 ( .A(n8), .B(regs[120]), .C(n48), .D(regs[56]), .Q(n1625) );
  AOI221 U551 ( .A(n12), .B(regs[335]), .C(n24), .D(regs[271]), .Q(n1416) );
  AOI221 U552 ( .A(n46), .B(regs[216]), .C(n50), .D(regs[152]), .Q(n1626) );
  AOI221 U553 ( .A(n8), .B(regs[632]), .C(n48), .D(regs[568]), .Q(n1621) );
  AOI221 U554 ( .A(n46), .B(regs[728]), .C(n50), .D(regs[664]), .Q(n1622) );
  OAI211 U555 ( .A(n120), .B(n49), .C(n1037), .Q(n1038) );
  AOI221 U556 ( .A(n46), .B(regs[729]), .C(n50), .D(regs[665]), .Q(n1644) );
  AOI221 U557 ( .A(n8), .B(regs[376]), .C(n48), .D(regs[312]), .Q(n1615) );
  AOI221 U558 ( .A(n8), .B(regs[633]), .C(n48), .D(regs[569]), .Q(n1643) );
  AOI221 U559 ( .A(n46), .B(regs[717]), .C(n52), .D(regs[653]), .Q(n1380) );
  OAI211 U560 ( .A(n151), .B(n49), .C(n652), .Q(n653) );
  AOI221 U561 ( .A(n12), .B(regs[856]), .C(n24), .D(regs[792]), .Q(n1610) );
  AOI221 U562 ( .A(n8), .B(regs[121]), .C(n48), .D(regs[57]), .Q(n1647) );
  OAI211 U563 ( .A(n148), .B(n49), .C(n622), .Q(n623) );
  AOI221 U564 ( .A(n12), .B(regs[86]), .C(n24), .D(regs[22]), .Q(n1580) );
  AOI221 U565 ( .A(n8), .B(regs[379]), .C(n48), .D(regs[315]), .Q(n1681) );
  AOI221 U566 ( .A(n12), .B(regs[347]), .C(n24), .D(regs[283]), .Q(n1680) );
  AOI221 U567 ( .A(n8), .B(regs[610]), .C(n48), .D(regs[546]), .Q(n1137) );
  AOI221 U568 ( .A(n46), .B(regs[716]), .C(n52), .D(regs[652]), .Q(n1358) );
  AOI221 U569 ( .A(n46), .B(regs[731]), .C(n1782), .D(regs[667]), .Q(n1688) );
  OAI211 U570 ( .A(n147), .B(n49), .C(n602), .Q(n603) );
  AOI221 U571 ( .A(n8), .B(regs[635]), .C(n48), .D(regs[571]), .Q(n1687) );
  OAI211 U572 ( .A(n163), .B(n49), .C(n802), .Q(n803) );
  AOI221 U573 ( .A(n12), .B(regs[342]), .C(n24), .D(regs[278]), .Q(n1570) );
  AOI221 U574 ( .A(n12), .B(regs[854]), .C(n24), .D(regs[790]), .Q(n1566) );
  AOI221 U575 ( .A(n46), .B(regs[219]), .C(n1782), .D(regs[155]), .Q(n1692) );
  AOI221 U576 ( .A(n12), .B(regs[332]), .C(n24), .D(regs[268]), .Q(n1350) );
  AOI221 U577 ( .A(n8), .B(regs[123]), .C(n1784), .D(regs[59]), .Q(n1691) );
  AOI221 U578 ( .A(n12), .B(regs[87]), .C(n24), .D(regs[23]), .Q(n1602) );
  AOI221 U579 ( .A(n46), .B(regs[973]), .C(n52), .D(regs[909]), .Q(n1370) );
  OAI211 U580 ( .A(n156), .B(n49), .C(n722), .Q(n723) );
  AOI221 U581 ( .A(n8), .B(regs[364]), .C(n48), .D(regs[300]), .Q(n1351) );
  AOI221 U582 ( .A(n46), .B(regs[986]), .C(n50), .D(regs[922]), .Q(n1656) );
  OAI211 U583 ( .A(n178), .B(n49), .C(n927), .Q(n928) );
  AOI221 U584 ( .A(n8), .B(regs[890]), .C(n48), .D(regs[826]), .Q(n1655) );
  OAI211 U585 ( .A(n157), .B(n49), .C(n727), .Q(n728) );
  AOI221 U586 ( .A(n8), .B(regs[98]), .C(n1784), .D(regs[34]), .Q(n1141) );
  OAI211 U587 ( .A(n94), .B(n49), .C(n592), .Q(n593) );
  AOI221 U588 ( .A(n12), .B(regs[343]), .C(n24), .D(regs[279]), .Q(n1592) );
  AOI221 U589 ( .A(n8), .B(regs[378]), .C(n48), .D(regs[314]), .Q(n1659) );
  AOI221 U590 ( .A(n12), .B(regs[346]), .C(n24), .D(regs[282]), .Q(n1658) );
  AOI221 U591 ( .A(n12), .B(regs[844]), .C(n24), .D(regs[780]), .Q(n1346) );
  OAI211 U592 ( .A(n115), .B(n49), .C(n912), .Q(n913) );
  OAI211 U593 ( .A(n173), .B(n49), .C(n892), .Q(n893) );
  AOI221 U594 ( .A(n12), .B(regs[331]), .C(n24), .D(regs[267]), .Q(n1328) );
  OAI211 U595 ( .A(n183), .B(n49), .C(n972), .Q(n973) );
  AOI221 U596 ( .A(n12), .B(regs[329]), .C(n24), .D(regs[265]), .Q(n1284) );
  OAI211 U597 ( .A(n78), .B(n49), .C(n392), .Q(n393) );
  AOI221 U598 ( .A(n46), .B(regs[977]), .C(n52), .D(regs[913]), .Q(n1458) );
  AOI221 U599 ( .A(n12), .B(regs[75]), .C(n24), .D(regs[11]), .Q(n1338) );
  OAI211 U600 ( .A(n82), .B(n49), .C(n442), .Q(n443) );
  AOI221 U601 ( .A(n8), .B(regs[106]), .C(n48), .D(regs[42]), .Q(n1317) );
  OAI211 U602 ( .A(n175), .B(n49), .C(n902), .Q(n903) );
  AOI221 U603 ( .A(n12), .B(regs[74]), .C(n24), .D(regs[10]), .Q(n1316) );
  AOI221 U604 ( .A(n8), .B(regs[363]), .C(n48), .D(regs[299]), .Q(n1329) );
  AOI221 U605 ( .A(n8), .B(regs[358]), .C(n48), .D(regs[294]), .Q(n1219) );
  OAI211 U606 ( .A(n81), .B(n49), .C(n437), .Q(n438) );
  AOI221 U607 ( .A(n12), .B(regs[330]), .C(n24), .D(regs[266]), .Q(n1306) );
  OAI211 U608 ( .A(n130), .B(n49), .C(n397), .Q(n398) );
  OAI211 U609 ( .A(n180), .B(n49), .C(n947), .Q(n948) );
  OAI211 U610 ( .A(n134), .B(n49), .C(n447), .Q(n448) );
  OAI211 U611 ( .A(n77), .B(n49), .C(n387), .Q(n388) );
  AOI221 U612 ( .A(n8), .B(regs[615]), .C(n48), .D(regs[551]), .Q(n1247) );
  AOI221 U613 ( .A(n8), .B(regs[104]), .C(n1784), .D(regs[40]), .Q(n1273) );
  OAI211 U614 ( .A(n86), .B(n49), .C(n492), .Q(n493) );
  AOI221 U615 ( .A(n8), .B(regs[361]), .C(n48), .D(regs[297]), .Q(n1285) );
  OAI211 U616 ( .A(n138), .B(n49), .C(n497), .Q(n498) );
  AOI221 U617 ( .A(n8), .B(regs[102]), .C(n1784), .D(regs[38]), .Q(n1229) );
  AOI221 U618 ( .A(n12), .B(regs[327]), .C(n24), .D(regs[263]), .Q(n1240) );
  AOI221 U619 ( .A(n12), .B(regs[70]), .C(n24), .D(regs[6]), .Q(n1228) );
  AOI221 U620 ( .A(n12), .B(regs[840]), .C(n24), .D(regs[776]), .Q(n1258) );
  OAI211 U621 ( .A(n187), .B(n49), .C(n1002), .Q(n1003) );
  OAI211 U622 ( .A(n83), .B(n49), .C(n462), .Q(n463) );
  AOI221 U623 ( .A(n8), .B(regs[107]), .C(n1784), .D(regs[43]), .Q(n1339) );
  OAI211 U624 ( .A(n76), .B(n49), .C(n367), .Q(n368) );
  OAI211 U625 ( .A(n135), .B(n49), .C(n452), .Q(n453) );
  AOI221 U626 ( .A(n46), .B(regs[465]), .C(n52), .D(regs[401]), .Q(n1462) );
  AOI221 U627 ( .A(n46), .B(regs[464]), .C(n52), .D(regs[400]), .Q(n1440) );
  OAI211 U628 ( .A(n75), .B(n49), .C(n362), .Q(n363) );
  AOI221 U629 ( .A(n46), .B(regs[721]), .C(n52), .D(regs[657]), .Q(n1468) );
  AOI221 U630 ( .A(n8), .B(regs[362]), .C(n48), .D(regs[298]), .Q(n1307) );
  AOI221 U631 ( .A(n8), .B(regs[614]), .C(n48), .D(regs[550]), .Q(n1225) );
  AOI221 U632 ( .A(n8), .B(regs[872]), .C(n48), .D(regs[808]), .Q(n1259) );
  AOI221 U633 ( .A(n8), .B(regs[105]), .C(n1784), .D(regs[41]), .Q(n1295) );
  OAI211 U634 ( .A(n131), .B(n49), .C(n402), .Q(n403) );
  OAI211 U635 ( .A(n84), .B(n49), .C(n467), .Q(n468) );
  OAI211 U636 ( .A(n137), .B(n49), .C(n477), .Q(n478) );
  AOI221 U637 ( .A(n8), .B(regs[377]), .C(n48), .D(regs[313]), .Q(n1637) );
  OAI211 U638 ( .A(n116), .B(n49), .C(n937), .Q(n938) );
  AOI221 U639 ( .A(n8), .B(regs[870]), .C(n48), .D(regs[806]), .Q(n1215) );
  OAI211 U640 ( .A(n85), .B(n49), .C(n487), .Q(n488) );
  OAI211 U641 ( .A(n133), .B(n49), .C(n427), .Q(n428) );
  OAI211 U642 ( .A(n136), .B(n49), .C(n472), .Q(n473) );
  OAI211 U643 ( .A(n80), .B(n49), .C(n417), .Q(n418) );
  OAI211 U644 ( .A(n171), .B(n49), .C(n872), .Q(n873) );
  OAI211 U645 ( .A(n128), .B(n49), .C(n372), .Q(n373) );
  AOI221 U646 ( .A(n12), .B(regs[328]), .C(n24), .D(regs[264]), .Q(n1262) );
  OAI211 U647 ( .A(n79), .B(n49), .C(n412), .Q(n413) );
  AOI221 U648 ( .A(n46), .B(regs[209]), .C(n52), .D(regs[145]), .Q(n1472) );
  AOI221 U649 ( .A(n46), .B(regs[720]), .C(n52), .D(regs[656]), .Q(n1446) );
  AOI221 U650 ( .A(n46), .B(regs[978]), .C(n52), .D(regs[914]), .Q(n1480) );
  OAI211 U651 ( .A(n181), .B(n49), .C(n952), .Q(n953) );
  OAI211 U652 ( .A(n117), .B(n49), .C(n962), .Q(n963) );
  AOI221 U653 ( .A(n12), .B(regs[843]), .C(n24), .D(regs[779]), .Q(n1324) );
  AOI221 U654 ( .A(n12), .B(regs[842]), .C(n24), .D(regs[778]), .Q(n1302) );
  OAI211 U655 ( .A(n184), .B(n49), .C(n977), .Q(n978) );
  AOI221 U656 ( .A(n12), .B(regs[841]), .C(n24), .D(regs[777]), .Q(n1280) );
  OAI211 U657 ( .A(n179), .B(n49), .C(n942), .Q(n943) );
  AOI221 U658 ( .A(n12), .B(regs[605]), .C(n24), .D(regs[541]), .Q(n1730) );
  AOI221 U659 ( .A(n12), .B(regs[349]), .C(n24), .D(regs[285]), .Q(n1724) );
  AOI221 U660 ( .A(n12), .B(regs[601]), .C(n24), .D(regs[537]), .Q(n1642) );
  AOI221 U661 ( .A(n47), .B(regs[60]), .C(n19), .D(regs[28]), .Q(n975) );
  AOI221 U662 ( .A(n14), .B(regs[767]), .C(n10), .D(regs[703]), .Q(n1779) );
  AOI221 U663 ( .A(n12), .B(regs[860]), .C(n24), .D(regs[796]), .Q(n1698) );
  AOI221 U664 ( .A(regs[736]), .B(n14), .C(regs[672]), .D(n10), .Q(n1095) );
  AOI221 U665 ( .A(n12), .B(regs[603]), .C(n24), .D(regs[539]), .Q(n1686) );
  AOI221 U666 ( .A(n12), .B(regs[93]), .C(n24), .D(regs[29]), .Q(n1734) );
  AOI221 U667 ( .A(n12), .B(regs[861]), .C(n24), .D(regs[797]), .Q(n1720) );
  AOI221 U668 ( .A(regs[576]), .B(n12), .C(regs[512]), .D(n24), .Q(n1092) );
  AOI221 U669 ( .A(n47), .B(regs[553]), .C(n19), .D(regs[521]), .Q(n505) );
  AOI221 U670 ( .A(n12), .B(regs[858]), .C(n24), .D(regs[794]), .Q(n1654) );
  AOI221 U671 ( .A(n12), .B(regs[91]), .C(n24), .D(regs[27]), .Q(n1690) );
  AOI221 U672 ( .A(n12), .B(regs[90]), .C(n24), .D(regs[26]), .Q(n1668) );
  AOI221 U673 ( .A(n47), .B(regs[554]), .C(n19), .D(regs[522]), .Q(n530) );
  AOI221 U674 ( .A(n12), .B(regs[92]), .C(n24), .D(regs[28]), .Q(n1712) );
  AOI221 U675 ( .A(n14), .B(regs[511]), .C(n10), .D(regs[447]), .Q(n1771) );
  AOI221 U676 ( .A(n12), .B(regs[859]), .C(n24), .D(regs[795]), .Q(n1676) );
  AOI221 U677 ( .A(n47), .B(regs[42]), .C(n19), .D(regs[10]), .Q(n525) );
  AOI221 U678 ( .A(n47), .B(regs[41]), .C(n19), .D(regs[9]), .Q(n500) );
  AOI221 U679 ( .A(n12), .B(regs[602]), .C(n24), .D(regs[538]), .Q(n1664) );
  AOI221 U680 ( .A(n12), .B(regs[857]), .C(n24), .D(regs[793]), .Q(n1632) );
  AOI221 U681 ( .A(n14), .B(regs[1023]), .C(n10), .D(regs[959]), .Q(n1767) );
  AOI221 U682 ( .A(n12), .B(regs[862]), .C(n24), .D(regs[798]), .Q(n1742) );
  AOI221 U683 ( .A(n14), .B(regs[510]), .C(n10), .D(regs[446]), .Q(n1749) );
  AOI221 U684 ( .A(n12), .B(regs[604]), .C(n24), .D(regs[540]), .Q(n1708) );
  AOI221 U685 ( .A(n14), .B(regs[766]), .C(n10), .D(regs[702]), .Q(n1755) );
  AOI221 U686 ( .A(n47), .B(regs[810]), .C(n19), .D(regs[778]), .Q(n520) );
  AOI221 U687 ( .A(n47), .B(regs[570]), .C(n19), .D(regs[538]), .Q(n930) );
  AOI221 U688 ( .A(n14), .B(regs[254]), .C(n10), .D(regs[190]), .Q(n1759) );
  AOI221 U689 ( .A(n47), .B(regs[315]), .C(n19), .D(regs[283]), .Q(n940) );
  AOI221 U690 ( .A(n12), .B(regs[348]), .C(n24), .D(regs[284]), .Q(n1702) );
  AOI221 U691 ( .A(n12), .B(regs[345]), .C(n24), .D(regs[281]), .Q(n1636) );
  AOI221 U692 ( .A(n47), .B(regs[809]), .C(n19), .D(regs[777]), .Q(n495) );
  AOI221 U693 ( .A(n8), .B(regs[119]), .C(n48), .D(regs[55]), .Q(n1603) );
  AOI221 U694 ( .A(n47), .B(regs[314]), .C(n19), .D(regs[282]), .Q(n915) );
  AOI221 U695 ( .A(n47), .B(regs[551]), .C(n19), .D(regs[519]), .Q(n455) );
  AOI221 U696 ( .A(n8), .B(regs[631]), .C(n48), .D(regs[567]), .Q(n1599) );
  AOI221 U697 ( .A(n47), .B(regs[39]), .C(n19), .D(regs[7]), .Q(n450) );
  AOI221 U698 ( .A(n47), .B(regs[811]), .C(n19), .D(regs[779]), .Q(n545) );
  AOI221 U699 ( .A(n47), .B(regs[807]), .C(n19), .D(regs[775]), .Q(n445) );
  AOI221 U700 ( .A(n47), .B(regs[813]), .C(n19), .D(regs[781]), .Q(n595) );
  AOI221 U701 ( .A(n8), .B(regs[375]), .C(n48), .D(regs[311]), .Q(n1593) );
  AOI221 U702 ( .A(n47), .B(regs[295]), .C(n19), .D(regs[263]), .Q(n440) );
  AOI221 U703 ( .A(n47), .B(regs[812]), .C(n19), .D(regs[780]), .Q(n570) );
  AOI221 U704 ( .A(n47), .B(regs[552]), .C(n19), .D(regs[520]), .Q(n480) );
  AOI221 U705 ( .A(n8), .B(regs[887]), .C(n48), .D(regs[823]), .Q(n1589) );
  AOI221 U706 ( .A(n47), .B(regs[301]), .C(n19), .D(regs[269]), .Q(n590) );
  AOI221 U707 ( .A(n8), .B(regs[372]), .C(n48), .D(regs[308]), .Q(n1527) );
  AOI221 U708 ( .A(n47), .B(regs[575]), .C(n19), .D(regs[543]), .Q(n1066) );
  AOI221 U709 ( .A(n8), .B(regs[885]), .C(n48), .D(regs[821]), .Q(n1545) );
  AOI221 U710 ( .A(n47), .B(regs[318]), .C(n19), .D(regs[286]), .Q(n1015) );
  AOI221 U711 ( .A(n47), .B(regs[573]), .C(n19), .D(regs[541]), .Q(n1005) );
  AOI221 U712 ( .A(n47), .B(regs[830]), .C(n19), .D(regs[798]), .Q(n1020) );
  AOI221 U713 ( .A(n8), .B(regs[373]), .C(n48), .D(regs[309]), .Q(n1549) );
  AOI221 U714 ( .A(n47), .B(regs[568]), .C(n19), .D(regs[536]), .Q(n880) );
  AOI221 U715 ( .A(n47), .B(regs[57]), .C(n19), .D(regs[25]), .Q(n900) );
  AOI221 U716 ( .A(n8), .B(regs[118]), .C(n48), .D(regs[54]), .Q(n1581) );
  AOI221 U717 ( .A(n47), .B(regs[300]), .C(n19), .D(regs[268]), .Q(n565) );
  AOI221 U718 ( .A(n8), .B(regs[629]), .C(n48), .D(regs[565]), .Q(n1555) );
  AOI221 U719 ( .A(n8), .B(regs[630]), .C(n48), .D(regs[566]), .Q(n1577) );
  AOI221 U720 ( .A(n8), .B(regs[374]), .C(n48), .D(regs[310]), .Q(n1571) );
  AOI221 U721 ( .A(n8), .B(regs[886]), .C(n48), .D(regs[822]), .Q(n1567) );
  AOI221 U722 ( .A(n8), .B(regs[117]), .C(n48), .D(regs[53]), .Q(n1559) );
  AOI221 U723 ( .A(n47), .B(regs[574]), .C(n19), .D(regs[542]), .Q(n1030) );
  AOI221 U724 ( .A(n47), .B(regs[296]), .C(n19), .D(regs[264]), .Q(n465) );
  AOI221 U725 ( .A(n47), .B(regs[61]), .C(n19), .D(regs[29]), .Q(n1000) );
  AOI221 U726 ( .A(n47), .B(regs[291]), .C(n19), .D(regs[259]), .Q(n340) );
  AOI221 U727 ( .A(n8), .B(regs[888]), .C(n48), .D(regs[824]), .Q(n1611) );
  AOI221 U728 ( .A(n47), .B(regs[825]), .C(n19), .D(regs[793]), .Q(n895) );
  AOI221 U729 ( .A(n12), .B(regs[344]), .C(n24), .D(regs[280]), .Q(n1614) );
  AOI221 U730 ( .A(n47), .B(regs[35]), .C(n19), .D(regs[3]), .Q(n350) );
  AOI221 U731 ( .A(n47), .B(regs[829]), .C(n19), .D(regs[797]), .Q(n995) );
  AOI221 U732 ( .A(n47), .B(regs[808]), .C(n19), .D(regs[776]), .Q(n470) );
  AOI221 U733 ( .A(n8), .B(regs[883]), .C(n48), .D(regs[819]), .Q(n1501) );
  AOI221 U734 ( .A(n8), .B(regs[628]), .C(n48), .D(regs[564]), .Q(n1533) );
  AOI221 U735 ( .A(n12), .B(regs[600]), .C(n24), .D(regs[536]), .Q(n1620) );
  AOI221 U736 ( .A(n47), .B(regs[547]), .C(n19), .D(regs[515]), .Q(n355) );
  AOI221 U737 ( .A(n47), .B(regs[44]), .C(n19), .D(regs[12]), .Q(n575) );
  AOI221 U738 ( .A(n8), .B(regs[116]), .C(n48), .D(regs[52]), .Q(n1537) );
  AOI221 U739 ( .A(n47), .B(regs[46]), .C(n19), .D(regs[14]), .Q(n625) );
  AOI221 U740 ( .A(n12), .B(regs[89]), .C(n24), .D(regs[25]), .Q(n1646) );
  AOI221 U741 ( .A(n14), .B(regs[992]), .C(n10), .D(regs[928]), .Q(n1083) );
  AOI221 U742 ( .A(n8), .B(regs[371]), .C(n48), .D(regs[307]), .Q(n1505) );
  AOI221 U743 ( .A(n47), .B(regs[555]), .C(n19), .D(regs[523]), .Q(n555) );
  AOI221 U744 ( .A(n47), .B(regs[59]), .C(n19), .D(regs[27]), .Q(n950) );
  AOI221 U745 ( .A(n47), .B(regs[556]), .C(n19), .D(regs[524]), .Q(n580) );
  AOI221 U746 ( .A(n12), .B(regs[88]), .C(n24), .D(regs[24]), .Q(n1624) );
  AOI221 U747 ( .A(n47), .B(regs[569]), .C(n19), .D(regs[537]), .Q(n905) );
  INV2 U748 ( .A(i_con_RegWr), .Q(n1811) );
  NAND33 U749 ( .A(i_con_RegWr), .B(i_addr_Rd[4]), .C(i_addr_Rd[3]), .Q(n1814)
         );
  AOI221 U750 ( .A(n45), .B(regs[352]), .C(n51), .D(regs[480]), .Q(n276) );
  AOI221 U751 ( .A(n14), .B(regs[1017]), .C(n10), .D(regs[953]), .Q(n1635) );
  AOI221 U752 ( .A(n14), .B(regs[495]), .C(n10), .D(regs[431]), .Q(n1419) );
  AOI221 U753 ( .A(n12), .B(regs[847]), .C(n24), .D(regs[783]), .Q(n1412) );
  AOI221 U754 ( .A(n14), .B(regs[1009]), .C(n10), .D(regs[945]), .Q(n1459) );
  AOI221 U755 ( .A(n12), .B(regs[848]), .C(n24), .D(regs[784]), .Q(n1434) );
  AOI221 U756 ( .A(n14), .B(regs[1008]), .C(n10), .D(regs[944]), .Q(n1437) );
  AOI221 U757 ( .A(n12), .B(regs[320]), .C(n24), .D(regs[256]), .Q(n1085) );
  AOI221 U758 ( .A(n46), .B(regs[467]), .C(n50), .D(regs[403]), .Q(n1506) );
  AOI221 U759 ( .A(n12), .B(regs[333]), .C(n24), .D(regs[269]), .Q(n1372) );
  AOI221 U760 ( .A(n12), .B(regs[845]), .C(n24), .D(regs[781]), .Q(n1368) );
  AOI221 U761 ( .A(n12), .B(regs[78]), .C(n24), .D(regs[14]), .Q(n1404) );
  AOI221 U762 ( .A(n12), .B(regs[584]), .C(n24), .D(regs[520]), .Q(n1268) );
  AOI221 U763 ( .A(n12), .B(regs[586]), .C(n24), .D(regs[522]), .Q(n1312) );
  AOI221 U764 ( .A(n14), .B(regs[1002]), .C(n10), .D(regs[938]), .Q(n1305) );
  AOI221 U765 ( .A(n12), .B(regs[73]), .C(n24), .D(regs[9]), .Q(n1294) );
  AOI221 U766 ( .A(n14), .B(regs[1001]), .C(n10), .D(regs[937]), .Q(n1283) );
  AOI221 U767 ( .A(n8), .B(regs[97]), .C(n48), .D(regs[33]), .Q(n1119) );
  AOI221 U768 ( .A(n12), .B(regs[321]), .C(n24), .D(regs[257]), .Q(n1108) );
  AOI221 U769 ( .A(n8), .B(regs[865]), .C(n48), .D(regs[801]), .Q(n1105) );
  AOI221 U770 ( .A(n12), .B(regs[587]), .C(n24), .D(regs[523]), .Q(n1334) );
  AOI221 U771 ( .A(n8), .B(regs[639]), .C(n48), .D(regs[575]), .Q(n1777) );
  AOI221 U772 ( .A(n8), .B(regs[895]), .C(n48), .D(regs[831]), .Q(n1765) );
  AOI221 U773 ( .A(n46), .B(regs[991]), .C(n50), .D(regs[927]), .Q(n1766) );
  AOI221 U774 ( .A(n8), .B(regs[101]), .C(n48), .D(regs[37]), .Q(n1207) );
  AOI221 U775 ( .A(n8), .B(regs[613]), .C(n48), .D(regs[549]), .Q(n1203) );
  AOI221 U776 ( .A(n8), .B(regs[869]), .C(n48), .D(regs[805]), .Q(n1193) );
  AOI221 U777 ( .A(n12), .B(regs[836]), .C(n24), .D(regs[772]), .Q(n1170) );
  AOI221 U778 ( .A(n14), .B(regs[504]), .C(n10), .D(regs[440]), .Q(n1617) );
  AOI221 U779 ( .A(n12), .B(regs[66]), .C(n24), .D(regs[2]), .Q(n1140) );
  AOI221 U780 ( .A(n12), .B(regs[322]), .C(n24), .D(regs[258]), .Q(n1130) );
  AOI221 U781 ( .A(n46), .B(regs[450]), .C(n52), .D(regs[386]), .Q(n1132) );
  AOI221 U782 ( .A(n12), .B(regs[834]), .C(n24), .D(regs[770]), .Q(n1126) );
  AOI221 U783 ( .A(n12), .B(regs[323]), .C(n24), .D(regs[259]), .Q(n1152) );
  AOI221 U784 ( .A(n12), .B(regs[835]), .C(n24), .D(regs[771]), .Q(n1148) );
  AOI221 U785 ( .A(n14), .B(regs[1018]), .C(n10), .D(regs[954]), .Q(n1657) );
  AOI221 U786 ( .A(n12), .B(regs[839]), .C(n24), .D(regs[775]), .Q(n1236) );
  AOI221 U787 ( .A(n46), .B(regs[454]), .C(n52), .D(regs[390]), .Q(n1220) );
  AOI221 U788 ( .A(n14), .B(regs[486]), .C(n10), .D(regs[422]), .Q(n1221) );
  AOI221 U789 ( .A(n47), .B(regs[804]), .C(n19), .D(regs[772]), .Q(n370) );
  AOI221 U790 ( .A(n47), .B(regs[292]), .C(n19), .D(regs[260]), .Q(n365) );
  AOI221 U791 ( .A(n33), .B(regs[193]), .C(n7), .D(regs[129]), .Q(n309) );
  AOI221 U792 ( .A(n45), .B(regs[97]), .C(n1), .D(regs[225]), .Q(n307) );
  AOI221 U793 ( .A(n33), .B(regs[705]), .C(n7), .D(regs[641]), .Q(n304) );
  AOI221 U794 ( .A(n33), .B(regs[449]), .C(n7), .D(regs[385]), .Q(n299) );
  AOI221 U795 ( .A(n33), .B(regs[961]), .C(n7), .D(regs[897]), .Q(n294) );
  AOI221 U796 ( .A(n8), .B(regs[638]), .C(n48), .D(regs[574]), .Q(n1753) );
  AOI221 U797 ( .A(n46), .B(regs[471]), .C(n50), .D(regs[407]), .Q(n1594) );
  AOI221 U798 ( .A(n46), .B(regs[470]), .C(n50), .D(regs[406]), .Q(n1572) );
  AOI221 U799 ( .A(n46), .B(regs[982]), .C(n50), .D(regs[918]), .Q(n1568) );
  AOI221 U800 ( .A(n33), .B(regs[723]), .C(n7), .D(regs[659]), .Q(n756) );
  AOI221 U801 ( .A(n47), .B(regs[312]), .C(n19), .D(regs[280]), .Q(n865) );
  AOI221 U802 ( .A(n47), .B(regs[55]), .C(n19), .D(regs[23]), .Q(n850) );
  AOI221 U803 ( .A(n47), .B(regs[823]), .C(n19), .D(regs[791]), .Q(n845) );
  AOI221 U804 ( .A(n47), .B(regs[311]), .C(n19), .D(regs[279]), .Q(n840) );
  AOI221 U805 ( .A(n47), .B(regs[58]), .C(n19), .D(regs[26]), .Q(n925) );
  AOI221 U806 ( .A(n47), .B(regs[826]), .C(n19), .D(regs[794]), .Q(n920) );
  AOI221 U807 ( .A(n47), .B(regs[546]), .C(n19), .D(regs[514]), .Q(n330) );
  AOI221 U808 ( .A(n47), .B(regs[34]), .C(n19), .D(regs[2]), .Q(n325) );
  AOI221 U809 ( .A(n47), .B(regs[802]), .C(n19), .D(regs[770]), .Q(n320) );
  AOI221 U810 ( .A(n47), .B(regs[290]), .C(n19), .D(regs[258]), .Q(n315) );
  AOI221 U811 ( .A(n45), .B(regs[638]), .C(n199), .D(regs[766]), .Q(n1027) );
  AOI221 U812 ( .A(n45), .B(regs[639]), .C(n199), .D(regs[767]), .Q(n1060) );
  AOI221 U813 ( .A(n47), .B(regs[313]), .C(n19), .D(regs[281]), .Q(n890) );
  AOI221 U814 ( .A(n47), .B(regs[45]), .C(n19), .D(regs[13]), .Q(n600) );
  AOI221 U815 ( .A(n47), .B(regs[43]), .C(n19), .D(regs[11]), .Q(n550) );
  AOI221 U816 ( .A(n47), .B(regs[297]), .C(n19), .D(regs[265]), .Q(n490) );
  AOI221 U817 ( .A(n47), .B(regs[817]), .C(n19), .D(regs[785]), .Q(n695) );
  AOI221 U818 ( .A(n47), .B(regs[305]), .C(n19), .D(regs[273]), .Q(n690) );
  AOI221 U819 ( .A(n14), .B(regs[1007]), .C(n10), .D(regs[943]), .Q(n1415) );
  AOI221 U820 ( .A(n12), .B(regs[337]), .C(n24), .D(regs[273]), .Q(n1460) );
  AOI221 U821 ( .A(n12), .B(regs[849]), .C(n24), .D(regs[785]), .Q(n1456) );
  AOI221 U822 ( .A(n12), .B(regs[336]), .C(n24), .D(regs[272]), .Q(n1438) );
  AOI221 U823 ( .A(n12), .B(regs[338]), .C(n24), .D(regs[274]), .Q(n1482) );
  AOI221 U824 ( .A(n12), .B(regs[850]), .C(n24), .D(regs[786]), .Q(n1478) );
  AOI221 U825 ( .A(n12), .B(regs[339]), .C(n24), .D(regs[275]), .Q(n1504) );
  AOI221 U826 ( .A(n12), .B(regs[851]), .C(n24), .D(regs[787]), .Q(n1500) );
  AOI221 U827 ( .A(n14), .B(regs[1005]), .C(n10), .D(regs[941]), .Q(n1371) );
  AOI221 U828 ( .A(n12), .B(regs[334]), .C(n24), .D(regs[270]), .Q(n1394) );
  AOI221 U829 ( .A(n12), .B(regs[846]), .C(n24), .D(regs[782]), .Q(n1390) );
  AOI221 U830 ( .A(n12), .B(regs[72]), .C(n24), .D(regs[8]), .Q(n1272) );
  AOI221 U831 ( .A(n14), .B(regs[234]), .C(n10), .D(regs[170]), .Q(n1319) );
  AOI221 U832 ( .A(n14), .B(regs[746]), .C(n10), .D(regs[682]), .Q(n1315) );
  AOI221 U833 ( .A(n14), .B(regs[490]), .C(n10), .D(regs[426]), .Q(n1309) );
  AOI221 U834 ( .A(n12), .B(regs[577]), .C(n24), .D(regs[513]), .Q(n1114) );
  AOI221 U835 ( .A(n14), .B(regs[748]), .C(n10), .D(regs[684]), .Q(n1359) );
  AOI221 U836 ( .A(n14), .B(regs[492]), .C(n10), .D(regs[428]), .Q(n1353) );
  AOI221 U837 ( .A(n14), .B(regs[1004]), .C(n10), .D(regs[940]), .Q(n1349) );
  AOI221 U838 ( .A(n14), .B(regs[235]), .C(n10), .D(regs[171]), .Q(n1341) );
  AOI221 U839 ( .A(n14), .B(regs[747]), .C(n10), .D(regs[683]), .Q(n1337) );
  AOI221 U840 ( .A(n14), .B(regs[491]), .C(n10), .D(regs[427]), .Q(n1331) );
  AOI221 U841 ( .A(n14), .B(regs[1003]), .C(n10), .D(regs[939]), .Q(n1327) );
  AOI221 U842 ( .A(n14), .B(regs[485]), .C(n10), .D(regs[421]), .Q(n1199) );
  AOI221 U843 ( .A(n14), .B(regs[997]), .C(n10), .D(regs[933]), .Q(n1195) );
  AOI221 U844 ( .A(n8), .B(regs[612]), .C(n48), .D(regs[548]), .Q(n1181) );
  AOI221 U845 ( .A(n14), .B(regs[248]), .C(n10), .D(regs[184]), .Q(n1627) );
  AOI221 U846 ( .A(n12), .B(regs[578]), .C(n24), .D(regs[514]), .Q(n1136) );
  AOI221 U847 ( .A(n12), .B(regs[67]), .C(n24), .D(regs[3]), .Q(n1162) );
  AOI221 U848 ( .A(n12), .B(regs[579]), .C(n24), .D(regs[515]), .Q(n1158) );
  AOI221 U849 ( .A(n14), .B(regs[762]), .C(n10), .D(regs[698]), .Q(n1667) );
  AOI221 U850 ( .A(n14), .B(regs[507]), .C(n10), .D(regs[443]), .Q(n1683) );
  AOI221 U851 ( .A(n14), .B(regs[1019]), .C(n10), .D(regs[955]), .Q(n1679) );
  AOI221 U852 ( .A(n12), .B(regs[582]), .C(n24), .D(regs[518]), .Q(n1224) );
  AOI221 U853 ( .A(n14), .B(regs[998]), .C(n10), .D(regs[934]), .Q(n1217) );
  AOI221 U854 ( .A(n12), .B(regs[852]), .C(n24), .D(regs[788]), .Q(n1522) );
  AOI221 U855 ( .A(n12), .B(regs[81]), .C(n24), .D(regs[17]), .Q(n1470) );
  AOI221 U856 ( .A(n12), .B(regs[80]), .C(n24), .D(regs[16]), .Q(n1448) );
  AOI221 U857 ( .A(n14), .B(regs[240]), .C(n10), .D(regs[176]), .Q(n1451) );
  AOI221 U858 ( .A(n12), .B(regs[82]), .C(n24), .D(regs[18]), .Q(n1492) );
  AOI221 U859 ( .A(n12), .B(regs[64]), .C(n24), .D(regs[0]), .Q(n1096) );
  AOI221 U860 ( .A(n46), .B(regs[712]), .C(n50), .D(regs[648]), .Q(n1270) );
  AOI221 U861 ( .A(n12), .B(regs[585]), .C(n24), .D(regs[521]), .Q(n1290) );
  AOI221 U862 ( .A(n14), .B(regs[489]), .C(n10), .D(regs[425]), .Q(n1287) );
  AOI221 U863 ( .A(n12), .B(regs[65]), .C(n24), .D(regs[1]), .Q(n1118) );
  AOI221 U864 ( .A(n12), .B(regs[833]), .C(n24), .D(regs[769]), .Q(n1104) );
  AOI221 U865 ( .A(n12), .B(regs[76]), .C(n24), .D(regs[12]), .Q(n1360) );
  AOI221 U866 ( .A(n12), .B(regs[69]), .C(n24), .D(regs[5]), .Q(n1206) );
  AOI221 U867 ( .A(n12), .B(regs[581]), .C(n24), .D(regs[517]), .Q(n1202) );
  AOI221 U868 ( .A(n12), .B(regs[325]), .C(n24), .D(regs[261]), .Q(n1196) );
  AOI221 U869 ( .A(n12), .B(regs[837]), .C(n24), .D(regs[773]), .Q(n1192) );
  AOI221 U870 ( .A(n12), .B(regs[68]), .C(n24), .D(regs[4]), .Q(n1184) );
  AOI221 U871 ( .A(n14), .B(regs[250]), .C(n10), .D(regs[186]), .Q(n1671) );
  AOI221 U872 ( .A(n12), .B(regs[71]), .C(n24), .D(regs[7]), .Q(n1250) );
  AOI221 U873 ( .A(n12), .B(regs[326]), .C(n24), .D(regs[262]), .Q(n1218) );
  AOI221 U874 ( .A(n12), .B(regs[838]), .C(n24), .D(regs[774]), .Q(n1214) );
  AOI221 U875 ( .A(n33), .B(regs[734]), .C(n7), .D(regs[670]), .Q(n1031) );
  AOI221 U876 ( .A(n14), .B(regs[241]), .C(n10), .D(regs[177]), .Q(n1473) );
  AOI221 U877 ( .A(n46), .B(regs[200]), .C(n50), .D(regs[136]), .Q(n1274) );
  AOI221 U878 ( .A(n46), .B(regs[196]), .C(n52), .D(regs[132]), .Q(n1186) );
  AOI221 U879 ( .A(n12), .B(regs[580]), .C(n24), .D(regs[516]), .Q(n1180) );
  AOI221 U880 ( .A(n14), .B(regs[760]), .C(n10), .D(regs[696]), .Q(n1623) );
  AOI221 U881 ( .A(n46), .B(regs[713]), .C(n50), .D(regs[649]), .Q(n1292) );
  AOI221 U882 ( .A(n14), .B(regs[225]), .C(n10), .D(regs[161]), .Q(n1121) );
  AOI221 U883 ( .A(n14), .B(regs[737]), .C(n10), .D(regs[673]), .Q(n1117) );
  AOI221 U884 ( .A(n12), .B(regs[588]), .C(n24), .D(regs[524]), .Q(n1356) );
  AOI221 U885 ( .A(n14), .B(regs[227]), .C(n10), .D(regs[163]), .Q(n1165) );
  AOI221 U886 ( .A(n46), .B(regs[711]), .C(n52), .D(regs[647]), .Q(n1248) );
  AOI221 U887 ( .A(n12), .B(regs[599]), .C(n24), .D(regs[535]), .Q(n1598) );
  AOI221 U888 ( .A(n8), .B(regs[96]), .C(n48), .D(regs[32]), .Q(n1097) );
  AOI221 U889 ( .A(n12), .B(regs[598]), .C(n24), .D(regs[534]), .Q(n1576) );
  AOI221 U890 ( .A(n1775), .B(n1377), .C(n1773), .D(n1376), .Q(n1389) );
  AOI221 U891 ( .A(n1775), .B(n1399), .C(n1773), .D(n1398), .Q(n1411) );
  AOI221 U892 ( .A(n1775), .B(n1311), .C(n1773), .D(n1310), .Q(n1323) );
  AOI221 U893 ( .A(n1775), .B(n1289), .C(n1773), .D(n1288), .Q(n1301) );
  AOI221 U894 ( .A(n1775), .B(n1113), .C(n1773), .D(n1112), .Q(n1125) );
  AOI221 U895 ( .A(n1775), .B(n1355), .C(n1773), .D(n1354), .Q(n1367) );
  AOI221 U896 ( .A(n1775), .B(n1333), .C(n1773), .D(n1332), .Q(n1345) );
  AOI221 U897 ( .A(n1775), .B(n1201), .C(n1773), .D(n1200), .Q(n1213) );
  AOI221 U898 ( .A(n1775), .B(n1135), .C(n1773), .D(n1134), .Q(n1147) );
  AOI221 U899 ( .A(n1775), .B(n1245), .C(n1773), .D(n1244), .Q(n1257) );
  AOI221 U900 ( .A(n45), .B(regs[353]), .C(n51), .D(regs[481]), .Q(n297) );
  AOI221 U901 ( .A(n45), .B(regs[865]), .C(n51), .D(regs[993]), .Q(n292) );
  AOI221 U902 ( .A(n45), .B(regs[635]), .C(n1), .D(regs[763]), .Q(n952) );
  AOI221 U903 ( .A(n45), .B(regs[123]), .C(n1), .D(regs[251]), .Q(n947) );
  AOI221 U904 ( .A(n45), .B(regs[891]), .C(n1), .D(regs[1019]), .Q(n942) );
  AOI221 U905 ( .A(n45), .B(regs[379]), .C(n1), .D(regs[507]), .Q(n937) );
  AOI221 U906 ( .A(n45), .B(regs[632]), .C(n1), .D(regs[760]), .Q(n877) );
  AOI221 U907 ( .A(n45), .B(regs[637]), .C(n1), .D(regs[765]), .Q(n1002) );
  AOI221 U908 ( .A(n45), .B(regs[125]), .C(n1), .D(regs[253]), .Q(n997) );
  AOI221 U909 ( .A(n45), .B(regs[893]), .C(n1), .D(regs[1021]), .Q(n992) );
  AOI221 U910 ( .A(n45), .B(regs[381]), .C(n1), .D(regs[509]), .Q(n987) );
  AOI221 U911 ( .A(n45), .B(regs[636]), .C(n1), .D(regs[764]), .Q(n977) );
  AOI221 U912 ( .A(n45), .B(regs[124]), .C(n1), .D(regs[252]), .Q(n972) );
  AOI221 U913 ( .A(n45), .B(regs[892]), .C(n1), .D(regs[1020]), .Q(n967) );
  AOI221 U914 ( .A(n45), .B(regs[380]), .C(n1), .D(regs[508]), .Q(n962) );
  AOI221 U915 ( .A(n45), .B(regs[383]), .C(n1), .D(regs[511]), .Q(n1037) );
  AOI221 U916 ( .A(n45), .B(regs[633]), .C(n1), .D(regs[761]), .Q(n902) );
  AOI221 U917 ( .A(n45), .B(regs[630]), .C(n1), .D(regs[758]), .Q(n827) );
  AOI221 U918 ( .A(n45), .B(regs[118]), .C(n1), .D(regs[246]), .Q(n822) );
  AOI221 U919 ( .A(n45), .B(regs[886]), .C(n1), .D(regs[1014]), .Q(n817) );
  AOI221 U920 ( .A(n1795), .B(n1651), .C(n1793), .D(n1650), .Q(n1652) );
  AOI221 U921 ( .A(n1795), .B(n1431), .C(n1793), .D(n1430), .Q(n1432) );
  AOI221 U922 ( .A(n1795), .B(n1475), .C(n1793), .D(n1474), .Q(n1476) );
  AOI221 U923 ( .A(n1795), .B(n1453), .C(n1793), .D(n1452), .Q(n1454) );
  AOI221 U924 ( .A(n1795), .B(n1497), .C(n1793), .D(n1496), .Q(n1498) );
  AOI220 U925 ( .A(n1781), .B(regs[498]), .C(n10), .D(regs[434]), .Q(n1485) );
  AOI221 U926 ( .A(n1795), .B(n1101), .C(n1793), .D(n1100), .Q(n1102) );
  AOI221 U927 ( .A(n1795), .B(n1519), .C(n1793), .D(n1518), .Q(n1520) );
  AOI220 U928 ( .A(n1781), .B(regs[499]), .C(n10), .D(regs[435]), .Q(n1507) );
  AOI221 U929 ( .A(n1795), .B(n1387), .C(n1793), .D(n1386), .Q(n1388) );
  AOI221 U930 ( .A(n1795), .B(n1409), .C(n1793), .D(n1408), .Q(n1410) );
  AOI221 U931 ( .A(n1795), .B(n1277), .C(n1793), .D(n1276), .Q(n1278) );
  AOI221 U932 ( .A(n1795), .B(n1321), .C(n1793), .D(n1320), .Q(n1322) );
  AOI221 U933 ( .A(n1795), .B(n1299), .C(n1793), .D(n1298), .Q(n1300) );
  AOI221 U934 ( .A(n1795), .B(n1123), .C(n1793), .D(n1122), .Q(n1124) );
  AOI221 U935 ( .A(n1795), .B(n1365), .C(n1793), .D(n1364), .Q(n1366) );
  AOI221 U936 ( .A(n1795), .B(n1343), .C(n1793), .D(n1342), .Q(n1344) );
  AOI221 U937 ( .A(n1795), .B(n1794), .C(n1793), .D(n1792), .Q(n1796) );
  AOI221 U938 ( .A(n1795), .B(n1211), .C(n1793), .D(n1210), .Q(n1212) );
  AOI221 U939 ( .A(n1795), .B(n1189), .C(n1793), .D(n1188), .Q(n1190) );
  AOI221 U940 ( .A(n1795), .B(n1629), .C(n1793), .D(n1628), .Q(n1630) );
  AOI221 U941 ( .A(n1795), .B(n1145), .C(n1793), .D(n1144), .Q(n1146) );
  AOI221 U942 ( .A(n1795), .B(n1167), .C(n1793), .D(n1166), .Q(n1168) );
  AOI221 U943 ( .A(n1795), .B(n1673), .C(n1793), .D(n1672), .Q(n1674) );
  AOI221 U944 ( .A(n1795), .B(n1695), .C(n1793), .D(n1694), .Q(n1696) );
  AOI221 U945 ( .A(n1795), .B(n1739), .C(n1793), .D(n1738), .Q(n1740) );
  AOI221 U946 ( .A(n1795), .B(n1717), .C(n1793), .D(n1716), .Q(n1718) );
  AOI221 U947 ( .A(n1795), .B(n1255), .C(n1793), .D(n1254), .Q(n1256) );
  AOI221 U948 ( .A(n1795), .B(n1233), .C(n1793), .D(n1232), .Q(n1234) );
  AOI221 U949 ( .A(n1074), .B(n1808), .C(n1073), .D(n1807), .Q(n1809) );
  AOI221 U950 ( .A(n198), .B(n1806), .C(n1075), .D(n1805), .Q(n1810) );
  AOI221 U951 ( .A(n1795), .B(n1541), .C(n1793), .D(n1540), .Q(n1542) );
  AOI221 U952 ( .A(n1795), .B(n1563), .C(n1793), .D(n1562), .Q(n1564) );
  AOI221 U953 ( .A(n1795), .B(n1761), .C(n1793), .D(n1760), .Q(n1762) );
  AOI221 U954 ( .A(n1795), .B(n1607), .C(n1793), .D(n1606), .Q(n1608) );
  AOI221 U955 ( .A(n1795), .B(n1585), .C(n1793), .D(n1584), .Q(n1586) );
  NAND22 U956 ( .A(n1804), .B(n1803), .Q(o_data_Rs[0]) );
  AOI221 U957 ( .A(n1074), .B(n1802), .C(n1073), .D(n1801), .Q(n1803) );
  NAND31 U958 ( .A(n291), .B(n290), .C(n289), .Q(n1801) );
  AOI221 U959 ( .A(n33), .B(regs[192]), .C(n7), .D(regs[128]), .Q(n289) );
  AOI211 U960 ( .A(n3), .B(regs[64]), .C(n288), .Q(n291) );
  AOI221 U961 ( .A(n45), .B(regs[96]), .C(n51), .D(regs[224]), .Q(n287) );
  NAND31 U962 ( .A(n286), .B(n285), .C(n284), .Q(n1802) );
  AOI221 U963 ( .A(n33), .B(regs[704]), .C(n7), .D(regs[640]), .Q(n284) );
  AOI211 U964 ( .A(n4), .B(regs[576]), .C(n283), .Q(n286) );
  AOI221 U965 ( .A(n45), .B(regs[608]), .C(n51), .D(regs[736]), .Q(n282) );
  AOI221 U966 ( .A(n198), .B(n1800), .C(n1075), .D(n1799), .Q(n1804) );
  NAND31 U967 ( .A(n280), .B(n279), .C(n278), .Q(n1799) );
  AOI221 U968 ( .A(n33), .B(regs[448]), .C(n7), .D(regs[384]), .Q(n278) );
  AOI211 U969 ( .A(n4), .B(regs[320]), .C(n277), .Q(n280) );
  NAND31 U970 ( .A(n274), .B(n273), .C(n272), .Q(n1800) );
  AOI221 U971 ( .A(n33), .B(regs[960]), .C(n7), .D(regs[896]), .Q(n272) );
  AOI211 U972 ( .A(n4), .B(regs[832]), .C(n265), .Q(n274) );
  AOI221 U973 ( .A(n45), .B(regs[864]), .C(n51), .D(regs[992]), .Q(n264) );
  NAND22 U974 ( .A(n1653), .B(n1652), .Q(o_data_Rt[25]) );
  NAND41 U975 ( .A(n1649), .B(n1648), .C(n1647), .D(n1646), .Q(n1650) );
  AOI221 U976 ( .A(n14), .B(regs[249]), .C(n10), .D(regs[185]), .Q(n1649) );
  NAND41 U977 ( .A(n1645), .B(n1644), .C(n1643), .D(n1642), .Q(n1651) );
  AOI221 U978 ( .A(n14), .B(regs[761]), .C(n10), .D(regs[697]), .Q(n1645) );
  AOI221 U979 ( .A(n1775), .B(n1641), .C(n1773), .D(n1640), .Q(n1653) );
  NAND41 U980 ( .A(n1639), .B(n1638), .C(n1637), .D(n1636), .Q(n1640) );
  NAND41 U981 ( .A(n1635), .B(n1634), .C(n1633), .D(n1632), .Q(n1641) );
  NAND22 U982 ( .A(n1433), .B(n1432), .Q(o_data_Rt[15]) );
  NAND41 U983 ( .A(n1429), .B(n1428), .C(n1427), .D(n1426), .Q(n1430) );
  AOI221 U984 ( .A(n12), .B(regs[79]), .C(n24), .D(regs[15]), .Q(n1426) );
  AOI221 U985 ( .A(n14), .B(regs[239]), .C(n10), .D(regs[175]), .Q(n1429) );
  NAND41 U986 ( .A(n1425), .B(n1424), .C(n1423), .D(n1422), .Q(n1431) );
  AOI221 U987 ( .A(n12), .B(regs[591]), .C(n24), .D(regs[527]), .Q(n1422) );
  AOI221 U988 ( .A(n14), .B(regs[751]), .C(n10), .D(regs[687]), .Q(n1425) );
  AOI221 U989 ( .A(n1775), .B(n1421), .C(n1773), .D(n1420), .Q(n1433) );
  NAND41 U990 ( .A(n1419), .B(n1418), .C(n1417), .D(n1416), .Q(n1420) );
  NAND41 U991 ( .A(n1415), .B(n1414), .C(n1413), .D(n1412), .Q(n1421) );
  NAND22 U992 ( .A(n1477), .B(n1476), .Q(o_data_Rt[17]) );
  NAND41 U993 ( .A(n1473), .B(n1472), .C(n1471), .D(n1470), .Q(n1474) );
  NAND41 U994 ( .A(n1469), .B(n1468), .C(n1467), .D(n1466), .Q(n1475) );
  AOI221 U995 ( .A(n12), .B(regs[593]), .C(n24), .D(regs[529]), .Q(n1466) );
  AOI221 U996 ( .A(n14), .B(regs[753]), .C(n10), .D(regs[689]), .Q(n1469) );
  AOI221 U997 ( .A(n1775), .B(n1465), .C(n1773), .D(n1464), .Q(n1477) );
  NAND41 U998 ( .A(n1463), .B(n1462), .C(n1461), .D(n1460), .Q(n1464) );
  NAND41 U999 ( .A(n1459), .B(n1458), .C(n1457), .D(n1456), .Q(n1465) );
  NAND22 U1000 ( .A(n1455), .B(n1454), .Q(o_data_Rt[16]) );
  NAND41 U1001 ( .A(n1451), .B(n1450), .C(n1449), .D(n1448), .Q(n1452) );
  NAND41 U1002 ( .A(n1447), .B(n1446), .C(n1445), .D(n1444), .Q(n1453) );
  AOI221 U1003 ( .A(n12), .B(regs[592]), .C(n24), .D(regs[528]), .Q(n1444) );
  AOI221 U1004 ( .A(n14), .B(regs[752]), .C(n10), .D(regs[688]), .Q(n1447) );
  AOI221 U1005 ( .A(n1775), .B(n1443), .C(n1773), .D(n1442), .Q(n1455) );
  NAND41 U1006 ( .A(n1441), .B(n1440), .C(n1439), .D(n1438), .Q(n1442) );
  NAND41 U1007 ( .A(n1437), .B(n1436), .C(n1435), .D(n1434), .Q(n1443) );
  NAND22 U1008 ( .A(n1499), .B(n1498), .Q(o_data_Rt[18]) );
  NAND41 U1009 ( .A(n1495), .B(n1494), .C(n1493), .D(n1492), .Q(n1496) );
  AOI221 U1010 ( .A(n8), .B(regs[114]), .C(n48), .D(regs[50]), .Q(n1493) );
  AOI221 U1011 ( .A(n14), .B(regs[242]), .C(n10), .D(regs[178]), .Q(n1495) );
  NAND41 U1012 ( .A(n1491), .B(n1490), .C(n1489), .D(n1488), .Q(n1497) );
  AOI221 U1013 ( .A(n12), .B(regs[594]), .C(n24), .D(regs[530]), .Q(n1488) );
  AOI221 U1014 ( .A(n8), .B(regs[626]), .C(n48), .D(regs[562]), .Q(n1489) );
  AOI221 U1015 ( .A(n46), .B(regs[722]), .C(n50), .D(regs[658]), .Q(n1490) );
  AOI221 U1016 ( .A(n14), .B(regs[754]), .C(n10), .D(regs[690]), .Q(n1491) );
  AOI221 U1017 ( .A(n1775), .B(n1487), .C(n1773), .D(n1486), .Q(n1499) );
  NAND41 U1018 ( .A(n1485), .B(n1484), .C(n1483), .D(n1482), .Q(n1486) );
  AOI221 U1019 ( .A(n46), .B(regs[466]), .C(n50), .D(regs[402]), .Q(n1484) );
  NAND41 U1020 ( .A(n1481), .B(n1480), .C(n1479), .D(n1478), .Q(n1487) );
  NAND22 U1021 ( .A(n1103), .B(n1102), .Q(o_data_Rt[0]) );
  NAND41 U1022 ( .A(n1099), .B(n1098), .C(n1097), .D(n1096), .Q(n1100) );
  AOI221 U1023 ( .A(n46), .B(regs[192]), .C(n52), .D(regs[128]), .Q(n1098) );
  AOI221 U1024 ( .A(n14), .B(regs[224]), .C(n10), .D(regs[160]), .Q(n1099) );
  NAND41 U1025 ( .A(n1095), .B(n1094), .C(n1093), .D(n1092), .Q(n1101) );
  AOI221 U1026 ( .A(n1775), .B(n1090), .C(n1773), .D(n1089), .Q(n1103) );
  NAND41 U1027 ( .A(n1088), .B(n1087), .C(n1086), .D(n1085), .Q(n1089) );
  AOI221 U1028 ( .A(n46), .B(regs[448]), .C(n52), .D(regs[384]), .Q(n1087) );
  AOI221 U1029 ( .A(n14), .B(regs[480]), .C(n10), .D(regs[416]), .Q(n1088) );
  NAND41 U1030 ( .A(n1083), .B(n1082), .C(n1081), .D(n1080), .Q(n1090) );
  AOI221 U1031 ( .A(n46), .B(regs[960]), .C(n50), .D(regs[896]), .Q(n1082) );
  NAND22 U1032 ( .A(n1521), .B(n1520), .Q(o_data_Rt[19]) );
  NAND41 U1033 ( .A(n1517), .B(n1516), .C(n1515), .D(n1514), .Q(n1518) );
  AOI221 U1034 ( .A(n12), .B(regs[83]), .C(n24), .D(regs[19]), .Q(n1514) );
  AOI221 U1035 ( .A(n8), .B(regs[115]), .C(n48), .D(regs[51]), .Q(n1515) );
  AOI221 U1036 ( .A(n14), .B(regs[243]), .C(n10), .D(regs[179]), .Q(n1517) );
  NAND41 U1037 ( .A(n1513), .B(n1512), .C(n1511), .D(n1510), .Q(n1519) );
  AOI221 U1038 ( .A(n12), .B(regs[595]), .C(n24), .D(regs[531]), .Q(n1510) );
  AOI221 U1039 ( .A(n8), .B(regs[627]), .C(n48), .D(regs[563]), .Q(n1511) );
  AOI221 U1040 ( .A(n46), .B(regs[723]), .C(n50), .D(regs[659]), .Q(n1512) );
  AOI221 U1041 ( .A(n14), .B(regs[755]), .C(n10), .D(regs[691]), .Q(n1513) );
  AOI221 U1042 ( .A(n1775), .B(n1509), .C(n1773), .D(n1508), .Q(n1521) );
  NAND41 U1043 ( .A(n1507), .B(n1506), .C(n1505), .D(n1504), .Q(n1508) );
  NAND41 U1044 ( .A(n1503), .B(n1502), .C(n1501), .D(n1500), .Q(n1509) );
  AOI221 U1045 ( .A(n46), .B(regs[979]), .C(n50), .D(regs[915]), .Q(n1502) );
  AOI221 U1046 ( .A(n14), .B(regs[1011]), .C(n10), .D(regs[947]), .Q(n1503) );
  NAND22 U1047 ( .A(n1389), .B(n1388), .Q(o_data_Rt[13]) );
  NAND41 U1048 ( .A(n1385), .B(n1384), .C(n1383), .D(n1382), .Q(n1386) );
  AOI221 U1049 ( .A(n12), .B(regs[77]), .C(n24), .D(regs[13]), .Q(n1382) );
  NAND41 U1050 ( .A(n1381), .B(n1380), .C(n1379), .D(n1378), .Q(n1387) );
  AOI221 U1051 ( .A(n12), .B(regs[589]), .C(n24), .D(regs[525]), .Q(n1378) );
  AOI221 U1052 ( .A(n14), .B(regs[749]), .C(n10), .D(regs[685]), .Q(n1381) );
  NAND41 U1053 ( .A(n1375), .B(n1374), .C(n1373), .D(n1372), .Q(n1376) );
  NAND41 U1054 ( .A(n1371), .B(n1370), .C(n1369), .D(n1368), .Q(n1377) );
  NAND22 U1055 ( .A(n1411), .B(n1410), .Q(o_data_Rt[14]) );
  NAND41 U1056 ( .A(n1407), .B(n1406), .C(n1405), .D(n1404), .Q(n1408) );
  AOI221 U1057 ( .A(n14), .B(regs[238]), .C(n10), .D(regs[174]), .Q(n1407) );
  NAND41 U1058 ( .A(n1403), .B(n1402), .C(n1401), .D(n1400), .Q(n1409) );
  AOI221 U1059 ( .A(n12), .B(regs[590]), .C(n24), .D(regs[526]), .Q(n1400) );
  AOI221 U1060 ( .A(n14), .B(regs[750]), .C(n10), .D(regs[686]), .Q(n1403) );
  NAND41 U1061 ( .A(n1397), .B(n1396), .C(n1395), .D(n1394), .Q(n1398) );
  NAND41 U1062 ( .A(n1393), .B(n1392), .C(n1391), .D(n1390), .Q(n1399) );
  AOI221 U1063 ( .A(n14), .B(regs[1006]), .C(n10), .D(regs[942]), .Q(n1393) );
  NAND22 U1064 ( .A(n1279), .B(n1278), .Q(o_data_Rt[8]) );
  NAND41 U1065 ( .A(n1275), .B(n1274), .C(n1273), .D(n1272), .Q(n1276) );
  AOI221 U1066 ( .A(n14), .B(regs[232]), .C(n10), .D(regs[168]), .Q(n1275) );
  NAND41 U1067 ( .A(n1271), .B(n1270), .C(n1269), .D(n1268), .Q(n1277) );
  AOI221 U1068 ( .A(n14), .B(regs[744]), .C(n10), .D(regs[680]), .Q(n1271) );
  AOI221 U1069 ( .A(n1775), .B(n1267), .C(n1773), .D(n1266), .Q(n1279) );
  NAND41 U1070 ( .A(n1265), .B(n1264), .C(n1263), .D(n1262), .Q(n1266) );
  AOI221 U1071 ( .A(n46), .B(regs[456]), .C(n52), .D(regs[392]), .Q(n1264) );
  NAND41 U1072 ( .A(n1261), .B(n1260), .C(n1259), .D(n1258), .Q(n1267) );
  AOI221 U1073 ( .A(n46), .B(regs[968]), .C(n52), .D(regs[904]), .Q(n1260) );
  NAND22 U1074 ( .A(n1323), .B(n1322), .Q(o_data_Rt[10]) );
  NAND41 U1075 ( .A(n1319), .B(n1318), .C(n1317), .D(n1316), .Q(n1320) );
  NAND41 U1076 ( .A(n1315), .B(n1314), .C(n1313), .D(n1312), .Q(n1321) );
  NAND41 U1077 ( .A(n1309), .B(n1308), .C(n1307), .D(n1306), .Q(n1310) );
  AOI221 U1078 ( .A(n46), .B(regs[458]), .C(n50), .D(regs[394]), .Q(n1308) );
  NAND41 U1079 ( .A(n1305), .B(n1304), .C(n1303), .D(n1302), .Q(n1311) );
  AOI221 U1080 ( .A(n46), .B(regs[970]), .C(n50), .D(regs[906]), .Q(n1304) );
  NAND22 U1081 ( .A(n1301), .B(n1300), .Q(o_data_Rt[9]) );
  NAND41 U1082 ( .A(n1297), .B(n1296), .C(n1295), .D(n1294), .Q(n1298) );
  AOI221 U1083 ( .A(n14), .B(regs[233]), .C(n10), .D(regs[169]), .Q(n1297) );
  NAND41 U1084 ( .A(n1293), .B(n1292), .C(n1291), .D(n1290), .Q(n1299) );
  AOI221 U1085 ( .A(n14), .B(regs[745]), .C(n10), .D(regs[681]), .Q(n1293) );
  NAND41 U1086 ( .A(n1287), .B(n1286), .C(n1285), .D(n1284), .Q(n1288) );
  AOI221 U1087 ( .A(n46), .B(regs[457]), .C(n50), .D(regs[393]), .Q(n1286) );
  NAND41 U1088 ( .A(n1283), .B(n1282), .C(n1281), .D(n1280), .Q(n1289) );
  AOI221 U1089 ( .A(n46), .B(regs[969]), .C(n50), .D(regs[905]), .Q(n1282) );
  NAND22 U1090 ( .A(n1125), .B(n1124), .Q(o_data_Rt[1]) );
  NAND41 U1091 ( .A(n1121), .B(n1120), .C(n1119), .D(n1118), .Q(n1122) );
  AOI221 U1092 ( .A(n46), .B(regs[193]), .C(n52), .D(regs[129]), .Q(n1120) );
  NAND41 U1093 ( .A(n1117), .B(n1116), .C(n1115), .D(n1114), .Q(n1123) );
  AOI221 U1094 ( .A(n8), .B(regs[609]), .C(n48), .D(regs[545]), .Q(n1115) );
  AOI221 U1095 ( .A(n46), .B(regs[705]), .C(n52), .D(regs[641]), .Q(n1116) );
  NAND41 U1096 ( .A(n1111), .B(n1110), .C(n1109), .D(n1108), .Q(n1112) );
  AOI221 U1097 ( .A(n46), .B(regs[449]), .C(n52), .D(regs[385]), .Q(n1110) );
  AOI221 U1098 ( .A(n14), .B(regs[481]), .C(n10), .D(regs[417]), .Q(n1111) );
  NAND41 U1099 ( .A(n1107), .B(n1106), .C(n1105), .D(n1104), .Q(n1113) );
  AOI221 U1100 ( .A(n46), .B(regs[961]), .C(n52), .D(regs[897]), .Q(n1106) );
  AOI221 U1101 ( .A(n14), .B(regs[993]), .C(n10), .D(regs[929]), .Q(n1107) );
  NAND22 U1102 ( .A(n1367), .B(n1366), .Q(o_data_Rt[12]) );
  NAND41 U1103 ( .A(n1363), .B(n1362), .C(n1361), .D(n1360), .Q(n1364) );
  NAND41 U1104 ( .A(n1359), .B(n1358), .C(n1357), .D(n1356), .Q(n1365) );
  NAND41 U1105 ( .A(n1353), .B(n1352), .C(n1351), .D(n1350), .Q(n1354) );
  AOI221 U1106 ( .A(n46), .B(regs[460]), .C(n50), .D(regs[396]), .Q(n1352) );
  NAND41 U1107 ( .A(n1349), .B(n1348), .C(n1347), .D(n1346), .Q(n1355) );
  AOI221 U1108 ( .A(n46), .B(regs[972]), .C(n50), .D(regs[908]), .Q(n1348) );
  NAND22 U1109 ( .A(n1345), .B(n1344), .Q(o_data_Rt[11]) );
  NAND41 U1110 ( .A(n1341), .B(n1340), .C(n1339), .D(n1338), .Q(n1342) );
  NAND41 U1111 ( .A(n1337), .B(n1336), .C(n1335), .D(n1334), .Q(n1343) );
  NAND41 U1112 ( .A(n1331), .B(n1330), .C(n1329), .D(n1328), .Q(n1332) );
  AOI221 U1113 ( .A(n46), .B(regs[459]), .C(n50), .D(regs[395]), .Q(n1330) );
  NAND41 U1114 ( .A(n1327), .B(n1326), .C(n1325), .D(n1324), .Q(n1333) );
  AOI221 U1115 ( .A(n46), .B(regs[971]), .C(n50), .D(regs[907]), .Q(n1326) );
  NAND22 U1116 ( .A(n1797), .B(n1796), .Q(o_data_Rt[31]) );
  NAND41 U1117 ( .A(n1791), .B(n1790), .C(n1789), .D(n1788), .Q(n1792) );
  AOI221 U1118 ( .A(n12), .B(regs[95]), .C(n24), .D(regs[31]), .Q(n1788) );
  AOI221 U1119 ( .A(n14), .B(regs[255]), .C(n10), .D(regs[191]), .Q(n1791) );
  NAND41 U1120 ( .A(n1779), .B(n1778), .C(n1777), .D(n1776), .Q(n1794) );
  AOI221 U1121 ( .A(n12), .B(regs[607]), .C(n24), .D(regs[543]), .Q(n1776) );
  AOI221 U1122 ( .A(n46), .B(regs[735]), .C(n50), .D(regs[671]), .Q(n1778) );
  AOI221 U1123 ( .A(n1775), .B(n1774), .C(n1773), .D(n1772), .Q(n1797) );
  NAND41 U1124 ( .A(n1771), .B(n1770), .C(n1769), .D(n1768), .Q(n1772) );
  NAND41 U1125 ( .A(n1767), .B(n1766), .C(n1765), .D(n1764), .Q(n1774) );
  AOI221 U1126 ( .A(n12), .B(regs[863]), .C(n24), .D(regs[799]), .Q(n1764) );
  NAND22 U1127 ( .A(n1213), .B(n1212), .Q(o_data_Rt[5]) );
  NAND41 U1128 ( .A(n1209), .B(n1208), .C(n1207), .D(n1206), .Q(n1210) );
  AOI221 U1129 ( .A(n14), .B(regs[229]), .C(n10), .D(regs[165]), .Q(n1209) );
  NAND41 U1130 ( .A(n1205), .B(n1204), .C(n1203), .D(n1202), .Q(n1211) );
  AOI221 U1131 ( .A(n46), .B(regs[709]), .C(n52), .D(regs[645]), .Q(n1204) );
  AOI221 U1132 ( .A(n14), .B(regs[741]), .C(n10), .D(regs[677]), .Q(n1205) );
  NAND41 U1133 ( .A(n1199), .B(n1198), .C(n1197), .D(n1196), .Q(n1200) );
  AOI221 U1134 ( .A(n46), .B(regs[453]), .C(n52), .D(regs[389]), .Q(n1198) );
  NAND41 U1135 ( .A(n1195), .B(n1194), .C(n1193), .D(n1192), .Q(n1201) );
  AOI221 U1136 ( .A(n46), .B(regs[965]), .C(n52), .D(regs[901]), .Q(n1194) );
  NAND22 U1137 ( .A(n1191), .B(n1190), .Q(o_data_Rt[4]) );
  NAND41 U1138 ( .A(n1187), .B(n1186), .C(n1185), .D(n1184), .Q(n1188) );
  AOI221 U1139 ( .A(n14), .B(regs[228]), .C(n10), .D(regs[164]), .Q(n1187) );
  NAND41 U1140 ( .A(n1183), .B(n1182), .C(n1181), .D(n1180), .Q(n1189) );
  AOI221 U1141 ( .A(n46), .B(regs[708]), .C(n52), .D(regs[644]), .Q(n1182) );
  AOI221 U1142 ( .A(n14), .B(regs[740]), .C(n10), .D(regs[676]), .Q(n1183) );
  AOI221 U1143 ( .A(n1775), .B(n1179), .C(n1773), .D(n1178), .Q(n1191) );
  NAND41 U1144 ( .A(n1177), .B(n1176), .C(n1175), .D(n1174), .Q(n1178) );
  AOI221 U1145 ( .A(n46), .B(regs[452]), .C(n52), .D(regs[388]), .Q(n1176) );
  AOI221 U1146 ( .A(n14), .B(regs[484]), .C(n10), .D(regs[420]), .Q(n1177) );
  NAND41 U1147 ( .A(n1173), .B(n1172), .C(n1171), .D(n1170), .Q(n1179) );
  AOI221 U1148 ( .A(n46), .B(regs[964]), .C(n52), .D(regs[900]), .Q(n1172) );
  AOI221 U1149 ( .A(n14), .B(regs[996]), .C(n10), .D(regs[932]), .Q(n1173) );
  NAND22 U1150 ( .A(n1631), .B(n1630), .Q(o_data_Rt[24]) );
  NAND41 U1151 ( .A(n1627), .B(n1626), .C(n1625), .D(n1624), .Q(n1628) );
  NAND41 U1152 ( .A(n1623), .B(n1622), .C(n1621), .D(n1620), .Q(n1629) );
  AOI221 U1153 ( .A(n1775), .B(n1619), .C(n1773), .D(n1618), .Q(n1631) );
  NAND41 U1154 ( .A(n1617), .B(n1616), .C(n1615), .D(n1614), .Q(n1618) );
  NAND41 U1155 ( .A(n1613), .B(n1612), .C(n1611), .D(n1610), .Q(n1619) );
  AOI221 U1156 ( .A(n46), .B(regs[984]), .C(n50), .D(regs[920]), .Q(n1612) );
  AOI221 U1157 ( .A(n14), .B(regs[1016]), .C(n10), .D(regs[952]), .Q(n1613) );
  NAND22 U1158 ( .A(n1147), .B(n1146), .Q(o_data_Rt[2]) );
  NAND41 U1159 ( .A(n1143), .B(n1142), .C(n1141), .D(n1140), .Q(n1144) );
  NAND41 U1160 ( .A(n1139), .B(n1138), .C(n1137), .D(n1136), .Q(n1145) );
  AOI221 U1161 ( .A(n46), .B(regs[706]), .C(n52), .D(regs[642]), .Q(n1138) );
  AOI221 U1162 ( .A(n14), .B(regs[738]), .C(n10), .D(regs[674]), .Q(n1139) );
  NAND41 U1163 ( .A(n1133), .B(n1132), .C(n1131), .D(n1130), .Q(n1134) );
  AOI221 U1164 ( .A(n14), .B(regs[482]), .C(n10), .D(regs[418]), .Q(n1133) );
  NAND41 U1165 ( .A(n1129), .B(n1128), .C(n1127), .D(n1126), .Q(n1135) );
  AOI221 U1166 ( .A(n46), .B(regs[962]), .C(n52), .D(regs[898]), .Q(n1128) );
  AOI221 U1167 ( .A(n14), .B(regs[994]), .C(n10), .D(regs[930]), .Q(n1129) );
  NAND22 U1168 ( .A(n1169), .B(n1168), .Q(o_data_Rt[3]) );
  NAND41 U1169 ( .A(n1165), .B(n1164), .C(n1163), .D(n1162), .Q(n1166) );
  AOI221 U1170 ( .A(n46), .B(regs[195]), .C(n52), .D(regs[131]), .Q(n1164) );
  NAND41 U1171 ( .A(n1161), .B(n1160), .C(n1159), .D(n1158), .Q(n1167) );
  AOI221 U1172 ( .A(n46), .B(regs[707]), .C(n52), .D(regs[643]), .Q(n1160) );
  AOI221 U1173 ( .A(n14), .B(regs[739]), .C(n10), .D(regs[675]), .Q(n1161) );
  AOI221 U1174 ( .A(n1775), .B(n1157), .C(n1773), .D(n1156), .Q(n1169) );
  NAND41 U1175 ( .A(n1155), .B(n1154), .C(n1153), .D(n1152), .Q(n1156) );
  AOI221 U1176 ( .A(n46), .B(regs[451]), .C(n52), .D(regs[387]), .Q(n1154) );
  AOI221 U1177 ( .A(n14), .B(regs[483]), .C(n10), .D(regs[419]), .Q(n1155) );
  NAND41 U1178 ( .A(n1151), .B(n1150), .C(n1149), .D(n1148), .Q(n1157) );
  AOI221 U1179 ( .A(n46), .B(regs[963]), .C(n52), .D(regs[899]), .Q(n1150) );
  AOI221 U1180 ( .A(n14), .B(regs[995]), .C(n10), .D(regs[931]), .Q(n1151) );
  NAND22 U1181 ( .A(n1675), .B(n1674), .Q(o_data_Rt[26]) );
  NAND41 U1182 ( .A(n1671), .B(n1670), .C(n1669), .D(n1668), .Q(n1672) );
  NAND41 U1183 ( .A(n1667), .B(n1666), .C(n1665), .D(n1664), .Q(n1673) );
  AOI221 U1184 ( .A(n1775), .B(n1663), .C(n1773), .D(n1662), .Q(n1675) );
  NAND41 U1185 ( .A(n1661), .B(n1660), .C(n1659), .D(n1658), .Q(n1662) );
  NAND41 U1186 ( .A(n1657), .B(n1656), .C(n1655), .D(n1654), .Q(n1663) );
  NAND22 U1187 ( .A(n1697), .B(n1696), .Q(o_data_Rt[27]) );
  NAND41 U1188 ( .A(n1693), .B(n1692), .C(n1691), .D(n1690), .Q(n1694) );
  AOI221 U1189 ( .A(n14), .B(regs[251]), .C(n10), .D(regs[187]), .Q(n1693) );
  NAND41 U1190 ( .A(n1689), .B(n1688), .C(n1687), .D(n1686), .Q(n1695) );
  AOI221 U1191 ( .A(n1775), .B(n1685), .C(n1773), .D(n1684), .Q(n1697) );
  NAND41 U1192 ( .A(n1683), .B(n1682), .C(n1681), .D(n1680), .Q(n1684) );
  NAND41 U1193 ( .A(n1679), .B(n1678), .C(n1677), .D(n1676), .Q(n1685) );
  NAND22 U1194 ( .A(n1741), .B(n1740), .Q(o_data_Rt[29]) );
  NAND41 U1195 ( .A(n1737), .B(n1736), .C(n1735), .D(n1734), .Q(n1738) );
  AOI221 U1196 ( .A(n14), .B(regs[253]), .C(n10), .D(regs[189]), .Q(n1737) );
  NAND41 U1197 ( .A(n1733), .B(n1732), .C(n1731), .D(n1730), .Q(n1739) );
  AOI221 U1198 ( .A(n14), .B(regs[765]), .C(n10), .D(regs[701]), .Q(n1733) );
  AOI221 U1199 ( .A(n1775), .B(n1729), .C(n1773), .D(n1728), .Q(n1741) );
  NAND41 U1200 ( .A(n1727), .B(n1726), .C(n1725), .D(n1724), .Q(n1728) );
  AOI221 U1201 ( .A(n14), .B(regs[509]), .C(n10), .D(regs[445]), .Q(n1727) );
  NAND41 U1202 ( .A(n1723), .B(n1722), .C(n1721), .D(n1720), .Q(n1729) );
  AOI221 U1203 ( .A(n14), .B(regs[1021]), .C(n10), .D(regs[957]), .Q(n1723) );
  NAND22 U1204 ( .A(n1719), .B(n1718), .Q(o_data_Rt[28]) );
  NAND41 U1205 ( .A(n1715), .B(n1714), .C(n1713), .D(n1712), .Q(n1716) );
  AOI221 U1206 ( .A(n14), .B(regs[252]), .C(n10), .D(regs[188]), .Q(n1715) );
  NAND41 U1207 ( .A(n1711), .B(n1710), .C(n1709), .D(n1708), .Q(n1717) );
  AOI221 U1208 ( .A(n14), .B(regs[764]), .C(n10), .D(regs[700]), .Q(n1711) );
  AOI221 U1209 ( .A(n1775), .B(n1707), .C(n1773), .D(n1706), .Q(n1719) );
  NAND41 U1210 ( .A(n1705), .B(n1704), .C(n1703), .D(n1702), .Q(n1706) );
  AOI221 U1211 ( .A(n14), .B(regs[508]), .C(n10), .D(regs[444]), .Q(n1705) );
  NAND41 U1212 ( .A(n1701), .B(n1700), .C(n1699), .D(n1698), .Q(n1707) );
  NAND22 U1213 ( .A(n1257), .B(n1256), .Q(o_data_Rt[7]) );
  NAND41 U1214 ( .A(n1253), .B(n1252), .C(n1251), .D(n1250), .Q(n1254) );
  NAND41 U1215 ( .A(n1249), .B(n1248), .C(n1247), .D(n1246), .Q(n1255) );
  AOI221 U1216 ( .A(n12), .B(regs[583]), .C(n24), .D(regs[519]), .Q(n1246) );
  NAND41 U1217 ( .A(n1243), .B(n1242), .C(n1241), .D(n1240), .Q(n1244) );
  AOI221 U1218 ( .A(n46), .B(regs[455]), .C(n52), .D(regs[391]), .Q(n1242) );
  NAND41 U1219 ( .A(n1239), .B(n1238), .C(n1237), .D(n1236), .Q(n1245) );
  AOI221 U1220 ( .A(n46), .B(regs[967]), .C(n52), .D(regs[903]), .Q(n1238) );
  NAND22 U1221 ( .A(n1235), .B(n1234), .Q(o_data_Rt[6]) );
  NAND41 U1222 ( .A(n1231), .B(n1230), .C(n1229), .D(n1228), .Q(n1232) );
  NAND41 U1223 ( .A(n1227), .B(n1226), .C(n1225), .D(n1224), .Q(n1233) );
  AOI221 U1224 ( .A(n1775), .B(n1223), .C(n1773), .D(n1222), .Q(n1235) );
  NAND41 U1225 ( .A(n1221), .B(n1220), .C(n1219), .D(n1218), .Q(n1222) );
  NAND41 U1226 ( .A(n1217), .B(n1216), .C(n1215), .D(n1214), .Q(n1223) );
  AOI221 U1227 ( .A(n46), .B(regs[966]), .C(n52), .D(regs[902]), .Q(n1216) );
  AOI311 U1228 ( .A(n381), .B(n380), .C(n379), .D(n1064), .Q(n382) );
  AOI211 U1229 ( .A(n3), .B(regs[580]), .C(n378), .Q(n379) );
  AOI221 U1230 ( .A(n45), .B(regs[612]), .C(n1), .D(regs[740]), .Q(n377) );
  AOI221 U1231 ( .A(n33), .B(regs[708]), .C(n7), .D(regs[644]), .Q(n381) );
  AOI311 U1232 ( .A(n376), .B(n375), .C(n374), .D(n1051), .Q(n383) );
  AOI211 U1233 ( .A(n3), .B(regs[68]), .C(n373), .Q(n374) );
  AOI221 U1234 ( .A(n45), .B(regs[100]), .C(n1), .D(regs[228]), .Q(n372) );
  AOI221 U1235 ( .A(n33), .B(regs[196]), .C(n7), .D(regs[132]), .Q(n376) );
  AOI311 U1236 ( .A(n371), .B(n370), .C(n369), .D(n1045), .Q(n384) );
  AOI211 U1237 ( .A(n4), .B(regs[836]), .C(n368), .Q(n369) );
  AOI221 U1238 ( .A(n45), .B(regs[868]), .C(n1), .D(regs[996]), .Q(n367) );
  AOI221 U1239 ( .A(n33), .B(regs[964]), .C(n7), .D(regs[900]), .Q(n371) );
  AOI311 U1240 ( .A(n366), .B(n365), .C(n364), .D(n1039), .Q(n385) );
  AOI211 U1241 ( .A(n3), .B(regs[324]), .C(n363), .Q(n364) );
  AOI221 U1242 ( .A(n45), .B(regs[356]), .C(n1), .D(regs[484]), .Q(n362) );
  AOI221 U1243 ( .A(n33), .B(regs[452]), .C(n7), .D(regs[388]), .Q(n366) );
  AOI311 U1244 ( .A(n456), .B(n455), .C(n454), .D(n1064), .Q(n457) );
  AOI211 U1245 ( .A(n4), .B(regs[583]), .C(n453), .Q(n454) );
  AOI221 U1246 ( .A(n45), .B(regs[615]), .C(n199), .D(regs[743]), .Q(n452) );
  AOI221 U1247 ( .A(n33), .B(regs[711]), .C(n7), .D(regs[647]), .Q(n456) );
  AOI311 U1248 ( .A(n451), .B(n450), .C(n449), .D(n1051), .Q(n458) );
  AOI211 U1249 ( .A(n4), .B(regs[71]), .C(n448), .Q(n449) );
  AOI221 U1250 ( .A(n45), .B(regs[103]), .C(n199), .D(regs[231]), .Q(n447) );
  AOI221 U1251 ( .A(n33), .B(regs[199]), .C(n7), .D(regs[135]), .Q(n451) );
  AOI311 U1252 ( .A(n446), .B(n445), .C(n444), .D(n1045), .Q(n459) );
  AOI211 U1253 ( .A(n3), .B(regs[839]), .C(n443), .Q(n444) );
  AOI221 U1254 ( .A(n45), .B(regs[871]), .C(n199), .D(regs[999]), .Q(n442) );
  AOI221 U1255 ( .A(n33), .B(regs[967]), .C(n7), .D(regs[903]), .Q(n446) );
  AOI311 U1256 ( .A(n441), .B(n440), .C(n439), .D(n1039), .Q(n460) );
  AOI211 U1257 ( .A(n4), .B(regs[327]), .C(n438), .Q(n439) );
  AOI221 U1258 ( .A(n45), .B(regs[359]), .C(n199), .D(regs[487]), .Q(n437) );
  AOI221 U1259 ( .A(n33), .B(regs[455]), .C(n7), .D(regs[391]), .Q(n441) );
  NAND22 U1260 ( .A(n1810), .B(n1809), .Q(o_data_Rs[1]) );
  NAND31 U1261 ( .A(n311), .B(n310), .C(n309), .Q(n1807) );
  NAND31 U1262 ( .A(n306), .B(n305), .C(n304), .Q(n1808) );
  NAND31 U1263 ( .A(n301), .B(n300), .C(n299), .Q(n1805) );
  NAND31 U1264 ( .A(n296), .B(n295), .C(n294), .Q(n1806) );
  AOI311 U1265 ( .A(n806), .B(n805), .C(n804), .D(n1064), .Q(n807) );
  AOI211 U1266 ( .A(n3), .B(regs[597]), .C(n803), .Q(n804) );
  AOI221 U1267 ( .A(n45), .B(regs[629]), .C(n199), .D(regs[757]), .Q(n802) );
  AOI221 U1268 ( .A(n33), .B(regs[725]), .C(n7), .D(regs[661]), .Q(n806) );
  AOI311 U1269 ( .A(n801), .B(n800), .C(n799), .D(n1051), .Q(n808) );
  AOI211 U1270 ( .A(n4), .B(regs[85]), .C(n798), .Q(n799) );
  AOI221 U1271 ( .A(n33), .B(regs[213]), .C(n7), .D(regs[149]), .Q(n801) );
  AOI311 U1272 ( .A(n796), .B(n795), .C(n794), .D(n1045), .Q(n809) );
  AOI211 U1273 ( .A(n3), .B(regs[853]), .C(n793), .Q(n794) );
  AOI221 U1274 ( .A(n45), .B(regs[885]), .C(n199), .D(regs[1013]), .Q(n792) );
  AOI221 U1275 ( .A(n33), .B(regs[981]), .C(n7), .D(regs[917]), .Q(n796) );
  AOI311 U1276 ( .A(n791), .B(n790), .C(n789), .D(n1039), .Q(n810) );
  AOI211 U1277 ( .A(n4), .B(regs[341]), .C(n788), .Q(n789) );
  AOI221 U1278 ( .A(n45), .B(regs[373]), .C(n199), .D(regs[501]), .Q(n787) );
  AOI221 U1279 ( .A(n33), .B(regs[469]), .C(n7), .D(regs[405]), .Q(n791) );
  NAND22 U1280 ( .A(n1543), .B(n1542), .Q(o_data_Rt[20]) );
  NAND41 U1281 ( .A(n1539), .B(n1538), .C(n1537), .D(n1536), .Q(n1540) );
  AOI221 U1282 ( .A(n46), .B(regs[212]), .C(n50), .D(regs[148]), .Q(n1538) );
  AOI221 U1283 ( .A(n14), .B(regs[244]), .C(n10), .D(regs[180]), .Q(n1539) );
  NAND41 U1284 ( .A(n1535), .B(n1534), .C(n1533), .D(n1532), .Q(n1541) );
  AOI221 U1285 ( .A(n46), .B(regs[724]), .C(n50), .D(regs[660]), .Q(n1534) );
  AOI221 U1286 ( .A(n14), .B(regs[756]), .C(n10), .D(regs[692]), .Q(n1535) );
  AOI221 U1287 ( .A(n1775), .B(n1531), .C(n1773), .D(n1530), .Q(n1543) );
  NAND41 U1288 ( .A(n1529), .B(n1528), .C(n1527), .D(n1526), .Q(n1530) );
  AOI221 U1289 ( .A(n46), .B(regs[468]), .C(n50), .D(regs[404]), .Q(n1528) );
  AOI221 U1290 ( .A(n14), .B(regs[500]), .C(n10), .D(regs[436]), .Q(n1529) );
  NAND41 U1291 ( .A(n1525), .B(n1524), .C(n1523), .D(n1522), .Q(n1531) );
  AOI221 U1292 ( .A(n8), .B(regs[884]), .C(n48), .D(regs[820]), .Q(n1523) );
  AOI221 U1293 ( .A(n46), .B(regs[980]), .C(n50), .D(regs[916]), .Q(n1524) );
  AOI221 U1294 ( .A(n14), .B(regs[1012]), .C(n10), .D(regs[948]), .Q(n1525) );
  NAND22 U1295 ( .A(n1565), .B(n1564), .Q(o_data_Rt[21]) );
  NAND41 U1296 ( .A(n1561), .B(n1560), .C(n1559), .D(n1558), .Q(n1562) );
  AOI221 U1297 ( .A(n46), .B(regs[213]), .C(n50), .D(regs[149]), .Q(n1560) );
  AOI221 U1298 ( .A(n14), .B(regs[245]), .C(n10), .D(regs[181]), .Q(n1561) );
  NAND41 U1299 ( .A(n1557), .B(n1556), .C(n1555), .D(n1554), .Q(n1563) );
  AOI221 U1300 ( .A(n46), .B(regs[725]), .C(n50), .D(regs[661]), .Q(n1556) );
  AOI221 U1301 ( .A(n14), .B(regs[757]), .C(n10), .D(regs[693]), .Q(n1557) );
  AOI221 U1302 ( .A(n1775), .B(n1553), .C(n1773), .D(n1552), .Q(n1565) );
  NAND41 U1303 ( .A(n1551), .B(n1550), .C(n1549), .D(n1548), .Q(n1552) );
  AOI221 U1304 ( .A(n46), .B(regs[469]), .C(n50), .D(regs[405]), .Q(n1550) );
  AOI221 U1305 ( .A(n14), .B(regs[501]), .C(n10), .D(regs[437]), .Q(n1551) );
  NAND41 U1306 ( .A(n1547), .B(n1546), .C(n1545), .D(n1544), .Q(n1553) );
  AOI221 U1307 ( .A(n46), .B(regs[981]), .C(n50), .D(regs[917]), .Q(n1546) );
  AOI221 U1308 ( .A(n14), .B(regs[1013]), .C(n10), .D(regs[949]), .Q(n1547) );
  AOI311 U1309 ( .A(n481), .B(n480), .C(n479), .D(n1064), .Q(n482) );
  AOI211 U1310 ( .A(n3), .B(regs[584]), .C(n478), .Q(n479) );
  AOI221 U1311 ( .A(n45), .B(regs[616]), .C(n1), .D(regs[744]), .Q(n477) );
  AOI221 U1312 ( .A(n33), .B(regs[712]), .C(n7), .D(regs[648]), .Q(n481) );
  AOI311 U1313 ( .A(n476), .B(n475), .C(n474), .D(n1051), .Q(n483) );
  AOI211 U1314 ( .A(n4), .B(regs[72]), .C(n473), .Q(n474) );
  AOI221 U1315 ( .A(n45), .B(regs[104]), .C(n1), .D(regs[232]), .Q(n472) );
  AOI221 U1316 ( .A(n33), .B(regs[200]), .C(n7), .D(regs[136]), .Q(n476) );
  AOI311 U1317 ( .A(n471), .B(n470), .C(n469), .D(n1045), .Q(n484) );
  AOI211 U1318 ( .A(n4), .B(regs[840]), .C(n468), .Q(n469) );
  AOI221 U1319 ( .A(n45), .B(regs[872]), .C(n199), .D(regs[1000]), .Q(n467) );
  AOI221 U1320 ( .A(n33), .B(regs[968]), .C(n7), .D(regs[904]), .Q(n471) );
  AOI311 U1321 ( .A(n466), .B(n465), .C(n464), .D(n1039), .Q(n485) );
  AOI211 U1322 ( .A(n4), .B(regs[328]), .C(n463), .Q(n464) );
  AOI221 U1323 ( .A(n45), .B(regs[360]), .C(n199), .D(regs[488]), .Q(n462) );
  AOI221 U1324 ( .A(n33), .B(regs[456]), .C(n7), .D(regs[392]), .Q(n466) );
  AOI311 U1325 ( .A(n781), .B(n780), .C(n779), .D(n1064), .Q(n782) );
  AOI211 U1326 ( .A(n3), .B(regs[596]), .C(n778), .Q(n779) );
  AOI221 U1327 ( .A(n45), .B(regs[628]), .C(n199), .D(regs[756]), .Q(n777) );
  AOI221 U1328 ( .A(n47), .B(regs[564]), .C(n19), .D(regs[532]), .Q(n780) );
  AOI221 U1329 ( .A(n33), .B(regs[724]), .C(n7), .D(regs[660]), .Q(n781) );
  AOI311 U1330 ( .A(n776), .B(n775), .C(n774), .D(n1051), .Q(n783) );
  AOI211 U1331 ( .A(n3), .B(regs[84]), .C(n773), .Q(n774) );
  AOI221 U1332 ( .A(n47), .B(regs[52]), .C(n19), .D(regs[20]), .Q(n775) );
  AOI221 U1333 ( .A(n33), .B(regs[212]), .C(n7), .D(regs[148]), .Q(n776) );
  AOI311 U1334 ( .A(n771), .B(n770), .C(n769), .D(n1045), .Q(n784) );
  AOI211 U1335 ( .A(n4), .B(regs[852]), .C(n768), .Q(n769) );
  AOI221 U1336 ( .A(n47), .B(regs[820]), .C(n19), .D(regs[788]), .Q(n770) );
  AOI221 U1337 ( .A(n33), .B(regs[980]), .C(n7), .D(regs[916]), .Q(n771) );
  AOI311 U1338 ( .A(n766), .B(n765), .C(n764), .D(n1039), .Q(n785) );
  AOI211 U1339 ( .A(n3), .B(regs[340]), .C(n763), .Q(n764) );
  AOI221 U1340 ( .A(n47), .B(regs[308]), .C(n19), .D(regs[276]), .Q(n765) );
  AOI221 U1341 ( .A(n33), .B(regs[468]), .C(n7), .D(regs[404]), .Q(n766) );
  AOI311 U1342 ( .A(n406), .B(n405), .C(n404), .D(n1064), .Q(n407) );
  AOI211 U1343 ( .A(n4), .B(regs[581]), .C(n403), .Q(n404) );
  AOI221 U1344 ( .A(n45), .B(regs[613]), .C(n1), .D(regs[741]), .Q(n402) );
  AOI221 U1345 ( .A(n33), .B(regs[709]), .C(n7), .D(regs[645]), .Q(n406) );
  AOI311 U1346 ( .A(n401), .B(n400), .C(n399), .D(n1051), .Q(n408) );
  AOI211 U1347 ( .A(n4), .B(regs[69]), .C(n398), .Q(n399) );
  AOI221 U1348 ( .A(n45), .B(regs[101]), .C(n1), .D(regs[229]), .Q(n397) );
  AOI221 U1349 ( .A(n33), .B(regs[197]), .C(n7), .D(regs[133]), .Q(n401) );
  AOI311 U1350 ( .A(n396), .B(n395), .C(n394), .D(n1045), .Q(n409) );
  AOI211 U1351 ( .A(n4), .B(regs[837]), .C(n393), .Q(n394) );
  AOI221 U1352 ( .A(n45), .B(regs[869]), .C(n1), .D(regs[997]), .Q(n392) );
  AOI221 U1353 ( .A(n33), .B(regs[965]), .C(n7), .D(regs[901]), .Q(n396) );
  AOI311 U1354 ( .A(n391), .B(n390), .C(n389), .D(n1039), .Q(n410) );
  AOI211 U1355 ( .A(n4), .B(regs[325]), .C(n388), .Q(n389) );
  AOI221 U1356 ( .A(n45), .B(regs[357]), .C(n1), .D(regs[485]), .Q(n387) );
  AOI221 U1357 ( .A(n47), .B(regs[293]), .C(n19), .D(regs[261]), .Q(n390) );
  AOI221 U1358 ( .A(n33), .B(regs[453]), .C(n7), .D(regs[389]), .Q(n391) );
  NAND22 U1359 ( .A(n1763), .B(n1762), .Q(o_data_Rt[30]) );
  NAND41 U1360 ( .A(n1759), .B(n1758), .C(n1757), .D(n1756), .Q(n1760) );
  AOI221 U1361 ( .A(n46), .B(regs[222]), .C(n50), .D(regs[158]), .Q(n1758) );
  NAND41 U1362 ( .A(n1755), .B(n1754), .C(n1753), .D(n1752), .Q(n1761) );
  AOI221 U1363 ( .A(n12), .B(regs[606]), .C(n24), .D(regs[542]), .Q(n1752) );
  AOI221 U1364 ( .A(n46), .B(regs[734]), .C(n50), .D(regs[670]), .Q(n1754) );
  AOI221 U1365 ( .A(n1775), .B(n1751), .C(n1773), .D(n1750), .Q(n1763) );
  NAND41 U1366 ( .A(n1749), .B(n1748), .C(n1747), .D(n1746), .Q(n1750) );
  NAND41 U1367 ( .A(n1745), .B(n1744), .C(n1743), .D(n1742), .Q(n1751) );
  AOI221 U1368 ( .A(n14), .B(regs[1022]), .C(n10), .D(regs[958]), .Q(n1745) );
  NAND22 U1369 ( .A(n1609), .B(n1608), .Q(o_data_Rt[23]) );
  NAND41 U1370 ( .A(n1605), .B(n1604), .C(n1603), .D(n1602), .Q(n1606) );
  AOI221 U1371 ( .A(n46), .B(regs[215]), .C(n50), .D(regs[151]), .Q(n1604) );
  AOI221 U1372 ( .A(n14), .B(regs[247]), .C(n10), .D(regs[183]), .Q(n1605) );
  NAND41 U1373 ( .A(n1601), .B(n1600), .C(n1599), .D(n1598), .Q(n1607) );
  AOI221 U1374 ( .A(n46), .B(regs[727]), .C(n50), .D(regs[663]), .Q(n1600) );
  AOI221 U1375 ( .A(n14), .B(regs[759]), .C(n10), .D(regs[695]), .Q(n1601) );
  AOI221 U1376 ( .A(n1775), .B(n1597), .C(n1773), .D(n1596), .Q(n1609) );
  NAND41 U1377 ( .A(n1595), .B(n1594), .C(n1593), .D(n1592), .Q(n1596) );
  AOI221 U1378 ( .A(n14), .B(regs[503]), .C(n10), .D(regs[439]), .Q(n1595) );
  NAND41 U1379 ( .A(n1591), .B(n1590), .C(n1589), .D(n1588), .Q(n1597) );
  AOI221 U1380 ( .A(n46), .B(regs[983]), .C(n50), .D(regs[919]), .Q(n1590) );
  AOI221 U1381 ( .A(n14), .B(regs[1015]), .C(n10), .D(regs[951]), .Q(n1591) );
  NAND22 U1382 ( .A(n1587), .B(n1586), .Q(o_data_Rt[22]) );
  NAND41 U1383 ( .A(n1583), .B(n1582), .C(n1581), .D(n1580), .Q(n1584) );
  AOI221 U1384 ( .A(n46), .B(regs[214]), .C(n50), .D(regs[150]), .Q(n1582) );
  AOI221 U1385 ( .A(n14), .B(regs[246]), .C(n10), .D(regs[182]), .Q(n1583) );
  NAND41 U1386 ( .A(n1579), .B(n1578), .C(n1577), .D(n1576), .Q(n1585) );
  AOI221 U1387 ( .A(n46), .B(regs[726]), .C(n50), .D(regs[662]), .Q(n1578) );
  AOI221 U1388 ( .A(n14), .B(regs[758]), .C(n10), .D(regs[694]), .Q(n1579) );
  AOI221 U1389 ( .A(n1775), .B(n1575), .C(n1773), .D(n1574), .Q(n1587) );
  NAND41 U1390 ( .A(n1573), .B(n1572), .C(n1571), .D(n1570), .Q(n1574) );
  AOI221 U1391 ( .A(n14), .B(regs[502]), .C(n10), .D(regs[438]), .Q(n1573) );
  NAND41 U1392 ( .A(n1569), .B(n1568), .C(n1567), .D(n1566), .Q(n1575) );
  AOI221 U1393 ( .A(n14), .B(regs[1014]), .C(n10), .D(regs[950]), .Q(n1569) );
  AOI311 U1394 ( .A(n356), .B(n355), .C(n354), .D(n1064), .Q(n357) );
  AOI221 U1395 ( .A(n45), .B(regs[611]), .C(n1), .D(regs[739]), .Q(n352) );
  AOI221 U1396 ( .A(n33), .B(regs[707]), .C(n7), .D(regs[643]), .Q(n356) );
  AOI311 U1397 ( .A(n351), .B(n350), .C(n349), .D(n1051), .Q(n358) );
  AOI211 U1398 ( .A(n3), .B(regs[67]), .C(n348), .Q(n349) );
  AOI221 U1399 ( .A(n45), .B(regs[99]), .C(n1), .D(regs[227]), .Q(n347) );
  AOI221 U1400 ( .A(n33), .B(regs[195]), .C(n7), .D(regs[131]), .Q(n351) );
  AOI311 U1401 ( .A(n346), .B(n345), .C(n344), .D(n1045), .Q(n359) );
  AOI211 U1402 ( .A(n3), .B(regs[835]), .C(n343), .Q(n344) );
  AOI221 U1403 ( .A(n45), .B(regs[867]), .C(n1), .D(regs[995]), .Q(n342) );
  AOI221 U1404 ( .A(n33), .B(regs[963]), .C(n7), .D(regs[899]), .Q(n346) );
  AOI311 U1405 ( .A(n341), .B(n340), .C(n339), .D(n1039), .Q(n360) );
  AOI211 U1406 ( .A(n3), .B(regs[323]), .C(n338), .Q(n339) );
  AOI221 U1407 ( .A(n45), .B(regs[355]), .C(n1), .D(regs[483]), .Q(n337) );
  AOI221 U1408 ( .A(n33), .B(regs[451]), .C(n7), .D(regs[387]), .Q(n341) );
  AOI311 U1409 ( .A(n431), .B(n430), .C(n429), .D(n1064), .Q(n432) );
  AOI211 U1410 ( .A(n3), .B(regs[582]), .C(n428), .Q(n429) );
  AOI221 U1411 ( .A(n45), .B(regs[614]), .C(n1), .D(regs[742]), .Q(n427) );
  AOI221 U1412 ( .A(n33), .B(regs[710]), .C(n7), .D(regs[646]), .Q(n431) );
  AOI311 U1413 ( .A(n426), .B(n425), .C(n424), .D(n1051), .Q(n433) );
  AOI211 U1414 ( .A(n4), .B(regs[70]), .C(n423), .Q(n424) );
  AOI221 U1415 ( .A(n45), .B(regs[102]), .C(n1), .D(regs[230]), .Q(n422) );
  AOI221 U1416 ( .A(n33), .B(regs[198]), .C(n7), .D(regs[134]), .Q(n426) );
  AOI311 U1417 ( .A(n421), .B(n420), .C(n419), .D(n1045), .Q(n434) );
  AOI211 U1418 ( .A(n3), .B(regs[838]), .C(n418), .Q(n419) );
  AOI221 U1419 ( .A(n45), .B(regs[870]), .C(n1), .D(regs[998]), .Q(n417) );
  AOI221 U1420 ( .A(n33), .B(regs[966]), .C(n7), .D(regs[902]), .Q(n421) );
  AOI311 U1421 ( .A(n416), .B(n415), .C(n414), .D(n1039), .Q(n435) );
  AOI211 U1422 ( .A(n3), .B(regs[326]), .C(n413), .Q(n414) );
  AOI221 U1423 ( .A(n45), .B(regs[358]), .C(n199), .D(regs[486]), .Q(n412) );
  AOI221 U1424 ( .A(n33), .B(regs[454]), .C(n7), .D(regs[390]), .Q(n416) );
  AOI311 U1425 ( .A(n756), .B(n755), .C(n754), .D(n1064), .Q(n757) );
  AOI211 U1426 ( .A(n4), .B(regs[595]), .C(n753), .Q(n754) );
  AOI221 U1427 ( .A(n45), .B(regs[627]), .C(n199), .D(regs[755]), .Q(n752) );
  AOI221 U1428 ( .A(n47), .B(regs[563]), .C(n19), .D(regs[531]), .Q(n755) );
  AOI311 U1429 ( .A(n751), .B(n750), .C(n749), .D(n1051), .Q(n758) );
  AOI211 U1430 ( .A(n3), .B(regs[83]), .C(n748), .Q(n749) );
  AOI221 U1431 ( .A(n47), .B(regs[51]), .C(n19), .D(regs[19]), .Q(n750) );
  AOI221 U1432 ( .A(n33), .B(regs[211]), .C(n7), .D(regs[147]), .Q(n751) );
  AOI311 U1433 ( .A(n746), .B(n745), .C(n744), .D(n1045), .Q(n759) );
  AOI211 U1434 ( .A(n4), .B(regs[851]), .C(n743), .Q(n744) );
  AOI221 U1435 ( .A(n45), .B(regs[883]), .C(n199), .D(regs[1011]), .Q(n742) );
  AOI221 U1436 ( .A(n47), .B(regs[819]), .C(n19), .D(regs[787]), .Q(n745) );
  AOI221 U1437 ( .A(n33), .B(regs[979]), .C(n7), .D(regs[915]), .Q(n746) );
  AOI311 U1438 ( .A(n741), .B(n740), .C(n739), .D(n1039), .Q(n760) );
  AOI211 U1439 ( .A(n4), .B(regs[339]), .C(n738), .Q(n739) );
  AOI221 U1440 ( .A(n47), .B(regs[307]), .C(n19), .D(regs[275]), .Q(n740) );
  AOI221 U1441 ( .A(n33), .B(regs[467]), .C(n7), .D(regs[403]), .Q(n741) );
  AOI311 U1442 ( .A(n956), .B(n955), .C(n954), .D(n1064), .Q(n957) );
  AOI211 U1443 ( .A(n3), .B(regs[603]), .C(n953), .Q(n954) );
  AOI311 U1444 ( .A(n951), .B(n950), .C(n949), .D(n1051), .Q(n958) );
  AOI211 U1445 ( .A(n4), .B(regs[91]), .C(n948), .Q(n949) );
  AOI311 U1446 ( .A(n946), .B(n945), .C(n944), .D(n1045), .Q(n959) );
  AOI211 U1447 ( .A(n3), .B(regs[859]), .C(n943), .Q(n944) );
  AOI311 U1448 ( .A(n941), .B(n940), .C(n939), .D(n1039), .Q(n960) );
  AOI211 U1449 ( .A(n3), .B(regs[347]), .C(n938), .Q(n939) );
  AOI311 U1450 ( .A(n881), .B(n880), .C(n879), .D(n1064), .Q(n882) );
  AOI211 U1451 ( .A(n3), .B(regs[600]), .C(n878), .Q(n879) );
  AOI221 U1452 ( .A(n33), .B(regs[728]), .C(n7), .D(regs[664]), .Q(n881) );
  AOI311 U1453 ( .A(n876), .B(n875), .C(n874), .D(n1051), .Q(n883) );
  AOI211 U1454 ( .A(n3), .B(regs[88]), .C(n873), .Q(n874) );
  AOI221 U1455 ( .A(n45), .B(regs[120]), .C(n199), .D(regs[248]), .Q(n872) );
  AOI221 U1456 ( .A(n33), .B(regs[216]), .C(n7), .D(regs[152]), .Q(n876) );
  AOI311 U1457 ( .A(n871), .B(n870), .C(n869), .D(n1045), .Q(n884) );
  AOI211 U1458 ( .A(n3), .B(regs[856]), .C(n868), .Q(n869) );
  AOI221 U1459 ( .A(n45), .B(regs[888]), .C(n199), .D(regs[1016]), .Q(n867) );
  AOI221 U1460 ( .A(n33), .B(regs[984]), .C(n7), .D(regs[920]), .Q(n871) );
  AOI311 U1461 ( .A(n866), .B(n865), .C(n864), .D(n1039), .Q(n885) );
  AOI211 U1462 ( .A(n4), .B(regs[344]), .C(n863), .Q(n864) );
  AOI221 U1463 ( .A(n45), .B(regs[376]), .C(n1), .D(regs[504]), .Q(n862) );
  AOI221 U1464 ( .A(n33), .B(regs[472]), .C(n7), .D(regs[408]), .Q(n866) );
  AOI311 U1465 ( .A(n856), .B(n855), .C(n854), .D(n1064), .Q(n857) );
  AOI211 U1466 ( .A(n3), .B(regs[599]), .C(n853), .Q(n854) );
  AOI221 U1467 ( .A(n45), .B(regs[631]), .C(n199), .D(regs[759]), .Q(n852) );
  AOI221 U1468 ( .A(n33), .B(regs[727]), .C(n7), .D(regs[663]), .Q(n856) );
  AOI311 U1469 ( .A(n851), .B(n850), .C(n849), .D(n1051), .Q(n858) );
  AOI211 U1470 ( .A(n4), .B(regs[87]), .C(n848), .Q(n849) );
  AOI221 U1471 ( .A(n45), .B(regs[119]), .C(n199), .D(regs[247]), .Q(n847) );
  AOI221 U1472 ( .A(n33), .B(regs[215]), .C(n7), .D(regs[151]), .Q(n851) );
  AOI311 U1473 ( .A(n846), .B(n845), .C(n844), .D(n1045), .Q(n859) );
  AOI211 U1474 ( .A(n4), .B(regs[855]), .C(n843), .Q(n844) );
  AOI221 U1475 ( .A(n45), .B(regs[887]), .C(n199), .D(regs[1015]), .Q(n842) );
  AOI221 U1476 ( .A(n33), .B(regs[983]), .C(n7), .D(regs[919]), .Q(n846) );
  AOI311 U1477 ( .A(n841), .B(n840), .C(n839), .D(n1039), .Q(n860) );
  AOI211 U1478 ( .A(n4), .B(regs[343]), .C(n838), .Q(n839) );
  AOI221 U1479 ( .A(n45), .B(regs[375]), .C(n1), .D(regs[503]), .Q(n837) );
  AOI221 U1480 ( .A(n33), .B(regs[471]), .C(n7), .D(regs[407]), .Q(n841) );
  AOI311 U1481 ( .A(n1006), .B(n1005), .C(n1004), .D(n1064), .Q(n1007) );
  AOI211 U1482 ( .A(n4), .B(regs[605]), .C(n1003), .Q(n1004) );
  AOI221 U1483 ( .A(n33), .B(regs[733]), .C(n7), .D(regs[669]), .Q(n1006) );
  AOI311 U1484 ( .A(n1001), .B(n1000), .C(n999), .D(n1051), .Q(n1008) );
  AOI211 U1485 ( .A(n3), .B(regs[93]), .C(n998), .Q(n999) );
  AOI221 U1486 ( .A(n33), .B(regs[221]), .C(n7), .D(regs[157]), .Q(n1001) );
  AOI311 U1487 ( .A(n996), .B(n995), .C(n994), .D(n1045), .Q(n1009) );
  AOI211 U1488 ( .A(n4), .B(regs[861]), .C(n993), .Q(n994) );
  AOI221 U1489 ( .A(n33), .B(regs[989]), .C(n7), .D(regs[925]), .Q(n996) );
  AOI311 U1490 ( .A(n991), .B(n990), .C(n989), .D(n1039), .Q(n1010) );
  AOI211 U1491 ( .A(n4), .B(regs[349]), .C(n988), .Q(n989) );
  AOI311 U1492 ( .A(n931), .B(n930), .C(n929), .D(n1064), .Q(n932) );
  AOI211 U1493 ( .A(n4), .B(regs[602]), .C(n928), .Q(n929) );
  AOI221 U1494 ( .A(n45), .B(regs[634]), .C(n199), .D(regs[762]), .Q(n927) );
  AOI221 U1495 ( .A(n33), .B(regs[730]), .C(n7), .D(regs[666]), .Q(n931) );
  AOI311 U1496 ( .A(n926), .B(n925), .C(n924), .D(n1051), .Q(n933) );
  AOI211 U1497 ( .A(n3), .B(regs[90]), .C(n923), .Q(n924) );
  AOI221 U1498 ( .A(n45), .B(regs[122]), .C(n1), .D(regs[250]), .Q(n922) );
  AOI221 U1499 ( .A(n33), .B(regs[218]), .C(n7), .D(regs[154]), .Q(n926) );
  AOI311 U1500 ( .A(n921), .B(n920), .C(n919), .D(n1045), .Q(n934) );
  AOI211 U1501 ( .A(n3), .B(regs[858]), .C(n918), .Q(n919) );
  AOI221 U1502 ( .A(n45), .B(regs[890]), .C(n1), .D(regs[1018]), .Q(n917) );
  AOI221 U1503 ( .A(n33), .B(regs[986]), .C(n7), .D(regs[922]), .Q(n921) );
  AOI311 U1504 ( .A(n916), .B(n915), .C(n914), .D(n1039), .Q(n935) );
  AOI211 U1505 ( .A(n3), .B(regs[346]), .C(n913), .Q(n914) );
  AOI221 U1506 ( .A(n45), .B(regs[378]), .C(n199), .D(regs[506]), .Q(n912) );
  AOI221 U1507 ( .A(n33), .B(regs[474]), .C(n7), .D(regs[410]), .Q(n916) );
  AOI311 U1508 ( .A(n331), .B(n330), .C(n329), .D(n1064), .Q(n332) );
  AOI211 U1509 ( .A(n3), .B(regs[578]), .C(n328), .Q(n329) );
  AOI221 U1510 ( .A(n45), .B(regs[610]), .C(n1), .D(regs[738]), .Q(n327) );
  AOI221 U1511 ( .A(n33), .B(regs[706]), .C(n7), .D(regs[642]), .Q(n331) );
  AOI311 U1512 ( .A(n326), .B(n325), .C(n324), .D(n1051), .Q(n333) );
  AOI211 U1513 ( .A(n4), .B(regs[66]), .C(n323), .Q(n324) );
  AOI221 U1514 ( .A(n45), .B(regs[98]), .C(n1), .D(regs[226]), .Q(n322) );
  AOI221 U1515 ( .A(n33), .B(regs[194]), .C(n7), .D(regs[130]), .Q(n326) );
  AOI311 U1516 ( .A(n321), .B(n320), .C(n319), .D(n1045), .Q(n334) );
  AOI211 U1517 ( .A(n4), .B(regs[834]), .C(n318), .Q(n319) );
  AOI221 U1518 ( .A(n45), .B(regs[866]), .C(n1), .D(regs[994]), .Q(n317) );
  AOI221 U1519 ( .A(n33), .B(regs[962]), .C(n7), .D(regs[898]), .Q(n321) );
  AOI311 U1520 ( .A(n316), .B(n315), .C(n314), .D(n1039), .Q(n335) );
  AOI211 U1521 ( .A(n3), .B(regs[322]), .C(n313), .Q(n314) );
  AOI221 U1522 ( .A(n45), .B(regs[354]), .C(n1), .D(regs[482]), .Q(n312) );
  AOI221 U1523 ( .A(n33), .B(regs[450]), .C(n7), .D(regs[386]), .Q(n316) );
  AOI311 U1524 ( .A(n1031), .B(n1030), .C(n1029), .D(n1064), .Q(n1032) );
  AOI211 U1525 ( .A(n4), .B(regs[606]), .C(n1028), .Q(n1029) );
  AOI311 U1526 ( .A(n1026), .B(n1025), .C(n1024), .D(n1051), .Q(n1033) );
  AOI211 U1527 ( .A(n4), .B(regs[94]), .C(n1023), .Q(n1024) );
  AOI221 U1528 ( .A(n45), .B(regs[126]), .C(n199), .D(regs[254]), .Q(n1022) );
  AOI221 U1529 ( .A(n33), .B(regs[222]), .C(n7), .D(regs[158]), .Q(n1026) );
  AOI311 U1530 ( .A(n1021), .B(n1020), .C(n1019), .D(n1045), .Q(n1034) );
  AOI211 U1531 ( .A(n4), .B(regs[862]), .C(n1018), .Q(n1019) );
  AOI221 U1532 ( .A(n45), .B(regs[894]), .C(n199), .D(regs[1022]), .Q(n1017)
         );
  AOI221 U1533 ( .A(n33), .B(regs[990]), .C(n7), .D(regs[926]), .Q(n1021) );
  AOI311 U1534 ( .A(n1016), .B(n1015), .C(n1014), .D(n1039), .Q(n1035) );
  AOI211 U1535 ( .A(n3), .B(regs[350]), .C(n1013), .Q(n1014) );
  AOI221 U1536 ( .A(n45), .B(regs[382]), .C(n1), .D(regs[510]), .Q(n1012) );
  AOI221 U1537 ( .A(n33), .B(regs[478]), .C(n7), .D(regs[414]), .Q(n1016) );
  AOI311 U1538 ( .A(n981), .B(n980), .C(n979), .D(n1064), .Q(n982) );
  AOI211 U1539 ( .A(n4), .B(regs[604]), .C(n978), .Q(n979) );
  AOI311 U1540 ( .A(n976), .B(n975), .C(n974), .D(n1051), .Q(n983) );
  AOI211 U1541 ( .A(n4), .B(regs[92]), .C(n973), .Q(n974) );
  AOI311 U1542 ( .A(n971), .B(n970), .C(n969), .D(n1045), .Q(n984) );
  AOI211 U1543 ( .A(n3), .B(regs[860]), .C(n968), .Q(n969) );
  AOI311 U1544 ( .A(n966), .B(n965), .C(n964), .D(n1039), .Q(n985) );
  AOI211 U1545 ( .A(n4), .B(regs[348]), .C(n963), .Q(n964) );
  AOI311 U1546 ( .A(n1067), .B(n1066), .C(n1065), .D(n1064), .Q(n1068) );
  AOI211 U1547 ( .A(n4), .B(regs[607]), .C(n1062), .Q(n1065) );
  AOI311 U1548 ( .A(n1054), .B(n1053), .C(n1052), .D(n1051), .Q(n1069) );
  AOI211 U1549 ( .A(n3), .B(regs[95]), .C(n1050), .Q(n1052) );
  AOI221 U1550 ( .A(n45), .B(regs[127]), .C(n199), .D(regs[255]), .Q(n1049) );
  AOI221 U1551 ( .A(n33), .B(regs[223]), .C(n7), .D(regs[159]), .Q(n1054) );
  AOI311 U1552 ( .A(n1048), .B(n1047), .C(n1046), .D(n1045), .Q(n1070) );
  AOI211 U1553 ( .A(n3), .B(regs[863]), .C(n1044), .Q(n1046) );
  AOI221 U1554 ( .A(n45), .B(regs[895]), .C(n199), .D(regs[1023]), .Q(n1043)
         );
  AOI221 U1555 ( .A(n33), .B(regs[991]), .C(n7), .D(regs[927]), .Q(n1048) );
  AOI311 U1556 ( .A(n1042), .B(n1041), .C(n1040), .D(n1039), .Q(n1071) );
  AOI211 U1557 ( .A(n3), .B(regs[351]), .C(n1038), .Q(n1040) );
  AOI221 U1558 ( .A(n33), .B(regs[479]), .C(n7), .D(regs[415]), .Q(n1042) );
  AOI311 U1559 ( .A(n906), .B(n905), .C(n904), .D(n1064), .Q(n907) );
  AOI211 U1560 ( .A(n3), .B(regs[601]), .C(n903), .Q(n904) );
  AOI221 U1561 ( .A(n33), .B(regs[729]), .C(n7), .D(regs[665]), .Q(n906) );
  AOI311 U1562 ( .A(n901), .B(n900), .C(n899), .D(n1051), .Q(n908) );
  AOI211 U1563 ( .A(n3), .B(regs[89]), .C(n898), .Q(n899) );
  AOI221 U1564 ( .A(n45), .B(regs[121]), .C(n199), .D(regs[249]), .Q(n897) );
  AOI221 U1565 ( .A(n33), .B(regs[217]), .C(n7), .D(regs[153]), .Q(n901) );
  AOI311 U1566 ( .A(n896), .B(n895), .C(n894), .D(n1045), .Q(n909) );
  AOI211 U1567 ( .A(n4), .B(regs[857]), .C(n893), .Q(n894) );
  AOI221 U1568 ( .A(n45), .B(regs[889]), .C(n199), .D(regs[1017]), .Q(n892) );
  AOI221 U1569 ( .A(n33), .B(regs[985]), .C(n7), .D(regs[921]), .Q(n896) );
  AOI311 U1570 ( .A(n891), .B(n890), .C(n889), .D(n1039), .Q(n910) );
  AOI211 U1571 ( .A(n4), .B(regs[345]), .C(n888), .Q(n889) );
  AOI221 U1572 ( .A(n45), .B(regs[377]), .C(n1), .D(regs[505]), .Q(n887) );
  AOI221 U1573 ( .A(n33), .B(regs[473]), .C(n7), .D(regs[409]), .Q(n891) );
  AOI311 U1574 ( .A(n831), .B(n830), .C(n829), .D(n1064), .Q(n832) );
  AOI211 U1575 ( .A(n3), .B(regs[598]), .C(n828), .Q(n829) );
  AOI311 U1576 ( .A(n826), .B(n825), .C(n824), .D(n1051), .Q(n833) );
  AOI211 U1577 ( .A(n4), .B(regs[86]), .C(n823), .Q(n824) );
  AOI221 U1578 ( .A(n33), .B(regs[214]), .C(n7), .D(regs[150]), .Q(n826) );
  AOI311 U1579 ( .A(n821), .B(n820), .C(n819), .D(n1045), .Q(n834) );
  AOI211 U1580 ( .A(n3), .B(regs[854]), .C(n818), .Q(n819) );
  AOI221 U1581 ( .A(n33), .B(regs[982]), .C(n7), .D(regs[918]), .Q(n821) );
  AOI311 U1582 ( .A(n816), .B(n815), .C(n814), .D(n1039), .Q(n835) );
  AOI211 U1583 ( .A(n4), .B(regs[342]), .C(n813), .Q(n814) );
  AOI221 U1584 ( .A(n33), .B(regs[470]), .C(n7), .D(regs[406]), .Q(n816) );
  AOI311 U1585 ( .A(n581), .B(n580), .C(n579), .D(n1064), .Q(n582) );
  AOI211 U1586 ( .A(n4), .B(regs[588]), .C(n578), .Q(n579) );
  AOI221 U1587 ( .A(n45), .B(regs[620]), .C(n1), .D(regs[748]), .Q(n577) );
  AOI221 U1588 ( .A(n33), .B(regs[716]), .C(n7), .D(regs[652]), .Q(n581) );
  AOI311 U1589 ( .A(n576), .B(n575), .C(n574), .D(n1051), .Q(n583) );
  AOI211 U1590 ( .A(n4), .B(regs[76]), .C(n573), .Q(n574) );
  AOI221 U1591 ( .A(n45), .B(regs[108]), .C(n1), .D(regs[236]), .Q(n572) );
  AOI221 U1592 ( .A(n33), .B(regs[204]), .C(n7), .D(regs[140]), .Q(n576) );
  AOI311 U1593 ( .A(n571), .B(n570), .C(n569), .D(n1045), .Q(n584) );
  AOI211 U1594 ( .A(n4), .B(regs[844]), .C(n568), .Q(n569) );
  AOI221 U1595 ( .A(n45), .B(regs[876]), .C(n1), .D(regs[1004]), .Q(n567) );
  AOI221 U1596 ( .A(n33), .B(regs[972]), .C(n7), .D(regs[908]), .Q(n571) );
  AOI311 U1597 ( .A(n566), .B(n565), .C(n564), .D(n1039), .Q(n585) );
  AOI211 U1598 ( .A(n3), .B(regs[332]), .C(n563), .Q(n564) );
  AOI221 U1599 ( .A(n45), .B(regs[364]), .C(n1), .D(regs[492]), .Q(n562) );
  AOI221 U1600 ( .A(n33), .B(regs[460]), .C(n7), .D(regs[396]), .Q(n566) );
  AOI311 U1601 ( .A(n631), .B(n630), .C(n629), .D(n1064), .Q(n632) );
  AOI211 U1602 ( .A(n4), .B(regs[590]), .C(n628), .Q(n629) );
  AOI221 U1603 ( .A(n45), .B(regs[622]), .C(n1), .D(regs[750]), .Q(n627) );
  AOI311 U1604 ( .A(n626), .B(n625), .C(n624), .D(n1051), .Q(n633) );
  AOI211 U1605 ( .A(n3), .B(regs[78]), .C(n623), .Q(n624) );
  AOI221 U1606 ( .A(n45), .B(regs[110]), .C(n1), .D(regs[238]), .Q(n622) );
  AOI221 U1607 ( .A(n33), .B(regs[206]), .C(n7), .D(regs[142]), .Q(n626) );
  AOI311 U1608 ( .A(n621), .B(n620), .C(n619), .D(n1045), .Q(n634) );
  AOI211 U1609 ( .A(n3), .B(regs[846]), .C(n618), .Q(n619) );
  AOI221 U1610 ( .A(n45), .B(regs[878]), .C(n51), .D(regs[1006]), .Q(n617) );
  AOI221 U1611 ( .A(n33), .B(regs[974]), .C(n7), .D(regs[910]), .Q(n621) );
  AOI311 U1612 ( .A(n616), .B(n615), .C(n614), .D(n1039), .Q(n635) );
  AOI211 U1613 ( .A(n3), .B(regs[334]), .C(n613), .Q(n614) );
  AOI221 U1614 ( .A(n45), .B(regs[366]), .C(n1), .D(regs[494]), .Q(n612) );
  AOI221 U1615 ( .A(n33), .B(regs[462]), .C(n7), .D(regs[398]), .Q(n616) );
  AOI311 U1616 ( .A(n606), .B(n605), .C(n604), .D(n1064), .Q(n607) );
  AOI211 U1617 ( .A(n3), .B(regs[589]), .C(n603), .Q(n604) );
  AOI311 U1618 ( .A(n601), .B(n600), .C(n599), .D(n1051), .Q(n608) );
  AOI211 U1619 ( .A(n4), .B(regs[77]), .C(n598), .Q(n599) );
  AOI221 U1620 ( .A(n45), .B(regs[109]), .C(n1), .D(regs[237]), .Q(n597) );
  AOI311 U1621 ( .A(n596), .B(n595), .C(n594), .D(n1045), .Q(n609) );
  AOI211 U1622 ( .A(n4), .B(regs[845]), .C(n593), .Q(n594) );
  AOI221 U1623 ( .A(n45), .B(regs[877]), .C(n199), .D(regs[1005]), .Q(n592) );
  AOI221 U1624 ( .A(n33), .B(regs[973]), .C(n7), .D(regs[909]), .Q(n596) );
  AOI311 U1625 ( .A(n591), .B(n590), .C(n589), .D(n1039), .Q(n610) );
  AOI211 U1626 ( .A(n3), .B(regs[333]), .C(n588), .Q(n589) );
  AOI221 U1627 ( .A(n45), .B(regs[365]), .C(n199), .D(regs[493]), .Q(n587) );
  AOI221 U1628 ( .A(n33), .B(regs[461]), .C(n7), .D(regs[397]), .Q(n591) );
  AOI311 U1629 ( .A(n731), .B(n730), .C(n729), .D(n1064), .Q(n732) );
  AOI211 U1630 ( .A(n4), .B(regs[594]), .C(n728), .Q(n729) );
  AOI221 U1631 ( .A(n47), .B(regs[562]), .C(n19), .D(regs[530]), .Q(n730) );
  AOI221 U1632 ( .A(n33), .B(regs[722]), .C(n7), .D(regs[658]), .Q(n731) );
  AOI311 U1633 ( .A(n726), .B(n725), .C(n724), .D(n1051), .Q(n733) );
  AOI211 U1634 ( .A(n4), .B(regs[82]), .C(n723), .Q(n724) );
  AOI221 U1635 ( .A(n45), .B(regs[114]), .C(n199), .D(regs[242]), .Q(n722) );
  AOI221 U1636 ( .A(n47), .B(regs[50]), .C(n19), .D(regs[18]), .Q(n725) );
  AOI221 U1637 ( .A(n33), .B(regs[210]), .C(n7), .D(regs[146]), .Q(n726) );
  AOI311 U1638 ( .A(n721), .B(n720), .C(n719), .D(n1045), .Q(n734) );
  AOI211 U1639 ( .A(n3), .B(regs[850]), .C(n718), .Q(n719) );
  AOI221 U1640 ( .A(n47), .B(regs[818]), .C(n19), .D(regs[786]), .Q(n720) );
  AOI221 U1641 ( .A(n33), .B(regs[978]), .C(n7), .D(regs[914]), .Q(n721) );
  AOI311 U1642 ( .A(n716), .B(n715), .C(n714), .D(n1039), .Q(n735) );
  AOI211 U1643 ( .A(n3), .B(regs[338]), .C(n713), .Q(n714) );
  AOI221 U1644 ( .A(n45), .B(regs[370]), .C(n199), .D(regs[498]), .Q(n712) );
  AOI221 U1645 ( .A(n47), .B(regs[306]), .C(n19), .D(regs[274]), .Q(n715) );
  AOI221 U1646 ( .A(n33), .B(regs[466]), .C(n7), .D(regs[402]), .Q(n716) );
  AOI311 U1647 ( .A(n556), .B(n555), .C(n554), .D(n1064), .Q(n557) );
  AOI211 U1648 ( .A(n3), .B(regs[587]), .C(n553), .Q(n554) );
  AOI221 U1649 ( .A(n45), .B(regs[619]), .C(n1), .D(regs[747]), .Q(n552) );
  AOI221 U1650 ( .A(n33), .B(regs[715]), .C(n7), .D(regs[651]), .Q(n556) );
  AOI311 U1651 ( .A(n551), .B(n550), .C(n549), .D(n1051), .Q(n558) );
  AOI211 U1652 ( .A(n3), .B(regs[75]), .C(n548), .Q(n549) );
  AOI221 U1653 ( .A(n45), .B(regs[107]), .C(n1), .D(regs[235]), .Q(n547) );
  AOI221 U1654 ( .A(n33), .B(regs[203]), .C(n7), .D(regs[139]), .Q(n551) );
  AOI311 U1655 ( .A(n546), .B(n545), .C(n544), .D(n1045), .Q(n559) );
  AOI211 U1656 ( .A(n4), .B(regs[843]), .C(n543), .Q(n544) );
  AOI221 U1657 ( .A(n45), .B(regs[875]), .C(n199), .D(regs[1003]), .Q(n542) );
  AOI221 U1658 ( .A(n33), .B(regs[971]), .C(n7), .D(regs[907]), .Q(n546) );
  AOI311 U1659 ( .A(n541), .B(n540), .C(n539), .D(n1039), .Q(n560) );
  AOI211 U1660 ( .A(n3), .B(regs[331]), .C(n538), .Q(n539) );
  AOI221 U1661 ( .A(n45), .B(regs[363]), .C(n199), .D(regs[491]), .Q(n537) );
  AOI221 U1662 ( .A(n33), .B(regs[459]), .C(n7), .D(regs[395]), .Q(n541) );
  AOI311 U1663 ( .A(n531), .B(n530), .C(n529), .D(n1064), .Q(n532) );
  AOI211 U1664 ( .A(n3), .B(regs[586]), .C(n528), .Q(n529) );
  AOI221 U1665 ( .A(n45), .B(regs[618]), .C(n199), .D(regs[746]), .Q(n527) );
  AOI221 U1666 ( .A(n33), .B(regs[714]), .C(n7), .D(regs[650]), .Q(n531) );
  AOI311 U1667 ( .A(n526), .B(n525), .C(n524), .D(n1051), .Q(n533) );
  AOI211 U1668 ( .A(n4), .B(regs[74]), .C(n523), .Q(n524) );
  AOI221 U1669 ( .A(n45), .B(regs[106]), .C(n199), .D(regs[234]), .Q(n522) );
  AOI221 U1670 ( .A(n33), .B(regs[202]), .C(n7), .D(regs[138]), .Q(n526) );
  AOI311 U1671 ( .A(n521), .B(n520), .C(n519), .D(n1045), .Q(n534) );
  AOI211 U1672 ( .A(n4), .B(regs[842]), .C(n518), .Q(n519) );
  AOI221 U1673 ( .A(n45), .B(regs[874]), .C(n199), .D(regs[1002]), .Q(n517) );
  AOI221 U1674 ( .A(n33), .B(regs[970]), .C(n7), .D(regs[906]), .Q(n521) );
  AOI311 U1675 ( .A(n516), .B(n515), .C(n514), .D(n1039), .Q(n535) );
  AOI211 U1676 ( .A(n3), .B(regs[330]), .C(n513), .Q(n514) );
  AOI221 U1677 ( .A(n45), .B(regs[362]), .C(n199), .D(regs[490]), .Q(n512) );
  AOI221 U1678 ( .A(n33), .B(regs[458]), .C(n7), .D(regs[394]), .Q(n516) );
  AOI311 U1679 ( .A(n506), .B(n505), .C(n504), .D(n1064), .Q(n507) );
  AOI211 U1680 ( .A(n4), .B(regs[585]), .C(n503), .Q(n504) );
  AOI221 U1681 ( .A(n45), .B(regs[617]), .C(n1), .D(regs[745]), .Q(n502) );
  AOI221 U1682 ( .A(n33), .B(regs[713]), .C(n7), .D(regs[649]), .Q(n506) );
  AOI311 U1683 ( .A(n501), .B(n500), .C(n499), .D(n1051), .Q(n508) );
  AOI211 U1684 ( .A(n4), .B(regs[73]), .C(n498), .Q(n499) );
  AOI221 U1685 ( .A(n45), .B(regs[105]), .C(n199), .D(regs[233]), .Q(n497) );
  AOI221 U1686 ( .A(n33), .B(regs[201]), .C(n7), .D(regs[137]), .Q(n501) );
  AOI311 U1687 ( .A(n496), .B(n495), .C(n494), .D(n1045), .Q(n509) );
  AOI211 U1688 ( .A(n3), .B(regs[841]), .C(n493), .Q(n494) );
  AOI221 U1689 ( .A(n45), .B(regs[873]), .C(n1), .D(regs[1001]), .Q(n492) );
  AOI221 U1690 ( .A(n33), .B(regs[969]), .C(n7), .D(regs[905]), .Q(n496) );
  AOI311 U1691 ( .A(n491), .B(n490), .C(n489), .D(n1039), .Q(n510) );
  AOI211 U1692 ( .A(n4), .B(regs[329]), .C(n488), .Q(n489) );
  AOI221 U1693 ( .A(n45), .B(regs[361]), .C(n1), .D(regs[489]), .Q(n487) );
  AOI221 U1694 ( .A(n33), .B(regs[457]), .C(n7), .D(regs[393]), .Q(n491) );
  AOI311 U1695 ( .A(n656), .B(n655), .C(n654), .D(n1064), .Q(n657) );
  AOI211 U1696 ( .A(n4), .B(regs[591]), .C(n653), .Q(n654) );
  AOI311 U1697 ( .A(n651), .B(n650), .C(n649), .D(n1051), .Q(n658) );
  AOI211 U1698 ( .A(n4), .B(regs[79]), .C(n648), .Q(n649) );
  AOI221 U1699 ( .A(n45), .B(regs[111]), .C(n1), .D(regs[239]), .Q(n647) );
  AOI311 U1700 ( .A(n646), .B(n645), .C(n644), .D(n1045), .Q(n659) );
  AOI211 U1701 ( .A(n3), .B(regs[847]), .C(n643), .Q(n644) );
  AOI221 U1702 ( .A(n45), .B(regs[879]), .C(n1), .D(regs[1007]), .Q(n642) );
  AOI221 U1703 ( .A(n33), .B(regs[975]), .C(n7), .D(regs[911]), .Q(n646) );
  AOI311 U1704 ( .A(n641), .B(n640), .C(n639), .D(n1039), .Q(n660) );
  AOI211 U1705 ( .A(n3), .B(regs[335]), .C(n638), .Q(n639) );
  AOI221 U1706 ( .A(n45), .B(regs[367]), .C(n1), .D(regs[495]), .Q(n637) );
  AOI311 U1707 ( .A(n706), .B(n705), .C(n704), .D(n1064), .Q(n707) );
  AOI311 U1708 ( .A(n701), .B(n700), .C(n699), .D(n1051), .Q(n708) );
  AOI211 U1709 ( .A(n3), .B(regs[81]), .C(n698), .Q(n699) );
  AOI311 U1710 ( .A(n696), .B(n695), .C(n694), .D(n1045), .Q(n709) );
  AOI211 U1711 ( .A(n4), .B(regs[849]), .C(n693), .Q(n694) );
  AOI311 U1712 ( .A(n691), .B(n690), .C(n689), .D(n1039), .Q(n710) );
  AOI211 U1713 ( .A(n4), .B(regs[337]), .C(n688), .Q(n689) );
  AOI311 U1714 ( .A(n681), .B(n680), .C(n679), .D(n1064), .Q(n682) );
  AOI211 U1715 ( .A(n3), .B(regs[592]), .C(n678), .Q(n679) );
  AOI311 U1716 ( .A(n676), .B(n675), .C(n674), .D(n1051), .Q(n683) );
  AOI211 U1717 ( .A(n3), .B(regs[80]), .C(n673), .Q(n674) );
  AOI311 U1718 ( .A(n671), .B(n670), .C(n669), .D(n1045), .Q(n684) );
  AOI211 U1719 ( .A(n4), .B(regs[848]), .C(n668), .Q(n669) );
  AOI311 U1720 ( .A(n666), .B(n665), .C(n664), .D(n1039), .Q(n685) );
  AOI211 U1721 ( .A(n3), .B(regs[336]), .C(n663), .Q(n664) );
  AOI221 U1722 ( .A(n33), .B(regs[464]), .C(n7), .D(regs[400]), .Q(n666) );
  NAND22 U1723 ( .A(n270), .B(i_addr_Rs[0]), .Q(n1061) );
  AOI210 U1724 ( .A(n3), .B(regs[321]), .C(n298), .Q(n301) );
  AOI220 U1725 ( .A(n1056), .B(regs[731]), .C(n7), .D(regs[667]), .Q(n956) );
  AOI220 U1726 ( .A(n1056), .B(regs[219]), .C(n7), .D(regs[155]), .Q(n951) );
  AOI220 U1727 ( .A(n1056), .B(regs[987]), .C(n7), .D(regs[923]), .Q(n946) );
  AOI220 U1728 ( .A(n1056), .B(regs[475]), .C(n7), .D(regs[411]), .Q(n941) );
  AOI220 U1729 ( .A(n1056), .B(regs[477]), .C(n7), .D(regs[413]), .Q(n991) );
  AOI220 U1730 ( .A(n1056), .B(regs[732]), .C(n7), .D(regs[668]), .Q(n981) );
  AOI220 U1731 ( .A(n1056), .B(regs[220]), .C(n7), .D(regs[156]), .Q(n976) );
  AOI220 U1732 ( .A(n1056), .B(regs[988]), .C(n7), .D(regs[924]), .Q(n971) );
  AOI220 U1733 ( .A(n1056), .B(regs[476]), .C(n7), .D(regs[412]), .Q(n966) );
  AOI220 U1734 ( .A(n1056), .B(regs[735]), .C(n7), .D(regs[671]), .Q(n1067) );
  AOI220 U1735 ( .A(n1056), .B(regs[718]), .C(n7), .D(regs[654]), .Q(n631) );
  AOI220 U1736 ( .A(n1056), .B(regs[717]), .C(n7), .D(regs[653]), .Q(n606) );
  AOI220 U1737 ( .A(n1056), .B(regs[205]), .C(n7), .D(regs[141]), .Q(n601) );
  AOI220 U1738 ( .A(n1056), .B(regs[719]), .C(n7), .D(regs[655]), .Q(n656) );
  AOI220 U1739 ( .A(n1056), .B(regs[207]), .C(n7), .D(regs[143]), .Q(n651) );
  AOI220 U1740 ( .A(n1056), .B(regs[463]), .C(n7), .D(regs[399]), .Q(n641) );
  AOI220 U1741 ( .A(n1056), .B(regs[721]), .C(n7), .D(regs[657]), .Q(n706) );
  AOI220 U1742 ( .A(n1056), .B(regs[209]), .C(n7), .D(regs[145]), .Q(n701) );
  AOI220 U1743 ( .A(n1056), .B(regs[977]), .C(n7), .D(regs[913]), .Q(n696) );
  AOI220 U1744 ( .A(n1056), .B(regs[465]), .C(n7), .D(regs[401]), .Q(n691) );
  AOI220 U1745 ( .A(n1056), .B(regs[720]), .C(n7), .D(regs[656]), .Q(n681) );
  AOI220 U1746 ( .A(n1056), .B(regs[208]), .C(n7), .D(regs[144]), .Q(n676) );
  AOI220 U1747 ( .A(n1056), .B(regs[976]), .C(n7), .D(regs[912]), .Q(n671) );
  AOI220 U1748 ( .A(n1785), .B(regs[864]), .C(n48), .D(regs[800]), .Q(n1081)
         );
  AOI220 U1749 ( .A(n1787), .B(regs[832]), .C(n24), .D(regs[768]), .Q(n1080)
         );
  AOI220 U1750 ( .A(regs[608]), .B(n1785), .C(regs[544]), .D(n48), .Q(n1093)
         );
  AOI220 U1751 ( .A(n1785), .B(regs[359]), .C(n48), .D(regs[295]), .Q(n1241)
         );
  AOI220 U1752 ( .A(n1785), .B(regs[103]), .C(n48), .D(regs[39]), .Q(n1251) );
  AOI220 U1753 ( .A(n1785), .B(regs[360]), .C(n48), .D(regs[296]), .Q(n1263)
         );
  AOI220 U1754 ( .A(n1785), .B(regs[382]), .C(n48), .D(regs[318]), .Q(n1747)
         );
  AOI220 U1755 ( .A(n1787), .B(regs[350]), .C(n24), .D(regs[286]), .Q(n1746)
         );
  AOI220 U1756 ( .A(n1785), .B(regs[126]), .C(n48), .D(regs[62]), .Q(n1757) );
  AOI220 U1757 ( .A(n1787), .B(regs[94]), .C(n24), .D(regs[30]), .Q(n1756) );
  AOI220 U1758 ( .A(n1785), .B(regs[383]), .C(n48), .D(regs[319]), .Q(n1769)
         );
  AOI220 U1759 ( .A(n1787), .B(regs[351]), .C(n24), .D(regs[287]), .Q(n1768)
         );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, id_con_Wregwrite, ex_con_Wregwrite, mem_con_Wregwrite,
         for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst, ex_con_Mmemread,
         ex_con_Mmemwrite, ex_con_Malupc8, ex_con_Wmemtoreg, mem_con_Malupc8,
         mem_con_Wmemtoreg, wb_con_Wmemtoreg, u_fetch_jmux_i_addr_pc4_3_,
         u_fetch_jmux_i_addr_pc4_4_, u_fetch_jmux_i_addr_pc4_5_,
         u_fetch_jmux_i_addr_pc4_6_, u_fetch_jmux_i_addr_pc4_7_,
         u_fetch_jmux_i_addr_pc4_8_, u_fetch_jmux_i_addr_pc4_9_,
         u_fetch_jmux_i_addr_pc4_10_, u_fetch_jmux_i_addr_pc4_11_,
         u_fetch_jmux_i_addr_pc4_12_, u_fetch_jmux_i_addr_pc4_13_,
         u_fetch_jmux_i_addr_pc4_14_, u_fetch_jmux_i_addr_pc4_15_,
         u_fetch_jmux_i_addr_pc4_16_, u_fetch_jmux_i_addr_pc4_17_,
         u_fetch_jmux_i_addr_pc4_18_, u_fetch_jmux_i_addr_pc4_19_,
         u_fetch_jmux_i_addr_pc4_20_, u_fetch_jmux_i_addr_pc4_21_,
         u_fetch_jmux_i_addr_pc4_22_, u_fetch_jmux_i_addr_pc4_23_,
         u_fetch_jmux_i_addr_pc4_24_, u_fetch_jmux_i_addr_pc4_25_,
         u_fetch_jmux_i_addr_pc4_26_, u_fetch_jmux_i_addr_pc4_27_,
         u_fetch_jmux_i_addr_pc4_28_, u_fetch_jmux_i_addr_pc4_29_,
         u_fetch_jmux_i_addr_pc4_30_, u_fetch_jmux_i_addr_pc4_31_, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, u_decode_n6,
         u_decode_n1, u_decode_for_o_con_fa_0_, u_decode_for_o_con_fa_1_,
         u_decode_for_o_con_fa_2_, u_decode_control_o_con_regwrite,
         u_decode_control_o_con_memwrite, u_decode_control_o_con_memread,
         u_decode_jbcon_o_con_aluPC4, u_decode_control_o_con_regdst,
         u_decode_control_o_con_alusrc, u_decode_control_o_con_aluop_0_,
         u_decode_control_o_con_aluop_1_, u_decode_control_o_con_aluop_2_,
         u_decode_control_o_con_aluop_3_, u_decode_control_o_con_aluop_4_,
         u_decode_control_o_con_aluop_5_, u_decode_add_x_16_n217,
         u_decode_add_x_16_n216, u_decode_add_x_16_n213,
         u_decode_add_x_16_n211, u_decode_add_x_16_n210,
         u_decode_add_x_16_n208, u_decode_add_x_16_n206,
         u_decode_add_x_16_n204, u_decode_add_x_16_n201,
         u_decode_add_x_16_n199, u_decode_add_x_16_n197,
         u_decode_add_x_16_n195, u_decode_add_x_16_n190,
         u_decode_add_x_16_n188, u_decode_add_x_16_n187,
         u_decode_add_x_16_n186, u_decode_add_x_16_n185,
         u_decode_add_x_16_n184, u_decode_add_x_16_n183,
         u_decode_add_x_16_n182, u_decode_add_x_16_n181,
         u_decode_add_x_16_n180, u_decode_add_x_16_n179,
         u_decode_add_x_16_n178, u_decode_add_x_16_n177,
         u_decode_add_x_16_n176, u_decode_add_x_16_n175,
         u_decode_add_x_16_n174, u_decode_add_x_16_n170,
         u_decode_add_x_16_n169, u_decode_add_x_16_n168,
         u_decode_add_x_16_n167, u_decode_add_x_16_n166,
         u_decode_add_x_16_n165, u_decode_add_x_16_n164,
         u_decode_add_x_16_n163, u_decode_add_x_16_n162,
         u_decode_add_x_16_n161, u_decode_add_x_16_n160,
         u_decode_add_x_16_n159, u_decode_add_x_16_n158,
         u_decode_add_x_16_n157, u_decode_add_x_16_n156,
         u_decode_add_x_16_n155, u_decode_add_x_16_n154,
         u_decode_add_x_16_n153, u_decode_add_x_16_n152,
         u_decode_add_x_16_n151, u_decode_add_x_16_n150,
         u_decode_add_x_16_n149, u_decode_add_x_16_n148,
         u_decode_add_x_16_n147, u_decode_add_x_16_n146,
         u_decode_add_x_16_n145, u_decode_add_x_16_n144,
         u_decode_add_x_16_n143, u_decode_add_x_16_n139,
         u_decode_add_x_16_n138, u_decode_add_x_16_n137,
         u_decode_add_x_16_n136, u_decode_add_x_16_n135,
         u_decode_add_x_16_n134, u_decode_add_x_16_n133,
         u_decode_add_x_16_n132, u_decode_add_x_16_n131,
         u_decode_add_x_16_n130, u_decode_add_x_16_n126,
         u_decode_add_x_16_n125, u_decode_add_x_16_n124,
         u_decode_add_x_16_n123, u_decode_add_x_16_n122,
         u_decode_add_x_16_n121, u_decode_add_x_16_n120,
         u_decode_add_x_16_n119, u_decode_add_x_16_n118,
         u_decode_add_x_16_n114, u_decode_add_x_16_n113,
         u_decode_add_x_16_n112, u_decode_add_x_16_n111,
         u_decode_add_x_16_n109, u_decode_add_x_16_n106,
         u_decode_add_x_16_n105, u_decode_add_x_16_n104,
         u_decode_add_x_16_n103, u_decode_add_x_16_n99, u_decode_add_x_16_n98,
         u_decode_add_x_16_n97, u_decode_add_x_16_n96, u_decode_add_x_16_n95,
         u_decode_add_x_16_n94, u_decode_add_x_16_n93, u_decode_add_x_16_n92,
         u_decode_add_x_16_n91, u_decode_add_x_16_n90, u_decode_add_x_16_n89,
         u_decode_add_x_16_n88, u_decode_add_x_16_n87, u_decode_add_x_16_n86,
         u_decode_add_x_16_n85, u_decode_add_x_16_n84, u_decode_add_x_16_n83,
         u_decode_add_x_16_n82, u_decode_add_x_16_n81, u_decode_add_x_16_n80,
         u_decode_add_x_16_n79, u_decode_add_x_16_n78, u_decode_add_x_16_n77,
         u_decode_add_x_16_n76, u_decode_add_x_16_n75, u_decode_add_x_16_n74,
         u_decode_add_x_16_n73, u_decode_add_x_16_n72, u_decode_add_x_16_n71,
         u_decode_add_x_16_n70, u_decode_add_x_16_n69, u_decode_add_x_16_n68,
         u_decode_add_x_16_n67, u_decode_add_x_16_n66, u_decode_add_x_16_n65,
         u_decode_add_x_16_n64, u_decode_add_x_16_n63, u_decode_add_x_16_n62,
         u_decode_add_x_16_n61, u_decode_add_x_16_n60, u_decode_add_x_16_n59,
         u_decode_add_x_16_n58, u_decode_add_x_16_n57, u_decode_add_x_16_n56,
         u_decode_add_x_16_n55, u_decode_add_x_16_n54, u_decode_add_x_16_n53,
         u_decode_add_x_16_n52, u_decode_add_x_16_n51, u_decode_add_x_16_n50,
         u_decode_add_x_16_n49, u_decode_add_x_16_n48, u_decode_add_x_16_n47,
         u_decode_add_x_16_n46, u_decode_add_x_16_n45, u_decode_add_x_16_n44,
         u_decode_add_x_16_n43, u_decode_add_x_16_n42, u_decode_add_x_16_n41,
         u_decode_add_x_16_n40, u_decode_add_x_16_n39, u_decode_add_x_16_n38,
         u_decode_add_x_16_n37, u_decode_add_x_16_n36, u_decode_add_x_16_n35,
         u_decode_add_x_16_n34, u_decode_add_x_16_n32, u_decode_add_x_16_n31,
         u_decode_add_x_16_n27, u_decode_add_x_16_n26, u_decode_add_x_16_n23,
         u_decode_add_x_16_n21, u_decode_add_x_16_n20, u_decode_add_x_16_n18,
         u_decode_add_x_16_n16, u_decode_add_x_16_n14, u_decode_add_x_16_n11,
         u_decode_add_x_16_n10, u_decode_add_x_16_n9, u_decode_add_x_16_n8,
         u_decode_add_x_16_n7, u_decode_add_x_16_n5, u_decode_add_x_16_n4,
         u_decode_add_x_16_n2, add_x_4_n121, add_x_4_n116, add_x_4_n115,
         add_x_4_n112, add_x_4_n109, add_x_4_n108, add_x_4_n107, add_x_4_n103,
         add_x_4_n100, add_x_4_n99, add_x_4_n96, add_x_4_n93, add_x_4_n92,
         add_x_4_n91, add_x_4_n90, add_x_4_n87, add_x_4_n84, add_x_4_n83,
         add_x_4_n82, add_x_4_n78, add_x_4_n75, add_x_4_n74, add_x_4_n73,
         add_x_4_n72, add_x_4_n68, add_x_4_n65, add_x_4_n64, add_x_4_n63,
         add_x_4_n59, add_x_4_n56, add_x_4_n55, add_x_4_n54, add_x_4_n53,
         add_x_4_n52, add_x_4_n48, add_x_4_n45, add_x_4_n44, add_x_4_n41,
         add_x_4_n38, add_x_4_n37, add_x_4_n36, add_x_4_n35, add_x_4_n34,
         add_x_4_n30, add_x_4_n27, add_x_4_n26, add_x_4_n25, add_x_4_n21,
         add_x_4_n16, add_x_4_n15, add_x_4_n12, add_x_4_n9, add_x_4_n8,
         add_x_4_n7, add_x_4_n5, add_x_4_n2, add_x_4_n1, add_x_1_n118,
         add_x_1_n113, add_x_1_n112, add_x_1_n106, add_x_1_n105, add_x_1_n104,
         add_x_1_n103, add_x_1_n97, add_x_1_n96, add_x_1_n90, add_x_1_n89,
         add_x_1_n88, add_x_1_n87, add_x_1_n81, add_x_1_n80, add_x_1_n79,
         add_x_1_n78, add_x_1_n72, add_x_1_n71, add_x_1_n70, add_x_1_n69,
         add_x_1_n68, add_x_1_n62, add_x_1_n61, add_x_1_n60, add_x_1_n59,
         add_x_1_n50, add_x_1_n49, add_x_1_n48, add_x_1_n42, add_x_1_n41,
         add_x_1_n35, add_x_1_n34, add_x_1_n33, add_x_1_n32, add_x_1_n31,
         add_x_1_n30, add_x_1_n24, add_x_1_n23, add_x_1_n22, add_x_1_n21,
         add_x_1_n13, add_x_1_n12, add_x_1_n6, add_x_1_n5, add_x_1_n4,
         add_x_1_n3, add_x_1_n2, add_x_1_n1, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588;
  wire   [31:2] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [27:2] id_addr_pc4;
  wire   [31:26] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] wb_data_memout;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] mem_data_alures;
  wire   [31:2] mem_data_pc4;
  wire   [31:0] u_mem_resmux_o_data_alu;
  wire   [31:0] u_mem_pc8;
  wire   [1:0] u_decode_jbcon_o_con_bop;
  wire   [31:0] u_decode_pcadd_o_addr_pcbranchE;
  wire   [2:0] u_decode_for_o_con_fb;
  wire   [31:0] u_decode_regbank_o_data_Rt;

  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext({n341, 
        n341, n341, n341, n341, n341, n341, n341, n341, n341, n341, n341, n341, 
        n341, n341, ex_data_immext[31], ex_addr_rd, ex_data_immext[10:0]}), 
        .i_addr_rt(ex_addr_rt), .i_addr_rd({n341, n341, n341, n341, n341}), 
        .i_data_FEalures(data_address), .i_data_FMalures(mem_data_alures), 
        .i_data_FMmemout(wb_data_memout), .i_data_FWmemout(for_memout), 
        .i_con_Efamux(for_o_con_Efamux), .i_con_Efbmux(for_o_con_Efbmux), 
        .i_con_Ealuop(ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), 
        .i_con_Mmemwrite(ex_con_Mmemwrite), .i_con_Malupc8(ex_con_Malupc8), 
        .i_con_Wmemtoreg(ex_con_Wmemtoreg), .i_con_Wregwrite(ex_con_Wregwrite), 
        .i_con_bop(ex_con_bop), .o_data_pc4({mem_data_pc4, u_mem_pc8[1:0]}), 
        .o_data_alures(data_address), .o_data_rt(write_data), .o_addr_regdst(
        mem_addr_regdst), .o_con_Mmemread(mem_read), .o_con_Mmemwrite(
        mem_write), .o_con_Malupc8(mem_con_Malupc8), .o_con_Wmemtoreg(
        mem_con_Wmemtoreg), .o_con_Wregwrite(mem_con_Wregwrite), .o_addr_Erd(
        for_o_addr_Erd), .o_addr_Mrt(for_addr_rtM), .o_con_ifbranch(if_con_b)
         );
  DFC1 u_fetch_pipe_pc4_reg_0_ ( .D(instruction_address[0]), .C(clk), .RN(
        rst_n), .Q(u_decode_pcadd_o_addr_pcbranchE[0]) );
  DFC1 u_fetch_pipe_pc4_reg_1_ ( .D(instruction_address[1]), .C(clk), .RN(
        rst_n), .Q(u_decode_pcadd_o_addr_pcbranchE[1]) );
  DFC1 u_fetch_pipe_pc4_reg_2_ ( .D(n276), .C(clk), .RN(rst_n), .Q(
        id_addr_pc4[2]) );
  DFC1 u_fetch_pipe_pc4_reg_3_ ( .D(u_fetch_jmux_i_addr_pc4_3_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[3]) );
  DFC1 u_fetch_pipe_pc4_reg_4_ ( .D(u_fetch_jmux_i_addr_pc4_4_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[4]) );
  DFC1 u_fetch_pipe_pc4_reg_5_ ( .D(u_fetch_jmux_i_addr_pc4_5_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[5]) );
  DFC1 u_fetch_pipe_pc4_reg_6_ ( .D(u_fetch_jmux_i_addr_pc4_6_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[6]) );
  DFC1 u_fetch_pipe_pc4_reg_7_ ( .D(u_fetch_jmux_i_addr_pc4_7_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[7]) );
  DFC1 u_fetch_pipe_pc4_reg_8_ ( .D(u_fetch_jmux_i_addr_pc4_8_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[8]) );
  DFC1 u_fetch_pipe_pc4_reg_9_ ( .D(u_fetch_jmux_i_addr_pc4_9_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[9]) );
  DFC1 u_fetch_pipe_pc4_reg_10_ ( .D(u_fetch_jmux_i_addr_pc4_10_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[10]) );
  DFC1 u_fetch_pipe_pc4_reg_11_ ( .D(u_fetch_jmux_i_addr_pc4_11_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[11]) );
  DFC1 u_fetch_pipe_pc4_reg_12_ ( .D(u_fetch_jmux_i_addr_pc4_12_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[12]) );
  DFC1 u_fetch_pipe_pc4_reg_13_ ( .D(u_fetch_jmux_i_addr_pc4_13_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[13]) );
  DFC1 u_fetch_pipe_pc4_reg_14_ ( .D(u_fetch_jmux_i_addr_pc4_14_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[14]) );
  DFC1 u_fetch_pipe_pc4_reg_15_ ( .D(u_fetch_jmux_i_addr_pc4_15_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[15]) );
  DFC1 u_fetch_pipe_pc4_reg_16_ ( .D(u_fetch_jmux_i_addr_pc4_16_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[16]) );
  DFC1 u_fetch_pipe_pc4_reg_17_ ( .D(u_fetch_jmux_i_addr_pc4_17_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[17]) );
  DFC1 u_fetch_pipe_pc4_reg_18_ ( .D(u_fetch_jmux_i_addr_pc4_18_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[18]) );
  DFC1 u_fetch_pipe_pc4_reg_19_ ( .D(u_fetch_jmux_i_addr_pc4_19_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[19]) );
  DFC1 u_fetch_pipe_pc4_reg_20_ ( .D(u_fetch_jmux_i_addr_pc4_20_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[20]) );
  DFC1 u_fetch_pipe_pc4_reg_21_ ( .D(u_fetch_jmux_i_addr_pc4_21_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[21]) );
  DFC1 u_fetch_pipe_pc4_reg_22_ ( .D(u_fetch_jmux_i_addr_pc4_22_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[22]) );
  DFC1 u_fetch_pipe_pc4_reg_23_ ( .D(u_fetch_jmux_i_addr_pc4_23_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[23]) );
  DFC1 u_fetch_pipe_pc4_reg_24_ ( .D(u_fetch_jmux_i_addr_pc4_24_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[24]) );
  DFC1 u_fetch_pipe_pc4_reg_25_ ( .D(u_fetch_jmux_i_addr_pc4_25_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[25]) );
  DFC1 u_fetch_pipe_pc4_reg_26_ ( .D(u_fetch_jmux_i_addr_pc4_26_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[26]) );
  DFC1 u_fetch_pipe_pc4_reg_27_ ( .D(u_fetch_jmux_i_addr_pc4_27_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[27]) );
  DFC1 u_fetch_pipe_pc4_reg_28_ ( .D(u_fetch_jmux_i_addr_pc4_28_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[28]), .QN(n281) );
  DFC1 u_fetch_pipe_pc4_reg_29_ ( .D(u_fetch_jmux_i_addr_pc4_29_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[29]), .QN(n280) );
  DFC1 u_fetch_pipe_pc4_reg_30_ ( .D(u_fetch_jmux_i_addr_pc4_30_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[30]), .QN(n279) );
  DFC1 u_fetch_pipe_pc4_reg_31_ ( .D(u_fetch_jmux_i_addr_pc4_31_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[31]), .QN(n278) );
  DFC1 u_fetch_pipe_instr_reg_0_ ( .D(read_instruction[0]), .C(clk), .RN(rst_n), .Q(if_addr_j[2]), .QN(n284) );
  DFC1 u_fetch_pipe_instr_reg_3_ ( .D(read_instruction[3]), .C(clk), .RN(rst_n), .Q(if_addr_j[5]), .QN(n283) );
  DFC1 u_fetch_pipe_instr_reg_4_ ( .D(read_instruction[4]), .C(clk), .RN(rst_n), .Q(if_addr_j[6]), .QN(n282) );
  DFC1 u_fetch_pipe_instr_reg_5_ ( .D(read_instruction[5]), .C(clk), .RN(rst_n), .Q(if_addr_j[7]), .QN(n285) );
  DFC1 u_fetch_pipe_instr_reg_6_ ( .D(read_instruction[6]), .C(clk), .RN(rst_n), .Q(if_addr_j[8]), .QN(n294) );
  DFC1 u_fetch_pipe_instr_reg_7_ ( .D(read_instruction[7]), .C(clk), .RN(rst_n), .Q(if_addr_j[9]), .QN(n293) );
  DFC1 u_fetch_pipe_instr_reg_8_ ( .D(read_instruction[8]), .C(clk), .RN(rst_n), .Q(if_addr_j[10]), .QN(n292) );
  DFC1 u_fetch_pipe_instr_reg_9_ ( .D(read_instruction[9]), .C(clk), .RN(rst_n), .Q(if_addr_j[11]), .QN(n291) );
  DFC1 u_fetch_pipe_instr_reg_10_ ( .D(read_instruction[10]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[12]), .QN(n286) );
  DFC1 u_fetch_pipe_instr_reg_11_ ( .D(read_instruction[11]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[13]), .QN(n290) );
  DFC1 u_fetch_pipe_instr_reg_12_ ( .D(read_instruction[12]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[14]), .QN(n289) );
  DFC1 u_fetch_pipe_instr_reg_13_ ( .D(read_instruction[13]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[15]), .QN(n288) );
  DFC1 u_fetch_pipe_instr_reg_14_ ( .D(read_instruction[14]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[16]), .QN(n287) );
  DFC1 u_fetch_pipe_instr_reg_26_ ( .D(read_instruction[26]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[26]), .QN(n264) );
  DFC1 u_fetch_pipe_instr_reg_29_ ( .D(read_instruction[29]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[29]), .QN(n342) );
  DFC1 u_mem_pipe_data_memout_reg_0_ ( .D(read_data[0]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[0]) );
  DFC1 u_mem_pipe_data_memout_reg_1_ ( .D(read_data[1]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[1]) );
  DFC1 u_mem_pipe_data_memout_reg_2_ ( .D(read_data[2]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[2]) );
  DFC1 u_mem_pipe_data_memout_reg_3_ ( .D(read_data[3]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[3]) );
  DFC1 u_mem_pipe_data_memout_reg_4_ ( .D(read_data[4]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[4]) );
  DFC1 u_mem_pipe_data_memout_reg_5_ ( .D(read_data[5]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[5]) );
  DFC1 u_mem_pipe_data_memout_reg_6_ ( .D(read_data[6]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[6]) );
  DFC1 u_mem_pipe_data_memout_reg_7_ ( .D(read_data[7]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[7]) );
  DFC1 u_mem_pipe_data_memout_reg_8_ ( .D(read_data[8]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[8]) );
  DFC1 u_mem_pipe_data_memout_reg_9_ ( .D(read_data[9]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[9]) );
  DFC1 u_mem_pipe_data_memout_reg_10_ ( .D(read_data[10]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[10]) );
  DFC1 u_mem_pipe_data_memout_reg_11_ ( .D(read_data[11]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[11]) );
  DFC1 u_mem_pipe_data_memout_reg_12_ ( .D(read_data[12]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[12]) );
  DFC1 u_mem_pipe_data_memout_reg_13_ ( .D(read_data[13]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[13]) );
  DFC1 u_mem_pipe_data_memout_reg_14_ ( .D(read_data[14]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[14]) );
  DFC1 u_mem_pipe_data_memout_reg_15_ ( .D(read_data[15]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[15]) );
  DFC1 u_mem_pipe_data_memout_reg_16_ ( .D(read_data[16]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[16]) );
  DFC1 u_mem_pipe_data_memout_reg_17_ ( .D(read_data[17]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[17]) );
  DFC1 u_mem_pipe_data_memout_reg_18_ ( .D(read_data[18]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[18]) );
  DFC1 u_mem_pipe_data_memout_reg_19_ ( .D(read_data[19]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[19]) );
  DFC1 u_mem_pipe_data_memout_reg_20_ ( .D(read_data[20]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[20]) );
  DFC1 u_mem_pipe_data_memout_reg_21_ ( .D(read_data[21]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[21]) );
  DFC1 u_mem_pipe_data_memout_reg_22_ ( .D(read_data[22]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[22]) );
  DFC1 u_mem_pipe_data_memout_reg_23_ ( .D(read_data[23]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[23]) );
  DFC1 u_mem_pipe_data_memout_reg_24_ ( .D(read_data[24]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[24]) );
  DFC1 u_mem_pipe_data_memout_reg_25_ ( .D(read_data[25]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[25]) );
  DFC1 u_mem_pipe_data_memout_reg_26_ ( .D(read_data[26]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[26]) );
  DFC1 u_mem_pipe_data_memout_reg_27_ ( .D(read_data[27]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[27]) );
  DFC1 u_mem_pipe_data_memout_reg_28_ ( .D(read_data[28]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[28]) );
  DFC1 u_mem_pipe_data_memout_reg_29_ ( .D(read_data[29]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[29]) );
  DFC1 u_mem_pipe_data_memout_reg_30_ ( .D(read_data[30]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[30]) );
  DFC1 u_mem_pipe_data_memout_reg_31_ ( .D(read_data[31]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[31]) );
  DFC1 u_mem_pipe_rt_reg_4_ ( .D(for_addr_rtM[4]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[4]), .QN(n265) );
  DFC1 u_mem_pipe_con_FWmemread_reg ( .D(ex_con_Mmemread), .C(clk), .RN(rst_n), 
        .Q(for_FWmemread) );
  DFC1 u_mem_pipe_rt_reg_0_ ( .D(for_addr_rtM[0]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[0]) );
  DFC1 u_mem_pipe_rt_reg_1_ ( .D(for_addr_rtM[1]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[1]) );
  DFC1 u_mem_pipe_rt_reg_2_ ( .D(for_addr_rtM[2]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[2]) );
  DFC1 u_mem_pipe_rt_reg_3_ ( .D(for_addr_rtM[3]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[3]) );
  DFC1 u_mem_pipe_con_Wregwrite_reg ( .D(mem_con_Wregwrite), .C(clk), .RN(
        rst_n), .Q(id_con_Wregwrite) );
  DFC1 u_mem_pipe_addr_regdst_reg_0_ ( .D(mem_addr_regdst[0]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[0]) );
  DFC1 u_mem_pipe_addr_regdst_reg_1_ ( .D(mem_addr_regdst[1]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[1]) );
  DFC1 u_mem_pipe_addr_regdst_reg_2_ ( .D(mem_addr_regdst[2]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[2]) );
  DFC1 u_mem_pipe_addr_regdst_reg_3_ ( .D(mem_addr_regdst[3]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[3]) );
  DFC1 u_mem_pipe_addr_regdst_reg_4_ ( .D(mem_addr_regdst[4]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[4]) );
  DFC1 u_mem_pipe_data_alures_reg_0_ ( .D(u_mem_resmux_o_data_alu[0]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[0]) );
  DFC1 u_mem_pipe_data_alures_reg_1_ ( .D(u_mem_resmux_o_data_alu[1]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[1]) );
  DFC1 u_mem_pipe_data_alures_reg_2_ ( .D(u_mem_resmux_o_data_alu[2]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[2]) );
  DFC1 u_mem_pipe_data_alures_reg_3_ ( .D(u_mem_resmux_o_data_alu[3]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[3]) );
  DFC1 u_mem_pipe_data_alures_reg_4_ ( .D(u_mem_resmux_o_data_alu[4]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[4]) );
  DFC1 u_mem_pipe_data_alures_reg_5_ ( .D(u_mem_resmux_o_data_alu[5]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[5]) );
  DFC1 u_mem_pipe_data_alures_reg_6_ ( .D(u_mem_resmux_o_data_alu[6]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[6]) );
  DFC1 u_mem_pipe_data_alures_reg_7_ ( .D(u_mem_resmux_o_data_alu[7]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[7]) );
  DFC1 u_mem_pipe_data_alures_reg_8_ ( .D(u_mem_resmux_o_data_alu[8]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[8]) );
  DFC1 u_mem_pipe_data_alures_reg_9_ ( .D(u_mem_resmux_o_data_alu[9]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[9]) );
  DFC1 u_mem_pipe_data_alures_reg_10_ ( .D(u_mem_resmux_o_data_alu[10]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[10]) );
  DFC1 u_mem_pipe_data_alures_reg_11_ ( .D(u_mem_resmux_o_data_alu[11]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[11]) );
  DFC1 u_mem_pipe_data_alures_reg_12_ ( .D(u_mem_resmux_o_data_alu[12]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[12]) );
  DFC1 u_mem_pipe_data_alures_reg_13_ ( .D(u_mem_resmux_o_data_alu[13]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[13]) );
  DFC1 u_mem_pipe_data_alures_reg_14_ ( .D(u_mem_resmux_o_data_alu[14]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[14]) );
  DFC1 u_mem_pipe_data_alures_reg_15_ ( .D(u_mem_resmux_o_data_alu[15]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[15]) );
  DFC1 u_mem_pipe_data_alures_reg_16_ ( .D(u_mem_resmux_o_data_alu[16]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[16]) );
  DFC1 u_mem_pipe_data_alures_reg_17_ ( .D(u_mem_resmux_o_data_alu[17]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[17]) );
  DFC1 u_mem_pipe_data_alures_reg_18_ ( .D(u_mem_resmux_o_data_alu[18]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[18]) );
  DFC1 u_mem_pipe_data_alures_reg_19_ ( .D(u_mem_resmux_o_data_alu[19]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[19]) );
  DFC1 u_mem_pipe_data_alures_reg_20_ ( .D(u_mem_resmux_o_data_alu[20]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[20]) );
  DFC1 u_mem_pipe_data_alures_reg_21_ ( .D(u_mem_resmux_o_data_alu[21]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[21]) );
  DFC1 u_mem_pipe_data_alures_reg_22_ ( .D(u_mem_resmux_o_data_alu[22]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[22]) );
  DFC1 u_mem_pipe_data_alures_reg_23_ ( .D(u_mem_resmux_o_data_alu[23]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[23]) );
  DFC1 u_mem_pipe_data_alures_reg_24_ ( .D(u_mem_resmux_o_data_alu[24]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[24]) );
  DFC1 u_mem_pipe_data_alures_reg_25_ ( .D(u_mem_resmux_o_data_alu[25]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[25]) );
  DFC1 u_mem_pipe_data_alures_reg_26_ ( .D(u_mem_resmux_o_data_alu[26]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[26]) );
  DFC1 u_mem_pipe_data_alures_reg_27_ ( .D(u_mem_resmux_o_data_alu[27]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[27]) );
  DFC1 u_mem_pipe_data_alures_reg_28_ ( .D(u_mem_resmux_o_data_alu[28]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[28]) );
  DFC1 u_mem_pipe_data_alures_reg_29_ ( .D(u_mem_resmux_o_data_alu[29]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[29]) );
  DFC1 u_mem_pipe_data_alures_reg_30_ ( .D(u_mem_resmux_o_data_alu[30]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[30]) );
  DFC1 u_mem_pipe_data_alures_reg_31_ ( .D(u_mem_resmux_o_data_alu[31]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[31]) );
  DFC1 u_fetch_u_pc_program_counter_reg_0_ ( .D(n137), .C(clk), .RN(rst_n), 
        .Q(instruction_address[0]), .QN(n328) );
  DFC1 u_fetch_u_pc_program_counter_reg_1_ ( .D(n136), .C(clk), .RN(rst_n), 
        .Q(instruction_address[1]) );
  DFC1 u_fetch_u_pc_program_counter_reg_2_ ( .D(n135), .C(clk), .RN(rst_n), 
        .Q(instruction_address[2]), .QN(n276) );
  DFC1 u_fetch_u_pc_program_counter_reg_3_ ( .D(n134), .C(clk), .RN(rst_n), 
        .Q(instruction_address[3]), .QN(n318) );
  DFC1 u_fetch_u_pc_program_counter_reg_4_ ( .D(n133), .C(clk), .RN(rst_n), 
        .Q(instruction_address[4]), .QN(n275) );
  DFC1 u_fetch_u_pc_program_counter_reg_5_ ( .D(n132), .C(clk), .RN(rst_n), 
        .Q(instruction_address[5]), .QN(n307) );
  DFC1 u_fetch_u_pc_program_counter_reg_6_ ( .D(n131), .C(clk), .RN(rst_n), 
        .Q(instruction_address[6]), .QN(n317) );
  DFC1 u_fetch_u_pc_program_counter_reg_7_ ( .D(n130), .C(clk), .RN(rst_n), 
        .Q(instruction_address[7]), .QN(n306) );
  DFC1 u_fetch_u_pc_program_counter_reg_8_ ( .D(n129), .C(clk), .RN(rst_n), 
        .Q(instruction_address[8]), .QN(n274) );
  DFC1 u_fetch_u_pc_program_counter_reg_9_ ( .D(n128), .C(clk), .RN(rst_n), 
        .Q(instruction_address[9]), .QN(n305) );
  DFC1 u_fetch_u_pc_program_counter_reg_10_ ( .D(n127), .C(clk), .RN(rst_n), 
        .Q(instruction_address[10]), .QN(n273) );
  DFC1 u_fetch_u_pc_program_counter_reg_11_ ( .D(n126), .C(clk), .RN(rst_n), 
        .Q(instruction_address[11]), .QN(n304) );
  DFC1 u_fetch_u_pc_program_counter_reg_12_ ( .D(n125), .C(clk), .RN(rst_n), 
        .Q(instruction_address[12]), .QN(n316) );
  DFC1 u_fetch_u_pc_program_counter_reg_13_ ( .D(n124), .C(clk), .RN(rst_n), 
        .Q(instruction_address[13]), .QN(n303) );
  DFC1 u_fetch_u_pc_program_counter_reg_14_ ( .D(n123), .C(clk), .RN(rst_n), 
        .Q(instruction_address[14]), .QN(n315) );
  DFC1 u_fetch_u_pc_program_counter_reg_15_ ( .D(n122), .C(clk), .RN(rst_n), 
        .Q(instruction_address[15]), .QN(n302) );
  DFC1 u_fetch_u_pc_program_counter_reg_16_ ( .D(n121), .C(clk), .RN(rst_n), 
        .Q(instruction_address[16]), .QN(n314) );
  DFC1 u_fetch_u_pc_program_counter_reg_17_ ( .D(n120), .C(clk), .RN(rst_n), 
        .Q(instruction_address[17]), .QN(n301) );
  DFC1 u_fetch_u_pc_program_counter_reg_18_ ( .D(n119), .C(clk), .RN(rst_n), 
        .Q(instruction_address[18]), .QN(n313) );
  DFC1 u_fetch_u_pc_program_counter_reg_19_ ( .D(n118), .C(clk), .RN(rst_n), 
        .Q(instruction_address[19]), .QN(n300) );
  DFC1 u_fetch_u_pc_program_counter_reg_20_ ( .D(n117), .C(clk), .RN(rst_n), 
        .Q(instruction_address[20]), .QN(n272) );
  DFC1 u_fetch_u_pc_program_counter_reg_21_ ( .D(n116), .C(clk), .RN(rst_n), 
        .Q(instruction_address[21]), .QN(n299) );
  DFC1 u_fetch_u_pc_program_counter_reg_22_ ( .D(n115), .C(clk), .RN(rst_n), 
        .Q(instruction_address[22]), .QN(n312) );
  DFC1 u_fetch_u_pc_program_counter_reg_23_ ( .D(n114), .C(clk), .RN(rst_n), 
        .Q(instruction_address[23]), .QN(n298) );
  DFC1 u_fetch_u_pc_program_counter_reg_24_ ( .D(n113), .C(clk), .RN(rst_n), 
        .Q(instruction_address[24]), .QN(n311) );
  DFC1 u_fetch_u_pc_program_counter_reg_25_ ( .D(n112), .C(clk), .RN(rst_n), 
        .Q(instruction_address[25]), .QN(n297) );
  DFC1 u_fetch_u_pc_program_counter_reg_26_ ( .D(n111), .C(clk), .RN(rst_n), 
        .Q(instruction_address[26]), .QN(n271) );
  DFC1 u_fetch_u_pc_program_counter_reg_27_ ( .D(n110), .C(clk), .RN(rst_n), 
        .Q(instruction_address[27]), .QN(n296) );
  DFC1 u_fetch_u_pc_program_counter_reg_28_ ( .D(n109), .C(clk), .RN(rst_n), 
        .Q(instruction_address[28]), .QN(n324) );
  DFC1 u_fetch_u_pc_program_counter_reg_29_ ( .D(n108), .C(clk), .RN(rst_n), 
        .Q(instruction_address[29]), .QN(n295) );
  DFC1 u_fetch_u_pc_program_counter_reg_30_ ( .D(n107), .C(clk), .RN(rst_n), 
        .Q(instruction_address[30]), .QN(n322) );
  DFC1 u_fetch_u_pc_program_counter_reg_31_ ( .D(n138), .C(clk), .RN(rst_n), 
        .Q(instruction_address[31]), .QN(n319) );
  DFC1 u_decode_pipe_addr_branch_reg_0_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[0]), .C(clk), .RN(rst_n), .Q(
        ex_data_pc4[0]) );
  DFC1 u_decode_pipe_addr_branch_reg_1_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[1]), .C(clk), .RN(rst_n), .Q(
        ex_data_pc4[1]) );
  DFC1 u_decode_pipe_addr_branch_reg_2_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[2]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[2]) );
  DFC1 u_decode_pipe_addr_branch_reg_3_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[3]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[3]) );
  DFC1 u_decode_pipe_addr_branch_reg_4_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[4]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[4]) );
  DFC1 u_decode_pipe_addr_branch_reg_5_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[5]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[5]) );
  DFC1 u_decode_pipe_addr_branch_reg_6_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[6]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[6]) );
  DFC1 u_decode_pipe_addr_branch_reg_7_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[7]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[7]) );
  DFC1 u_decode_pipe_addr_branch_reg_8_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[8]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[8]) );
  DFC1 u_decode_pipe_addr_branch_reg_9_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[9]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[9]) );
  DFC1 u_decode_pipe_addr_branch_reg_10_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[10]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[10]) );
  DFC1 u_decode_pipe_addr_branch_reg_11_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[11]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[11]) );
  DFC1 u_decode_pipe_addr_branch_reg_12_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[12]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[12]) );
  DFC1 u_decode_pipe_addr_branch_reg_13_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[13]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[13]) );
  DFC1 u_decode_pipe_addr_branch_reg_14_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[14]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[14]) );
  DFC1 u_decode_pipe_addr_branch_reg_15_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[15]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[15]) );
  DFC1 u_decode_pipe_addr_branch_reg_16_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[16]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[16]) );
  DFC1 u_decode_pipe_addr_branch_reg_17_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[17]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[17]) );
  DFC1 u_decode_pipe_addr_branch_reg_18_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[18]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[18]) );
  DFC1 u_decode_pipe_addr_branch_reg_19_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[19]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[19]) );
  DFC1 u_decode_pipe_addr_branch_reg_20_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[20]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[20]) );
  DFC1 u_decode_pipe_addr_branch_reg_21_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[21]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[21]) );
  DFC1 u_decode_pipe_addr_branch_reg_22_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[22]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[22]) );
  DFC1 u_decode_pipe_addr_branch_reg_23_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[23]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[23]) );
  DFC1 u_decode_pipe_addr_branch_reg_24_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[24]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[24]) );
  DFC1 u_decode_pipe_addr_branch_reg_25_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[25]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[25]) );
  DFC1 u_decode_pipe_addr_branch_reg_26_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[26]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[26]) );
  DFC1 u_decode_pipe_addr_branch_reg_27_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[27]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[27]) );
  DFC1 u_decode_pipe_addr_branch_reg_28_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[28]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[28]) );
  DFC1 u_decode_pipe_addr_branch_reg_29_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[29]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[29]) );
  DFC1 u_decode_pipe_addr_branch_reg_30_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[30]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[30]) );
  DFC1 u_decode_pipe_addr_branch_reg_31_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[31]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[31]) );
  DFC1 u_decode_pipe_FWmemout_reg_0_ ( .D(wb_data_memout[0]), .C(clk), .RN(
        rst_n), .Q(for_memout[0]) );
  DFC1 u_decode_pipe_FWmemout_reg_1_ ( .D(wb_data_memout[1]), .C(clk), .RN(
        rst_n), .Q(for_memout[1]) );
  DFC1 u_decode_pipe_FWmemout_reg_2_ ( .D(wb_data_memout[2]), .C(clk), .RN(
        rst_n), .Q(for_memout[2]) );
  DFC1 u_decode_pipe_FWmemout_reg_3_ ( .D(wb_data_memout[3]), .C(clk), .RN(
        rst_n), .Q(for_memout[3]) );
  DFC1 u_decode_pipe_FWmemout_reg_4_ ( .D(wb_data_memout[4]), .C(clk), .RN(
        rst_n), .Q(for_memout[4]) );
  DFC1 u_decode_pipe_FWmemout_reg_5_ ( .D(wb_data_memout[5]), .C(clk), .RN(
        rst_n), .Q(for_memout[5]) );
  DFC1 u_decode_pipe_FWmemout_reg_6_ ( .D(wb_data_memout[6]), .C(clk), .RN(
        rst_n), .Q(for_memout[6]) );
  DFC1 u_decode_pipe_FWmemout_reg_7_ ( .D(wb_data_memout[7]), .C(clk), .RN(
        rst_n), .Q(for_memout[7]) );
  DFC1 u_decode_pipe_FWmemout_reg_8_ ( .D(wb_data_memout[8]), .C(clk), .RN(
        rst_n), .Q(for_memout[8]) );
  DFC1 u_decode_pipe_FWmemout_reg_9_ ( .D(wb_data_memout[9]), .C(clk), .RN(
        rst_n), .Q(for_memout[9]) );
  DFC1 u_decode_pipe_FWmemout_reg_10_ ( .D(wb_data_memout[10]), .C(clk), .RN(
        rst_n), .Q(for_memout[10]) );
  DFC1 u_decode_pipe_FWmemout_reg_11_ ( .D(wb_data_memout[11]), .C(clk), .RN(
        rst_n), .Q(for_memout[11]) );
  DFC1 u_decode_pipe_FWmemout_reg_12_ ( .D(wb_data_memout[12]), .C(clk), .RN(
        rst_n), .Q(for_memout[12]) );
  DFC1 u_decode_pipe_FWmemout_reg_13_ ( .D(wb_data_memout[13]), .C(clk), .RN(
        rst_n), .Q(for_memout[13]) );
  DFC1 u_decode_pipe_FWmemout_reg_14_ ( .D(wb_data_memout[14]), .C(clk), .RN(
        rst_n), .Q(for_memout[14]) );
  DFC1 u_decode_pipe_FWmemout_reg_15_ ( .D(wb_data_memout[15]), .C(clk), .RN(
        rst_n), .Q(for_memout[15]) );
  DFC1 u_decode_pipe_FWmemout_reg_16_ ( .D(wb_data_memout[16]), .C(clk), .RN(
        rst_n), .Q(for_memout[16]) );
  DFC1 u_decode_pipe_FWmemout_reg_17_ ( .D(wb_data_memout[17]), .C(clk), .RN(
        rst_n), .Q(for_memout[17]) );
  DFC1 u_decode_pipe_FWmemout_reg_18_ ( .D(wb_data_memout[18]), .C(clk), .RN(
        rst_n), .Q(for_memout[18]) );
  DFC1 u_decode_pipe_FWmemout_reg_19_ ( .D(wb_data_memout[19]), .C(clk), .RN(
        rst_n), .Q(for_memout[19]) );
  DFC1 u_decode_pipe_FWmemout_reg_20_ ( .D(wb_data_memout[20]), .C(clk), .RN(
        rst_n), .Q(for_memout[20]) );
  DFC1 u_decode_pipe_FWmemout_reg_21_ ( .D(wb_data_memout[21]), .C(clk), .RN(
        rst_n), .Q(for_memout[21]) );
  DFC1 u_decode_pipe_FWmemout_reg_22_ ( .D(wb_data_memout[22]), .C(clk), .RN(
        rst_n), .Q(for_memout[22]) );
  DFC1 u_decode_pipe_FWmemout_reg_23_ ( .D(wb_data_memout[23]), .C(clk), .RN(
        rst_n), .Q(for_memout[23]) );
  DFC1 u_decode_pipe_FWmemout_reg_24_ ( .D(wb_data_memout[24]), .C(clk), .RN(
        rst_n), .Q(for_memout[24]) );
  DFC1 u_decode_pipe_FWmemout_reg_25_ ( .D(wb_data_memout[25]), .C(clk), .RN(
        rst_n), .Q(for_memout[25]) );
  DFC1 u_decode_pipe_FWmemout_reg_26_ ( .D(wb_data_memout[26]), .C(clk), .RN(
        rst_n), .Q(for_memout[26]) );
  DFC1 u_decode_pipe_FWmemout_reg_28_ ( .D(wb_data_memout[28]), .C(clk), .RN(
        rst_n), .Q(for_memout[28]) );
  DFC1 u_decode_pipe_FWmemout_reg_29_ ( .D(wb_data_memout[29]), .C(clk), .RN(
        rst_n), .Q(for_memout[29]) );
  DFC1 u_decode_pipe_FWmemout_reg_30_ ( .D(wb_data_memout[30]), .C(clk), .RN(
        rst_n), .Q(for_memout[30]) );
  DFC1 u_decode_pipe_FWmemout_reg_31_ ( .D(wb_data_memout[31]), .C(clk), .RN(
        rst_n), .Q(for_memout[31]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_11_ ( .D(if_addr_j[13]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[0]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_12_ ( .D(if_addr_j[14]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[1]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_13_ ( .D(if_addr_j[15]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[2]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_14_ ( .D(if_addr_j[16]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[3]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_15_ ( .D(if_addr_j[17]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[4]) );
  DFC1 u_decode_pipe_con_Wregwrite_reg ( .D(u_decode_control_o_con_regwrite), 
        .C(clk), .RN(rst_n), .Q(ex_con_Wregwrite) );
  DFC1 u_decode_pipe_con_Wmemtoreg_reg ( .D(n512), .C(clk), .RN(rst_n), .Q(
        ex_con_Wmemtoreg) );
  DFC1 u_decode_pipe_con_Mmemwrite_reg ( .D(u_decode_control_o_con_memwrite), 
        .C(clk), .RN(rst_n), .Q(ex_con_Mmemwrite) );
  DFC1 u_decode_pipe_con_Mmemread_reg ( .D(u_decode_control_o_con_memread), 
        .C(clk), .RN(rst_n), .Q(ex_con_Mmemread) );
  DFC1 u_decode_pipe_con_MaluPC4_reg ( .D(u_decode_jbcon_o_con_aluPC4), .C(clk), .RN(rst_n), .Q(ex_con_Malupc8) );
  DFC1 u_decode_pipe_con_Eregdst_reg ( .D(u_decode_control_o_con_regdst), .C(
        clk), .RN(rst_n), .Q(ex_con_Eregdst) );
  DFC1 u_decode_pipe_con_Ealuop_reg_0_ ( .D(u_decode_control_o_con_aluop_0_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[0]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_2_ ( .D(u_decode_control_o_con_aluop_2_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[2]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_5_ ( .D(u_decode_control_o_con_aluop_5_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[5]) );
  DFC1 u_decode_pipe_addr_pc4_reg_2_ ( .D(id_addr_pc4[2]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[2]) );
  DFC1 u_decode_pipe_addr_pc4_reg_3_ ( .D(id_addr_pc4[3]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[3]) );
  DFC1 u_decode_pipe_addr_pc4_reg_4_ ( .D(id_addr_pc4[4]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[4]) );
  DFC1 u_decode_pipe_addr_pc4_reg_5_ ( .D(id_addr_pc4[5]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[5]) );
  DFC1 u_decode_pipe_addr_pc4_reg_6_ ( .D(id_addr_pc4[6]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[6]) );
  DFC1 u_decode_pipe_addr_pc4_reg_7_ ( .D(id_addr_pc4[7]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[7]) );
  DFC1 u_decode_pipe_addr_pc4_reg_8_ ( .D(id_addr_pc4[8]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[8]) );
  DFC1 u_decode_pipe_addr_pc4_reg_9_ ( .D(id_addr_pc4[9]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[9]) );
  DFC1 u_decode_pipe_addr_pc4_reg_10_ ( .D(id_addr_pc4[10]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[10]) );
  DFC1 u_decode_pipe_addr_pc4_reg_11_ ( .D(id_addr_pc4[11]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[11]) );
  DFC1 u_decode_pipe_addr_pc4_reg_12_ ( .D(id_addr_pc4[12]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[12]) );
  DFC1 u_decode_pipe_addr_pc4_reg_13_ ( .D(id_addr_pc4[13]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[13]) );
  DFC1 u_decode_pipe_addr_pc4_reg_14_ ( .D(id_addr_pc4[14]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[14]) );
  DFC1 u_decode_pipe_addr_pc4_reg_15_ ( .D(id_addr_pc4[15]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[15]) );
  DFC1 u_decode_pipe_addr_pc4_reg_16_ ( .D(id_addr_pc4[16]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[16]) );
  DFC1 u_decode_pipe_addr_pc4_reg_17_ ( .D(id_addr_pc4[17]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[17]) );
  DFC1 u_decode_pipe_addr_pc4_reg_18_ ( .D(id_addr_pc4[18]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[18]) );
  DFC1 u_decode_pipe_addr_pc4_reg_19_ ( .D(id_addr_pc4[19]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[19]) );
  DFC1 u_decode_pipe_addr_pc4_reg_20_ ( .D(id_addr_pc4[20]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[20]) );
  DFC1 u_decode_pipe_addr_pc4_reg_21_ ( .D(id_addr_pc4[21]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[21]) );
  DFC1 u_decode_pipe_addr_pc4_reg_22_ ( .D(id_addr_pc4[22]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[22]) );
  DFC1 u_decode_pipe_addr_pc4_reg_23_ ( .D(id_addr_pc4[23]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[23]) );
  DFC1 u_decode_pipe_addr_pc4_reg_24_ ( .D(id_addr_pc4[24]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[24]) );
  DFC1 u_decode_pipe_addr_pc4_reg_25_ ( .D(id_addr_pc4[25]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[25]) );
  DFC1 u_decode_pipe_addr_pc4_reg_26_ ( .D(id_addr_pc4[26]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[26]) );
  DFC1 u_decode_pipe_addr_pc4_reg_27_ ( .D(id_addr_pc4[27]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[27]) );
  DFC1 u_decode_pipe_addr_pc4_reg_28_ ( .D(if_addr_j[28]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[28]) );
  DFC1 u_decode_pipe_addr_pc4_reg_29_ ( .D(if_addr_j[29]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[29]) );
  DFC1 u_decode_pipe_addr_pc4_reg_30_ ( .D(if_addr_j[30]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[30]) );
  DFC1 u_decode_pipe_addr_pc4_reg_31_ ( .D(if_addr_j[31]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[31]) );
  DFC1 u_decode_pipe_addr_rt_reg_0_ ( .D(if_addr_j[18]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[0]) );
  DFC1 u_decode_pipe_addr_rt_reg_1_ ( .D(if_addr_j[19]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[1]) );
  DFC1 u_decode_pipe_addr_rt_reg_2_ ( .D(if_addr_j[20]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[2]) );
  DFC1 u_decode_pipe_addr_rt_reg_3_ ( .D(if_addr_j[21]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[3]) );
  DFC1 u_decode_pipe_addr_rt_reg_4_ ( .D(if_addr_j[22]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[4]) );
  DFC1 u_decode_pipe_data_rt_reg_0_ ( .D(u_decode_regbank_o_data_Rt[0]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[0]) );
  DFC1 u_decode_pipe_data_rt_reg_1_ ( .D(u_decode_regbank_o_data_Rt[1]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[1]) );
  DFC1 u_decode_pipe_data_rt_reg_2_ ( .D(u_decode_regbank_o_data_Rt[2]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[2]) );
  DFC1 u_decode_pipe_data_rt_reg_3_ ( .D(u_decode_regbank_o_data_Rt[3]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[3]) );
  DFC1 u_decode_pipe_data_rt_reg_4_ ( .D(u_decode_regbank_o_data_Rt[4]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[4]) );
  DFC1 u_decode_pipe_data_rt_reg_5_ ( .D(u_decode_regbank_o_data_Rt[5]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[5]) );
  DFC1 u_decode_pipe_data_rt_reg_6_ ( .D(u_decode_regbank_o_data_Rt[6]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[6]) );
  DFC1 u_decode_pipe_data_rt_reg_7_ ( .D(u_decode_regbank_o_data_Rt[7]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[7]) );
  DFC1 u_decode_pipe_data_rt_reg_8_ ( .D(u_decode_regbank_o_data_Rt[8]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[8]) );
  DFC1 u_decode_pipe_data_rt_reg_9_ ( .D(u_decode_regbank_o_data_Rt[9]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[9]) );
  DFC1 u_decode_pipe_data_rt_reg_10_ ( .D(u_decode_regbank_o_data_Rt[10]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[10]) );
  DFC1 u_decode_pipe_data_rt_reg_11_ ( .D(u_decode_regbank_o_data_Rt[11]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[11]) );
  DFC1 u_decode_pipe_data_rt_reg_12_ ( .D(u_decode_regbank_o_data_Rt[12]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[12]) );
  DFC1 u_decode_pipe_data_rt_reg_13_ ( .D(u_decode_regbank_o_data_Rt[13]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[13]) );
  DFC1 u_decode_pipe_data_rt_reg_14_ ( .D(u_decode_regbank_o_data_Rt[14]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[14]) );
  DFC1 u_decode_pipe_data_rt_reg_15_ ( .D(u_decode_regbank_o_data_Rt[15]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[15]) );
  DFC1 u_decode_pipe_data_rt_reg_16_ ( .D(u_decode_regbank_o_data_Rt[16]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[16]) );
  DFC1 u_decode_pipe_data_rt_reg_17_ ( .D(u_decode_regbank_o_data_Rt[17]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[17]) );
  DFC1 u_decode_pipe_data_rt_reg_18_ ( .D(u_decode_regbank_o_data_Rt[18]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[18]) );
  DFC1 u_decode_pipe_data_rt_reg_19_ ( .D(u_decode_regbank_o_data_Rt[19]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[19]) );
  DFC1 u_decode_pipe_data_rt_reg_20_ ( .D(u_decode_regbank_o_data_Rt[20]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[20]) );
  DFC1 u_decode_pipe_data_rt_reg_21_ ( .D(u_decode_regbank_o_data_Rt[21]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[21]) );
  DFC1 u_decode_pipe_data_rt_reg_22_ ( .D(u_decode_regbank_o_data_Rt[22]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[22]) );
  DFC1 u_decode_pipe_data_rt_reg_23_ ( .D(u_decode_regbank_o_data_Rt[23]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[23]) );
  DFC1 u_decode_pipe_data_rt_reg_24_ ( .D(u_decode_regbank_o_data_Rt[24]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[24]) );
  DFC1 u_decode_pipe_data_rt_reg_25_ ( .D(u_decode_regbank_o_data_Rt[25]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[25]) );
  DFC1 u_decode_pipe_data_rt_reg_26_ ( .D(u_decode_regbank_o_data_Rt[26]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[26]) );
  DFC1 u_decode_pipe_data_rt_reg_27_ ( .D(u_decode_regbank_o_data_Rt[27]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[27]) );
  DFC1 u_decode_pipe_data_rt_reg_28_ ( .D(u_decode_regbank_o_data_Rt[28]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[28]) );
  DFC1 u_decode_pipe_data_rt_reg_29_ ( .D(u_decode_regbank_o_data_Rt[29]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[29]) );
  DFC1 u_decode_pipe_data_rt_reg_30_ ( .D(u_decode_regbank_o_data_Rt[30]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[30]) );
  DFC1 u_decode_pipe_data_rt_reg_31_ ( .D(u_decode_regbank_o_data_Rt[31]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[31]) );
  DFC1 u_decode_pipe_data_rs_reg_0_ ( .D(id_data_jr[0]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[0]) );
  DFC1 u_decode_pipe_data_rs_reg_1_ ( .D(id_data_jr[1]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[1]) );
  DFC1 u_decode_pipe_data_rs_reg_2_ ( .D(id_data_jr[2]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[2]) );
  DFC1 u_decode_pipe_data_rs_reg_3_ ( .D(id_data_jr[3]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[3]) );
  DFC1 u_decode_pipe_data_rs_reg_4_ ( .D(id_data_jr[4]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[4]) );
  DFC1 u_decode_pipe_data_rs_reg_5_ ( .D(id_data_jr[5]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[5]) );
  DFC1 u_decode_pipe_data_rs_reg_6_ ( .D(id_data_jr[6]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[6]) );
  DFC1 u_decode_pipe_data_rs_reg_7_ ( .D(id_data_jr[7]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[7]) );
  DFC1 u_decode_pipe_data_rs_reg_8_ ( .D(id_data_jr[8]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[8]) );
  DFC1 u_decode_pipe_data_rs_reg_9_ ( .D(id_data_jr[9]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[9]) );
  DFC1 u_decode_pipe_data_rs_reg_10_ ( .D(id_data_jr[10]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[10]) );
  DFC1 u_decode_pipe_data_rs_reg_11_ ( .D(id_data_jr[11]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[11]) );
  DFC1 u_decode_pipe_data_rs_reg_12_ ( .D(id_data_jr[12]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[12]) );
  DFC1 u_decode_pipe_data_rs_reg_13_ ( .D(id_data_jr[13]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[13]) );
  DFC1 u_decode_pipe_data_rs_reg_14_ ( .D(id_data_jr[14]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[14]) );
  DFC1 u_decode_pipe_data_rs_reg_15_ ( .D(id_data_jr[15]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[15]) );
  DFC1 u_decode_pipe_data_rs_reg_16_ ( .D(id_data_jr[16]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[16]) );
  DFC1 u_decode_pipe_data_rs_reg_17_ ( .D(id_data_jr[17]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[17]) );
  DFC1 u_decode_pipe_data_rs_reg_18_ ( .D(id_data_jr[18]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[18]) );
  DFC1 u_decode_pipe_data_rs_reg_19_ ( .D(id_data_jr[19]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[19]) );
  DFC1 u_decode_pipe_data_rs_reg_20_ ( .D(id_data_jr[20]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[20]) );
  DFC1 u_decode_pipe_data_rs_reg_21_ ( .D(id_data_jr[21]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[21]) );
  DFC1 u_decode_pipe_data_rs_reg_22_ ( .D(id_data_jr[22]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[22]) );
  DFC1 u_decode_pipe_data_rs_reg_23_ ( .D(id_data_jr[23]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[23]) );
  DFC1 u_decode_pipe_data_rs_reg_24_ ( .D(id_data_jr[24]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[24]) );
  DFC1 u_decode_pipe_data_rs_reg_25_ ( .D(id_data_jr[25]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[25]) );
  DFC1 u_decode_pipe_data_rs_reg_26_ ( .D(id_data_jr[26]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[26]) );
  DFC1 u_decode_pipe_data_rs_reg_27_ ( .D(id_data_jr[27]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[27]) );
  DFC1 u_decode_pipe_data_rs_reg_28_ ( .D(id_data_jr[28]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[28]) );
  DFC1 u_decode_pipe_data_rs_reg_29_ ( .D(id_data_jr[29]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[29]) );
  DFC1 u_decode_pipe_data_rs_reg_30_ ( .D(id_data_jr[30]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[30]) );
  DFC1 u_decode_pipe_data_rs_reg_31_ ( .D(id_data_jr[31]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[31]) );
  DFC1 u_decode_pipe_bop_reg_0_ ( .D(u_decode_jbcon_o_con_bop[0]), .C(clk), 
        .RN(rst_n), .Q(ex_con_bop[0]) );
  DFC1 u_decode_pipe_bop_reg_1_ ( .D(u_decode_jbcon_o_con_bop[1]), .C(clk), 
        .RN(rst_n), .Q(ex_con_bop[1]) );
  DFC1 u_decode_pipe_bop_reg_2_ ( .D(u_decode_n6), .C(clk), .RN(rst_n), .Q(
        ex_con_bop[2]) );
  D_register_bank u_decode_u_regbank ( .i_clk(clk), .i_rst_n(rst_n), 
        .i_addr_Rs(if_addr_j[27:23]), .i_con_RegWr(id_con_Wregwrite), 
        .i_addr_Rd(id_addr_Wregwrite), .i_data_Rd(id_data_Wregwrite), 
        .o_data_Rs(id_data_jr), .o_data_Rt(u_decode_regbank_o_data_Rt), 
        .i_addr_Rt_4_(if_addr_j[22]), .i_addr_Rt_3_(if_addr_j[21]), 
        .i_addr_Rt_2_(if_addr_j[20]), .i_addr_Rt_1_(if_addr_j[19]), 
        .i_addr_Rt_0_(if_addr_j[18]) );
  OAI212 u_decode_add_x_16_U193 ( .A(u_decode_add_x_16_n157), .B(
        u_decode_add_x_16_n177), .C(u_decode_add_x_16_n158), .Q(
        u_decode_add_x_16_n156) );
  DFC3 u_fetch_pipe_instr_reg_16_ ( .D(read_instruction[16]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[18]), .QN(n251) );
  DFC3 u_fetch_pipe_instr_reg_17_ ( .D(read_instruction[17]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[19]), .QN(n329) );
  DFC3 u_fetch_pipe_instr_reg_18_ ( .D(read_instruction[18]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[20]), .QN(n330) );
  DFC3 u_fetch_pipe_instr_reg_19_ ( .D(read_instruction[19]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[21]), .QN(n325) );
  DFC3 u_fetch_pipe_instr_reg_28_ ( .D(read_instruction[28]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[28]), .QN(n270) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_16_ ( .D(u_decode_n1), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[31]) );
  DFC3 u_fetch_pipe_instr_reg_21_ ( .D(read_instruction[21]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[23]), .QN(n309) );
  DFC3 u_fetch_pipe_instr_reg_22_ ( .D(read_instruction[22]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[24]), .QN(n321) );
  DFC3 u_decode_pipe_con_Efbmux_reg_1_ ( .D(u_decode_for_o_con_fb[1]), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[1]) );
  DFC3 u_decode_pipe_con_Efbmux_reg_2_ ( .D(u_decode_for_o_con_fb[2]), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[2]) );
  DFC3 u_decode_pipe_con_Efbmux_reg_0_ ( .D(u_decode_for_o_con_fb[0]), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[0]) );
  DFC3 u_decode_pipe_con_Efamux_reg_2_ ( .D(u_decode_for_o_con_fa_2_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[2]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_10_ ( .D(if_addr_j[12]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[10]) );
  DFC3 u_fetch_pipe_instr_reg_23_ ( .D(read_instruction[23]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[25]), .QN(n323) );
  DFC3 u_decode_pipe_con_Efamux_reg_1_ ( .D(u_decode_for_o_con_fa_1_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[1]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_1_ ( .D(if_addr_j[3]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[1]) );
  DFC3 u_fetch_pipe_instr_reg_1_ ( .D(read_instruction[1]), .C(clk), .RN(rst_n), .Q(if_addr_j[3]), .QN(n327) );
  DFC3 u_decode_pipe_con_Efamux_reg_0_ ( .D(u_decode_for_o_con_fa_0_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[0]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_5_ ( .D(if_addr_j[7]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[5]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_3_ ( .D(if_addr_j[5]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[3]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_2_ ( .D(if_addr_j[4]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[2]) );
  DFC3 u_fetch_pipe_instr_reg_2_ ( .D(read_instruction[2]), .C(clk), .RN(rst_n), .Q(if_addr_j[4]), .QN(n326) );
  DFC3 u_decode_pipe_con_Ealusrc_reg ( .D(u_decode_control_o_con_alusrc), .C(
        clk), .RN(rst_n), .Q(ex_con_Ealusrc) );
  DFC3 u_fetch_pipe_instr_reg_24_ ( .D(read_instruction[24]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[26]), .QN(n320) );
  DFC3 u_fetch_pipe_instr_reg_25_ ( .D(read_instruction[25]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[27]), .QN(n308) );
  DFC3 u_mem_pipe_con_Wmemtoreg_reg ( .D(mem_con_Wmemtoreg), .C(clk), .RN(
        rst_n), .Q(wb_con_Wmemtoreg) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_6_ ( .D(if_addr_j[8]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[6]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_9_ ( .D(if_addr_j[11]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[9]) );
  XNR21 add_x_4_U79 ( .A(n302), .B(add_x_4_n68), .Q(
        u_fetch_jmux_i_addr_pc4_15_) );
  XNR21 add_x_4_U90 ( .A(n303), .B(add_x_4_n78), .Q(
        u_fetch_jmux_i_addr_pc4_13_) );
  NAND22 add_x_4_U12 ( .A(add_x_4_n8), .B(add_x_4_n53), .Q(add_x_4_n7) );
  NAND22 add_x_4_U5 ( .A(add_x_4_n5), .B(instruction_address[29]), .Q(
        add_x_4_n2) );
  XNR21 add_x_4_U56 ( .A(n300), .B(add_x_4_n48), .Q(
        u_fetch_jmux_i_addr_pc4_19_) );
  XNR21 add_x_4_U119 ( .A(n274), .B(add_x_4_n99), .Q(
        u_fetch_jmux_i_addr_pc4_8_) );
  XNR21 add_x_4_U123 ( .A(n306), .B(add_x_4_n103), .Q(
        u_fetch_jmux_i_addr_pc4_7_) );
  OAI210 u_decode_add_x_16_U51 ( .A(u_decode_add_x_16_n69), .B(
        u_decode_add_x_16_n63), .C(u_decode_add_x_16_n64), .Q(
        u_decode_add_x_16_n62) );
  NAND22 add_x_1_U140 ( .A(mem_data_pc4[2]), .B(mem_data_pc4[3]), .Q(
        add_x_1_n113) );
  XNR21 add_x_1_U80 ( .A(add_x_1_n68), .B(add_x_1_n69), .Q(u_mem_pc8[14]) );
  XNR21 u_decode_add_x_16_U6 ( .A(u_decode_add_x_16_n2), .B(
        u_decode_add_x_16_n38), .Q(u_decode_pcadd_o_addr_pcbranchE[30]) );
  XNR21 u_decode_add_x_16_U56 ( .A(u_decode_add_x_16_n8), .B(
        u_decode_add_x_16_n70), .Q(u_decode_pcadd_o_addr_pcbranchE[24]) );
  XNR21 u_decode_add_x_16_U82 ( .A(u_decode_add_x_16_n11), .B(
        u_decode_add_x_16_n92), .Q(u_decode_pcadd_o_addr_pcbranchE[21]) );
  XNR21 u_decode_add_x_16_U28 ( .A(u_decode_add_x_16_n5), .B(
        u_decode_add_x_16_n53), .Q(u_decode_pcadd_o_addr_pcbranchE[27]) );
  XNR21 u_decode_add_x_16_U74 ( .A(u_decode_add_x_16_n10), .B(
        u_decode_add_x_16_n82), .Q(u_decode_pcadd_o_addr_pcbranchE[22]) );
  XNR21 u_decode_add_x_16_U130 ( .A(u_decode_add_x_16_n16), .B(
        u_decode_add_x_16_n120), .Q(u_decode_pcadd_o_addr_pcbranchE[16]) );
  XNR21 u_decode_add_x_16_U20 ( .A(u_decode_add_x_16_n4), .B(
        u_decode_add_x_16_n46), .Q(u_decode_pcadd_o_addr_pcbranchE[28]) );
  XNR21 u_decode_add_x_16_U109 ( .A(u_decode_add_x_16_n14), .B(
        u_decode_add_x_16_n105), .Q(u_decode_pcadd_o_addr_pcbranchE[18]) );
  XNR21 u_decode_add_x_16_U167 ( .A(u_decode_add_x_16_n20), .B(
        u_decode_add_x_16_n145), .Q(u_decode_pcadd_o_addr_pcbranchE[12]) );
  XNR21 u_decode_add_x_16_U175 ( .A(u_decode_add_x_16_n21), .B(
        u_decode_add_x_16_n152), .Q(u_decode_pcadd_o_addr_pcbranchE[11]) );
  XNR21 u_decode_add_x_16_U191 ( .A(u_decode_add_x_16_n23), .B(
        u_decode_add_x_16_n163), .Q(u_decode_pcadd_o_addr_pcbranchE[9]) );
  XNR21 u_decode_add_x_16_U216 ( .A(u_decode_add_x_16_n26), .B(
        u_decode_add_x_16_n176), .Q(u_decode_pcadd_o_addr_pcbranchE[6]) );
  XNR21 u_decode_add_x_16_U224 ( .A(u_decode_add_x_16_n27), .B(
        u_decode_add_x_16_n182), .Q(u_decode_pcadd_o_addr_pcbranchE[5]) );
  XNR21 add_x_4_U108 ( .A(n273), .B(add_x_4_n90), .Q(
        u_fetch_jmux_i_addr_pc4_10_) );
  XNR21 add_x_4_U85 ( .A(n315), .B(add_x_4_n72), .Q(
        u_fetch_jmux_i_addr_pc4_14_) );
  XNR21 add_x_4_U143 ( .A(instruction_address[2]), .B(n318), .Q(
        u_fetch_jmux_i_addr_pc4_3_) );
  XNR21 add_x_4_U139 ( .A(n275), .B(add_x_4_n115), .Q(
        u_fetch_jmux_i_addr_pc4_4_) );
  NOR20 u_decode_add_x_16_U4 ( .A(if_addr_j[31]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n31) );
  NAND22 add_x_4_U145 ( .A(instruction_address[3]), .B(instruction_address[2]), 
        .Q(add_x_4_n116) );
  NAND22 u_decode_add_x_16_U48 ( .A(u_decode_add_x_16_n73), .B(
        u_decode_add_x_16_n61), .Q(u_decode_add_x_16_n59) );
  NAND22 u_decode_add_x_16_U87 ( .A(u_decode_add_x_16_n96), .B(
        u_decode_add_x_16_n88), .Q(u_decode_add_x_16_n86) );
  NAND22 u_decode_add_x_16_U30 ( .A(u_decode_add_x_16_n57), .B(
        u_decode_add_x_16_n49), .Q(u_decode_add_x_16_n47) );
  NAND22 u_decode_add_x_16_U194 ( .A(u_decode_add_x_16_n167), .B(
        u_decode_add_x_16_n159), .Q(u_decode_add_x_16_n157) );
  OAI212 u_decode_add_x_16_U241 ( .A(u_decode_add_x_16_n190), .B(
        u_decode_add_x_16_n187), .C(u_decode_add_x_16_n188), .Q(
        u_decode_add_x_16_n186) );
  OAI212 u_decode_add_x_16_U211 ( .A(u_decode_add_x_16_n175), .B(
        u_decode_add_x_16_n169), .C(u_decode_add_x_16_n170), .Q(
        u_decode_add_x_16_n168) );
  NAND22 u_decode_add_x_16_U159 ( .A(u_decode_add_x_16_n148), .B(
        u_decode_add_x_16_n136), .Q(u_decode_add_x_16_n134) );
  NAND22 u_decode_add_x_16_U122 ( .A(u_decode_add_x_16_n111), .B(
        u_decode_add_x_16_n123), .Q(u_decode_add_x_16_n109) );
  AOI211 u_decode_add_x_16_U49 ( .A(u_decode_add_x_16_n74), .B(
        u_decode_add_x_16_n61), .C(u_decode_add_x_16_n62), .Q(
        u_decode_add_x_16_n60) );
  OAI212 u_decode_add_x_16_U29 ( .A(u_decode_add_x_16_n47), .B(
        u_decode_add_x_16_n106), .C(u_decode_add_x_16_n48), .Q(
        u_decode_add_x_16_n46) );
  OAI212 u_decode_add_x_16_U15 ( .A(u_decode_add_x_16_n39), .B(
        u_decode_add_x_16_n41), .C(u_decode_add_x_16_n40), .Q(
        u_decode_add_x_16_n38) );
  NAND22 add_x_1_U31 ( .A(mem_data_pc4[22]), .B(mem_data_pc4[23]), .Q(
        add_x_1_n24) );
  NOR21 add_x_1_U8 ( .A(add_x_1_n6), .B(add_x_1_n13), .Q(add_x_1_n5) );
  NAND22 add_x_1_U120 ( .A(mem_data_pc4[6]), .B(mem_data_pc4[7]), .Q(
        add_x_1_n97) );
  NAND22 add_x_1_U131 ( .A(mem_data_pc4[4]), .B(mem_data_pc4[5]), .Q(
        add_x_1_n106) );
  NAND22 add_x_1_U100 ( .A(mem_data_pc4[10]), .B(mem_data_pc4[11]), .Q(
        add_x_1_n81) );
  XOR21 add_x_1_U1 ( .A(mem_data_pc4[31]), .B(add_x_1_n1), .Q(u_mem_pc8[31])
         );
  NAND22 add_x_1_U87 ( .A(add_x_1_n87), .B(add_x_1_n71), .Q(add_x_1_n70) );
  NAND22 add_x_1_U75 ( .A(add_x_1_n69), .B(add_x_1_n61), .Q(add_x_1_n60) );
  XOR21 add_x_1_U69 ( .A(add_x_1_n59), .B(add_x_1_n60), .Q(u_mem_pc8[16]) );
  NAND22 add_x_1_U98 ( .A(add_x_1_n87), .B(add_x_1_n80), .Q(add_x_1_n79) );
  XOR21 add_x_1_U92 ( .A(add_x_1_n78), .B(add_x_1_n79), .Q(u_mem_pc8[12]) );
  NAND22 u_decode_add_x_16_U10 ( .A(u_decode_add_x_16_n34), .B(
        u_decode_add_x_16_n37), .Q(u_decode_add_x_16_n2) );
  OAI212 u_decode_add_x_16_U65 ( .A(u_decode_add_x_16_n71), .B(
        u_decode_add_x_16_n83), .C(u_decode_add_x_16_n72), .Q(
        u_decode_add_x_16_n70) );
  XOR21 u_decode_add_x_16_U44 ( .A(u_decode_add_x_16_n7), .B(
        u_decode_add_x_16_n65), .Q(u_decode_pcadd_o_addr_pcbranchE[25]) );
  XOR21 u_decode_add_x_16_U64 ( .A(u_decode_add_x_16_n9), .B(
        u_decode_add_x_16_n77), .Q(u_decode_pcadd_o_addr_pcbranchE[23]) );
  OAI212 u_decode_add_x_16_U158 ( .A(u_decode_add_x_16_n134), .B(
        u_decode_add_x_16_n155), .C(u_decode_add_x_16_n135), .Q(
        u_decode_add_x_16_n133) );
  OAI212 u_decode_add_x_16_U139 ( .A(u_decode_add_x_16_n121), .B(
        u_decode_add_x_16_n132), .C(u_decode_add_x_16_n122), .Q(
        u_decode_add_x_16_n120) );
  XOR21 add_x_1_U34 ( .A(add_x_1_n30), .B(add_x_1_n31), .Q(u_mem_pc8[22]) );
  OAI212 u_decode_add_x_16_U176 ( .A(u_decode_add_x_16_n146), .B(
        u_decode_add_x_16_n155), .C(u_decode_add_x_16_n147), .Q(
        u_decode_add_x_16_n145) );
  NAND22 add_x_1_U29 ( .A(add_x_1_n32), .B(add_x_1_n23), .Q(add_x_1_n22) );
  XOR21 add_x_1_U23 ( .A(add_x_1_n21), .B(add_x_1_n22), .Q(u_mem_pc8[24]) );
  ADD22 add_x_1_U3 ( .A(add_x_1_n3), .B(mem_data_pc4[29]), .CO(add_x_1_n2), 
        .S(u_mem_pc8[29]) );
  NAND22 add_x_4_U116 ( .A(instruction_address[8]), .B(instruction_address[9]), 
        .Q(add_x_4_n93) );
  NAND22 add_x_4_U125 ( .A(instruction_address[6]), .B(instruction_address[7]), 
        .Q(add_x_4_n100) );
  NAND22 add_x_4_U136 ( .A(instruction_address[4]), .B(instruction_address[5]), 
        .Q(add_x_4_n109) );
  NAND22 add_x_4_U94 ( .A(instruction_address[12]), .B(instruction_address[13]), .Q(add_x_4_n75) );
  NAND22 add_x_4_U105 ( .A(instruction_address[10]), .B(
        instruction_address[11]), .Q(add_x_4_n84) );
  NAND22 add_x_4_U82 ( .A(instruction_address[14]), .B(instruction_address[15]), .Q(add_x_4_n65) );
  XOR21 add_x_4_U74 ( .A(n314), .B(add_x_4_n63), .Q(
        u_fetch_jmux_i_addr_pc4_16_) );
  NAND22 add_x_4_U71 ( .A(instruction_address[16]), .B(instruction_address[17]), .Q(add_x_4_n56) );
  NOR21 add_x_4_U98 ( .A(n316), .B(add_x_4_n82), .Q(add_x_4_n78) );
  NAND22 add_x_4_U49 ( .A(instruction_address[20]), .B(instruction_address[21]), .Q(add_x_4_n38) );
  NAND22 add_x_4_U58 ( .A(instruction_address[18]), .B(instruction_address[19]), .Q(add_x_4_n45) );
  NAND22 add_x_4_U36 ( .A(instruction_address[22]), .B(instruction_address[23]), .Q(add_x_4_n27) );
  NAND22 add_x_4_U14 ( .A(instruction_address[26]), .B(instruction_address[27]), .Q(add_x_4_n9) );
  NAND22 add_x_4_U18 ( .A(add_x_4_n15), .B(instruction_address[26]), .Q(
        add_x_4_n12) );
  NAND22 add_x_4_U53 ( .A(add_x_4_n44), .B(instruction_address[20]), .Q(
        add_x_4_n41) );
  NOR21 u_decode_add_x_16_U222 ( .A(id_addr_pc4[6]), .B(if_addr_j[6]), .Q(
        u_decode_add_x_16_n174) );
  NAND22 u_decode_add_x_16_U250 ( .A(if_addr_j[2]), .B(id_addr_pc4[2]), .Q(
        u_decode_add_x_16_n190) );
  NAND22 u_decode_add_x_16_U238 ( .A(if_addr_j[4]), .B(id_addr_pc4[4]), .Q(
        u_decode_add_x_16_n184) );
  NAND22 u_decode_add_x_16_U223 ( .A(if_addr_j[6]), .B(id_addr_pc4[6]), .Q(
        u_decode_add_x_16_n175) );
  NAND22 u_decode_add_x_16_U207 ( .A(if_addr_j[8]), .B(id_addr_pc4[8]), .Q(
        u_decode_add_x_16_n165) );
  NAND22 u_decode_add_x_16_U190 ( .A(if_addr_j[10]), .B(id_addr_pc4[10]), .Q(
        u_decode_add_x_16_n154) );
  NAND22 u_decode_add_x_16_U174 ( .A(if_addr_j[12]), .B(id_addr_pc4[12]), .Q(
        u_decode_add_x_16_n144) );
  NAND22 u_decode_add_x_16_U155 ( .A(if_addr_j[14]), .B(id_addr_pc4[14]), .Q(
        u_decode_add_x_16_n131) );
  NAND22 u_decode_add_x_16_U116 ( .A(n346), .B(id_addr_pc4[18]), .Q(
        u_decode_add_x_16_n104) );
  NAND22 u_decode_add_x_16_U100 ( .A(n346), .B(id_addr_pc4[20]), .Q(
        u_decode_add_x_16_n94) );
  NAND22 u_decode_add_x_16_U81 ( .A(n346), .B(id_addr_pc4[22]), .Q(
        u_decode_add_x_16_n81) );
  NAND22 u_decode_add_x_16_U63 ( .A(n346), .B(id_addr_pc4[24]), .Q(
        u_decode_add_x_16_n69) );
  NOR21 u_decode_add_x_16_U26 ( .A(if_addr_j[28]), .B(n346), .Q(
        u_decode_add_x_16_n44) );
  NAND22 u_decode_add_x_16_U27 ( .A(n346), .B(if_addr_j[28]), .Q(
        u_decode_add_x_16_n45) );
  NAND22 add_x_1_U44 ( .A(mem_data_pc4[20]), .B(mem_data_pc4[21]), .Q(
        add_x_1_n35) );
  NAND22 add_x_1_U53 ( .A(mem_data_pc4[18]), .B(mem_data_pc4[19]), .Q(
        add_x_1_n42) );
  NAND22 add_x_1_U111 ( .A(mem_data_pc4[8]), .B(mem_data_pc4[9]), .Q(
        add_x_1_n90) );
  NAND22 add_x_1_U89 ( .A(mem_data_pc4[12]), .B(mem_data_pc4[13]), .Q(
        add_x_1_n72) );
  NAND22 add_x_1_U77 ( .A(mem_data_pc4[14]), .B(mem_data_pc4[15]), .Q(
        add_x_1_n62) );
  ADD22 add_x_1_U2 ( .A(add_x_1_n2), .B(mem_data_pc4[30]), .CO(add_x_1_n1), 
        .S(u_mem_pc8[30]) );
  NAND22 u_decode_add_x_16_U52 ( .A(u_decode_add_x_16_n197), .B(
        u_decode_add_x_16_n64), .Q(u_decode_add_x_16_n7) );
  NAND22 u_decode_add_x_16_U60 ( .A(u_decode_add_x_16_n66), .B(
        u_decode_add_x_16_n69), .Q(u_decode_add_x_16_n8) );
  NAND22 u_decode_add_x_16_U70 ( .A(u_decode_add_x_16_n199), .B(
        u_decode_add_x_16_n76), .Q(u_decode_add_x_16_n9) );
  NAND22 u_decode_add_x_16_U91 ( .A(u_decode_add_x_16_n201), .B(
        u_decode_add_x_16_n91), .Q(u_decode_add_x_16_n11) );
  NAND22 u_decode_add_x_16_U34 ( .A(u_decode_add_x_16_n195), .B(
        u_decode_add_x_16_n52), .Q(u_decode_add_x_16_n5) );
  DFC3 u_decode_pipe_con_Ealuop_reg_3_ ( .D(u_decode_control_o_con_aluop_3_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[3]) );
  DFC3 u_decode_pipe_con_Ealuop_reg_1_ ( .D(u_decode_control_o_con_aluop_1_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[1]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_4_ ( .D(if_addr_j[6]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[4]) );
  DFC3 u_decode_pipe_FWmemout_reg_27_ ( .D(wb_data_memout[27]), .C(clk), .RN(
        rst_n), .Q(for_memout[27]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_0_ ( .D(if_addr_j[2]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[0]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_8_ ( .D(if_addr_j[10]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[8]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_7_ ( .D(if_addr_j[9]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[7]) );
  DFC3 u_fetch_pipe_instr_reg_20_ ( .D(read_instruction[20]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[22]), .QN(n277) );
  NAND22 u_decode_add_x_16_U245 ( .A(if_addr_j[3]), .B(id_addr_pc4[3]), .Q(
        u_decode_add_x_16_n188) );
  NAND21 u_decode_add_x_16_U166 ( .A(if_addr_j[13]), .B(id_addr_pc4[13]), .Q(
        u_decode_add_x_16_n139) );
  NAND21 u_decode_add_x_16_U147 ( .A(if_addr_j[15]), .B(id_addr_pc4[15]), .Q(
        u_decode_add_x_16_n126) );
  NAND22 u_decode_add_x_16_U137 ( .A(if_addr_j[16]), .B(id_addr_pc4[16]), .Q(
        u_decode_add_x_16_n119) );
  NAND21 u_decode_add_x_16_U201 ( .A(if_addr_j[9]), .B(id_addr_pc4[9]), .Q(
        u_decode_add_x_16_n162) );
  OAI211 u_decode_add_x_16_U197 ( .A(u_decode_add_x_16_n165), .B(
        u_decode_add_x_16_n161), .C(u_decode_add_x_16_n162), .Q(
        u_decode_add_x_16_n160) );
  NAND22 u_decode_add_x_16_U73 ( .A(n346), .B(id_addr_pc4[23]), .Q(
        u_decode_add_x_16_n76) );
  NAND22 u_decode_add_x_16_U13 ( .A(n346), .B(if_addr_j[30]), .Q(
        u_decode_add_x_16_n37) );
  NAND22 u_decode_add_x_16_U19 ( .A(n346), .B(if_addr_j[29]), .Q(
        u_decode_add_x_16_n40) );
  NAND21 u_decode_add_x_16_U129 ( .A(n346), .B(id_addr_pc4[17]), .Q(
        u_decode_add_x_16_n114) );
  NAND22 u_decode_add_x_16_U108 ( .A(n346), .B(id_addr_pc4[19]), .Q(
        u_decode_add_x_16_n99) );
  NAND22 u_decode_add_x_16_U43 ( .A(n346), .B(id_addr_pc4[26]), .Q(
        u_decode_add_x_16_n55) );
  NOR21 u_decode_add_x_16_U12 ( .A(if_addr_j[30]), .B(n346), .Q(
        u_decode_add_x_16_n36) );
  NAND21 u_decode_add_x_16_U5 ( .A(n346), .B(if_addr_j[31]), .Q(
        u_decode_add_x_16_n32) );
  OAI211 u_decode_add_x_16_U162 ( .A(u_decode_add_x_16_n144), .B(
        u_decode_add_x_16_n138), .C(u_decode_add_x_16_n139), .Q(
        u_decode_add_x_16_n137) );
  OAI211 u_decode_add_x_16_U90 ( .A(u_decode_add_x_16_n94), .B(
        u_decode_add_x_16_n90), .C(u_decode_add_x_16_n91), .Q(
        u_decode_add_x_16_n89) );
  OAI211 u_decode_add_x_16_U234 ( .A(u_decode_add_x_16_n183), .B(
        u_decode_add_x_16_n185), .C(u_decode_add_x_16_n184), .Q(
        u_decode_add_x_16_n182) );
  XOR21 add_x_4_U133 ( .A(n307), .B(add_x_4_n112), .Q(
        u_fetch_jmux_i_addr_pc4_5_) );
  XOR21 add_x_4_U128 ( .A(n317), .B(add_x_4_n107), .Q(
        u_fetch_jmux_i_addr_pc4_6_) );
  NOR21 add_x_4_U129 ( .A(n317), .B(add_x_4_n107), .Q(add_x_4_n103) );
  XOR21 add_x_4_U61 ( .A(n313), .B(add_x_4_n52), .Q(
        u_fetch_jmux_i_addr_pc4_18_) );
  NOR21 add_x_4_U62 ( .A(n313), .B(add_x_4_n52), .Q(add_x_4_n48) );
  XOR21 add_x_4_U8 ( .A(n324), .B(add_x_4_n7), .Q(u_fetch_jmux_i_addr_pc4_28_)
         );
  NOR21 add_x_4_U86 ( .A(n315), .B(add_x_4_n73), .Q(add_x_4_n68) );
  XOR21 add_x_4_U97 ( .A(n316), .B(add_x_4_n82), .Q(
        u_fetch_jmux_i_addr_pc4_12_) );
  ADD22 add_x_1_U4 ( .A(add_x_1_n118), .B(mem_data_pc4[28]), .CO(add_x_1_n3), 
        .S(u_mem_pc8[28]) );
  ADD22 add_x_4_U2 ( .A(add_x_4_n121), .B(instruction_address[30]), .CO(
        add_x_4_n1), .S(u_fetch_jmux_i_addr_pc4_30_) );
  OAI211 u_decode_add_x_16_U33 ( .A(u_decode_add_x_16_n55), .B(
        u_decode_add_x_16_n51), .C(u_decode_add_x_16_n52), .Q(
        u_decode_add_x_16_n50) );
  XOR21 u_decode_add_x_16_U148 ( .A(u_decode_add_x_16_n18), .B(
        u_decode_add_x_16_n132), .Q(u_decode_pcadd_o_addr_pcbranchE[14]) );
  NOR21 u_decode_add_x_16_U244 ( .A(id_addr_pc4[3]), .B(if_addr_j[3]), .Q(
        u_decode_add_x_16_n187) );
  NAND22 u_decode_add_x_16_U232 ( .A(if_addr_j[5]), .B(id_addr_pc4[5]), .Q(
        u_decode_add_x_16_n181) );
  NAND22 u_decode_add_x_16_U37 ( .A(n346), .B(id_addr_pc4[27]), .Q(
        u_decode_add_x_16_n52) );
  NAND22 u_decode_add_x_16_U94 ( .A(n346), .B(id_addr_pc4[21]), .Q(
        u_decode_add_x_16_n91) );
  NOR21 u_decode_add_x_16_U50 ( .A(u_decode_add_x_16_n63), .B(
        u_decode_add_x_16_n68), .Q(u_decode_add_x_16_n61) );
  NOR21 add_x_1_U119 ( .A(add_x_1_n97), .B(add_x_1_n104), .Q(add_x_1_n96) );
  NAND22 add_x_4_U103 ( .A(add_x_4_n90), .B(add_x_4_n83), .Q(add_x_4_n82) );
  AOI211 u_decode_add_x_16_U31 ( .A(u_decode_add_x_16_n58), .B(
        u_decode_add_x_16_n49), .C(u_decode_add_x_16_n50), .Q(
        u_decode_add_x_16_n48) );
  XOR21 add_x_4_U102 ( .A(n304), .B(add_x_4_n87), .Q(
        u_fetch_jmux_i_addr_pc4_11_) );
  XOR21 add_x_4_U112 ( .A(n305), .B(add_x_4_n96), .Q(
        u_fetch_jmux_i_addr_pc4_9_) );
  XNR21 add_x_4_U52 ( .A(n272), .B(add_x_4_n44), .Q(
        u_fetch_jmux_i_addr_pc4_20_) );
  XNR21 add_x_4_U17 ( .A(n271), .B(add_x_4_n15), .Q(
        u_fetch_jmux_i_addr_pc4_26_) );
  XNR21 add_x_4_U4 ( .A(n295), .B(add_x_4_n5), .Q(u_fetch_jmux_i_addr_pc4_29_)
         );
  XOR21 add_x_4_U44 ( .A(n299), .B(add_x_4_n41), .Q(
        u_fetch_jmux_i_addr_pc4_21_) );
  XNR21 add_x_4_U66 ( .A(n301), .B(add_x_4_n59), .Q(
        u_fetch_jmux_i_addr_pc4_17_) );
  NOR21 u_decode_add_x_16_U136 ( .A(id_addr_pc4[16]), .B(if_addr_j[16]), .Q(
        u_decode_add_x_16_n118) );
  NAND22 add_x_1_U9 ( .A(mem_data_pc4[26]), .B(mem_data_pc4[27]), .Q(
        add_x_1_n6) );
  NAND22 u_decode_add_x_16_U215 ( .A(if_addr_j[7]), .B(id_addr_pc4[7]), .Q(
        u_decode_add_x_16_n170) );
  NAND22 u_decode_add_x_16_U184 ( .A(if_addr_j[11]), .B(id_addr_pc4[11]), .Q(
        u_decode_add_x_16_n151) );
  NOR21 u_decode_add_x_16_U62 ( .A(id_addr_pc4[24]), .B(n346), .Q(
        u_decode_add_x_16_n68) );
  NOR21 u_decode_add_x_16_U18 ( .A(if_addr_j[29]), .B(n346), .Q(
        u_decode_add_x_16_n39) );
  NOR21 u_decode_add_x_16_U227 ( .A(u_decode_add_x_16_n180), .B(
        u_decode_add_x_16_n183), .Q(u_decode_add_x_16_n178) );
  NOR21 u_decode_add_x_16_U210 ( .A(u_decode_add_x_16_n169), .B(
        u_decode_add_x_16_n174), .Q(u_decode_add_x_16_n167) );
  NOR21 u_decode_add_x_16_U124 ( .A(u_decode_add_x_16_n118), .B(
        u_decode_add_x_16_n113), .Q(u_decode_add_x_16_n111) );
  NOR21 u_decode_add_x_16_U32 ( .A(u_decode_add_x_16_n51), .B(
        u_decode_add_x_16_n54), .Q(u_decode_add_x_16_n49) );
  NOR21 add_x_4_U13 ( .A(add_x_4_n9), .B(add_x_4_n16), .Q(add_x_4_n8) );
  NOR21 add_x_1_U17 ( .A(add_x_1_n13), .B(add_x_1_n49), .Q(add_x_1_n12) );
  NOR21 add_x_1_U52 ( .A(add_x_1_n42), .B(add_x_1_n49), .Q(add_x_1_n41) );
  NAND22 add_x_4_U34 ( .A(add_x_4_n35), .B(add_x_4_n26), .Q(add_x_4_n25) );
  XOR21 add_x_4_U11 ( .A(n296), .B(add_x_4_n12), .Q(
        u_fetch_jmux_i_addr_pc4_27_) );
  NOR21 add_x_4_U75 ( .A(n314), .B(add_x_4_n63), .Q(add_x_4_n59) );
  XOR21 add_x_4_U28 ( .A(n311), .B(add_x_4_n25), .Q(
        u_fetch_jmux_i_addr_pc4_24_) );
  XOR21 add_x_4_U39 ( .A(n312), .B(add_x_4_n34), .Q(
        u_fetch_jmux_i_addr_pc4_22_) );
  XNR21 add_x_4_U21 ( .A(n297), .B(add_x_4_n21), .Q(
        u_fetch_jmux_i_addr_pc4_25_) );
  XNR21 add_x_4_U33 ( .A(n298), .B(add_x_4_n30), .Q(
        u_fetch_jmux_i_addr_pc4_23_) );
  XOR21 add_x_4_U1 ( .A(instruction_address[31]), .B(add_x_4_n1), .Q(
        u_fetch_jmux_i_addr_pc4_31_) );
  NOR21 u_decode_add_x_16_U173 ( .A(id_addr_pc4[12]), .B(if_addr_j[12]), .Q(
        u_decode_add_x_16_n143) );
  NOR21 u_decode_add_x_16_U154 ( .A(id_addr_pc4[14]), .B(if_addr_j[14]), .Q(
        u_decode_add_x_16_n130) );
  NOR21 add_x_1_U110 ( .A(add_x_1_n90), .B(add_x_1_n97), .Q(add_x_1_n89) );
  NOR21 u_decode_add_x_16_U179 ( .A(u_decode_add_x_16_n150), .B(
        u_decode_add_x_16_n153), .Q(u_decode_add_x_16_n148) );
  NOR21 add_x_1_U88 ( .A(add_x_1_n72), .B(add_x_1_n81), .Q(add_x_1_n71) );
  NAND22 u_decode_add_x_16_U55 ( .A(n346), .B(id_addr_pc4[25]), .Q(
        u_decode_add_x_16_n64) );
  NOR21 add_x_4_U70 ( .A(add_x_4_n56), .B(add_x_4_n65), .Q(add_x_4_n55) );
  NOR21 add_x_1_U43 ( .A(add_x_1_n35), .B(add_x_1_n42), .Q(add_x_1_n34) );
  NOR21 u_decode_add_x_16_U142 ( .A(u_decode_add_x_16_n125), .B(
        u_decode_add_x_16_n130), .Q(u_decode_add_x_16_n123) );
  NOR21 u_decode_add_x_16_U161 ( .A(u_decode_add_x_16_n138), .B(
        u_decode_add_x_16_n143), .Q(u_decode_add_x_16_n136) );
  NOR21 u_decode_add_x_16_U68 ( .A(u_decode_add_x_16_n75), .B(
        u_decode_add_x_16_n80), .Q(u_decode_add_x_16_n73) );
  NAND22 add_x_4_U69 ( .A(add_x_4_n74), .B(add_x_4_n55), .Q(add_x_4_n54) );
  NAND22 add_x_1_U109 ( .A(add_x_1_n89), .B(add_x_1_n105), .Q(add_x_1_n88) );
  AOI211 u_decode_add_x_16_U195 ( .A(u_decode_add_x_16_n168), .B(
        u_decode_add_x_16_n159), .C(u_decode_add_x_16_n160), .Q(
        u_decode_add_x_16_n158) );
  NAND21 add_x_4_U140 ( .A(add_x_4_n115), .B(instruction_address[4]), .Q(
        add_x_4_n112) );
  AOI211 u_decode_add_x_16_U160 ( .A(u_decode_add_x_16_n149), .B(
        u_decode_add_x_16_n136), .C(u_decode_add_x_16_n137), .Q(
        u_decode_add_x_16_n135) );
  NOR21 add_x_4_U124 ( .A(add_x_4_n100), .B(add_x_4_n107), .Q(add_x_4_n99) );
  NOR21 u_decode_add_x_16_U46 ( .A(u_decode_add_x_16_n59), .B(
        u_decode_add_x_16_n86), .Q(u_decode_add_x_16_n57) );
  NAND22 add_x_4_U92 ( .A(add_x_4_n90), .B(add_x_4_n74), .Q(add_x_4_n73) );
  OAI211 u_decode_add_x_16_U203 ( .A(u_decode_add_x_16_n164), .B(
        u_decode_add_x_16_n166), .C(u_decode_add_x_16_n165), .Q(
        u_decode_add_x_16_n163) );
  NAND22 add_x_4_U80 ( .A(add_x_4_n72), .B(add_x_4_n64), .Q(add_x_4_n63) );
  NOR21 add_x_4_U29 ( .A(n311), .B(add_x_4_n25), .Q(add_x_4_n21) );
  NOR21 add_x_4_U40 ( .A(n312), .B(add_x_4_n34), .Q(add_x_4_n30) );
  NOR21 u_decode_add_x_16_U196 ( .A(u_decode_add_x_16_n161), .B(
        u_decode_add_x_16_n164), .Q(u_decode_add_x_16_n159) );
  NOR21 u_decode_add_x_16_U80 ( .A(id_addr_pc4[22]), .B(n346), .Q(
        u_decode_add_x_16_n80) );
  NOR21 add_x_4_U115 ( .A(add_x_4_n93), .B(add_x_4_n100), .Q(add_x_4_n92) );
  NOR21 add_x_4_U48 ( .A(add_x_4_n38), .B(add_x_4_n45), .Q(add_x_4_n37) );
  NAND22 add_x_4_U114 ( .A(add_x_4_n92), .B(add_x_4_n108), .Q(add_x_4_n91) );
  NOR21 u_decode_add_x_16_U103 ( .A(u_decode_add_x_16_n98), .B(
        u_decode_add_x_16_n103), .Q(u_decode_add_x_16_n96) );
  NOR21 add_x_4_U22 ( .A(add_x_4_n16), .B(add_x_4_n52), .Q(add_x_4_n15) );
  NOR21 add_x_1_U41 ( .A(add_x_1_n33), .B(add_x_1_n49), .Q(add_x_1_n32) );
  NOR21 add_x_4_U57 ( .A(add_x_4_n45), .B(add_x_4_n52), .Q(add_x_4_n44) );
  OAI211 u_decode_add_x_16_U186 ( .A(u_decode_add_x_16_n153), .B(
        u_decode_add_x_16_n155), .C(u_decode_add_x_16_n154), .Q(
        u_decode_add_x_16_n152) );
  AOI211 u_decode_add_x_16_U57 ( .A(u_decode_add_x_16_n70), .B(
        u_decode_add_x_16_n66), .C(u_decode_add_x_16_n67), .Q(
        u_decode_add_x_16_n65) );
  AOI211 u_decode_add_x_16_U75 ( .A(u_decode_add_x_16_n82), .B(
        u_decode_add_x_16_n78), .C(u_decode_add_x_16_n79), .Q(
        u_decode_add_x_16_n77) );
  NOR21 u_decode_add_x_16_U200 ( .A(id_addr_pc4[9]), .B(if_addr_j[9]), .Q(
        u_decode_add_x_16_n161) );
  NOR21 u_decode_add_x_16_U115 ( .A(id_addr_pc4[18]), .B(n346), .Q(
        u_decode_add_x_16_n103) );
  NOR21 add_x_4_U93 ( .A(add_x_4_n75), .B(add_x_4_n84), .Q(add_x_4_n74) );
  NOR21 u_decode_add_x_16_U89 ( .A(u_decode_add_x_16_n90), .B(
        u_decode_add_x_16_n93), .Q(u_decode_add_x_16_n88) );
  AOI211 u_decode_add_x_16_U226 ( .A(u_decode_add_x_16_n186), .B(
        u_decode_add_x_16_n178), .C(u_decode_add_x_16_n179), .Q(
        u_decode_add_x_16_n177) );
  AOI211 u_decode_add_x_16_U88 ( .A(u_decode_add_x_16_n97), .B(
        u_decode_add_x_16_n88), .C(u_decode_add_x_16_n89), .Q(
        u_decode_add_x_16_n87) );
  AOI211 u_decode_add_x_16_U209 ( .A(u_decode_add_x_16_n176), .B(
        u_decode_add_x_16_n167), .C(u_decode_add_x_16_n168), .Q(
        u_decode_add_x_16_n166) );
  NOR21 add_x_4_U9 ( .A(n324), .B(add_x_4_n7), .Q(add_x_4_n5) );
  NOR21 add_x_4_U46 ( .A(add_x_4_n36), .B(add_x_4_n52), .Q(add_x_4_n35) );
  NOR21 u_decode_add_x_16_U165 ( .A(id_addr_pc4[13]), .B(if_addr_j[13]), .Q(
        u_decode_add_x_16_n138) );
  NOR21 u_decode_add_x_16_U231 ( .A(id_addr_pc4[5]), .B(if_addr_j[5]), .Q(
        u_decode_add_x_16_n180) );
  NOR21 u_decode_add_x_16_U206 ( .A(id_addr_pc4[8]), .B(if_addr_j[8]), .Q(
        u_decode_add_x_16_n164) );
  NOR21 u_decode_add_x_16_U189 ( .A(id_addr_pc4[10]), .B(if_addr_j[10]), .Q(
        u_decode_add_x_16_n153) );
  OAI211 u_decode_add_x_16_U228 ( .A(u_decode_add_x_16_n184), .B(
        u_decode_add_x_16_n180), .C(u_decode_add_x_16_n181), .Q(
        u_decode_add_x_16_n179) );
  NOR21 add_x_1_U130 ( .A(add_x_1_n113), .B(add_x_1_n106), .Q(add_x_1_n105) );
  NAND21 add_x_4_U109 ( .A(add_x_4_n90), .B(instruction_address[10]), .Q(
        add_x_4_n87) );
  XOR20 add_x_1_U56 ( .A(add_x_1_n48), .B(add_x_1_n49), .Q(u_mem_pc8[18]) );
  NOR21 u_decode_add_x_16_U183 ( .A(id_addr_pc4[11]), .B(if_addr_j[11]), .Q(
        u_decode_add_x_16_n150) );
  NOR21 u_decode_add_x_16_U237 ( .A(id_addr_pc4[4]), .B(if_addr_j[4]), .Q(
        u_decode_add_x_16_n183) );
  NOR21 u_decode_add_x_16_U214 ( .A(id_addr_pc4[7]), .B(if_addr_j[7]), .Q(
        u_decode_add_x_16_n169) );
  NOR21 u_decode_add_x_16_U146 ( .A(id_addr_pc4[15]), .B(if_addr_j[15]), .Q(
        u_decode_add_x_16_n125) );
  NOR21 u_decode_add_x_16_U54 ( .A(id_addr_pc4[25]), .B(n346), .Q(
        u_decode_add_x_16_n63) );
  NOR21 add_x_4_U135 ( .A(add_x_4_n116), .B(add_x_4_n109), .Q(add_x_4_n108) );
  OAI211 u_decode_add_x_16_U143 ( .A(u_decode_add_x_16_n131), .B(
        u_decode_add_x_16_n125), .C(u_decode_add_x_16_n126), .Q(
        u_decode_add_x_16_n124) );
  NOR21 add_x_4_U68 ( .A(add_x_4_n91), .B(add_x_4_n54), .Q(add_x_4_n53) );
  AOI211 u_decode_add_x_16_U102 ( .A(u_decode_add_x_16_n105), .B(
        u_decode_add_x_16_n96), .C(u_decode_add_x_16_n97), .Q(
        u_decode_add_x_16_n95) );
  AOI211 u_decode_add_x_16_U84 ( .A(u_decode_add_x_16_n105), .B(
        u_decode_add_x_16_n84), .C(u_decode_add_x_16_n85), .Q(
        u_decode_add_x_16_n83) );
  AOI211 u_decode_add_x_16_U45 ( .A(u_decode_add_x_16_n105), .B(
        u_decode_add_x_16_n57), .C(u_decode_add_x_16_n58), .Q(
        u_decode_add_x_16_n56) );
  OAI211 u_decode_add_x_16_U96 ( .A(u_decode_add_x_16_n93), .B(
        u_decode_add_x_16_n95), .C(u_decode_add_x_16_n94), .Q(
        u_decode_add_x_16_n92) );
  OAI211 u_decode_add_x_16_U39 ( .A(u_decode_add_x_16_n54), .B(
        u_decode_add_x_16_n56), .C(u_decode_add_x_16_n55), .Q(
        u_decode_add_x_16_n53) );
  NOR21 u_decode_add_x_16_U36 ( .A(id_addr_pc4[27]), .B(n346), .Q(
        u_decode_add_x_16_n51) );
  NOR21 u_decode_add_x_16_U42 ( .A(id_addr_pc4[26]), .B(n346), .Q(
        u_decode_add_x_16_n54) );
  NOR21 u_decode_add_x_16_U72 ( .A(id_addr_pc4[23]), .B(n346), .Q(
        u_decode_add_x_16_n75) );
  NOR21 u_decode_add_x_16_U128 ( .A(id_addr_pc4[17]), .B(n346), .Q(
        u_decode_add_x_16_n113) );
  NOR21 u_decode_add_x_16_U93 ( .A(id_addr_pc4[21]), .B(n346), .Q(
        u_decode_add_x_16_n90) );
  NOR21 u_decode_add_x_16_U99 ( .A(id_addr_pc4[20]), .B(n346), .Q(
        u_decode_add_x_16_n93) );
  NOR21 u_decode_add_x_16_U107 ( .A(id_addr_pc4[19]), .B(n346), .Q(
        u_decode_add_x_16_n98) );
  NAND21 u_decode_add_x_16_U229 ( .A(u_decode_add_x_16_n217), .B(
        u_decode_add_x_16_n181), .Q(u_decode_add_x_16_n27) );
  OAI210 u_decode_add_x_16_U125 ( .A(u_decode_add_x_16_n119), .B(
        u_decode_add_x_16_n113), .C(u_decode_add_x_16_n114), .Q(
        u_decode_add_x_16_n112) );
  OAI211 u_decode_add_x_16_U69 ( .A(u_decode_add_x_16_n81), .B(
        u_decode_add_x_16_n75), .C(u_decode_add_x_16_n76), .Q(
        u_decode_add_x_16_n74) );
  NAND21 u_decode_add_x_16_U24 ( .A(u_decode_add_x_16_n42), .B(
        u_decode_add_x_16_n45), .Q(u_decode_add_x_16_n4) );
  NAND21 add_x_4_U120 ( .A(add_x_4_n99), .B(instruction_address[8]), .Q(
        add_x_4_n96) );
  AOI211 u_decode_add_x_16_U21 ( .A(u_decode_add_x_16_n46), .B(
        u_decode_add_x_16_n42), .C(u_decode_add_x_16_n43), .Q(
        u_decode_add_x_16_n41) );
  OAI211 u_decode_add_x_16_U180 ( .A(u_decode_add_x_16_n154), .B(
        u_decode_add_x_16_n150), .C(u_decode_add_x_16_n151), .Q(
        u_decode_add_x_16_n149) );
  NAND21 u_decode_add_x_16_U220 ( .A(u_decode_add_x_16_n216), .B(
        u_decode_add_x_16_n175), .Q(u_decode_add_x_16_n26) );
  NAND21 u_decode_add_x_16_U198 ( .A(u_decode_add_x_16_n213), .B(
        u_decode_add_x_16_n162), .Q(u_decode_add_x_16_n23) );
  NAND21 u_decode_add_x_16_U152 ( .A(u_decode_add_x_16_n208), .B(
        u_decode_add_x_16_n131), .Q(u_decode_add_x_16_n18) );
  NAND21 u_decode_add_x_16_U113 ( .A(u_decode_add_x_16_n204), .B(
        u_decode_add_x_16_n104), .Q(u_decode_add_x_16_n14) );
  XOR20 add_x_1_U123 ( .A(add_x_1_n103), .B(add_x_1_n104), .Q(u_mem_pc8[6]) );
  NAND22 add_x_1_U7 ( .A(add_x_1_n5), .B(add_x_1_n50), .Q(add_x_1_n4) );
  OAI212 u_decode_add_x_16_U47 ( .A(u_decode_add_x_16_n59), .B(
        u_decode_add_x_16_n87), .C(u_decode_add_x_16_n60), .Q(
        u_decode_add_x_16_n58) );
  OAI212 u_decode_add_x_16_U104 ( .A(u_decode_add_x_16_n104), .B(
        u_decode_add_x_16_n98), .C(u_decode_add_x_16_n99), .Q(
        u_decode_add_x_16_n97) );
  NAND21 u_decode_add_x_16_U134 ( .A(u_decode_add_x_16_n206), .B(
        u_decode_add_x_16_n119), .Q(u_decode_add_x_16_n16) );
  NAND21 u_decode_add_x_16_U171 ( .A(u_decode_add_x_16_n210), .B(
        u_decode_add_x_16_n144), .Q(u_decode_add_x_16_n20) );
  NAND21 u_decode_add_x_16_U181 ( .A(u_decode_add_x_16_n211), .B(
        u_decode_add_x_16_n151), .Q(u_decode_add_x_16_n21) );
  NAND21 u_decode_add_x_16_U78 ( .A(u_decode_add_x_16_n78), .B(
        u_decode_add_x_16_n81), .Q(u_decode_add_x_16_n10) );
  DFC3 u_fetch_pipe_instr_reg_31_ ( .D(read_instruction[31]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[31]), .QN(n269) );
  DFC3 u_fetch_pipe_instr_reg_27_ ( .D(read_instruction[27]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[27]), .QN(n268) );
  DFC3 u_decode_pipe_con_Ealuop_reg_4_ ( .D(u_decode_control_o_con_aluop_4_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[4]) );
  DFC3 u_fetch_pipe_instr_reg_15_ ( .D(read_instruction[15]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[17]), .QN(n266) );
  DFC3 u_fetch_pipe_instr_reg_30_ ( .D(read_instruction[30]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[30]), .QN(n310) );
  NAND28 U204 ( .A(n452), .B(u_fetch_jmux_i_addr_pc4_18_), .Q(n260) );
  NAND22 U205 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_28_), .Q(n378) );
  NAND33 U206 ( .A(n371), .B(n369), .C(n370), .Q(n107) );
  NAND33 U207 ( .A(n456), .B(n455), .C(n454), .Q(n125) );
  NAND33 U208 ( .A(n395), .B(n393), .C(n394), .Q(n112) );
  NAND33 U209 ( .A(n461), .B(n460), .C(n459), .Q(n126) );
  NAND33 U210 ( .A(n420), .B(n419), .C(n418), .Q(n117) );
  NAND33 U211 ( .A(n488), .B(n487), .C(n486), .Q(n132) );
  AOI211 U212 ( .A(id_data_jr[27]), .B(n255), .C(n381), .Q(n385) );
  AOI211 U213 ( .A(id_data_jr[24]), .B(n255), .C(n396), .Q(n400) );
  AOI211 U214 ( .A(id_data_jr[31]), .B(n255), .C(n360), .Q(n366) );
  AOI212 U215 ( .A(u_fetch_jmux_i_addr_pc4_13_), .B(n452), .C(n446), .Q(n450)
         );
  AOI212 U216 ( .A(u_fetch_jmux_i_addr_pc4_15_), .B(n452), .C(n436), .Q(n440)
         );
  AOI212 U217 ( .A(u_fetch_jmux_i_addr_pc4_8_), .B(n452), .C(n471), .Q(n475)
         );
  AOI212 U218 ( .A(u_fetch_jmux_i_addr_pc4_3_), .B(n452), .C(n494), .Q(n498)
         );
  INV12 U219 ( .A(n343), .Q(n256) );
  AOI212 U220 ( .A(n452), .B(u_fetch_jmux_i_addr_pc4_16_), .C(n152), .Q(n435)
         );
  CLKBU15 U221 ( .A(n332), .Q(n253) );
  IMUX20 U222 ( .A(if_addr_j[26]), .B(n320), .S(for_addr_rtM[3]), .Q(n140) );
  IMUX20 U223 ( .A(if_addr_j[25]), .B(n323), .S(for_addr_rtM[2]), .Q(n141) );
  XNR20 U224 ( .A(if_addr_j[27]), .B(for_addr_rtM[4]), .Q(n142) );
  NAND40 U225 ( .A(mem_read), .B(n140), .C(n141), .D(n142), .Q(n143) );
  IMUX20 U226 ( .A(n321), .B(if_addr_j[24]), .S(for_addr_rtM[1]), .Q(n144) );
  IMUX20 U227 ( .A(n309), .B(if_addr_j[23]), .S(for_addr_rtM[0]), .Q(n145) );
  CLKIN0 U228 ( .A(n559), .Q(n146) );
  NOR40 U229 ( .A(n143), .B(n144), .C(n145), .D(n146), .Q(n558) );
  NOR21 U230 ( .A(n280), .B(n345), .Q(n147) );
  AOI211 U231 ( .A(n255), .B(id_data_jr[29]), .C(n147), .Q(n375) );
  CLKIN0 U232 ( .A(add_x_1_n24), .Q(n148) );
  NAND40 U233 ( .A(mem_data_pc4[24]), .B(mem_data_pc4[25]), .C(add_x_1_n34), 
        .D(n148), .Q(add_x_1_n13) );
  NOR21 U234 ( .A(n329), .B(n345), .Q(n149) );
  AOI211 U235 ( .A(n452), .B(u_fetch_jmux_i_addr_pc4_19_), .C(n149), .Q(n424)
         );
  NAND31 U236 ( .A(mem_data_pc4[16]), .B(mem_data_pc4[17]), .C(add_x_1_n71), 
        .Q(n150) );
  NOR30 U237 ( .A(add_x_1_n88), .B(add_x_1_n62), .C(n150), .Q(add_x_1_n50) );
  NOR21 U238 ( .A(n266), .B(n345), .Q(n151) );
  AOI211 U239 ( .A(n452), .B(u_fetch_jmux_i_addr_pc4_17_), .C(n151), .Q(n431)
         );
  NOR21 U240 ( .A(n287), .B(n345), .Q(n152) );
  NOR21 U241 ( .A(n292), .B(n344), .Q(n153) );
  AOI211 U242 ( .A(n452), .B(u_fetch_jmux_i_addr_pc4_10_), .C(n153), .Q(n465)
         );
  NAND20 U243 ( .A(add_x_1_n12), .B(mem_data_pc4[26]), .Q(n154) );
  XNR20 U244 ( .A(mem_data_pc4[27]), .B(n154), .Q(n155) );
  MUX21 U245 ( .A(data_address[27]), .B(n155), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[27]) );
  AOI210 U246 ( .A(u_decode_add_x_16_n124), .B(u_decode_add_x_16_n111), .C(
        u_decode_add_x_16_n112), .Q(n156) );
  OAI212 U247 ( .A(u_decode_add_x_16_n109), .B(u_decode_add_x_16_n135), .C(
        n156), .Q(n157) );
  NOR20 U248 ( .A(u_decode_add_x_16_n134), .B(u_decode_add_x_16_n109), .Q(n158) );
  AOI211 U249 ( .A(n158), .B(u_decode_add_x_16_n156), .C(n157), .Q(
        u_decode_add_x_16_n106) );
  NOR21 U250 ( .A(n285), .B(n344), .Q(n159) );
  AOI211 U251 ( .A(n452), .B(u_fetch_jmux_i_addr_pc4_7_), .C(n159), .Q(n479)
         );
  CLKIN0 U252 ( .A(data_address[26]), .Q(n160) );
  XNR20 U253 ( .A(add_x_1_n12), .B(mem_data_pc4[26]), .Q(n161) );
  IMUX20 U254 ( .A(n160), .B(n161), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[26]) );
  CLKIN0 U255 ( .A(data_address[15]), .Q(n162) );
  NOR20 U256 ( .A(add_x_1_n70), .B(add_x_1_n68), .Q(n163) );
  XNR20 U257 ( .A(mem_data_pc4[15]), .B(n163), .Q(n164) );
  IMUX20 U258 ( .A(n162), .B(n164), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[15]) );
  NOR22 U259 ( .A(n284), .B(n252), .Q(n165) );
  AOI211 U260 ( .A(n257), .B(if_addr_b[2]), .C(n165), .Q(n501) );
  CLKIN0 U261 ( .A(u_decode_add_x_16_n55), .Q(n166) );
  NOR20 U262 ( .A(u_decode_add_x_16_n54), .B(n166), .Q(n167) );
  XNR20 U263 ( .A(u_decode_add_x_16_n56), .B(n167), .Q(
        u_decode_pcadd_o_addr_pcbranchE[26]) );
  CLKIN0 U264 ( .A(u_decode_add_x_16_n131), .Q(n168) );
  AOI210 U265 ( .A(u_decode_add_x_16_n133), .B(u_decode_add_x_16_n208), .C(
        n168), .Q(n169) );
  CLKIN0 U266 ( .A(u_decode_add_x_16_n126), .Q(n170) );
  NOR20 U267 ( .A(u_decode_add_x_16_n125), .B(n170), .Q(n171) );
  XNR20 U268 ( .A(n169), .B(n171), .Q(u_decode_pcadd_o_addr_pcbranchE[15]) );
  NAND20 U269 ( .A(add_x_1_n41), .B(mem_data_pc4[20]), .Q(n172) );
  XNR20 U270 ( .A(mem_data_pc4[21]), .B(n172), .Q(n173) );
  MUX21 U271 ( .A(data_address[21]), .B(n173), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[21]) );
  CLKIN0 U272 ( .A(data_address[13]), .Q(n174) );
  NOR20 U273 ( .A(add_x_1_n79), .B(add_x_1_n78), .Q(n175) );
  XNR20 U274 ( .A(mem_data_pc4[13]), .B(n175), .Q(n176) );
  IMUX20 U275 ( .A(n174), .B(n176), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[13]) );
  NAND20 U276 ( .A(add_x_1_n96), .B(mem_data_pc4[8]), .Q(n177) );
  XNR20 U277 ( .A(mem_data_pc4[9]), .B(n177), .Q(n178) );
  MUX21 U278 ( .A(data_address[9]), .B(n178), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[9]) );
  NOR22 U279 ( .A(n282), .B(n252), .Q(n179) );
  AOI211 U280 ( .A(n452), .B(u_fetch_jmux_i_addr_pc4_6_), .C(n179), .Q(n483)
         );
  NAND30 U281 ( .A(n264), .B(id_data_instr[27]), .C(id_data_instr[28]), .Q(
        n180) );
  OAI210 U282 ( .A(if_addr_j[18]), .B(id_data_instr[28]), .C(n354), .Q(n181)
         );
  AOI210 U283 ( .A(n180), .B(n181), .C(n581), .Q(u_decode_jbcon_o_con_bop[1])
         );
  AOI211 U284 ( .A(u_decode_add_x_16_n38), .B(u_decode_add_x_16_n34), .C(
        u_decode_add_x_16_n35), .Q(n182) );
  CLKIN0 U285 ( .A(u_decode_add_x_16_n32), .Q(n183) );
  NOR20 U286 ( .A(u_decode_add_x_16_n31), .B(n183), .Q(n184) );
  XNR21 U287 ( .A(n182), .B(n184), .Q(u_decode_pcadd_o_addr_pcbranchE[31]) );
  CLKIN0 U288 ( .A(u_decode_add_x_16_n94), .Q(n185) );
  NOR20 U289 ( .A(u_decode_add_x_16_n93), .B(n185), .Q(n186) );
  XNR20 U290 ( .A(u_decode_add_x_16_n95), .B(n186), .Q(
        u_decode_pcadd_o_addr_pcbranchE[20]) );
  CLKIN0 U291 ( .A(u_decode_add_x_16_n144), .Q(n187) );
  AOI210 U292 ( .A(u_decode_add_x_16_n145), .B(u_decode_add_x_16_n210), .C(
        n187), .Q(n188) );
  CLKIN0 U293 ( .A(u_decode_add_x_16_n139), .Q(n189) );
  NOR20 U294 ( .A(u_decode_add_x_16_n138), .B(n189), .Q(n190) );
  XNR20 U295 ( .A(n188), .B(n190), .Q(u_decode_pcadd_o_addr_pcbranchE[13]) );
  CLKIN0 U296 ( .A(u_decode_add_x_16_n165), .Q(n191) );
  NOR20 U297 ( .A(u_decode_add_x_16_n164), .B(n191), .Q(n192) );
  XNR20 U298 ( .A(u_decode_add_x_16_n166), .B(n192), .Q(
        u_decode_pcadd_o_addr_pcbranchE[8]) );
  CLKIN0 U299 ( .A(u_decode_add_x_16_n188), .Q(n193) );
  NOR20 U300 ( .A(u_decode_add_x_16_n187), .B(n193), .Q(n194) );
  XNR20 U301 ( .A(u_decode_add_x_16_n190), .B(n194), .Q(
        u_decode_pcadd_o_addr_pcbranchE[3]) );
  CLKIN0 U302 ( .A(data_address[25]), .Q(n195) );
  NOR20 U303 ( .A(add_x_1_n22), .B(add_x_1_n21), .Q(n196) );
  XNR20 U304 ( .A(mem_data_pc4[25]), .B(n196), .Q(n197) );
  IMUX20 U305 ( .A(n195), .B(n197), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[25]) );
  CLKIN0 U306 ( .A(data_address[20]), .Q(n198) );
  XNR20 U307 ( .A(add_x_1_n41), .B(mem_data_pc4[20]), .Q(n199) );
  IMUX20 U308 ( .A(n198), .B(n199), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[20]) );
  NAND20 U309 ( .A(add_x_1_n87), .B(mem_data_pc4[10]), .Q(n200) );
  XNR20 U310 ( .A(mem_data_pc4[11]), .B(n200), .Q(n201) );
  MUX21 U311 ( .A(data_address[11]), .B(n201), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[11]) );
  CLKIN0 U312 ( .A(data_address[8]), .Q(n202) );
  XNR20 U313 ( .A(add_x_1_n96), .B(mem_data_pc4[8]), .Q(n203) );
  IMUX20 U314 ( .A(n202), .B(n203), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[8]) );
  NAND20 U315 ( .A(add_x_1_n112), .B(mem_data_pc4[4]), .Q(n204) );
  XNR20 U316 ( .A(mem_data_pc4[5]), .B(n204), .Q(n205) );
  MUX21 U317 ( .A(data_address[5]), .B(n205), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[5]) );
  CLKIN0 U318 ( .A(data_address[3]), .Q(n206) );
  XNR20 U319 ( .A(mem_data_pc4[2]), .B(mem_data_pc4[3]), .Q(n207) );
  IMUX20 U320 ( .A(n206), .B(n207), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[3]) );
  CLKIN0 U321 ( .A(add_x_4_n27), .Q(n208) );
  NAND40 U322 ( .A(instruction_address[24]), .B(instruction_address[25]), .C(
        add_x_4_n37), .D(n208), .Q(add_x_4_n16) );
  NOR40 U323 ( .A(n569), .B(n570), .C(n571), .D(n547), .Q(n209) );
  IMUX20 U324 ( .A(n560), .B(if_addr_j[24]), .S(mem_addr_regdst[1]), .Q(n210)
         );
  IMUX20 U325 ( .A(n323), .B(if_addr_j[25]), .S(mem_addr_regdst[2]), .Q(n211)
         );
  NOR30 U326 ( .A(n211), .B(n555), .C(n210), .Q(n212) );
  NAND20 U327 ( .A(n209), .B(n212), .Q(n213) );
  AOI210 U328 ( .A(n557), .B(n213), .C(n558), .Q(u_decode_for_o_con_fa_0_) );
  NAND20 U329 ( .A(n513), .B(n352), .Q(n214) );
  CLKIN0 U330 ( .A(n214), .Q(u_decode_jbcon_o_con_aluPC4) );
  CLKIN0 U331 ( .A(u_decode_add_x_16_n40), .Q(n215) );
  NOR20 U332 ( .A(u_decode_add_x_16_n39), .B(n215), .Q(n216) );
  XNR20 U333 ( .A(u_decode_add_x_16_n41), .B(n216), .Q(
        u_decode_pcadd_o_addr_pcbranchE[29]) );
  CLKIN0 U334 ( .A(u_decode_add_x_16_n104), .Q(n217) );
  AOI210 U335 ( .A(u_decode_add_x_16_n105), .B(u_decode_add_x_16_n204), .C(
        n217), .Q(n218) );
  CLKIN0 U336 ( .A(u_decode_add_x_16_n99), .Q(n219) );
  NOR20 U337 ( .A(u_decode_add_x_16_n98), .B(n219), .Q(n220) );
  XNR20 U338 ( .A(n218), .B(n220), .Q(u_decode_pcadd_o_addr_pcbranchE[19]) );
  CLKIN0 U339 ( .A(u_decode_add_x_16_n119), .Q(n221) );
  AOI210 U340 ( .A(u_decode_add_x_16_n120), .B(u_decode_add_x_16_n206), .C(
        n221), .Q(n222) );
  CLKIN0 U341 ( .A(u_decode_add_x_16_n114), .Q(n223) );
  NOR20 U342 ( .A(u_decode_add_x_16_n113), .B(n223), .Q(n224) );
  XNR20 U343 ( .A(n222), .B(n224), .Q(u_decode_pcadd_o_addr_pcbranchE[17]) );
  CLKIN0 U344 ( .A(u_decode_add_x_16_n154), .Q(n225) );
  NOR20 U345 ( .A(u_decode_add_x_16_n153), .B(n225), .Q(n226) );
  XNR20 U346 ( .A(u_decode_add_x_16_n155), .B(n226), .Q(
        u_decode_pcadd_o_addr_pcbranchE[10]) );
  CLKIN0 U347 ( .A(u_decode_add_x_16_n175), .Q(n227) );
  AOI210 U348 ( .A(u_decode_add_x_16_n176), .B(u_decode_add_x_16_n216), .C(
        n227), .Q(n228) );
  CLKIN0 U349 ( .A(u_decode_add_x_16_n170), .Q(n229) );
  NOR20 U350 ( .A(u_decode_add_x_16_n169), .B(n229), .Q(n230) );
  XNR20 U351 ( .A(n228), .B(n230), .Q(u_decode_pcadd_o_addr_pcbranchE[7]) );
  CLKIN0 U352 ( .A(u_decode_add_x_16_n184), .Q(n231) );
  NOR20 U353 ( .A(u_decode_add_x_16_n183), .B(n231), .Q(n232) );
  XNR20 U354 ( .A(u_decode_add_x_16_n185), .B(n232), .Q(
        u_decode_pcadd_o_addr_pcbranchE[4]) );
  OAI210 U355 ( .A(if_addr_j[2]), .B(id_addr_pc4[2]), .C(
        u_decode_add_x_16_n190), .Q(n233) );
  CLKIN0 U356 ( .A(n233), .Q(u_decode_pcadd_o_addr_pcbranchE[2]) );
  CLKIN0 U357 ( .A(data_address[23]), .Q(n234) );
  NOR20 U358 ( .A(add_x_1_n31), .B(add_x_1_n30), .Q(n235) );
  XNR20 U359 ( .A(mem_data_pc4[23]), .B(n235), .Q(n236) );
  IMUX20 U360 ( .A(n234), .B(n236), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[23]) );
  CLKIN0 U361 ( .A(data_address[19]), .Q(n237) );
  NOR20 U362 ( .A(add_x_1_n49), .B(add_x_1_n48), .Q(n238) );
  XNR20 U363 ( .A(mem_data_pc4[19]), .B(n238), .Q(n239) );
  IMUX20 U364 ( .A(n237), .B(n239), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[19]) );
  CLKIN0 U365 ( .A(data_address[17]), .Q(n240) );
  NOR20 U366 ( .A(add_x_1_n60), .B(add_x_1_n59), .Q(n241) );
  XNR20 U367 ( .A(mem_data_pc4[17]), .B(n241), .Q(n242) );
  IMUX20 U368 ( .A(n240), .B(n242), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[17]) );
  CLKIN0 U369 ( .A(data_address[10]), .Q(n243) );
  XNR20 U370 ( .A(add_x_1_n87), .B(mem_data_pc4[10]), .Q(n244) );
  IMUX20 U371 ( .A(n243), .B(n244), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[10]) );
  CLKIN0 U372 ( .A(data_address[7]), .Q(n245) );
  NOR20 U373 ( .A(add_x_1_n104), .B(add_x_1_n103), .Q(n246) );
  XNR20 U374 ( .A(mem_data_pc4[7]), .B(n246), .Q(n247) );
  IMUX20 U375 ( .A(n245), .B(n247), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[7]) );
  CLKIN0 U376 ( .A(data_address[4]), .Q(n248) );
  XNR20 U377 ( .A(add_x_1_n112), .B(mem_data_pc4[4]), .Q(n249) );
  IMUX20 U378 ( .A(n248), .B(n249), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[4]) );
  CLKIN0 U379 ( .A(data_address[2]), .Q(n250) );
  IMUX20 U380 ( .A(n250), .B(mem_data_pc4[2]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[2]) );
  NAND28 U381 ( .A(n426), .B(n359), .Q(n344) );
  NAND20 U382 ( .A(n338), .B(n508), .Q(n511) );
  NOR21 U383 ( .A(n279), .B(n252), .Q(n367) );
  NOR21 U384 ( .A(n320), .B(n252), .Q(n386) );
  NOR21 U385 ( .A(n323), .B(n252), .Q(n391) );
  INV3 U386 ( .A(n260), .Q(n259) );
  INV15 U387 ( .A(n343), .Q(n255) );
  NAND23 U388 ( .A(n258), .B(n427), .Q(n119) );
  NAND33 U389 ( .A(n410), .B(n409), .C(n408), .Q(n115) );
  AOI212 U390 ( .A(id_data_jr[22]), .B(n256), .C(n406), .Q(n410) );
  NAND33 U391 ( .A(n405), .B(n404), .C(n403), .Q(n114) );
  AOI212 U392 ( .A(id_data_jr[23]), .B(n256), .C(n401), .Q(n405) );
  NAND33 U393 ( .A(n380), .B(n379), .C(n378), .Q(n109) );
  AOI212 U394 ( .A(id_data_jr[28]), .B(n256), .C(n376), .Q(n380) );
  NAND33 U395 ( .A(n400), .B(n399), .C(n398), .Q(n113) );
  NAND33 U396 ( .A(n375), .B(n373), .C(n374), .Q(n108) );
  NAND33 U397 ( .A(n366), .B(n365), .C(n364), .Q(n138) );
  NAND33 U398 ( .A(n385), .B(n384), .C(n383), .Q(n110) );
  NAND33 U399 ( .A(n500), .B(n501), .C(n499), .Q(n135) );
  IMUX21 U400 ( .A(n253), .B(n502), .S(instruction_address[2]), .Q(n500) );
  NAND28 U401 ( .A(n426), .B(n359), .Q(n252) );
  OAI212 U402 ( .A(n502), .B(n452), .C(instruction_address[1]), .Q(n505) );
  INV15 U403 ( .A(n338), .Q(n257) );
  INV15 U404 ( .A(n338), .Q(n254) );
  NAND26 U405 ( .A(if_con_b), .B(n506), .Q(n338) );
  AOI211 U406 ( .A(u_fetch_jmux_i_addr_pc4_4_), .B(n452), .C(n489), .Q(n493)
         );
  AOI211 U407 ( .A(u_fetch_jmux_i_addr_pc4_14_), .B(n452), .C(n441), .Q(n445)
         );
  AOI211 U408 ( .A(u_fetch_jmux_i_addr_pc4_9_), .B(n452), .C(n466), .Q(n470)
         );
  AOI211 U409 ( .A(u_fetch_jmux_i_addr_pc4_21_), .B(n452), .C(n411), .Q(n415)
         );
  AOI211 U410 ( .A(u_fetch_jmux_i_addr_pc4_11_), .B(n452), .C(n457), .Q(n461)
         );
  INV15 U411 ( .A(if_con_b), .Q(n426) );
  NAND33 U412 ( .A(n475), .B(n474), .C(n473), .Q(n129) );
  NAND33 U413 ( .A(n479), .B(n478), .C(n477), .Q(n130) );
  INV15 U414 ( .A(n339), .Q(n452) );
  NAND26 U415 ( .A(n426), .B(n340), .Q(n339) );
  NOR33 U416 ( .A(id_data_instr[29]), .B(id_data_instr[31]), .C(
        id_data_instr[30]), .Q(n513) );
  NAND28 U417 ( .A(n426), .B(n263), .Q(n343) );
  NAND33 U418 ( .A(n498), .B(n497), .C(n496), .Q(n134) );
  NAND33 U419 ( .A(n465), .B(n464), .C(n463), .Q(n127) );
  NAND33 U420 ( .A(n435), .B(n434), .C(n433), .Q(n121) );
  NAND33 U421 ( .A(n424), .B(n423), .C(n422), .Q(n118) );
  NAND28 U422 ( .A(n426), .B(n359), .Q(n345) );
  AOI212 U423 ( .A(id_data_jr[30]), .B(n256), .C(n367), .Q(n371) );
  AOI212 U424 ( .A(id_data_jr[25]), .B(n255), .C(n391), .Q(n395) );
  NAND33 U425 ( .A(n493), .B(n492), .C(n491), .Q(n133) );
  NOR22 U426 ( .A(n283), .B(n252), .Q(n484) );
  NOR22 U427 ( .A(n330), .B(n252), .Q(n416) );
  NAND33 U428 ( .A(n390), .B(n389), .C(n388), .Q(n111) );
  AOI212 U429 ( .A(id_data_jr[26]), .B(n255), .C(n386), .Q(n390) );
  NAND33 U430 ( .A(n482), .B(n483), .C(n481), .Q(n131) );
  NAND33 U431 ( .A(n450), .B(n449), .C(n448), .Q(n124) );
  NAND33 U432 ( .A(n440), .B(n439), .C(n438), .Q(n122) );
  NAND33 U433 ( .A(n445), .B(n444), .C(n443), .Q(n123) );
  NAND33 U434 ( .A(n431), .B(n430), .C(n429), .Q(n120) );
  NAND33 U435 ( .A(n470), .B(n469), .C(n468), .Q(n128) );
  NAND33 U436 ( .A(n415), .B(n414), .C(n413), .Q(n116) );
  AOI2112 U437 ( .A(n255), .B(id_data_jr[18]), .C(n261), .D(n259), .Q(n258) );
  NOR22 U438 ( .A(n291), .B(n252), .Q(n457) );
  NOR22 U439 ( .A(n286), .B(n252), .Q(n451) );
  OAI212 U440 ( .A(n344), .B(n251), .C(n262), .Q(n261) );
  NAND22 U441 ( .A(n254), .B(if_addr_b[17]), .Q(n429) );
  NAND21 U442 ( .A(n257), .B(if_addr_b[9]), .Q(n468) );
  NAND21 U443 ( .A(n254), .B(if_addr_b[15]), .Q(n438) );
  NAND21 U444 ( .A(n257), .B(if_addr_b[16]), .Q(n433) );
  NAND21 U445 ( .A(n254), .B(if_addr_b[14]), .Q(n443) );
  NAND21 U446 ( .A(n257), .B(if_addr_b[4]), .Q(n491) );
  NAND21 U447 ( .A(n257), .B(if_addr_b[13]), .Q(n448) );
  NAND22 U448 ( .A(n257), .B(if_addr_b[12]), .Q(n454) );
  NAND22 U449 ( .A(n257), .B(if_addr_b[5]), .Q(n486) );
  NAND21 U450 ( .A(n254), .B(if_addr_b[7]), .Q(n477) );
  NAND21 U451 ( .A(n257), .B(if_addr_b[10]), .Q(n463) );
  NAND22 U452 ( .A(n254), .B(if_addr_b[20]), .Q(n418) );
  MUX21 U453 ( .A(data_address[30]), .B(u_mem_pc8[30]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[30]) );
  INV3 U454 ( .A(n362), .Q(n356) );
  INV2 U455 ( .A(u_decode_add_x_16_n86), .Q(u_decode_add_x_16_n84) );
  OAI210 U456 ( .A(n268), .B(n583), .C(n584), .Q(
        u_decode_control_o_con_memread) );
  INV1 U457 ( .A(u_decode_control_o_con_aluop_5_), .Q(n587) );
  INV1 U458 ( .A(u_decode_add_x_16_n124), .Q(u_decode_add_x_16_n122) );
  INV2 U459 ( .A(u_decode_add_x_16_n69), .Q(u_decode_add_x_16_n67) );
  INV3 U460 ( .A(n588), .Q(n586) );
  INV2 U461 ( .A(mem_data_pc4[24]), .Q(add_x_1_n21) );
  NAND21 U462 ( .A(n254), .B(if_addr_b[11]), .Q(n459) );
  NOR21 U463 ( .A(n502), .B(n363), .Q(n359) );
  INV2 U464 ( .A(add_x_4_n91), .Q(add_x_4_n90) );
  INV3 U465 ( .A(n352), .Q(n350) );
  NOR21 U466 ( .A(n355), .B(n581), .Q(n502) );
  INV1 U467 ( .A(u_decode_add_x_16_n149), .Q(u_decode_add_x_16_n147) );
  INV1 U468 ( .A(add_x_4_n65), .Q(add_x_4_n64) );
  INV2 U469 ( .A(add_x_4_n27), .Q(add_x_4_n26) );
  INV1 U470 ( .A(add_x_1_n62), .Q(add_x_1_n61) );
  INV3 U471 ( .A(mem_con_Wregwrite), .Q(n547) );
  NAND21 U472 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_23_), .Q(n403) );
  NAND21 U473 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_25_), .Q(n393) );
  NAND21 U474 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_27_), .Q(n383) );
  NAND21 U475 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_26_), .Q(n388) );
  NAND21 U476 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_22_), .Q(n408) );
  NAND21 U477 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_24_), .Q(n398) );
  NAND21 U478 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_30_), .Q(n369) );
  NAND21 U479 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_31_), .Q(n364) );
  NOR22 U480 ( .A(n507), .B(if_con_b), .Q(n332) );
  INV2 U481 ( .A(n507), .Q(n340) );
  CLKIN3 U482 ( .A(add_x_1_n32), .Q(add_x_1_n31) );
  NAND31 U483 ( .A(n363), .B(n362), .C(n506), .Q(n507) );
  INV2 U484 ( .A(u_decode_add_x_16_n87), .Q(u_decode_add_x_16_n85) );
  INV2 U485 ( .A(u_decode_add_x_16_n74), .Q(u_decode_add_x_16_n72) );
  INV2 U486 ( .A(add_x_1_n88), .Q(add_x_1_n87) );
  INV6 U487 ( .A(n502), .Q(n506) );
  INV1 U488 ( .A(u_decode_add_x_16_n51), .Q(u_decode_add_x_16_n195) );
  INV1 U489 ( .A(u_decode_add_x_16_n123), .Q(u_decode_add_x_16_n121) );
  INV1 U490 ( .A(u_decode_add_x_16_n148), .Q(u_decode_add_x_16_n146) );
  INV2 U491 ( .A(add_x_1_n24), .Q(add_x_1_n23) );
  NOR21 U492 ( .A(n517), .B(id_data_instr[28]), .Q(n352) );
  INV2 U493 ( .A(mem_addr_regdst[4]), .Q(n331) );
  NAND21 U494 ( .A(n253), .B(u_fetch_jmux_i_addr_pc4_29_), .Q(n373) );
  MUX21 U495 ( .A(data_address[31]), .B(u_mem_pc8[31]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[31]) );
  MUX21 U496 ( .A(data_address[28]), .B(u_mem_pc8[28]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[28]) );
  CLKIN3 U497 ( .A(add_x_4_n35), .Q(add_x_4_n34) );
  INV2 U498 ( .A(n524), .Q(n526) );
  NAND31 U499 ( .A(for_FWmemread), .B(n548), .C(n549), .Q(n524) );
  NOR40 U500 ( .A(n550), .B(n551), .C(n552), .D(n553), .Q(n548) );
  INV2 U501 ( .A(add_x_4_n108), .Q(add_x_4_n107) );
  INV1 U502 ( .A(u_decode_add_x_16_n75), .Q(u_decode_add_x_16_n199) );
  INV1 U503 ( .A(u_decode_add_x_16_n63), .Q(u_decode_add_x_16_n197) );
  INV1 U504 ( .A(add_x_4_n84), .Q(add_x_4_n83) );
  NOR21 U505 ( .A(n264), .B(id_data_instr[27]), .Q(n354) );
  BUF6 U506 ( .A(if_addr_j[17]), .Q(n346) );
  NAND21 U507 ( .A(id_data_jr[0]), .B(n256), .Q(n509) );
  NAND21 U508 ( .A(id_data_jr[1]), .B(n255), .Q(n504) );
  NAND21 U509 ( .A(n257), .B(ex_data_pc4[0]), .Q(n510) );
  MUX21 U510 ( .A(data_address[16]), .B(u_mem_pc8[16]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[16]) );
  INV3 U511 ( .A(add_x_4_n53), .Q(add_x_4_n52) );
  INV2 U512 ( .A(u_decode_add_x_16_n177), .Q(u_decode_add_x_16_n176) );
  INV2 U513 ( .A(u_decode_add_x_16_n68), .Q(u_decode_add_x_16_n66) );
  INV1 U514 ( .A(u_decode_add_x_16_n90), .Q(u_decode_add_x_16_n201) );
  INV2 U515 ( .A(u_decode_add_x_16_n186), .Q(u_decode_add_x_16_n185) );
  INV1 U516 ( .A(add_x_1_n81), .Q(add_x_1_n80) );
  NOR21 U517 ( .A(id_data_instr[28]), .B(n354), .Q(n355) );
  INV3 U518 ( .A(n513), .Q(n581) );
  INV2 U519 ( .A(mem_data_pc4[16]), .Q(add_x_1_n59) );
  INV2 U520 ( .A(mem_data_pc4[22]), .Q(add_x_1_n30) );
  INV3 U521 ( .A(n357), .Q(n263) );
  MUX21 U522 ( .A(data_address[14]), .B(u_mem_pc8[14]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[14]) );
  INV3 U523 ( .A(u_decode_add_x_16_n106), .Q(u_decode_add_x_16_n105) );
  MUX21 U524 ( .A(data_address[18]), .B(u_mem_pc8[18]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[18]) );
  MUX21 U525 ( .A(data_address[12]), .B(u_mem_pc8[12]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[12]) );
  INV2 U526 ( .A(if_con_j[1]), .Q(n358) );
  INV2 U527 ( .A(u_decode_add_x_16_n103), .Q(u_decode_add_x_16_n204) );
  INV2 U528 ( .A(add_x_1_n105), .Q(add_x_1_n104) );
  INV2 U529 ( .A(u_decode_add_x_16_n81), .Q(u_decode_add_x_16_n79) );
  INV2 U530 ( .A(add_x_4_n37), .Q(add_x_4_n36) );
  INV1 U531 ( .A(u_decode_add_x_16_n150), .Q(u_decode_add_x_16_n211) );
  INV1 U532 ( .A(u_decode_add_x_16_n180), .Q(u_decode_add_x_16_n217) );
  INV1 U533 ( .A(u_decode_add_x_16_n161), .Q(u_decode_add_x_16_n213) );
  NAND22 U534 ( .A(n356), .B(n506), .Q(n357) );
  INV2 U535 ( .A(n555), .Q(n554) );
  OAI210 U536 ( .A(n585), .B(n586), .C(n515), .Q(
        u_decode_control_o_con_aluop_3_) );
  NOR21 U537 ( .A(n333), .B(n564), .Q(n555) );
  NAND22 U538 ( .A(n353), .B(if_con_j[1]), .Q(n362) );
  NOR20 U539 ( .A(n312), .B(n506), .Q(n407) );
  INV3 U540 ( .A(u_decode_add_x_16_n156), .Q(u_decode_add_x_16_n155) );
  INV3 U541 ( .A(add_x_1_n50), .Q(add_x_1_n49) );
  AOI211 U542 ( .A(n583), .B(n348), .C(n268), .Q(
        u_decode_control_o_con_aluop_4_) );
  NAND22 U543 ( .A(n358), .B(if_con_j[0]), .Q(n363) );
  NOR21 U544 ( .A(n296), .B(n506), .Q(n382) );
  INV2 U545 ( .A(u_decode_add_x_16_n80), .Q(u_decode_add_x_16_n78) );
  INV2 U546 ( .A(mem_data_pc4[12]), .Q(add_x_1_n78) );
  AOI211 U547 ( .A(n254), .B(if_addr_b[25]), .C(n392), .Q(n394) );
  AOI211 U548 ( .A(n257), .B(if_addr_b[31]), .C(n361), .Q(n365) );
  AOI211 U549 ( .A(n254), .B(if_addr_b[30]), .C(n368), .Q(n370) );
  AOI211 U550 ( .A(n254), .B(if_addr_b[28]), .C(n377), .Q(n379) );
  AOI211 U551 ( .A(n257), .B(if_addr_b[22]), .C(n407), .Q(n409) );
  NOR21 U552 ( .A(n271), .B(n506), .Q(n387) );
  NOR21 U553 ( .A(n298), .B(n506), .Q(n402) );
  NOR20 U554 ( .A(n311), .B(n506), .Q(n397) );
  INV2 U555 ( .A(u_decode_add_x_16_n73), .Q(u_decode_add_x_16_n71) );
  OAI211 U556 ( .A(for_o_addr_Erd[2]), .B(n567), .C(n323), .Q(n566) );
  INV2 U557 ( .A(add_x_1_n34), .Q(add_x_1_n33) );
  INV2 U558 ( .A(u_decode_add_x_16_n130), .Q(u_decode_add_x_16_n208) );
  MUX21 U559 ( .A(data_address[0]), .B(u_mem_pc8[0]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[0]) );
  INV2 U560 ( .A(u_decode_add_x_16_n118), .Q(u_decode_add_x_16_n206) );
  MUX21 U561 ( .A(data_address[1]), .B(u_mem_pc8[1]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[1]) );
  INV2 U562 ( .A(u_decode_add_x_16_n143), .Q(u_decode_add_x_16_n210) );
  INV2 U563 ( .A(mem_data_pc4[14]), .Q(add_x_1_n68) );
  AOI211 U564 ( .A(n257), .B(if_addr_b[27]), .C(n382), .Q(n384) );
  AOI211 U565 ( .A(n257), .B(if_addr_b[24]), .C(n397), .Q(n399) );
  INV3 U566 ( .A(u_decode_add_x_16_n133), .Q(u_decode_add_x_16_n132) );
  INV3 U567 ( .A(add_x_4_n73), .Q(add_x_4_n72) );
  NOR20 U568 ( .A(n304), .B(n506), .Q(n458) );
  NOR20 U569 ( .A(n273), .B(n506), .Q(n462) );
  NOR20 U570 ( .A(n307), .B(n506), .Q(n485) );
  NOR20 U571 ( .A(n306), .B(n506), .Q(n476) );
  NOR20 U572 ( .A(n275), .B(n506), .Q(n490) );
  NOR20 U573 ( .A(n303), .B(n506), .Q(n447) );
  NOR20 U574 ( .A(n302), .B(n506), .Q(n437) );
  NOR20 U575 ( .A(n274), .B(n506), .Q(n472) );
  NOR20 U576 ( .A(n318), .B(n506), .Q(n495) );
  NOR20 U577 ( .A(n305), .B(n506), .Q(n467) );
  NOR20 U578 ( .A(n272), .B(n506), .Q(n417) );
  NOR20 U579 ( .A(n300), .B(n506), .Q(n421) );
  NOR20 U580 ( .A(n299), .B(n506), .Q(n412) );
  OAI210 U581 ( .A(n354), .B(n586), .C(n587), .Q(
        u_decode_control_o_con_aluop_2_) );
  NOR20 U582 ( .A(n301), .B(n506), .Q(n428) );
  NOR40 U583 ( .A(n531), .B(n533), .C(n337), .D(n532), .Q(n336) );
  NOR40 U584 ( .A(n576), .B(n577), .C(n578), .D(n579), .Q(n573) );
  IMUX21 U585 ( .A(if_addr_j[22]), .B(n277), .S(for_addr_rtW[4]), .Q(n549) );
  AOI211 U586 ( .A(n256), .B(id_data_jr[3]), .C(n495), .Q(n497) );
  AOI211 U587 ( .A(n255), .B(id_data_jr[16]), .C(n432), .Q(n434) );
  AOI211 U588 ( .A(n255), .B(id_data_jr[8]), .C(n472), .Q(n474) );
  AOI211 U589 ( .A(n256), .B(id_data_jr[6]), .C(n480), .Q(n482) );
  AOI211 U590 ( .A(n256), .B(id_data_jr[9]), .C(n467), .Q(n469) );
  AOI211 U591 ( .A(n255), .B(id_data_jr[13]), .C(n447), .Q(n449) );
  AOI211 U592 ( .A(n255), .B(id_data_jr[17]), .C(n428), .Q(n430) );
  AOI211 U593 ( .A(n255), .B(id_data_jr[14]), .C(n442), .Q(n444) );
  AOI211 U594 ( .A(n256), .B(id_data_jr[5]), .C(n485), .Q(n487) );
  AOI211 U595 ( .A(n255), .B(id_data_jr[10]), .C(n462), .Q(n464) );
  AOI211 U596 ( .A(n255), .B(id_data_jr[20]), .C(n417), .Q(n419) );
  AOI211 U597 ( .A(n256), .B(id_data_jr[21]), .C(n412), .Q(n414) );
  AOI211 U598 ( .A(n256), .B(id_data_jr[4]), .C(n490), .Q(n492) );
  AOI211 U599 ( .A(n255), .B(id_data_jr[19]), .C(n421), .Q(n423) );
  AOI211 U600 ( .A(n255), .B(id_data_jr[7]), .C(n476), .Q(n478) );
  AOI211 U601 ( .A(n255), .B(id_data_jr[15]), .C(n437), .Q(n439) );
  AOI211 U602 ( .A(n255), .B(id_data_jr[11]), .C(n458), .Q(n460) );
  AOI211 U603 ( .A(n257), .B(if_addr_b[23]), .C(n402), .Q(n404) );
  AOI211 U604 ( .A(n257), .B(if_addr_b[26]), .C(n387), .Q(n389) );
  AOI211 U605 ( .A(n254), .B(if_addr_b[29]), .C(n372), .Q(n374) );
  NOR21 U606 ( .A(n554), .B(u_decode_for_o_con_fa_2_), .Q(
        u_decode_for_o_con_fa_1_) );
  AOI211 U607 ( .A(n528), .B(n524), .C(n523), .Q(u_decode_for_o_con_fb[0]) );
  NAND41 U608 ( .A(for_FWmemread), .B(n573), .C(n574), .D(n559), .Q(n557) );
  IMUX21 U609 ( .A(if_addr_j[20]), .B(n330), .S(for_o_addr_Erd[2]), .Q(n539)
         );
  IMUX21 U610 ( .A(n251), .B(if_addr_j[18]), .S(for_addr_rtW[0]), .Q(n553) );
  INV2 U611 ( .A(add_x_4_n116), .Q(add_x_4_n115) );
  INV3 U612 ( .A(n516), .Q(n582) );
  AOI311 U613 ( .A(if_addr_j[5]), .B(n522), .C(n285), .D(id_data_instr[26]), 
        .Q(n521) );
  INV2 U614 ( .A(mem_data_pc4[18]), .Q(add_x_1_n48) );
  NAND22 U615 ( .A(id_data_instr[26]), .B(id_data_instr[27]), .Q(n517) );
  NAND31 U616 ( .A(n505), .B(n504), .C(n503), .Q(n136) );
  AOI211 U617 ( .A(n256), .B(id_data_jr[12]), .C(n453), .Q(n455) );
  AOI211 U618 ( .A(n514), .B(n515), .C(n266), .Q(u_decode_n1) );
  NOR21 U619 ( .A(n297), .B(n506), .Q(n392) );
  IMUX21 U620 ( .A(n329), .B(if_addr_j[19]), .S(for_addr_rtW[1]), .Q(n552) );
  NAND31 U621 ( .A(n509), .B(n510), .C(n511), .Q(n137) );
  AOI211 U622 ( .A(u_fetch_jmux_i_addr_pc4_12_), .B(n452), .C(n451), .Q(n456)
         );
  AOI211 U623 ( .A(u_fetch_jmux_i_addr_pc4_5_), .B(n452), .C(n484), .Q(n488)
         );
  NOR21 U624 ( .A(n309), .B(n344), .Q(n401) );
  MUX22 U625 ( .A(data_address[29]), .B(u_mem_pc8[29]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[29]) );
  OAI211 U626 ( .A(n523), .B(n524), .C(n525), .Q(u_decode_for_o_con_fb[2]) );
  INV2 U627 ( .A(n425), .Q(n262) );
  NOR21 U628 ( .A(n295), .B(n506), .Q(n372) );
  INV2 U629 ( .A(n558), .Q(n556) );
  INV2 U630 ( .A(n351), .Q(u_decode_control_o_con_regwrite) );
  AOI211 U631 ( .A(n350), .B(n342), .C(n349), .Q(n512) );
  OAI211 U632 ( .A(n350), .B(n349), .C(n582), .Q(u_decode_control_o_con_alusrc) );
  NOR21 U633 ( .A(id_data_instr[31]), .B(n582), .Q(
        u_decode_control_o_con_aluop_0_) );
  NOR21 U634 ( .A(n269), .B(n582), .Q(u_decode_control_o_con_memwrite) );
  INV2 U635 ( .A(add_x_1_n113), .Q(add_x_1_n112) );
  NAND21 U636 ( .A(id_data_instr[26]), .B(n588), .Q(n583) );
  INV2 U637 ( .A(u_decode_add_x_16_n174), .Q(u_decode_add_x_16_n216) );
  XNR20 U638 ( .A(n331), .B(if_addr_j[27]), .Q(n571) );
  NAND21 U639 ( .A(n310), .B(id_data_instr[31]), .Q(n349) );
  INV2 U640 ( .A(mem_data_pc4[6]), .Q(add_x_1_n103) );
  NOR21 U641 ( .A(n342), .B(id_data_instr[30]), .Q(n516) );
  NOR21 U642 ( .A(n293), .B(n344), .Q(n466) );
  NAND31 U643 ( .A(n264), .B(n270), .C(u_decode_control_o_con_aluop_0_), .Q(
        n348) );
  NAND22 U644 ( .A(n534), .B(n277), .Q(n529) );
  NOR21 U645 ( .A(n322), .B(n506), .Q(n368) );
  NOR21 U646 ( .A(n319), .B(n506), .Q(n361) );
  NOR21 U647 ( .A(id_data_instr[26]), .B(id_data_instr[27]), .Q(n585) );
  NOR21 U648 ( .A(n277), .B(n344), .Q(n406) );
  NOR20 U649 ( .A(n581), .B(n519), .Q(u_decode_control_o_con_regdst) );
  XOR21 U650 ( .A(n308), .B(for_o_addr_Erd[4]), .Q(n568) );
  AOI211 U651 ( .A(u_fetch_jmux_i_addr_pc4_20_), .B(n452), .C(n416), .Q(n420)
         );
  NOR21 U652 ( .A(id_data_instr[27]), .B(n521), .Q(n520) );
  AOI211 U653 ( .A(n580), .B(n352), .C(u_decode_control_o_con_aluop_1_), .Q(
        n351) );
  INV3 U654 ( .A(u_decode_control_o_con_aluop_4_), .Q(n515) );
  NOR40 U655 ( .A(id_data_instr[30]), .B(id_data_instr[31]), .C(n342), .D(n270), .Q(n588) );
  NOR31 U656 ( .A(n523), .B(n527), .C(n526), .Q(u_decode_for_o_con_fb[1]) );
  INV3 U657 ( .A(add_x_1_n70), .Q(add_x_1_n69) );
  INV3 U658 ( .A(add_x_1_n4), .Q(add_x_1_n118) );
  NAND22 U659 ( .A(n336), .B(n529), .Q(n525) );
  NAND31 U660 ( .A(n267), .B(n530), .C(mem_read), .Q(n337) );
  NAND41 U661 ( .A(n535), .B(n527), .C(n536), .D(n537), .Q(n528) );
  NAND31 U662 ( .A(ex_con_Wregwrite), .B(n538), .C(n539), .Q(n527) );
  INV3 U663 ( .A(u_decode_add_x_16_n37), .Q(u_decode_add_x_16_n35) );
  INV3 U664 ( .A(u_decode_add_x_16_n45), .Q(u_decode_add_x_16_n43) );
  NAND22 U665 ( .A(n556), .B(n557), .Q(u_decode_for_o_con_fa_2_) );
  NAND22 U666 ( .A(n575), .B(n308), .Q(n559) );
  OAI2111 U667 ( .A(for_o_addr_Erd[2]), .B(n323), .C(n565), .D(n566), .Q(n564)
         );
  NAND22 U668 ( .A(n335), .B(n334), .Q(n333) );
  NOR21 U669 ( .A(n561), .B(n562), .Q(n334) );
  INV3 U670 ( .A(n563), .Q(n335) );
  NAND22 U671 ( .A(ex_con_Wregwrite), .B(n568), .Q(n563) );
  MUX22 U672 ( .A(mem_data_alures[23]), .B(wb_data_memout[23]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[23]) );
  MUX22 U673 ( .A(mem_data_alures[7]), .B(wb_data_memout[7]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[7]) );
  MUX22 U674 ( .A(mem_data_alures[8]), .B(wb_data_memout[8]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[8]) );
  MUX22 U675 ( .A(mem_data_alures[5]), .B(wb_data_memout[5]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[5]) );
  MUX22 U676 ( .A(mem_data_alures[4]), .B(wb_data_memout[4]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[4]) );
  MUX22 U677 ( .A(mem_data_alures[9]), .B(wb_data_memout[9]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[9]) );
  MUX22 U678 ( .A(mem_data_alures[2]), .B(wb_data_memout[2]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[2]) );
  MUX22 U679 ( .A(mem_data_alures[29]), .B(wb_data_memout[29]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[29]) );
  MUX22 U680 ( .A(mem_data_alures[30]), .B(wb_data_memout[30]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[30]) );
  MUX22 U681 ( .A(mem_data_alures[28]), .B(wb_data_memout[28]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[28]) );
  MUX22 U682 ( .A(mem_data_alures[31]), .B(wb_data_memout[31]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[31]) );
  MUX22 U683 ( .A(mem_data_alures[18]), .B(wb_data_memout[18]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[18]) );
  MUX22 U684 ( .A(mem_data_alures[17]), .B(wb_data_memout[17]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[17]) );
  MUX22 U685 ( .A(mem_data_alures[11]), .B(wb_data_memout[11]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[11]) );
  MUX22 U686 ( .A(mem_data_alures[27]), .B(wb_data_memout[27]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[27]) );
  MUX22 U687 ( .A(mem_data_alures[10]), .B(wb_data_memout[10]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[10]) );
  MUX22 U688 ( .A(mem_data_alures[26]), .B(wb_data_memout[26]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[26]) );
  MUX22 U689 ( .A(mem_data_alures[12]), .B(wb_data_memout[12]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[12]) );
  MUX22 U690 ( .A(mem_data_alures[24]), .B(wb_data_memout[24]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[24]) );
  MUX22 U691 ( .A(mem_data_alures[15]), .B(wb_data_memout[15]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[15]) );
  MUX22 U692 ( .A(mem_data_alures[22]), .B(wb_data_memout[22]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[22]) );
  MUX22 U693 ( .A(mem_data_alures[0]), .B(wb_data_memout[0]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[0]) );
  MUX22 U694 ( .A(mem_data_alures[21]), .B(wb_data_memout[21]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[21]) );
  MUX22 U695 ( .A(mem_data_alures[25]), .B(wb_data_memout[25]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[25]) );
  MUX22 U696 ( .A(mem_data_alures[13]), .B(wb_data_memout[13]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[13]) );
  MUX22 U697 ( .A(mem_data_alures[20]), .B(wb_data_memout[20]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[20]) );
  MUX22 U698 ( .A(mem_data_alures[19]), .B(wb_data_memout[19]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[19]) );
  MUX22 U699 ( .A(mem_data_alures[3]), .B(wb_data_memout[3]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[3]) );
  MUX22 U700 ( .A(mem_data_alures[6]), .B(wb_data_memout[6]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[6]) );
  MUX22 U701 ( .A(mem_data_alures[1]), .B(wb_data_memout[1]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[1]) );
  MUX22 U702 ( .A(mem_data_alures[16]), .B(wb_data_memout[16]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[16]) );
  MUX22 U703 ( .A(mem_data_alures[14]), .B(wb_data_memout[14]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[14]) );
  NOR21 U704 ( .A(n326), .B(n344), .Q(n489) );
  NAND22 U705 ( .A(n257), .B(ex_data_pc4[1]), .Q(n503) );
  NAND22 U706 ( .A(n257), .B(if_addr_b[21]), .Q(n413) );
  NOR21 U707 ( .A(n325), .B(n344), .Q(n411) );
  NAND22 U708 ( .A(n254), .B(if_addr_b[8]), .Q(n473) );
  NOR21 U709 ( .A(n294), .B(n345), .Q(n471) );
  NAND22 U710 ( .A(n254), .B(if_addr_b[3]), .Q(n496) );
  NOR21 U711 ( .A(n327), .B(n345), .Q(n494) );
  NAND22 U712 ( .A(n257), .B(if_addr_b[6]), .Q(n481) );
  NAND22 U713 ( .A(n254), .B(if_addr_b[19]), .Q(n422) );
  NOR21 U714 ( .A(n308), .B(n345), .Q(n381) );
  NOR21 U715 ( .A(n321), .B(n345), .Q(n396) );
  NAND22 U716 ( .A(n255), .B(id_data_jr[2]), .Q(n499) );
  NOR21 U717 ( .A(n281), .B(n344), .Q(n376) );
  NOR21 U718 ( .A(n278), .B(n345), .Q(n360) );
  NOR21 U719 ( .A(n289), .B(n344), .Q(n441) );
  NOR21 U720 ( .A(n290), .B(n345), .Q(n446) );
  NAND22 U721 ( .A(n257), .B(if_addr_b[18]), .Q(n427) );
  NOR21 U722 ( .A(n288), .B(n345), .Q(n436) );
  INV3 U723 ( .A(if_con_j[0]), .Q(n353) );
  OAI212 U724 ( .A(id_data_instr[28]), .B(n520), .C(n513), .Q(if_con_j[0]) );
  NOR20 U725 ( .A(id_data_instr[30]), .B(id_data_instr[29]), .Q(n580) );
  MUX21 U726 ( .A(data_address[24]), .B(u_mem_pc8[24]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[24]) );
  MUX21 U727 ( .A(data_address[22]), .B(u_mem_pc8[22]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[22]) );
  MUX21 U728 ( .A(data_address[6]), .B(u_mem_pc8[6]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[6]) );
  NAND22 U729 ( .A(n513), .B(n519), .Q(if_con_j[1]) );
  NAND22 U730 ( .A(n585), .B(n270), .Q(n519) );
  AOI2110 U731 ( .A(id_data_instr[28]), .B(id_data_instr[26]), .C(n347), .D(
        n581), .Q(u_decode_jbcon_o_con_bop[0]) );
  AOI210 U732 ( .A(n354), .B(n251), .C(id_data_instr[28]), .Q(n347) );
  NAND30 U733 ( .A(n352), .B(id_data_instr[31]), .C(n580), .Q(n584) );
  INV3 U734 ( .A(u_decode_add_x_16_n83), .Q(u_decode_add_x_16_n82) );
  NAND22 U735 ( .A(n525), .B(n529), .Q(n523) );
  MUX21 U736 ( .A(n325), .B(if_addr_j[21]), .S(for_addr_rtM[3]), .Q(n267) );
  INV3 U737 ( .A(u_decode_add_x_16_n36), .Q(u_decode_add_x_16_n34) );
  INV3 U738 ( .A(u_decode_add_x_16_n44), .Q(u_decode_add_x_16_n42) );
  XNR21 U739 ( .A(n265), .B(if_addr_j[27]), .Q(n578) );
  NOR40 U740 ( .A(for_o_addr_Erd[1]), .B(for_o_addr_Erd[3]), .C(
        for_o_addr_Erd[0]), .D(if_addr_j[27]), .Q(n567) );
  AOI210 U741 ( .A(n507), .B(n506), .C(n328), .Q(n508) );
  NOR20 U742 ( .A(n317), .B(n506), .Q(n480) );
  NOR20 U743 ( .A(n324), .B(n506), .Q(n377) );
  INV3 U744 ( .A(add_x_4_n2), .Q(add_x_4_n121) );
  NOR20 U745 ( .A(n316), .B(n506), .Q(n453) );
  NOR20 U746 ( .A(n315), .B(n506), .Q(n442) );
  NOR20 U747 ( .A(n313), .B(n506), .Q(n425) );
  NOR20 U748 ( .A(n314), .B(n506), .Q(n432) );
  LOGIC0 U749 ( .Q(n341) );
  AOI310 U750 ( .A(n516), .B(n270), .C(n517), .D(n512), .Q(n514) );
  AOI210 U751 ( .A(n270), .B(id_data_instr[27]), .C(n518), .Q(u_decode_n6) );
  OAI2110 U752 ( .A(n270), .B(id_data_instr[27]), .C(n513), .D(
        id_data_instr[26]), .Q(n518) );
  NOR40 U753 ( .A(if_addr_j[2]), .B(if_addr_j[3]), .C(if_addr_j[4]), .D(
        if_addr_j[6]), .Q(n522) );
  IMUX20 U754 ( .A(if_addr_j[20]), .B(n330), .S(for_addr_rtM[2]), .Q(n530) );
  IMUX20 U755 ( .A(n329), .B(if_addr_j[19]), .S(for_addr_rtM[1]), .Q(n533) );
  IMUX20 U756 ( .A(n277), .B(if_addr_j[22]), .S(for_addr_rtM[4]), .Q(n532) );
  IMUX20 U757 ( .A(n251), .B(if_addr_j[18]), .S(for_addr_rtM[0]), .Q(n531) );
  NOR40 U758 ( .A(if_addr_j[19]), .B(if_addr_j[21]), .C(if_addr_j[18]), .D(
        if_addr_j[20]), .Q(n534) );
  IMUX20 U759 ( .A(if_addr_j[18]), .B(n251), .S(mem_addr_regdst[0]), .Q(n537)
         );
  IMUX20 U760 ( .A(if_addr_j[19]), .B(n329), .S(mem_addr_regdst[1]), .Q(n536)
         );
  NOR40 U761 ( .A(n540), .B(n541), .C(n542), .D(n543), .Q(n538) );
  IMUX20 U762 ( .A(n251), .B(if_addr_j[18]), .S(for_o_addr_Erd[0]), .Q(n543)
         );
  IMUX20 U763 ( .A(n325), .B(if_addr_j[21]), .S(for_o_addr_Erd[3]), .Q(n542)
         );
  IMUX20 U764 ( .A(n329), .B(if_addr_j[19]), .S(for_o_addr_Erd[1]), .Q(n541)
         );
  IMUX20 U765 ( .A(n277), .B(if_addr_j[22]), .S(for_o_addr_Erd[4]), .Q(n540)
         );
  NOR40 U766 ( .A(n544), .B(n545), .C(n546), .D(n547), .Q(n535) );
  IMUX20 U767 ( .A(n325), .B(if_addr_j[21]), .S(mem_addr_regdst[3]), .Q(n546)
         );
  IMUX20 U768 ( .A(n330), .B(if_addr_j[20]), .S(mem_addr_regdst[2]), .Q(n545)
         );
  IMUX20 U769 ( .A(n277), .B(if_addr_j[22]), .S(mem_addr_regdst[4]), .Q(n544)
         );
  IMUX20 U770 ( .A(n330), .B(if_addr_j[20]), .S(for_addr_rtW[2]), .Q(n551) );
  IMUX20 U771 ( .A(n325), .B(if_addr_j[21]), .S(for_addr_rtW[3]), .Q(n550) );
  IMUX20 U772 ( .A(if_addr_j[23]), .B(n309), .S(for_o_addr_Erd[0]), .Q(n565)
         );
  IMUX20 U773 ( .A(n320), .B(if_addr_j[26]), .S(for_o_addr_Erd[3]), .Q(n562)
         );
  IMUX20 U774 ( .A(n321), .B(if_addr_j[24]), .S(for_o_addr_Erd[1]), .Q(n561)
         );
  IMUX20 U775 ( .A(n320), .B(if_addr_j[26]), .S(mem_addr_regdst[3]), .Q(n570)
         );
  IMUX20 U776 ( .A(n309), .B(if_addr_j[23]), .S(mem_addr_regdst[0]), .Q(n569)
         );
  NOR20 U777 ( .A(if_addr_j[24]), .B(n572), .Q(n560) );
  NOR40 U778 ( .A(mem_addr_regdst[0]), .B(mem_addr_regdst[4]), .C(
        mem_addr_regdst[2]), .D(mem_addr_regdst[3]), .Q(n572) );
  NOR40 U779 ( .A(if_addr_j[23]), .B(if_addr_j[25]), .C(if_addr_j[26]), .D(
        if_addr_j[24]), .Q(n575) );
  IMUX20 U780 ( .A(if_addr_j[26]), .B(n320), .S(for_addr_rtW[3]), .Q(n574) );
  IMUX20 U781 ( .A(n323), .B(if_addr_j[25]), .S(for_addr_rtW[2]), .Q(n579) );
  IMUX20 U782 ( .A(n309), .B(if_addr_j[23]), .S(for_addr_rtW[0]), .Q(n577) );
  IMUX20 U783 ( .A(n321), .B(if_addr_j[24]), .S(for_addr_rtW[1]), .Q(n576) );
  AOI2110 U784 ( .A(n342), .B(n519), .C(id_data_instr[30]), .D(
        id_data_instr[31]), .Q(u_decode_control_o_con_aluop_1_) );
  NOR40 U785 ( .A(id_data_instr[28]), .B(id_data_instr[31]), .C(n517), .D(n582), .Q(u_decode_control_o_con_aluop_5_) );
endmodule

