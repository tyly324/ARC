// Verilog simulation library for c35_IOLIBC_ANA_3B_4M
// Owner: austriamicrosystems AG  HIT-Kit: Digital
module APRIO1K5C_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO200C_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO50C_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module APRIO500C_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module AVSUBC_3B (A);
  input A ;
endmodule
module APRIOWC_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
module AGNDALLC_3B (A);
  input A ;
endmodule
module AVDDALLC_3B (A);
  input A ;
endmodule
module APRIOC_3B (PAD,Z);
  inout PAD ;
  inout Z ;
endmodule
