
module F_jumpmux ( i_addr_j, i_addr_jr, i_addr_pc4, i_con_jump, o_addr_jumpmux
 );
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [31:0] i_addr_pc4;
  input [1:0] i_con_jump;
  output [31:0] o_addr_jumpmux;
  wire   n3, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n23,
         n24, n45, n46, n67, n68, n1, n2, n5, n6, n19, n20, n21, n22, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n69, n70, n71, n72,
         n73, n74, n75, n76, n77;

  NAND22 U1 ( .A(n66), .B(n65), .Q(o_addr_jumpmux[28]) );
  BUF6 U2 ( .A(n75), .Q(n1) );
  AOI221 U3 ( .A(i_addr_pc4[3]), .B(n6), .C(i_addr_jr[3]), .D(n75), .Q(n17) );
  NAND22 U4 ( .A(n62), .B(n61), .Q(o_addr_jumpmux[26]) );
  NAND22 U5 ( .A(n11), .B(n12), .Q(o_addr_jumpmux[6]) );
  AOI221 U6 ( .A(i_addr_pc4[6]), .B(n5), .C(i_addr_jr[6]), .D(n75), .Q(n11) );
  NAND22 U7 ( .A(n34), .B(n33), .Q(o_addr_jumpmux[13]) );
  NAND22 U8 ( .A(i_addr_jr[13]), .B(n75), .Q(n33) );
  NAND22 U9 ( .A(n48), .B(n47), .Q(o_addr_jumpmux[19]) );
  NAND22 U10 ( .A(i_addr_jr[19]), .B(n1), .Q(n47) );
  AOI221 U11 ( .A(i_addr_j[22]), .B(n19), .C(i_addr_pc4[22]), .D(n2), .Q(n54)
         );
  AOI221 U12 ( .A(i_addr_j[26]), .B(n19), .C(i_addr_pc4[26]), .D(n5), .Q(n62)
         );
  AOI221 U13 ( .A(i_addr_j[31]), .B(n20), .C(i_addr_pc4[31]), .D(n5), .Q(n74)
         );
  INV2 U14 ( .A(i_con_jump[0]), .Q(n25) );
  NAND20 U15 ( .A(i_con_jump[0]), .B(n21), .Q(n22) );
  AOI220 U16 ( .A(i_addr_j[15]), .B(n19), .C(i_addr_pc4[15]), .D(n2), .Q(n38)
         );
  INV2 U17 ( .A(i_con_jump[1]), .Q(n21) );
  AOI220 U18 ( .A(i_addr_j[25]), .B(n19), .C(i_addr_pc4[25]), .D(n5), .Q(n60)
         );
  NAND22 U19 ( .A(n17), .B(n18), .Q(o_addr_jumpmux[3]) );
  NAND22 U20 ( .A(n7), .B(n8), .Q(o_addr_jumpmux[8]) );
  NAND20 U21 ( .A(i_addr_j[8]), .B(n20), .Q(n8) );
  NAND22 U22 ( .A(n15), .B(n16), .Q(o_addr_jumpmux[4]) );
  NAND20 U23 ( .A(i_addr_j[4]), .B(n20), .Q(n16) );
  NAND22 U24 ( .A(n9), .B(n10), .Q(o_addr_jumpmux[7]) );
  NAND20 U25 ( .A(i_addr_j[7]), .B(n20), .Q(n10) );
  NAND22 U26 ( .A(n3), .B(n4), .Q(o_addr_jumpmux[9]) );
  NAND20 U27 ( .A(i_addr_j[9]), .B(n20), .Q(n4) );
  NAND20 U28 ( .A(i_addr_j[6]), .B(n20), .Q(n12) );
  NAND22 U29 ( .A(n13), .B(n14), .Q(o_addr_jumpmux[5]) );
  NAND22 U30 ( .A(n67), .B(n68), .Q(o_addr_jumpmux[0]) );
  NAND20 U31 ( .A(i_addr_j[0]), .B(n20), .Q(n68) );
  NAND22 U32 ( .A(n45), .B(n46), .Q(o_addr_jumpmux[1]) );
  NAND20 U33 ( .A(i_addr_j[1]), .B(n19), .Q(n46) );
  NAND22 U34 ( .A(n23), .B(n24), .Q(o_addr_jumpmux[2]) );
  AOI220 U35 ( .A(i_addr_j[18]), .B(n19), .C(i_addr_pc4[18]), .D(n2), .Q(n44)
         );
  AOI220 U36 ( .A(i_addr_j[23]), .B(n19), .C(i_addr_pc4[23]), .D(n5), .Q(n56)
         );
  AOI220 U37 ( .A(i_addr_pc4[7]), .B(n5), .C(i_addr_jr[7]), .D(n75), .Q(n9) );
  AOI220 U38 ( .A(i_addr_pc4[8]), .B(n5), .C(i_addr_jr[8]), .D(n75), .Q(n7) );
  AOI220 U39 ( .A(i_addr_pc4[9]), .B(n5), .C(i_addr_jr[9]), .D(n75), .Q(n3) );
  AOI220 U40 ( .A(i_addr_pc4[2]), .B(n6), .C(i_addr_jr[2]), .D(n75), .Q(n23)
         );
  AOI220 U41 ( .A(i_addr_pc4[4]), .B(n6), .C(i_addr_jr[4]), .D(n75), .Q(n15)
         );
  AOI220 U42 ( .A(i_addr_pc4[5]), .B(n6), .C(i_addr_jr[5]), .D(n75), .Q(n13)
         );
  AOI220 U43 ( .A(i_addr_j[28]), .B(n19), .C(i_addr_pc4[28]), .D(n5), .Q(n66)
         );
  AOI220 U44 ( .A(i_addr_j[29]), .B(n20), .C(i_addr_pc4[29]), .D(n5), .Q(n70)
         );
  AOI220 U45 ( .A(i_addr_j[30]), .B(n20), .C(i_addr_pc4[30]), .D(n5), .Q(n72)
         );
  AOI220 U46 ( .A(i_addr_j[12]), .B(n19), .C(i_addr_pc4[12]), .D(n2), .Q(n32)
         );
  AOI220 U47 ( .A(i_addr_j[13]), .B(n19), .C(i_addr_pc4[13]), .D(n2), .Q(n34)
         );
  AOI220 U48 ( .A(i_addr_j[14]), .B(n19), .C(i_addr_pc4[14]), .D(n2), .Q(n36)
         );
  AOI220 U49 ( .A(i_addr_j[16]), .B(n19), .C(i_addr_pc4[16]), .D(n2), .Q(n40)
         );
  AOI220 U50 ( .A(i_addr_j[17]), .B(n19), .C(i_addr_pc4[17]), .D(n2), .Q(n42)
         );
  AOI220 U51 ( .A(i_addr_j[19]), .B(n19), .C(i_addr_pc4[19]), .D(n2), .Q(n48)
         );
  AOI220 U52 ( .A(i_addr_j[21]), .B(n19), .C(i_addr_pc4[21]), .D(n2), .Q(n52)
         );
  AOI220 U53 ( .A(i_addr_j[24]), .B(n19), .C(i_addr_pc4[24]), .D(n5), .Q(n58)
         );
  AOI220 U54 ( .A(i_addr_pc4[1]), .B(n6), .C(i_addr_jr[1]), .D(n75), .Q(n45)
         );
  AOI220 U55 ( .A(i_addr_pc4[0]), .B(n6), .C(i_addr_jr[0]), .D(n75), .Q(n67)
         );
  AOI220 U56 ( .A(i_addr_j[10]), .B(n20), .C(i_addr_pc4[10]), .D(n2), .Q(n28)
         );
  AOI220 U57 ( .A(i_addr_j[11]), .B(n20), .C(i_addr_pc4[11]), .D(n2), .Q(n30)
         );
  NAND20 U58 ( .A(i_addr_j[3]), .B(n20), .Q(n18) );
  NAND20 U59 ( .A(i_addr_j[5]), .B(n20), .Q(n14) );
  NAND20 U60 ( .A(i_addr_j[2]), .B(n20), .Q(n24) );
  BUF2 U61 ( .A(n77), .Q(n19) );
  BUF2 U62 ( .A(n76), .Q(n2) );
  BUF2 U63 ( .A(n76), .Q(n5) );
  BUF2 U64 ( .A(n76), .Q(n6) );
  BUF2 U65 ( .A(n77), .Q(n20) );
  INV3 U66 ( .A(n26), .Q(n75) );
  AOI220 U67 ( .A(i_addr_j[20]), .B(n19), .C(i_addr_pc4[20]), .D(n2), .Q(n50)
         );
  AOI220 U68 ( .A(i_addr_j[27]), .B(n19), .C(i_addr_pc4[27]), .D(n5), .Q(n64)
         );
  CLKIN3 U69 ( .A(n22), .Q(n77) );
  XNR21 U70 ( .A(i_con_jump[0]), .B(i_con_jump[1]), .Q(n76) );
  NAND22 U71 ( .A(i_con_jump[1]), .B(n25), .Q(n26) );
  NAND22 U72 ( .A(i_addr_jr[10]), .B(n75), .Q(n27) );
  NAND22 U73 ( .A(n28), .B(n27), .Q(o_addr_jumpmux[10]) );
  NAND22 U74 ( .A(i_addr_jr[11]), .B(n75), .Q(n29) );
  NAND22 U75 ( .A(n30), .B(n29), .Q(o_addr_jumpmux[11]) );
  NAND22 U76 ( .A(i_addr_jr[12]), .B(n75), .Q(n31) );
  NAND22 U77 ( .A(n32), .B(n31), .Q(o_addr_jumpmux[12]) );
  NAND22 U78 ( .A(i_addr_jr[14]), .B(n75), .Q(n35) );
  NAND22 U79 ( .A(n36), .B(n35), .Q(o_addr_jumpmux[14]) );
  NAND22 U80 ( .A(i_addr_jr[15]), .B(n1), .Q(n37) );
  NAND22 U81 ( .A(n38), .B(n37), .Q(o_addr_jumpmux[15]) );
  NAND22 U82 ( .A(i_addr_jr[16]), .B(n1), .Q(n39) );
  NAND22 U83 ( .A(n40), .B(n39), .Q(o_addr_jumpmux[16]) );
  NAND22 U84 ( .A(i_addr_jr[17]), .B(n1), .Q(n41) );
  NAND22 U85 ( .A(n42), .B(n41), .Q(o_addr_jumpmux[17]) );
  NAND22 U86 ( .A(i_addr_jr[18]), .B(n1), .Q(n43) );
  NAND22 U87 ( .A(n44), .B(n43), .Q(o_addr_jumpmux[18]) );
  NAND22 U88 ( .A(i_addr_jr[20]), .B(n1), .Q(n49) );
  NAND22 U89 ( .A(n50), .B(n49), .Q(o_addr_jumpmux[20]) );
  NAND22 U90 ( .A(i_addr_jr[21]), .B(n1), .Q(n51) );
  NAND22 U91 ( .A(n52), .B(n51), .Q(o_addr_jumpmux[21]) );
  NAND22 U92 ( .A(i_addr_jr[22]), .B(n1), .Q(n53) );
  NAND22 U93 ( .A(n54), .B(n53), .Q(o_addr_jumpmux[22]) );
  NAND22 U94 ( .A(i_addr_jr[23]), .B(n1), .Q(n55) );
  NAND22 U95 ( .A(n56), .B(n55), .Q(o_addr_jumpmux[23]) );
  NAND22 U96 ( .A(i_addr_jr[24]), .B(n1), .Q(n57) );
  NAND22 U97 ( .A(n58), .B(n57), .Q(o_addr_jumpmux[24]) );
  NAND22 U98 ( .A(i_addr_jr[25]), .B(n1), .Q(n59) );
  NAND22 U99 ( .A(n60), .B(n59), .Q(o_addr_jumpmux[25]) );
  NAND22 U100 ( .A(i_addr_jr[26]), .B(n1), .Q(n61) );
  NAND22 U101 ( .A(i_addr_jr[27]), .B(n1), .Q(n63) );
  NAND22 U102 ( .A(n64), .B(n63), .Q(o_addr_jumpmux[27]) );
  NAND22 U103 ( .A(i_addr_jr[28]), .B(n1), .Q(n65) );
  NAND22 U104 ( .A(i_addr_jr[29]), .B(n1), .Q(n69) );
  NAND22 U105 ( .A(n70), .B(n69), .Q(o_addr_jumpmux[29]) );
  NAND22 U106 ( .A(i_addr_jr[30]), .B(n1), .Q(n71) );
  NAND22 U107 ( .A(n72), .B(n71), .Q(o_addr_jumpmux[30]) );
  NAND22 U108 ( .A(i_addr_jr[31]), .B(n1), .Q(n73) );
  NAND22 U109 ( .A(n74), .B(n73), .Q(o_addr_jumpmux[31]) );
endmodule


module F_branchmux ( i_addr_jumpmux, i_addr_b, i_con_ifbranch, o_addr_nextpc
 );
  input [31:0] i_addr_jumpmux;
  input [31:0] i_addr_b;
  output [31:0] o_addr_nextpc;
  input i_con_ifbranch;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23;

  MUX22 U1 ( .A(i_addr_jumpmux[28]), .B(i_addr_b[28]), .S(n22), .Q(
        o_addr_nextpc[28]) );
  CLKBU15 U2 ( .A(i_con_ifbranch), .Q(n21) );
  MUX24 U3 ( .A(i_addr_jumpmux[8]), .B(i_addr_b[8]), .S(n22), .Q(
        o_addr_nextpc[8]) );
  BUF12 U4 ( .A(i_con_ifbranch), .Q(n23) );
  CLKBU15 U5 ( .A(i_con_ifbranch), .Q(n22) );
  INV3 U6 ( .A(i_addr_b[22]), .Q(n4) );
  INV3 U7 ( .A(i_addr_jumpmux[22]), .Q(n3) );
  INV3 U8 ( .A(i_addr_b[26]), .Q(n20) );
  INV3 U9 ( .A(i_addr_jumpmux[26]), .Q(n19) );
  INV3 U10 ( .A(i_addr_b[9]), .Q(n8) );
  INV3 U11 ( .A(i_addr_jumpmux[9]), .Q(n7) );
  INV3 U12 ( .A(i_addr_b[5]), .Q(n2) );
  INV3 U13 ( .A(i_addr_jumpmux[5]), .Q(n1) );
  INV3 U14 ( .A(i_addr_b[1]), .Q(n6) );
  INV3 U15 ( .A(i_addr_jumpmux[1]), .Q(n5) );
  INV3 U16 ( .A(i_addr_b[31]), .Q(n18) );
  INV3 U17 ( .A(i_addr_b[2]), .Q(n14) );
  INV3 U18 ( .A(i_addr_jumpmux[2]), .Q(n13) );
  INV3 U19 ( .A(i_addr_b[3]), .Q(n12) );
  INV3 U20 ( .A(i_addr_jumpmux[3]), .Q(n11) );
  INV3 U21 ( .A(i_addr_b[10]), .Q(n10) );
  INV3 U22 ( .A(i_addr_jumpmux[10]), .Q(n9) );
  INV3 U23 ( .A(i_addr_b[11]), .Q(n16) );
  INV3 U24 ( .A(i_addr_jumpmux[11]), .Q(n15) );
  INV3 U25 ( .A(i_addr_jumpmux[31]), .Q(n17) );
  IMUX22 U26 ( .A(n1), .B(n2), .S(n23), .Q(o_addr_nextpc[5]) );
  IMUX22 U27 ( .A(n3), .B(n4), .S(n23), .Q(o_addr_nextpc[22]) );
  IMUX22 U28 ( .A(n5), .B(n6), .S(n23), .Q(o_addr_nextpc[1]) );
  IMUX21 U29 ( .A(n19), .B(n20), .S(n22), .Q(o_addr_nextpc[26]) );
  IMUX21 U30 ( .A(n17), .B(n18), .S(n22), .Q(o_addr_nextpc[31]) );
  IMUX22 U31 ( .A(n7), .B(n8), .S(n22), .Q(o_addr_nextpc[9]) );
  IMUX22 U32 ( .A(n9), .B(n10), .S(n22), .Q(o_addr_nextpc[10]) );
  IMUX22 U33 ( .A(n11), .B(n12), .S(n22), .Q(o_addr_nextpc[3]) );
  IMUX22 U34 ( .A(n13), .B(n14), .S(n22), .Q(o_addr_nextpc[2]) );
  IMUX22 U35 ( .A(n15), .B(n16), .S(n22), .Q(o_addr_nextpc[11]) );
  MUX24 U36 ( .A(i_addr_jumpmux[29]), .B(i_addr_b[29]), .S(n23), .Q(
        o_addr_nextpc[29]) );
  MUX24 U37 ( .A(i_addr_jumpmux[30]), .B(i_addr_b[30]), .S(n23), .Q(
        o_addr_nextpc[30]) );
  MUX24 U38 ( .A(i_addr_jumpmux[20]), .B(i_addr_b[20]), .S(n23), .Q(
        o_addr_nextpc[20]) );
  MUX24 U39 ( .A(i_addr_jumpmux[17]), .B(i_addr_b[17]), .S(n23), .Q(
        o_addr_nextpc[17]) );
  MUX24 U40 ( .A(i_addr_jumpmux[18]), .B(i_addr_b[18]), .S(n21), .Q(
        o_addr_nextpc[18]) );
  MUX24 U41 ( .A(i_addr_jumpmux[21]), .B(i_addr_b[21]), .S(n21), .Q(
        o_addr_nextpc[21]) );
  MUX24 U42 ( .A(i_addr_jumpmux[19]), .B(i_addr_b[19]), .S(n21), .Q(
        o_addr_nextpc[19]) );
  MUX24 U43 ( .A(i_addr_jumpmux[25]), .B(i_addr_b[25]), .S(n21), .Q(
        o_addr_nextpc[25]) );
  MUX24 U44 ( .A(i_addr_jumpmux[15]), .B(i_addr_b[15]), .S(n21), .Q(
        o_addr_nextpc[15]) );
  MUX24 U45 ( .A(i_addr_jumpmux[24]), .B(i_addr_b[24]), .S(n23), .Q(
        o_addr_nextpc[24]) );
  MUX24 U46 ( .A(i_addr_jumpmux[23]), .B(i_addr_b[23]), .S(n21), .Q(
        o_addr_nextpc[23]) );
  MUX24 U47 ( .A(i_addr_jumpmux[16]), .B(i_addr_b[16]), .S(n21), .Q(
        o_addr_nextpc[16]) );
  MUX24 U48 ( .A(i_addr_jumpmux[27]), .B(i_addr_b[27]), .S(n21), .Q(
        o_addr_nextpc[27]) );
  MUX24 U49 ( .A(i_addr_jumpmux[14]), .B(i_addr_b[14]), .S(n21), .Q(
        o_addr_nextpc[14]) );
  MUX24 U50 ( .A(i_addr_jumpmux[13]), .B(i_addr_b[13]), .S(n23), .Q(
        o_addr_nextpc[13]) );
  MUX24 U51 ( .A(i_addr_jumpmux[0]), .B(i_addr_b[0]), .S(n21), .Q(
        o_addr_nextpc[0]) );
  MUX24 U52 ( .A(i_addr_jumpmux[4]), .B(i_addr_b[4]), .S(n23), .Q(
        o_addr_nextpc[4]) );
  MUX24 U53 ( .A(i_addr_jumpmux[6]), .B(i_addr_b[6]), .S(n21), .Q(
        o_addr_nextpc[6]) );
  MUX24 U54 ( .A(i_addr_jumpmux[7]), .B(i_addr_b[7]), .S(n21), .Q(
        o_addr_nextpc[7]) );
  MUX24 U55 ( .A(i_addr_jumpmux[12]), .B(i_addr_b[12]), .S(n22), .Q(
        o_addr_nextpc[12]) );
endmodule


module F_pc ( i_clk, i_rst_n, i_con_stall, i_addr_next_pc, o_addr_pc );
  input [31:0] i_addr_next_pc;
  output [31:0] o_addr_pc;
  input i_clk, i_rst_n, i_con_stall;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  DFC1 program_counter_reg_21_ ( .D(n20), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[21]) );
  DFC1 program_counter_reg_19_ ( .D(n19), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[19]) );
  DFC1 program_counter_reg_18_ ( .D(n18), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[18]) );
  DFC1 program_counter_reg_16_ ( .D(n17), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[16]) );
  DFC1 program_counter_reg_13_ ( .D(n16), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[13]) );
  DFC1 program_counter_reg_12_ ( .D(n15), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[12]) );
  DFC1 program_counter_reg_11_ ( .D(n14), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[11]) );
  DFC1 program_counter_reg_10_ ( .D(n13), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[10]) );
  DFC1 program_counter_reg_9_ ( .D(n12), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[9]) );
  DFC1 program_counter_reg_6_ ( .D(n10), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[6]) );
  DFC1 program_counter_reg_4_ ( .D(n9), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[4]) );
  DFC1 program_counter_reg_3_ ( .D(n8), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[3]) );
  DFC1 program_counter_reg_2_ ( .D(n7), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[2]) );
  DFC1 program_counter_reg_0_ ( .D(n6), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[0]) );
  DFEC3 program_counter_reg_27_ ( .D(i_addr_next_pc[27]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[27]) );
  DFEC3 program_counter_reg_29_ ( .D(i_addr_next_pc[29]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[29]) );
  DFEC3 program_counter_reg_26_ ( .D(i_addr_next_pc[26]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[26]) );
  DFEC3 program_counter_reg_30_ ( .D(i_addr_next_pc[30]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[30]) );
  DFEC3 program_counter_reg_31_ ( .D(i_addr_next_pc[31]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[31]) );
  DFC1 program_counter_reg_8_ ( .D(n11), .C(i_clk), .RN(i_rst_n), .Q(
        o_addr_pc[8]) );
  DFEC3 program_counter_reg_1_ ( .D(i_addr_next_pc[1]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[1]) );
  DFEC3 program_counter_reg_25_ ( .D(i_addr_next_pc[25]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[25]) );
  DFEC3 program_counter_reg_22_ ( .D(i_addr_next_pc[22]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[22]) );
  DFEC3 program_counter_reg_23_ ( .D(i_addr_next_pc[23]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[23]) );
  DFEC3 program_counter_reg_7_ ( .D(i_addr_next_pc[7]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[7]) );
  DFEC3 program_counter_reg_5_ ( .D(i_addr_next_pc[5]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[5]) );
  DFEC3 program_counter_reg_24_ ( .D(i_addr_next_pc[24]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[24]) );
  DFEC3 program_counter_reg_15_ ( .D(i_addr_next_pc[15]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[15]) );
  DFEC3 program_counter_reg_17_ ( .D(i_addr_next_pc[17]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[17]) );
  DFEC3 program_counter_reg_20_ ( .D(i_addr_next_pc[20]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[20]) );
  DFEC3 program_counter_reg_14_ ( .D(i_addr_next_pc[14]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[14]) );
  DFEC1 program_counter_reg_28_ ( .D(i_addr_next_pc[28]), .E(n21), .C(i_clk), 
        .RN(i_rst_n), .Q(o_addr_pc[28]) );
  NAND26 U2 ( .A(i_addr_next_pc[4]), .B(n1), .Q(n2) );
  NAND20 U3 ( .A(o_addr_pc[4]), .B(n5), .Q(n3) );
  NAND26 U4 ( .A(n2), .B(n3), .Q(n9) );
  INV12 U5 ( .A(n5), .Q(n1) );
  INV3 U6 ( .A(i_con_stall), .Q(n5) );
  INV3 U7 ( .A(i_con_stall), .Q(n4) );
  MUX24 U8 ( .A(i_addr_next_pc[11]), .B(o_addr_pc[11]), .S(n4), .Q(n14) );
  MUX24 U9 ( .A(i_addr_next_pc[9]), .B(o_addr_pc[9]), .S(n4), .Q(n12) );
  MUX24 U10 ( .A(i_addr_next_pc[10]), .B(o_addr_pc[10]), .S(n5), .Q(n13) );
  MUX24 U11 ( .A(i_addr_next_pc[3]), .B(o_addr_pc[3]), .S(n4), .Q(n8) );
  MUX24 U12 ( .A(i_addr_next_pc[2]), .B(o_addr_pc[2]), .S(n5), .Q(n7) );
  MUX24 U13 ( .A(i_addr_next_pc[13]), .B(o_addr_pc[13]), .S(n5), .Q(n16) );
  MUX24 U14 ( .A(i_addr_next_pc[12]), .B(o_addr_pc[12]), .S(n4), .Q(n15) );
  MUX24 U15 ( .A(i_addr_next_pc[6]), .B(o_addr_pc[6]), .S(n5), .Q(n10) );
  MUX24 U16 ( .A(i_addr_next_pc[16]), .B(o_addr_pc[16]), .S(n4), .Q(n17) );
  MUX24 U17 ( .A(i_addr_next_pc[21]), .B(o_addr_pc[21]), .S(n4), .Q(n20) );
  MUX24 U18 ( .A(i_addr_next_pc[18]), .B(o_addr_pc[18]), .S(n5), .Q(n18) );
  MUX24 U19 ( .A(i_addr_next_pc[19]), .B(o_addr_pc[19]), .S(n5), .Q(n19) );
  MUX24 U20 ( .A(i_addr_next_pc[0]), .B(o_addr_pc[0]), .S(n4), .Q(n6) );
  MUX26 U21 ( .A(o_addr_pc[8]), .B(i_addr_next_pc[8]), .S(n21), .Q(n11) );
  BUF2 U22 ( .A(i_con_stall), .Q(n21) );
endmodule


module F_add4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  NAND31 U2 ( .A(A[24]), .B(n23), .C(n32), .Q(n36) );
  INV3 U3 ( .A(n26), .Q(n32) );
  NAND22 U4 ( .A(n49), .B(A[21]), .Q(n48) );
  NAND22 U5 ( .A(A[8]), .B(n90), .Q(n1) );
  NAND22 U6 ( .A(n79), .B(n90), .Q(n80) );
  NAND22 U7 ( .A(n78), .B(n90), .Q(n77) );
  NAND22 U8 ( .A(A[16]), .B(n32), .Q(n63) );
  NAND22 U9 ( .A(n60), .B(n32), .Q(n61) );
  NAND22 U10 ( .A(n39), .B(n32), .Q(n52) );
  NAND22 U11 ( .A(n23), .B(n32), .Q(n37) );
  NAND22 U12 ( .A(n35), .B(A[25]), .Q(n34) );
  NAND22 U13 ( .A(n16), .B(n22), .Q(n17) );
  NAND31 U14 ( .A(n23), .B(n24), .C(n25), .Q(n18) );
  INV3 U15 ( .A(n18), .Q(n22) );
  INV2 U16 ( .A(n26), .Q(n25) );
  NAND30 U17 ( .A(n31), .B(n32), .C(n23), .Q(n30) );
  NAND30 U18 ( .A(n47), .B(n32), .C(n46), .Q(n45) );
  XOR21 U19 ( .A(n50), .B(n42), .Q(SUM[21]) );
  NOR20 U20 ( .A(SUM[2]), .B(n14), .Q(n12) );
  INV2 U21 ( .A(A[10]), .Q(n87) );
  XNR20 U22 ( .A(n71), .B(n72), .Q(SUM[14]) );
  INV0 U23 ( .A(n75), .Q(n78) );
  INV0 U24 ( .A(A[5]), .Q(n9) );
  INV0 U25 ( .A(A[7]), .Q(n5) );
  INV0 U26 ( .A(A[11]), .Q(n84) );
  CLKIN3 U27 ( .A(A[2]), .Q(SUM[2]) );
  XNR20 U28 ( .A(A[3]), .B(SUM[2]), .Q(SUM[3]) );
  INV0 U29 ( .A(A[9]), .Q(n3) );
  NAND20 U30 ( .A(n60), .B(n32), .Q(n59) );
  XOR20 U31 ( .A(n36), .B(n28), .Q(SUM[25]) );
  NAND21 U32 ( .A(n46), .B(n32), .Q(n50) );
  XOR21 U33 ( .A(n55), .B(n63), .Q(SUM[17]) );
  XOR21 U34 ( .A(n56), .B(n61), .Q(SUM[18]) );
  INV0 U35 ( .A(n69), .Q(n79) );
  XOR21 U36 ( .A(n29), .B(n34), .Q(SUM[26]) );
  XOR20 U37 ( .A(n32), .B(A[16]), .Q(SUM[16]) );
  XNR20 U38 ( .A(A[15]), .B(n70), .Q(SUM[15]) );
  XNR21 U39 ( .A(A[23]), .B(n45), .Q(SUM[23]) );
  XNR21 U40 ( .A(A[27]), .B(n30), .Q(SUM[27]) );
  NAND20 U41 ( .A(A[4]), .B(n12), .Q(n11) );
  CLKIN3 U42 ( .A(n91), .Q(n68) );
  XNR20 U43 ( .A(A[12]), .B(n80), .Q(SUM[12]) );
  XOR20 U44 ( .A(A[4]), .B(n12), .Q(SUM[4]) );
  XNR20 U45 ( .A(A[8]), .B(n4), .Q(SUM[8]) );
  INV0 U46 ( .A(A[8]), .Q(n2) );
  INV3 U47 ( .A(n36), .Q(n35) );
  INV3 U48 ( .A(n50), .Q(n49) );
  XNR21 U49 ( .A(n86), .B(n87), .Q(SUM[10]) );
  XNR21 U50 ( .A(A[13]), .B(n77), .Q(SUM[13]) );
  XNR21 U51 ( .A(A[22]), .B(n48), .Q(SUM[22]) );
  XNR21 U52 ( .A(A[9]), .B(n1), .Q(SUM[9]) );
  INV3 U53 ( .A(n38), .Q(n23) );
  NAND22 U54 ( .A(n39), .B(n40), .Q(n38) );
  NOR31 U55 ( .A(n41), .B(n42), .C(n43), .Q(n40) );
  INV3 U56 ( .A(n90), .Q(n4) );
  NOR31 U57 ( .A(n68), .B(n14), .C(SUM[2]), .Q(n90) );
  INV3 U58 ( .A(n88), .Q(n86) );
  NAND22 U59 ( .A(n89), .B(n90), .Q(n88) );
  NOR21 U60 ( .A(n3), .B(n2), .Q(n89) );
  INV3 U61 ( .A(n73), .Q(n71) );
  NAND22 U62 ( .A(n74), .B(n90), .Q(n73) );
  NOR21 U63 ( .A(n75), .B(n76), .Q(n74) );
  XNR21 U64 ( .A(n10), .B(n9), .Q(SUM[5]) );
  XNR21 U65 ( .A(n7), .B(n8), .Q(SUM[6]) );
  NOR21 U66 ( .A(n9), .B(n11), .Q(n7) );
  NOR21 U67 ( .A(n55), .B(n62), .Q(n60) );
  NAND41 U68 ( .A(A[14]), .B(A[13]), .C(A[12]), .D(A[15]), .Q(n66) );
  NOR31 U69 ( .A(n29), .B(n27), .C(n28), .Q(n24) );
  NAND22 U70 ( .A(A[27]), .B(A[24]), .Q(n27) );
  XNR21 U71 ( .A(A[20]), .B(n52), .Q(SUM[20]) );
  XNR21 U72 ( .A(A[24]), .B(n37), .Q(SUM[24]) );
  XOR21 U73 ( .A(n84), .B(n85), .Q(SUM[11]) );
  NAND22 U74 ( .A(n86), .B(A[10]), .Q(n85) );
  XOR21 U75 ( .A(A[19]), .B(n58), .Q(SUM[19]) );
  NOR21 U76 ( .A(n56), .B(n59), .Q(n58) );
  NAND22 U77 ( .A(n71), .B(A[14]), .Q(n70) );
  NOR21 U78 ( .A(n43), .B(n42), .Q(n47) );
  XOR21 U79 ( .A(n22), .B(A[28]), .Q(SUM[28]) );
  XOR21 U80 ( .A(n20), .B(n21), .Q(SUM[29]) );
  NAND22 U81 ( .A(A[28]), .B(n22), .Q(n21) );
  XNR21 U82 ( .A(A[30]), .B(n17), .Q(SUM[30]) );
  NOR31 U83 ( .A(n33), .B(n29), .C(n28), .Q(n31) );
  INV3 U84 ( .A(A[3]), .Q(n14) );
  NAND22 U85 ( .A(A[23]), .B(A[20]), .Q(n41) );
  XNR21 U86 ( .A(A[31]), .B(n15), .Q(SUM[31]) );
  NAND31 U87 ( .A(n22), .B(n16), .C(A[30]), .Q(n15) );
  NAND22 U88 ( .A(n64), .B(n65), .Q(n26) );
  NOR21 U89 ( .A(n68), .B(n69), .Q(n64) );
  NOR21 U90 ( .A(n66), .B(n67), .Q(n65) );
  NAND22 U91 ( .A(A[3]), .B(A[2]), .Q(n67) );
  INV3 U92 ( .A(A[17]), .Q(n55) );
  INV3 U93 ( .A(A[18]), .Q(n56) );
  NAND22 U94 ( .A(n79), .B(A[12]), .Q(n75) );
  NOR21 U95 ( .A(n92), .B(n93), .Q(n91) );
  NAND22 U96 ( .A(A[6]), .B(A[7]), .Q(n93) );
  NAND22 U97 ( .A(A[4]), .B(A[5]), .Q(n92) );
  INV3 U98 ( .A(n81), .Q(n69) );
  NOR21 U99 ( .A(n82), .B(n83), .Q(n81) );
  NAND22 U100 ( .A(A[10]), .B(A[11]), .Q(n83) );
  NAND22 U101 ( .A(A[8]), .B(A[9]), .Q(n82) );
  NAND22 U102 ( .A(n53), .B(n54), .Q(n44) );
  NOR21 U103 ( .A(n55), .B(n56), .Q(n54) );
  NOR21 U104 ( .A(n62), .B(n57), .Q(n53) );
  INV3 U105 ( .A(A[19]), .Q(n57) );
  NOR21 U106 ( .A(n51), .B(n44), .Q(n46) );
  INV3 U107 ( .A(A[20]), .Q(n51) );
  INV3 U108 ( .A(A[24]), .Q(n33) );
  INV3 U109 ( .A(A[16]), .Q(n62) );
  INV3 U110 ( .A(A[25]), .Q(n28) );
  INV3 U111 ( .A(A[21]), .Q(n42) );
  INV3 U112 ( .A(A[14]), .Q(n72) );
  INV3 U113 ( .A(A[13]), .Q(n76) );
  INV3 U114 ( .A(A[6]), .Q(n8) );
  INV3 U115 ( .A(A[22]), .Q(n43) );
  INV3 U116 ( .A(A[26]), .Q(n29) );
  NOR21 U117 ( .A(n19), .B(n20), .Q(n16) );
  INV3 U118 ( .A(A[29]), .Q(n20) );
  XOR21 U119 ( .A(n5), .B(n6), .Q(SUM[7]) );
  NAND22 U120 ( .A(n7), .B(A[6]), .Q(n6) );
  INV3 U121 ( .A(A[28]), .Q(n19) );
  INV3 U122 ( .A(n11), .Q(n10) );
  CLKIN3 U123 ( .A(n44), .Q(n39) );
endmodule


module F_add4 ( i_addr_pc, o_addr_pcadd4 );
  input [31:0] i_addr_pc;
  output [31:0] o_addr_pcadd4;
  wire   n2, n1;

  F_add4_DW01_add_1 add_5 ( .A(i_addr_pc), .B({n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n2, n1, n1}), .CI(n1), .SUM(o_addr_pcadd4) );
  LOGIC0 U3 ( .Q(n1) );
  LOGIC1 U4 ( .Q(n2) );
endmodule


module fetch ( i_clk, i_nrst, i_addr_b, i_addr_j, i_addr_jr, i_con_b, i_con_j, 
        i_data_instr, i_con_ifstall, o_addr_pc, o_addr_pc4, o_data_instr );
  input [31:0] i_addr_b;
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [1:0] i_con_j;
  input [31:0] i_data_instr;
  output [31:0] o_addr_pc;
  output [31:0] o_addr_pc4;
  output [31:0] o_data_instr;
  input i_clk, i_nrst, i_con_b, i_con_ifstall;

  wire   [31:0] jmux_i_addr_pc4;
  wire   [31:0] bmux_i_addr_jumpmux;
  wire   [31:0] pc_i_addr_next_pc;

  DFC3 pipe_instr_reg_31_ ( .D(i_data_instr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[31]) );
  DFC3 pipe_instr_reg_30_ ( .D(i_data_instr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[30]) );
  DFC3 pipe_instr_reg_29_ ( .D(i_data_instr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[29]) );
  DFC3 pipe_instr_reg_28_ ( .D(i_data_instr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[28]) );
  DFC3 pipe_instr_reg_27_ ( .D(i_data_instr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[27]) );
  DFC3 pipe_instr_reg_26_ ( .D(i_data_instr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[26]) );
  DFC3 pipe_instr_reg_25_ ( .D(i_data_instr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[25]) );
  DFC3 pipe_instr_reg_24_ ( .D(i_data_instr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[24]) );
  DFC3 pipe_instr_reg_23_ ( .D(i_data_instr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[23]) );
  DFC3 pipe_instr_reg_22_ ( .D(i_data_instr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[22]) );
  DFC3 pipe_instr_reg_21_ ( .D(i_data_instr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[21]) );
  DFC3 pipe_instr_reg_20_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[20]) );
  DFC3 pipe_instr_reg_19_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[19]) );
  DFC3 pipe_instr_reg_18_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[18]) );
  DFC3 pipe_instr_reg_17_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[17]) );
  DFC3 pipe_instr_reg_16_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[16]) );
  DFC3 pipe_instr_reg_15_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[15]) );
  DFC3 pipe_instr_reg_14_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[14]) );
  DFC3 pipe_instr_reg_13_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[13]) );
  DFC3 pipe_instr_reg_12_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[12]) );
  DFC3 pipe_instr_reg_11_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[11]) );
  DFC3 pipe_instr_reg_10_ ( .D(i_data_instr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[10]) );
  DFC3 pipe_instr_reg_9_ ( .D(i_data_instr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[9]) );
  DFC3 pipe_instr_reg_8_ ( .D(i_data_instr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[8]) );
  DFC3 pipe_instr_reg_7_ ( .D(i_data_instr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[7]) );
  DFC3 pipe_instr_reg_6_ ( .D(i_data_instr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[6]) );
  DFC3 pipe_instr_reg_5_ ( .D(i_data_instr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[5]) );
  DFC3 pipe_instr_reg_4_ ( .D(i_data_instr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[4]) );
  DFC3 pipe_instr_reg_3_ ( .D(i_data_instr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[3]) );
  DFC3 pipe_instr_reg_2_ ( .D(i_data_instr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[2]) );
  DFC3 pipe_instr_reg_1_ ( .D(i_data_instr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[1]) );
  DFC3 pipe_instr_reg_0_ ( .D(i_data_instr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(jmux_i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(jmux_i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(jmux_i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(jmux_i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(jmux_i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(jmux_i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(jmux_i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(jmux_i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(jmux_i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_pc4_reg_21_ ( .D(jmux_i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(jmux_i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_pc4_reg_18_ ( .D(jmux_i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(jmux_i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(jmux_i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(jmux_i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(jmux_i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(jmux_i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(jmux_i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(jmux_i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(jmux_i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(jmux_i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(jmux_i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(jmux_i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(jmux_i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(jmux_i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(jmux_i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(jmux_i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(jmux_i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(jmux_i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(jmux_i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  F_jumpmux u_jumpmux ( .i_addr_j(i_addr_j), .i_addr_jr(i_addr_jr), 
        .i_addr_pc4(jmux_i_addr_pc4), .i_con_jump(i_con_j), .o_addr_jumpmux(
        bmux_i_addr_jumpmux) );
  F_branchmux u_branchmux ( .i_addr_jumpmux(bmux_i_addr_jumpmux), .i_addr_b(
        i_addr_b), .i_con_ifbranch(i_con_b), .o_addr_nextpc(pc_i_addr_next_pc)
         );
  F_pc u_pc ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_con_stall(i_con_ifstall), 
        .i_addr_next_pc(pc_i_addr_next_pc), .o_addr_pc(o_addr_pc) );
  F_add4 u_add4 ( .i_addr_pc(o_addr_pc), .o_addr_pcadd4(jmux_i_addr_pc4) );
  DFC1 pipe_pc4_reg_22_ ( .D(jmux_i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC1 pipe_pc4_reg_19_ ( .D(jmux_i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
endmodule


module D_control ( o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite, 
        o_con_alusrc, o_con_regwrite, o_con_ifsign, o_con_aluop, i_con_instru
 );
  output [5:0] o_con_aluop;
  input [5:0] i_con_instru;
  output o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite,
         o_con_alusrc, o_con_regwrite, o_con_ifsign;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n1, n2, n3, n5, n6, n7, n8, n9, n10;

  OAI212 U3 ( .A(n5), .B(n13), .C(n3), .Q(n12) );
  NAND21 U2 ( .A(i_con_instru[5]), .B(n7), .Q(n15) );
  NOR30 U4 ( .A(i_con_instru[2]), .B(i_con_instru[4]), .C(n27), .Q(n13) );
  NAND20 U5 ( .A(i_con_instru[3]), .B(n6), .Q(n20) );
  INV0 U6 ( .A(i_con_instru[4]), .Q(n6) );
  NAND20 U7 ( .A(i_con_instru[0]), .B(i_con_instru[1]), .Q(n24) );
  NAND20 U8 ( .A(i_con_instru[5]), .B(n5), .Q(n16) );
  OAI220 U9 ( .A(i_con_instru[3]), .B(n15), .C(i_con_instru[4]), .D(n17), .Q(
        o_con_memread) );
  NOR20 U10 ( .A(i_con_instru[3]), .B(n14), .Q(o_con_regdst) );
  OAI210 U11 ( .A(i_con_instru[3]), .B(n11), .C(n12), .Q(o_con_regwrite) );
  OAI210 U12 ( .A(i_con_instru[5]), .B(n20), .C(n14), .Q(o_con_aluop[1]) );
  INV0 U13 ( .A(i_con_instru[2]), .Q(n8) );
  NAND30 U14 ( .A(n2), .B(n9), .C(i_con_instru[2]), .Q(n17) );
  NAND30 U15 ( .A(i_con_instru[1]), .B(n10), .C(n2), .Q(n23) );
  NAND20 U16 ( .A(i_con_instru[3]), .B(n3), .Q(n21) );
  AOI2110 U17 ( .A(n24), .B(n26), .C(n21), .D(i_con_instru[4]), .Q(
        o_con_aluop[2]) );
  NAND20 U18 ( .A(i_con_instru[2]), .B(n10), .Q(n26) );
  AOI210 U19 ( .A(n23), .B(n25), .C(i_con_instru[4]), .Q(o_con_aluop[3]) );
  NAND30 U20 ( .A(n2), .B(i_con_instru[0]), .C(i_con_instru[2]), .Q(n25) );
  NOR20 U21 ( .A(i_con_instru[4]), .B(n21), .Q(o_con_aluop[0]) );
  INV0 U22 ( .A(i_con_instru[5]), .Q(n3) );
  AOI210 U23 ( .A(n17), .B(n22), .C(i_con_instru[4]), .Q(o_con_aluop[4]) );
  NAND31 U24 ( .A(n24), .B(n3), .C(n13), .Q(n14) );
  NAND22 U25 ( .A(n9), .B(n13), .Q(n11) );
  AOI211 U26 ( .A(n5), .B(n8), .C(o_con_memwrite), .Q(n18) );
  INV3 U27 ( .A(n20), .Q(n5) );
  INV3 U28 ( .A(n24), .Q(n9) );
  NAND22 U29 ( .A(n20), .B(n15), .Q(o_con_alusrc) );
  NAND22 U30 ( .A(n15), .B(n16), .Q(o_con_memtoreg) );
  NOR21 U31 ( .A(n11), .B(n21), .Q(o_con_aluop[5]) );
  INV3 U32 ( .A(n16), .Q(o_con_memwrite) );
  INV3 U33 ( .A(n21), .Q(n2) );
  XNR21 U34 ( .A(i_con_instru[1]), .B(n10), .Q(n27) );
  INV3 U35 ( .A(n11), .Q(n7) );
  OAI2111 U36 ( .A(n9), .B(n18), .C(n19), .D(n15), .Q(o_con_ifsign) );
  NAND31 U37 ( .A(n9), .B(n5), .C(i_con_instru[2]), .Q(n19) );
  INV3 U38 ( .A(i_con_instru[0]), .Q(n10) );
  NAND22 U39 ( .A(n1), .B(n8), .Q(n22) );
  INV3 U40 ( .A(n23), .Q(n1) );
endmodule


module D_jb_control ( o_con_jump, o_con_bop, o_con_aluPC4, o_con_ifstall, 
        i_con_instru, i_con_func, i_con_rt );
  output [1:0] o_con_jump;
  output [2:0] o_con_bop;
  input [5:0] i_con_instru;
  input [5:0] i_con_func;
  input i_con_rt;
  output o_con_aluPC4, o_con_ifstall;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n2, n3, n4,
         n5, n6;

  OAI222 U13 ( .A(n5), .B(n16), .C(n14), .D(n17), .Q(o_con_bop[1]) );
  NOR32 U3 ( .A(i_con_instru[3]), .B(i_con_instru[5]), .C(i_con_instru[4]), 
        .Q(n7) );
  INV3 U4 ( .A(i_con_instru[2]), .Q(n3) );
  NAND21 U5 ( .A(n7), .B(n8), .Q(o_con_jump[1]) );
  INV0 U6 ( .A(n7), .Q(n2) );
  NAND20 U7 ( .A(n7), .B(n4), .Q(n17) );
  CLKIN3 U8 ( .A(i_con_instru[1]), .Q(n5) );
  NAND20 U9 ( .A(i_con_instru[0]), .B(n5), .Q(n14) );
  NAND30 U10 ( .A(n7), .B(n6), .C(i_con_instru[2]), .Q(n16) );
  XNR20 U11 ( .A(n5), .B(i_con_instru[2]), .Q(n15) );
  NOR20 U12 ( .A(i_con_instru[2]), .B(i_con_rt), .Q(n18) );
  NAND31 U14 ( .A(n5), .B(n3), .C(n6), .Q(n8) );
  INV3 U15 ( .A(n13), .Q(o_con_ifstall) );
  AOI211 U16 ( .A(n3), .B(n14), .C(n2), .Q(n13) );
  OAI311 U17 ( .A(n4), .B(n2), .C(n14), .D(n16), .Q(o_con_bop[0]) );
  OAI2111 U18 ( .A(n9), .B(n8), .C(n10), .D(n7), .Q(o_con_jump[0]) );
  NOR40 U19 ( .A(n11), .B(i_con_func[2]), .C(i_con_func[5]), .D(i_con_func[4]), 
        .Q(n9) );
  NAND22 U20 ( .A(i_con_instru[1]), .B(n3), .Q(n10) );
  NAND22 U21 ( .A(n12), .B(i_con_func[3]), .Q(n11) );
  INV3 U22 ( .A(i_con_instru[0]), .Q(n6) );
  NOR21 U23 ( .A(i_con_func[1]), .B(i_con_func[0]), .Q(n12) );
  NOR40 U24 ( .A(i_con_instru[2]), .B(n2), .C(n5), .D(n6), .Q(o_con_aluPC4) );
  NOR31 U25 ( .A(n15), .B(n2), .C(n6), .Q(o_con_bop[2]) );
  INV3 U26 ( .A(n18), .Q(n4) );
endmodule


module D_pcadd_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300;

  NAND22 U2 ( .A(n89), .B(n102), .Q(n103) );
  NAND22 U3 ( .A(n27), .B(n29), .Q(n30) );
  NAND22 U4 ( .A(n16), .B(n17), .Q(n14) );
  NAND22 U5 ( .A(n244), .B(n204), .Q(n245) );
  NAND22 U6 ( .A(n165), .B(n169), .Q(n187) );
  NAND22 U7 ( .A(n167), .B(n163), .Q(n183) );
  NAND22 U8 ( .A(n131), .B(n144), .Q(n145) );
  MUX22 U9 ( .A(B[0]), .B(n300), .S(A[0]), .Q(SUM[0]) );
  INV3 U10 ( .A(n233), .Q(n225) );
  NOR21 U11 ( .A(A[5]), .B(B[5]), .Q(n35) );
  NAND22 U12 ( .A(n185), .B(n165), .Q(n184) );
  NAND24 U13 ( .A(n118), .B(n119), .Q(n65) );
  AOI212 U14 ( .A(n124), .B(n125), .C(n126), .Q(n118) );
  INV3 U15 ( .A(A[3]), .Q(n292) );
  INV1 U16 ( .A(B[3]), .Q(n293) );
  NOR20 U17 ( .A(A[3]), .B(B[3]), .Q(n297) );
  OAI2111 U18 ( .A(n225), .B(n224), .C(n220), .D(n221), .Q(n255) );
  AOI211 U19 ( .A(n181), .B(n167), .C(n182), .Q(n180) );
  INV2 U20 ( .A(B[15]), .Q(n205) );
  CLKIN2 U21 ( .A(B[19]), .Q(n8) );
  NOR20 U22 ( .A(n272), .B(n217), .Q(n273) );
  INV3 U23 ( .A(n226), .Q(n222) );
  AOI310 U24 ( .A(n259), .B(n17), .C(n215), .D(n217), .Q(n258) );
  NAND21 U25 ( .A(B[10]), .B(A[10]), .Q(n215) );
  CLKIN1 U26 ( .A(B[18]), .Q(n7) );
  NOR20 U27 ( .A(A[11]), .B(B[11]), .Q(n218) );
  NOR20 U28 ( .A(A[8]), .B(B[8]), .Q(n275) );
  AOI220 U29 ( .A(B[15]), .B(A[15]), .C(n199), .D(n200), .Q(n198) );
  NAND21 U30 ( .A(B[11]), .B(A[11]), .Q(n212) );
  XNR20 U31 ( .A(B[15]), .B(A[15]), .Q(n236) );
  IMUX20 U32 ( .A(n190), .B(n191), .S(n121), .Q(SUM[16]) );
  NOR20 U33 ( .A(A[10]), .B(B[10]), .Q(n264) );
  NAND20 U34 ( .A(A[12]), .B(B[12]), .Q(n202) );
  INV0 U35 ( .A(B[8]), .Q(n214) );
  INV0 U36 ( .A(A[8]), .Q(n213) );
  NOR20 U37 ( .A(A[12]), .B(B[12]), .Q(n251) );
  NAND20 U38 ( .A(B[8]), .B(A[8]), .Q(n23) );
  NAND20 U39 ( .A(B[12]), .B(A[12]), .Q(n248) );
  XNR20 U40 ( .A(B[8]), .B(A[8]), .Q(n19) );
  NOR20 U41 ( .A(B[8]), .B(A[8]), .Q(n21) );
  XNR20 U42 ( .A(B[12]), .B(A[12]), .Q(n253) );
  AOI210 U43 ( .A(n222), .B(n255), .C(n249), .Q(n254) );
  NAND20 U44 ( .A(B[8]), .B(A[8]), .Q(n259) );
  NOR30 U45 ( .A(n296), .B(n51), .C(n297), .Q(n295) );
  NOR20 U46 ( .A(n162), .B(n8), .Q(n161) );
  AOI210 U47 ( .A(n113), .B(n65), .C(n106), .Q(n112) );
  XOR20 U48 ( .A(n148), .B(n146), .Q(SUM[21]) );
  NAND20 U49 ( .A(n169), .B(n184), .Q(n181) );
  XNR20 U50 ( .A(n145), .B(n143), .Q(SUM[22]) );
  XNR20 U51 ( .A(n103), .B(n101), .Q(SUM[26]) );
  INV0 U52 ( .A(n122), .Q(n158) );
  NOR30 U53 ( .A(n153), .B(n122), .C(n151), .Q(n149) );
  CLKIN0 U54 ( .A(B[17]), .Q(n6) );
  INV0 U55 ( .A(B[22]), .Q(n10) );
  OAI2110 U56 ( .A(A[6]), .B(B[6]), .C(A[5]), .D(B[5]), .Q(n280) );
  NAND21 U57 ( .A(B[18]), .B(A[18]), .Q(n163) );
  XNR21 U58 ( .A(n2), .B(n142), .Q(SUM[23]) );
  XOR21 U59 ( .A(B[23]), .B(A[23]), .Q(n2) );
  NAND20 U60 ( .A(B[22]), .B(A[22]), .Q(n144) );
  NAND20 U61 ( .A(A[2]), .B(B[2]), .Q(n299) );
  NAND20 U62 ( .A(B[27]), .B(A[27]), .Q(n87) );
  NOR20 U63 ( .A(A[27]), .B(B[27]), .Q(n86) );
  NOR20 U64 ( .A(A[19]), .B(B[19]), .Q(n170) );
  OAI220 U65 ( .A(A[5]), .B(B[5]), .C(A[6]), .D(B[6]), .Q(n278) );
  XNR20 U66 ( .A(n3), .B(n54), .Q(SUM[30]) );
  XNR21 U67 ( .A(B[30]), .B(A[30]), .Q(n3) );
  XNR20 U68 ( .A(B[27]), .B(A[27]), .Q(n99) );
  XNR20 U69 ( .A(B[28]), .B(A[28]), .Q(n83) );
  AOI210 U70 ( .A(n81), .B(n65), .C(n79), .Q(n84) );
  XNR21 U71 ( .A(n4), .B(n52), .Q(SUM[31]) );
  XOR21 U72 ( .A(B[31]), .B(A[31]), .Q(n4) );
  AOI210 U73 ( .A(n76), .B(n65), .C(n61), .Q(n75) );
  XOR20 U74 ( .A(n74), .B(n75), .Q(SUM[29]) );
  XNR20 U75 ( .A(B[19]), .B(A[19]), .Q(n179) );
  AOI210 U76 ( .A(n158), .B(n121), .C(n125), .Q(n157) );
  NAND20 U77 ( .A(B[28]), .B(A[28]), .Q(n78) );
  NOR20 U78 ( .A(A[28]), .B(B[28]), .Q(n82) );
  NOR20 U79 ( .A(B[27]), .B(A[27]), .Q(n98) );
  NOR20 U80 ( .A(A[2]), .B(B[2]), .Q(n51) );
  NAND20 U81 ( .A(B[5]), .B(A[5]), .Q(n31) );
  XNR21 U82 ( .A(n46), .B(n5), .Q(SUM[3]) );
  XNR20 U83 ( .A(B[3]), .B(A[3]), .Q(n5) );
  NAND20 U84 ( .A(B[2]), .B(A[2]), .Q(n47) );
  INV3 U85 ( .A(n153), .Q(n121) );
  INV3 U86 ( .A(n152), .Q(n125) );
  INV3 U87 ( .A(B[30]), .Q(n13) );
  OAI2111 U88 ( .A(n20), .B(n246), .C(n247), .D(n248), .Q(n243) );
  NAND22 U89 ( .A(n249), .B(n250), .Q(n247) );
  NAND22 U90 ( .A(n250), .B(n222), .Q(n246) );
  INV3 U91 ( .A(n251), .Q(n250) );
  AOI2111 U92 ( .A(n192), .B(n193), .C(n194), .D(n195), .Q(n153) );
  INV3 U93 ( .A(n224), .Q(n193) );
  NOR31 U94 ( .A(n225), .B(n197), .C(n226), .Q(n192) );
  NAND22 U95 ( .A(n120), .B(n121), .Q(n119) );
  NAND31 U96 ( .A(n287), .B(n288), .C(n286), .Q(n233) );
  INV3 U97 ( .A(n295), .Q(n287) );
  AOI211 U98 ( .A(n289), .B(n290), .C(n291), .Q(n288) );
  INV3 U99 ( .A(n298), .Q(n286) );
  NAND22 U100 ( .A(n222), .B(n223), .Q(n219) );
  AOI311 U101 ( .A(n208), .B(n209), .C(n210), .D(n211), .Q(n196) );
  INV3 U102 ( .A(n212), .Q(n211) );
  NAND22 U103 ( .A(n216), .B(n215), .Q(n209) );
  OAI2111 U104 ( .A(n213), .B(n214), .C(n17), .D(n215), .Q(n210) );
  NAND31 U105 ( .A(n165), .B(n166), .C(n167), .Q(n164) );
  NAND22 U106 ( .A(n168), .B(n169), .Q(n166) );
  NAND22 U107 ( .A(n274), .B(n17), .Q(n270) );
  NAND22 U108 ( .A(n16), .B(n15), .Q(n274) );
  NAND22 U109 ( .A(n204), .B(n242), .Q(n238) );
  NAND22 U110 ( .A(n243), .B(n244), .Q(n242) );
  XNR21 U111 ( .A(n183), .B(n181), .Q(SUM[18]) );
  XOR21 U112 ( .A(n111), .B(n112), .Q(SUM[25]) );
  NAND22 U113 ( .A(n95), .B(n92), .Q(n111) );
  INV3 U114 ( .A(n109), .Q(n113) );
  NAND22 U115 ( .A(n104), .B(n105), .Q(n101) );
  NAND22 U116 ( .A(n106), .B(n95), .Q(n105) );
  AOI211 U117 ( .A(n107), .B(n65), .C(n108), .Q(n104) );
  INV3 U118 ( .A(n92), .Q(n108) );
  NOR21 U119 ( .A(n122), .B(n123), .Q(n120) );
  NOR21 U120 ( .A(n217), .B(n218), .Q(n208) );
  AOI211 U121 ( .A(n159), .B(n160), .C(n161), .Q(n152) );
  INV3 U122 ( .A(n170), .Q(n159) );
  NAND22 U123 ( .A(n163), .B(n164), .Q(n160) );
  NOR21 U124 ( .A(n292), .B(n293), .Q(n291) );
  NAND22 U125 ( .A(n81), .B(n80), .Q(n66) );
  NAND22 U126 ( .A(n212), .B(n256), .Q(n249) );
  NAND22 U127 ( .A(n257), .B(n258), .Q(n256) );
  AOI211 U128 ( .A(n216), .B(n215), .C(n218), .Q(n257) );
  XOR21 U129 ( .A(n270), .B(n273), .Q(SUM[10]) );
  XOR21 U130 ( .A(n238), .B(n241), .Q(SUM[14]) );
  NOR21 U131 ( .A(n240), .B(n207), .Q(n241) );
  XNR21 U132 ( .A(n14), .B(n15), .Q(SUM[9]) );
  XNR21 U133 ( .A(n245), .B(n243), .Q(SUM[13]) );
  XNR21 U134 ( .A(n187), .B(n185), .Q(SUM[17]) );
  NAND22 U135 ( .A(n136), .B(n135), .Q(n148) );
  NAND22 U136 ( .A(n31), .B(n32), .Q(n26) );
  NAND22 U137 ( .A(n33), .B(n34), .Q(n32) );
  INV3 U138 ( .A(n35), .Q(n34) );
  XNR21 U139 ( .A(n30), .B(n26), .Q(SUM[6]) );
  XNR21 U140 ( .A(n37), .B(n38), .Q(SUM[5]) );
  NOR21 U141 ( .A(n35), .B(n39), .Q(n38) );
  INV3 U142 ( .A(n33), .Q(n37) );
  INV3 U143 ( .A(n31), .Q(n39) );
  NOR21 U144 ( .A(n66), .B(n63), .Q(n64) );
  NOR21 U145 ( .A(n109), .B(n93), .Q(n107) );
  INV3 U146 ( .A(n63), .Q(n62) );
  XOR21 U147 ( .A(n49), .B(n67), .Q(SUM[2]) );
  NOR21 U148 ( .A(n68), .B(n51), .Q(n67) );
  XOR21 U149 ( .A(n71), .B(n176), .Q(SUM[1]) );
  NOR21 U150 ( .A(n177), .B(n73), .Q(n176) );
  INV3 U151 ( .A(n201), .Q(n244) );
  INV3 U152 ( .A(n216), .Q(n16) );
  INV3 U153 ( .A(n36), .Q(n27) );
  INV3 U154 ( .A(n168), .Q(n235) );
  NAND22 U155 ( .A(n69), .B(n70), .Q(n49) );
  NAND22 U156 ( .A(n71), .B(n72), .Q(n70) );
  INV3 U157 ( .A(n73), .Q(n72) );
  AOI211 U158 ( .A(n293), .B(n292), .C(n73), .Q(n289) );
  INV3 U159 ( .A(n51), .Q(n50) );
  NAND31 U160 ( .A(n167), .B(n165), .C(n171), .Q(n122) );
  NOR21 U161 ( .A(n172), .B(n173), .Q(n171) );
  NOR21 U162 ( .A(B[16]), .B(A[16]), .Q(n172) );
  NOR21 U163 ( .A(B[19]), .B(A[19]), .Q(n173) );
  NAND22 U164 ( .A(B[9]), .B(A[9]), .Q(n17) );
  NOR21 U165 ( .A(A[10]), .B(B[10]), .Q(n217) );
  NAND22 U166 ( .A(B[16]), .B(A[16]), .Q(n168) );
  NAND31 U167 ( .A(n58), .B(n59), .C(n60), .Q(n54) );
  NAND22 U168 ( .A(B[29]), .B(A[29]), .Q(n59) );
  NAND22 U169 ( .A(n61), .B(n62), .Q(n60) );
  NAND22 U170 ( .A(n64), .B(n65), .Q(n58) );
  NAND22 U171 ( .A(B[17]), .B(A[17]), .Q(n169) );
  NAND22 U172 ( .A(B[6]), .B(A[6]), .Q(n29) );
  NAND22 U173 ( .A(n227), .B(n228), .Q(n197) );
  NOR21 U174 ( .A(n231), .B(n232), .Q(n227) );
  NOR21 U175 ( .A(n229), .B(n230), .Q(n228) );
  NOR21 U176 ( .A(A[14]), .B(B[14]), .Q(n232) );
  NOR21 U177 ( .A(B[4]), .B(A[4]), .Q(n284) );
  NOR21 U178 ( .A(B[8]), .B(A[8]), .Q(n263) );
  AOI211 U179 ( .A(n205), .B(n206), .C(n207), .Q(n199) );
  OAI2111 U180 ( .A(n201), .B(n202), .C(n203), .D(n204), .Q(n200) );
  INV3 U181 ( .A(A[15]), .Q(n206) );
  NOR21 U182 ( .A(B[12]), .B(A[12]), .Q(n229) );
  NAND22 U183 ( .A(B[23]), .B(A[23]), .Q(n129) );
  NOR21 U184 ( .A(A[23]), .B(B[23]), .Q(n128) );
  AOI211 U185 ( .A(n130), .B(n131), .C(n132), .Q(n127) );
  AOI211 U186 ( .A(n88), .B(n89), .C(n90), .Q(n85) );
  NOR21 U187 ( .A(A[6]), .B(B[6]), .Q(n36) );
  NAND22 U188 ( .A(n282), .B(n283), .Q(n224) );
  NOR21 U189 ( .A(n284), .B(n285), .Q(n282) );
  NOR21 U190 ( .A(n35), .B(n36), .Q(n283) );
  NOR21 U191 ( .A(B[7]), .B(A[7]), .Q(n285) );
  NAND22 U192 ( .A(n260), .B(n261), .Q(n226) );
  NOR21 U193 ( .A(n264), .B(n265), .Q(n260) );
  NOR21 U194 ( .A(n262), .B(n263), .Q(n261) );
  NOR21 U195 ( .A(A[9]), .B(B[9]), .Q(n265) );
  AOI211 U196 ( .A(n91), .B(n92), .C(n93), .Q(n88) );
  NAND22 U197 ( .A(B[24]), .B(A[24]), .Q(n91) );
  NOR21 U198 ( .A(n149), .B(n150), .Q(n146) );
  NOR21 U199 ( .A(A[20]), .B(B[20]), .Q(n151) );
  NAND22 U200 ( .A(n276), .B(n277), .Q(n221) );
  INV3 U201 ( .A(n281), .Q(n276) );
  OAI2111 U202 ( .A(n278), .B(n279), .C(n280), .D(n29), .Q(n277) );
  NOR21 U203 ( .A(A[7]), .B(B[7]), .Q(n281) );
  NAND22 U204 ( .A(n77), .B(n78), .Q(n61) );
  NAND22 U205 ( .A(n79), .B(n80), .Q(n77) );
  NAND22 U206 ( .A(n188), .B(n168), .Q(n185) );
  NOR21 U207 ( .A(B[15]), .B(A[15]), .Q(n230) );
  NOR21 U208 ( .A(B[11]), .B(A[11]), .Q(n262) );
  NAND22 U209 ( .A(B[4]), .B(A[4]), .Q(n279) );
  NOR21 U210 ( .A(n297), .B(n299), .Q(n298) );
  XOR21 U211 ( .A(n268), .B(n269), .Q(SUM[11]) );
  XNR21 U212 ( .A(B[11]), .B(A[11]), .Q(n268) );
  AOI211 U213 ( .A(n270), .B(n271), .C(n272), .Q(n269) );
  INV3 U214 ( .A(n217), .Q(n271) );
  XOR21 U215 ( .A(n236), .B(n237), .Q(SUM[15]) );
  AOI211 U216 ( .A(n238), .B(n239), .C(n240), .Q(n237) );
  INV3 U217 ( .A(n207), .Q(n239) );
  AOI211 U218 ( .A(n143), .B(n131), .C(n132), .Q(n142) );
  XOR21 U219 ( .A(n99), .B(n100), .Q(SUM[27]) );
  AOI211 U220 ( .A(n101), .B(n89), .C(n90), .Q(n100) );
  XOR21 U221 ( .A(n83), .B(n84), .Q(SUM[28]) );
  XNR21 U222 ( .A(B[29]), .B(A[29]), .Q(n74) );
  AOI211 U223 ( .A(n53), .B(n54), .C(n55), .Q(n52) );
  NOR21 U224 ( .A(n56), .B(n13), .Q(n55) );
  XOR21 U225 ( .A(n179), .B(n180), .Q(SUM[19]) );
  NOR21 U226 ( .A(A[13]), .B(B[13]), .Q(n231) );
  IMUX21 U227 ( .A(n115), .B(n116), .S(n117), .Q(SUM[24]) );
  XNR21 U228 ( .A(B[24]), .B(A[24]), .Q(n116) );
  NOR21 U229 ( .A(n140), .B(n106), .Q(n115) );
  NAND31 U230 ( .A(n131), .B(n136), .C(n137), .Q(n123) );
  NOR21 U231 ( .A(n138), .B(n139), .Q(n137) );
  NOR21 U232 ( .A(B[23]), .B(A[23]), .Q(n139) );
  NOR21 U233 ( .A(B[20]), .B(A[20]), .Q(n138) );
  NAND22 U234 ( .A(n6), .B(n189), .Q(n165) );
  INV3 U235 ( .A(A[17]), .Q(n189) );
  NAND22 U236 ( .A(n7), .B(n186), .Q(n167) );
  INV3 U237 ( .A(A[18]), .Q(n186) );
  NAND22 U238 ( .A(n9), .B(n154), .Q(n136) );
  INV3 U239 ( .A(A[21]), .Q(n154) );
  INV3 U240 ( .A(B[21]), .Q(n9) );
  NAND22 U241 ( .A(n11), .B(n114), .Q(n95) );
  INV3 U242 ( .A(A[25]), .Q(n114) );
  INV3 U243 ( .A(B[25]), .Q(n11) );
  NOR21 U244 ( .A(A[4]), .B(B[4]), .Q(n40) );
  IMUX21 U245 ( .A(n252), .B(n253), .S(n254), .Q(SUM[12]) );
  NOR21 U246 ( .A(n266), .B(n267), .Q(n252) );
  NAND22 U247 ( .A(B[24]), .B(A[24]), .Q(n141) );
  NAND22 U248 ( .A(n10), .B(n147), .Q(n131) );
  INV3 U249 ( .A(A[22]), .Q(n147) );
  NAND22 U250 ( .A(B[25]), .B(A[25]), .Q(n92) );
  NAND22 U251 ( .A(B[13]), .B(A[13]), .Q(n204) );
  XOR21 U252 ( .A(n24), .B(n25), .Q(SUM[7]) );
  XNR21 U253 ( .A(B[7]), .B(A[7]), .Q(n24) );
  AOI211 U254 ( .A(n26), .B(n27), .C(n28), .Q(n25) );
  NOR21 U255 ( .A(A[14]), .B(B[14]), .Q(n207) );
  NOR21 U256 ( .A(A[24]), .B(B[24]), .Q(n109) );
  NOR21 U257 ( .A(A[9]), .B(B[9]), .Q(n216) );
  NAND22 U258 ( .A(B[20]), .B(A[20]), .Q(n134) );
  NAND22 U259 ( .A(B[21]), .B(A[21]), .Q(n135) );
  NOR21 U260 ( .A(A[29]), .B(B[29]), .Q(n63) );
  NAND22 U261 ( .A(B[4]), .B(A[4]), .Q(n41) );
  NAND22 U262 ( .A(B[26]), .B(A[26]), .Q(n102) );
  NOR21 U263 ( .A(A[13]), .B(B[13]), .Q(n201) );
  NAND22 U264 ( .A(B[7]), .B(A[7]), .Q(n220) );
  NOR21 U265 ( .A(B[24]), .B(A[24]), .Q(n97) );
  NAND22 U266 ( .A(B[14]), .B(A[14]), .Q(n203) );
  NAND31 U267 ( .A(n89), .B(n95), .C(n96), .Q(n94) );
  NOR21 U268 ( .A(n97), .B(n98), .Q(n96) );
  XNR21 U269 ( .A(B[16]), .B(A[16]), .Q(n190) );
  NOR21 U270 ( .A(n234), .B(n235), .Q(n191) );
  NOR21 U271 ( .A(B[16]), .B(A[16]), .Q(n234) );
  IMUX21 U272 ( .A(n18), .B(n19), .S(n20), .Q(SUM[8]) );
  NOR21 U273 ( .A(n21), .B(n22), .Q(n18) );
  IMUX21 U274 ( .A(n155), .B(n156), .S(n157), .Q(SUM[20]) );
  XNR21 U275 ( .A(B[20]), .B(A[20]), .Q(n156) );
  NOR21 U276 ( .A(n174), .B(n175), .Q(n155) );
  INV3 U277 ( .A(n82), .Q(n80) );
  INV3 U278 ( .A(A[19]), .Q(n162) );
  INV3 U279 ( .A(n57), .Q(n53) );
  NOR21 U280 ( .A(A[30]), .B(B[30]), .Q(n57) );
  NAND22 U281 ( .A(n12), .B(n110), .Q(n89) );
  INV3 U282 ( .A(A[26]), .Q(n110) );
  INV3 U283 ( .A(B[26]), .Q(n12) );
  NAND22 U284 ( .A(n47), .B(n48), .Q(n46) );
  NAND22 U285 ( .A(n49), .B(n50), .Q(n48) );
  NOR21 U286 ( .A(A[1]), .B(B[1]), .Q(n73) );
  NOR21 U287 ( .A(B[12]), .B(A[12]), .Q(n266) );
  NOR21 U288 ( .A(B[24]), .B(A[24]), .Q(n140) );
  NOR21 U289 ( .A(B[20]), .B(A[20]), .Q(n174) );
  IMUX21 U290 ( .A(n42), .B(n43), .S(n225), .Q(SUM[4]) );
  NOR21 U291 ( .A(n44), .B(n45), .Q(n42) );
  XNR21 U292 ( .A(B[4]), .B(A[4]), .Q(n43) );
  NOR21 U293 ( .A(B[4]), .B(A[4]), .Q(n44) );
  INV3 U294 ( .A(A[30]), .Q(n56) );
  INV3 U295 ( .A(B[0]), .Q(n300) );
  NAND22 U296 ( .A(B[1]), .B(A[1]), .Q(n296) );
  NAND22 U297 ( .A(B[1]), .B(A[1]), .Q(n69) );
  NOR21 U298 ( .A(n51), .B(n294), .Q(n290) );
  NAND22 U299 ( .A(B[0]), .B(A[0]), .Q(n294) );
  INV3 U300 ( .A(n178), .Q(n71) );
  NAND22 U301 ( .A(B[0]), .B(A[0]), .Q(n178) );
  CLKIN3 U302 ( .A(n23), .Q(n22) );
  CLKIN3 U303 ( .A(n29), .Q(n28) );
  OAI212 U304 ( .A(n225), .B(n40), .C(n41), .Q(n33) );
  CLKIN3 U305 ( .A(n41), .Q(n45) );
  CLKIN3 U306 ( .A(n47), .Q(n68) );
  CLKIN3 U307 ( .A(n66), .Q(n76) );
  OAI212 U308 ( .A(n85), .B(n86), .C(n87), .Q(n79) );
  CLKIN3 U309 ( .A(n94), .Q(n81) );
  CLKIN3 U310 ( .A(n102), .Q(n90) );
  CLKIN3 U311 ( .A(n95), .Q(n93) );
  CLKIN3 U312 ( .A(n65), .Q(n117) );
  OAI212 U313 ( .A(n127), .B(n128), .C(n129), .Q(n126) );
  OAI212 U314 ( .A(n133), .B(n134), .C(n135), .Q(n130) );
  CLKIN3 U315 ( .A(n123), .Q(n124) );
  CLKIN3 U316 ( .A(n141), .Q(n106) );
  CLKIN3 U317 ( .A(n144), .Q(n132) );
  OAI212 U318 ( .A(n133), .B(n146), .C(n135), .Q(n143) );
  CLKIN3 U319 ( .A(n136), .Q(n133) );
  OAI212 U320 ( .A(n151), .B(n152), .C(n134), .Q(n150) );
  CLKIN3 U321 ( .A(n134), .Q(n175) );
  CLKIN3 U322 ( .A(n69), .Q(n177) );
  CLKIN3 U323 ( .A(n163), .Q(n182) );
  OAI212 U324 ( .A(A[16]), .B(B[16]), .C(n121), .Q(n188) );
  OAI212 U325 ( .A(n196), .B(n197), .C(n198), .Q(n195) );
  OAI222 U326 ( .A(n219), .B(n220), .C(n219), .D(n221), .Q(n194) );
  CLKIN3 U327 ( .A(n197), .Q(n223) );
  CLKIN3 U328 ( .A(n203), .Q(n240) );
  CLKIN3 U329 ( .A(n248), .Q(n267) );
  CLKIN3 U330 ( .A(n215), .Q(n272) );
  OAI212 U331 ( .A(n20), .B(n275), .C(n23), .Q(n15) );
  CLKIN3 U332 ( .A(n255), .Q(n20) );
endmodule


module D_pcadd ( i_addr_pcadd4E, i_data_immshiftl, o_addr_pcbranchE );
  input [31:0] i_addr_pcadd4E;
  input [31:0] i_data_immshiftl;
  output [31:0] o_addr_pcbranchE;
  wire   n1;

  D_pcadd_DW01_add_1 add_5 ( .A(i_addr_pcadd4E), .B(i_data_immshiftl), .CI(n1), 
        .SUM(o_addr_pcbranchE) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_addr_Rt, i_con_RegWr, 
        i_addr_Rd, i_data_Rd, o_data_Rs, o_data_Rt );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rt;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr;
  wire   n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907;
  wire   [1023:0] regs;

  DFEC1 regs_reg_30__31_ ( .D(i_data_Rd[31]), .E(n871), .C(i_clk), .RN(n862), 
        .Q(regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(i_data_Rd[30]), .E(n871), .C(i_clk), .RN(n862), 
        .Q(regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(i_data_Rd[29]), .E(n871), .C(i_clk), .RN(n862), 
        .Q(regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(i_data_Rd[28]), .E(n871), .C(i_clk), .RN(n862), 
        .Q(regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(i_data_Rd[27]), .E(n871), .C(i_clk), .RN(n863), 
        .Q(regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(i_data_Rd[26]), .E(n871), .C(i_clk), .RN(n863), 
        .Q(regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(i_data_Rd[25]), .E(n871), .C(i_clk), .RN(n863), 
        .Q(regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(n856), .E(n871), .C(i_clk), .RN(n863), .Q(
        regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(i_data_Rd[23]), .E(n871), .C(i_clk), .RN(n863), 
        .Q(regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(n852), .E(n871), .C(i_clk), .RN(n863), .Q(
        regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(i_data_Rd[21]), .E(n871), .C(i_clk), .RN(n863), 
        .Q(regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(n848), .E(n871), .C(i_clk), .RN(n863), .Q(
        regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n871), .C(i_clk), .RN(n863), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(n844), .E(n871), .C(i_clk), .RN(n864), .Q(
        regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(i_data_Rd[17]), .E(n871), .C(i_clk), .RN(n864), 
        .Q(regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(n840), .E(n871), .C(i_clk), .RN(n864), .Q(
        regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(i_data_Rd[15]), .E(n871), .C(i_clk), .RN(n864), 
        .Q(regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(n836), .E(n871), .C(i_clk), .RN(n864), .Q(
        regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(i_data_Rd[13]), .E(n871), .C(i_clk), .RN(n864), 
        .Q(regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(n832), .E(n871), .C(i_clk), .RN(n864), .Q(
        regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(i_data_Rd[11]), .E(n871), .C(i_clk), .RN(n864), 
        .Q(regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(n828), .E(n871), .C(i_clk), .RN(n864), .Q(
        regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(n826), .E(n871), .C(i_clk), .RN(n865), .Q(
        regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(n824), .E(n871), .C(i_clk), .RN(n865), .Q(
        regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(i_data_Rd[7]), .E(n871), .C(i_clk), .RN(n865), 
        .Q(regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n871), .C(i_clk), .RN(n865), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(n818), .E(n871), .C(i_clk), .RN(n865), .Q(
        regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(n816), .E(n871), .C(i_clk), .RN(n865), .Q(
        regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(i_data_Rd[3]), .E(n871), .C(i_clk), .RN(n865), 
        .Q(regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(n811), .E(n871), .C(i_clk), .RN(n865), .Q(
        regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n871), .C(i_clk), .RN(n865), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(i_data_Rd[0]), .E(n871), .C(i_clk), .RN(n866), 
        .Q(regs[960]) );
  DFEC1 regs_reg_26__31_ ( .D(i_data_Rd[31]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(i_data_Rd[30]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(i_data_Rd[29]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(i_data_Rd[28]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(i_data_Rd[27]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(i_data_Rd[26]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(i_data_Rd[25]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(n856), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(i_data_Rd[23]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(n852), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(i_data_Rd[21]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(n848), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(n844), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(i_data_Rd[17]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(n840), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(i_data_Rd[15]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(n836), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(i_data_Rd[13]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(n832), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(i_data_Rd[11]), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(n828), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(n826), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(n824), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(i_data_Rd[7]), .E(n875), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n875), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(n818), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(n816), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(i_data_Rd[3]), .E(n875), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(n811), .E(n875), .C(i_clk), .RN(i_rst_n), .Q(
        regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n875), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(i_data_Rd[0]), .E(n875), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[832]) );
  DFEC1 regs_reg_22__31_ ( .D(i_data_Rd[31]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(i_data_Rd[30]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(i_data_Rd[29]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(i_data_Rd[28]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(i_data_Rd[27]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(i_data_Rd[26]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(i_data_Rd[25]), .E(n879), .C(i_clk), .RN(n869), 
        .Q(regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(i_data_Rd[24]), .E(n879), .C(i_clk), .RN(n864), 
        .Q(regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(i_data_Rd[23]), .E(n879), .C(i_clk), .RN(n861), 
        .Q(regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(i_data_Rd[22]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(i_data_Rd[21]), .E(n879), .C(i_clk), .RN(n867), 
        .Q(regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(i_data_Rd[20]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(i_data_Rd[19]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(i_data_Rd[18]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(i_data_Rd[17]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(i_data_Rd[16]), .E(n879), .C(i_clk), .RN(n866), 
        .Q(regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(i_data_Rd[15]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(i_data_Rd[14]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(i_data_Rd[13]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(i_data_Rd[12]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(i_data_Rd[11]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(i_data_Rd[10]), .E(n879), .C(i_clk), .RN(i_rst_n), .Q(regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(i_data_Rd[9]), .E(n879), .C(i_clk), .RN(n869), 
        .Q(regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(i_data_Rd[8]), .E(n879), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(i_data_Rd[7]), .E(n879), .C(i_clk), .RN(n861), 
        .Q(regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(i_data_Rd[6]), .E(n879), .C(i_clk), .RN(n862), 
        .Q(regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(i_data_Rd[5]), .E(n879), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(i_data_Rd[4]), .E(n879), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(i_data_Rd[3]), .E(n879), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(i_data_Rd[2]), .E(n879), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(i_data_Rd[1]), .E(n879), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(i_data_Rd[0]), .E(n879), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[704]) );
  DFEC1 regs_reg_18__31_ ( .D(i_data_Rd[31]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(i_data_Rd[30]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(i_data_Rd[29]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(i_data_Rd[28]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(i_data_Rd[27]), .E(n883), .C(i_clk), .RN(n863), 
        .Q(regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(i_data_Rd[26]), .E(n883), .C(i_clk), .RN(n868), 
        .Q(regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(i_data_Rd[25]), .E(n883), .C(i_clk), .RN(n861), 
        .Q(regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(i_data_Rd[24]), .E(n883), .C(i_clk), .RN(n863), 
        .Q(regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(i_data_Rd[23]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(i_data_Rd[22]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(i_data_Rd[21]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(i_data_Rd[20]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(i_data_Rd[19]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(i_data_Rd[18]), .E(n883), .C(i_clk), .RN(n865), 
        .Q(regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(i_data_Rd[17]), .E(n883), .C(i_clk), .RN(n866), 
        .Q(regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(i_data_Rd[16]), .E(n883), .C(i_clk), .RN(n862), 
        .Q(regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(i_data_Rd[15]), .E(n883), .C(i_clk), .RN(n869), 
        .Q(regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(i_data_Rd[14]), .E(n883), .C(i_clk), .RN(n865), 
        .Q(regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(i_data_Rd[13]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(i_data_Rd[12]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(i_data_Rd[11]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(i_data_Rd[10]), .E(n883), .C(i_clk), .RN(i_rst_n), .Q(regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(i_data_Rd[9]), .E(n883), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(i_data_Rd[8]), .E(n883), .C(i_clk), .RN(n865), 
        .Q(regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(i_data_Rd[7]), .E(n883), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(i_data_Rd[6]), .E(n883), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(i_data_Rd[5]), .E(n883), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(i_data_Rd[4]), .E(n883), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(i_data_Rd[3]), .E(n883), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(i_data_Rd[2]), .E(n883), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(i_data_Rd[1]), .E(n883), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(i_data_Rd[0]), .E(n883), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[576]) );
  DFEC1 regs_reg_14__31_ ( .D(n860), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(i_data_Rd[30]), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(i_data_Rd[29]), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(i_data_Rd[28]), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(i_data_Rd[27]), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(i_data_Rd[26]), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(n858), .E(n888), .C(i_clk), .RN(n867), .Q(
        regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(i_data_Rd[24]), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(n854), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(i_data_Rd[22]), .E(n888), .C(i_clk), .RN(n863), 
        .Q(regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(n850), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(i_data_Rd[20]), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(n846), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(i_data_Rd[18]), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(n842), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(i_data_Rd[16]), .E(n888), .C(i_clk), .RN(n868), 
        .Q(regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(n838), .E(n888), .C(i_clk), .RN(n863), .Q(
        regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n888), .C(i_clk), .RN(n864), 
        .Q(regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(n834), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(i_data_Rd[12]), .E(n888), .C(i_clk), .RN(n864), 
        .Q(regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(n830), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(i_data_Rd[9]), .E(n888), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(i_data_Rd[8]), .E(n888), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(n822), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(n820), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(i_data_Rd[5]), .E(n888), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(n815), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(n813), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(i_data_Rd[2]), .E(n888), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(n809), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(n807), .E(n888), .C(i_clk), .RN(i_rst_n), .Q(
        regs[448]) );
  DFEC1 regs_reg_10__31_ ( .D(n860), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(i_data_Rd[30]), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(i_data_Rd[29]), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(i_data_Rd[28]), .E(n892), .C(i_clk), .RN(n863), 
        .Q(regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(i_data_Rd[27]), .E(n892), .C(i_clk), .RN(n864), 
        .Q(regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(i_data_Rd[26]), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(n858), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(i_data_Rd[24]), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(n854), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(i_data_Rd[22]), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(n850), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(i_data_Rd[20]), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(n846), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(i_data_Rd[18]), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(n842), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(i_data_Rd[16]), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(n838), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(n834), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(i_data_Rd[12]), .E(n892), .C(i_clk), .RN(n865), 
        .Q(regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(n830), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n892), .C(i_clk), .RN(n861), 
        .Q(regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(i_data_Rd[9]), .E(n892), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(i_data_Rd[8]), .E(n892), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(n822), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(n820), .E(n892), .C(i_clk), .RN(n868), .Q(
        regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(i_data_Rd[5]), .E(n892), .C(i_clk), .RN(n869), 
        .Q(regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(n815), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(n813), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(i_data_Rd[2]), .E(n892), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(n809), .E(n892), .C(i_clk), .RN(i_rst_n), .Q(
        regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(n807), .E(n892), .C(i_clk), .RN(n867), .Q(
        regs[320]) );
  DFEC1 regs_reg_6__31_ ( .D(n859), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(i_data_Rd[30]), .E(n896), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(i_data_Rd[29]), .E(n896), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(i_data_Rd[28]), .E(n896), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(i_data_Rd[27]), .E(n896), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(i_data_Rd[26]), .E(n896), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(n857), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(n855), .E(n896), .C(i_clk), .RN(n861), .Q(
        regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(n853), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(n851), .E(n896), .C(i_clk), .RN(n863), .Q(
        regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(n849), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(n847), .E(n896), .C(i_clk), .RN(n868), .Q(
        regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(n845), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(n843), .E(n896), .C(i_clk), .RN(n863), .Q(
        regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(n841), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(n839), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(n837), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(n835), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(n833), .E(n896), .C(i_clk), .RN(n869), .Q(
        regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(n831), .E(n896), .C(i_clk), .RN(n861), .Q(
        regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(n829), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(n827), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(n825), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(n823), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(n821), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(n819), .E(n896), .C(i_clk), .RN(n867), .Q(
        regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(n817), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(n814), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(n812), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(n810), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(n808), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(n806), .E(n896), .C(i_clk), .RN(i_rst_n), .Q(
        regs[192]) );
  DFEC1 regs_reg_2__31_ ( .D(n859), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(i_data_Rd[30]), .E(n900), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(i_data_Rd[29]), .E(n900), .C(i_clk), .RN(n861), 
        .Q(regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(i_data_Rd[28]), .E(n900), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(i_data_Rd[27]), .E(n900), .C(i_clk), .RN(n867), 
        .Q(regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(i_data_Rd[26]), .E(n900), .C(i_clk), .RN(n861), 
        .Q(regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(n857), .E(n900), .C(i_clk), .RN(n865), .Q(
        regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(n855), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(n853), .E(n900), .C(i_clk), .RN(n866), .Q(
        regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(n851), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(n849), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(n847), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(n845), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(n843), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(n841), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(n839), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(n837), .E(n900), .C(i_clk), .RN(n869), .Q(
        regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(n835), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(n833), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(n831), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(n829), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(n827), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(n825), .E(n900), .C(i_clk), .RN(n862), .Q(regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(n823), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(n821), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(n819), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(n817), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(n814), .E(n900), .C(i_clk), .RN(n867), .Q(regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(n812), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(n810), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(n808), .E(n900), .C(i_clk), .RN(i_rst_n), .Q(
        regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(n806), .E(n900), .C(i_clk), .RN(n869), .Q(regs[64]) );
  DFEC1 regs_reg_31__31_ ( .D(i_data_Rd[31]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1023]) );
  DFEC1 regs_reg_31__30_ ( .D(i_data_Rd[30]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(i_data_Rd[29]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(i_data_Rd[28]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(i_data_Rd[27]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(i_data_Rd[26]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(i_data_Rd[25]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(n856), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(i_data_Rd[23]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(n852), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(i_data_Rd[21]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(n848), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(n844), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(i_data_Rd[17]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(n840), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(i_data_Rd[15]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(n836), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(i_data_Rd[13]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(n832), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(i_data_Rd[11]), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(n828), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(n826), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(n824), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(i_data_Rd[7]), .E(n870), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n870), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(n818), .E(n870), .C(i_clk), .RN(i_rst_n), .Q(
        regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(n816), .E(n870), .C(i_clk), .RN(n862), .Q(
        regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(i_data_Rd[3]), .E(n870), .C(i_clk), .RN(n862), 
        .Q(regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(n811), .E(n870), .C(i_clk), .RN(n862), .Q(
        regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n870), .C(i_clk), .RN(n862), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(i_data_Rd[0]), .E(n870), .C(i_clk), .RN(n862), 
        .Q(regs[992]) );
  DFEC1 regs_reg_29__31_ ( .D(i_data_Rd[31]), .E(n872), .C(i_clk), .RN(n866), 
        .Q(regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(i_data_Rd[30]), .E(n872), .C(i_clk), .RN(n866), 
        .Q(regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(i_data_Rd[29]), .E(n872), .C(i_clk), .RN(n866), 
        .Q(regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(i_data_Rd[28]), .E(n872), .C(i_clk), .RN(n866), 
        .Q(regs[956]) );
  DFEC1 regs_reg_29__27_ ( .D(i_data_Rd[27]), .E(n872), .C(i_clk), .RN(n866), 
        .Q(regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(i_data_Rd[26]), .E(n872), .C(i_clk), .RN(n866), 
        .Q(regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(i_data_Rd[25]), .E(n872), .C(i_clk), .RN(n866), 
        .Q(regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(n856), .E(n872), .C(i_clk), .RN(n866), .Q(
        regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(i_data_Rd[23]), .E(n872), .C(i_clk), .RN(n867), 
        .Q(regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(n852), .E(n872), .C(i_clk), .RN(n867), .Q(
        regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(i_data_Rd[21]), .E(n872), .C(i_clk), .RN(n867), 
        .Q(regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(n848), .E(n872), .C(i_clk), .RN(n867), .Q(
        regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n872), .C(i_clk), .RN(n867), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(n844), .E(n872), .C(i_clk), .RN(n867), .Q(
        regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(i_data_Rd[17]), .E(n872), .C(i_clk), .RN(n867), 
        .Q(regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(n840), .E(n872), .C(i_clk), .RN(n867), .Q(
        regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(i_data_Rd[15]), .E(n872), .C(i_clk), .RN(n867), 
        .Q(regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(n836), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(i_data_Rd[13]), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(n832), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(i_data_Rd[11]), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(n828), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(n826), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(n824), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(i_data_Rd[7]), .E(n872), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n872), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(n818), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(n816), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(i_data_Rd[3]), .E(n872), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(n811), .E(n872), .C(i_clk), .RN(i_rst_n), .Q(
        regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n872), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(i_data_Rd[0]), .E(n872), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[928]) );
  DFEC1 regs_reg_28__31_ ( .D(i_data_Rd[31]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(i_data_Rd[30]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(i_data_Rd[29]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(i_data_Rd[28]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(i_data_Rd[27]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(i_data_Rd[26]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(i_data_Rd[25]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(n856), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(i_data_Rd[23]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(n852), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(i_data_Rd[21]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(n848), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(n844), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(i_data_Rd[17]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(n840), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(i_data_Rd[15]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(n836), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(i_data_Rd[13]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(n832), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(i_data_Rd[11]), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(n828), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(n826), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(n824), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(i_data_Rd[7]), .E(n873), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n873), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(n818), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(n816), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(i_data_Rd[3]), .E(n873), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(n811), .E(n873), .C(i_clk), .RN(i_rst_n), .Q(
        regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n873), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(i_data_Rd[0]), .E(n873), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(i_data_Rd[31]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(i_data_Rd[30]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(i_data_Rd[29]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(i_data_Rd[28]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(i_data_Rd[27]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(i_data_Rd[26]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(i_data_Rd[25]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(n856), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(i_data_Rd[23]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(n852), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(i_data_Rd[21]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(n848), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(n844), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(i_data_Rd[17]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(n840), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(i_data_Rd[15]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(n836), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(i_data_Rd[13]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(n832), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(i_data_Rd[11]), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(n828), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(n826), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(n824), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(i_data_Rd[7]), .E(n874), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n874), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(n818), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(n816), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(i_data_Rd[3]), .E(n874), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(n811), .E(n874), .C(i_clk), .RN(i_rst_n), .Q(
        regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(i_data_Rd[1]), .E(n874), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(i_data_Rd[0]), .E(n874), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[864]) );
  DFEC1 regs_reg_25__31_ ( .D(n860), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(i_data_Rd[30]), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(i_data_Rd[29]), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(i_data_Rd[28]), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(i_data_Rd[27]), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(i_data_Rd[26]), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(n858), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(n856), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(n854), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(n852), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(n850), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(n848), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(n846), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(n844), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(n842), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(n840), .E(n876), .C(i_clk), .RN(n863), .Q(
        regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(n838), .E(n876), .C(i_clk), .RN(n864), .Q(
        regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(n836), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(n834), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(n832), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(n830), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(n828), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(n826), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(n824), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(n822), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(n820), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(n818), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(n816), .E(n876), .C(i_clk), .RN(n868), .Q(
        regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(n813), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(n811), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(n809), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(n807), .E(n876), .C(i_clk), .RN(i_rst_n), .Q(
        regs[800]) );
  DFEC1 regs_reg_24__31_ ( .D(n859), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(i_data_Rd[30]), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(i_data_Rd[29]), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(i_data_Rd[28]), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(i_data_Rd[27]), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(i_data_Rd[26]), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(n857), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(n856), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(n853), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(n852), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(n849), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(n848), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(n845), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(n844), .E(n877), .C(i_clk), .RN(n869), .Q(
        regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(n841), .E(n877), .C(i_clk), .RN(n867), .Q(
        regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(n840), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(n837), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(n836), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(n833), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(n832), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(n829), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(n828), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(n826), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(n824), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(n821), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(n819), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(n818), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(n816), .E(n877), .C(i_clk), .RN(n869), .Q(
        regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(n812), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(n811), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(n808), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(n806), .E(n877), .C(i_clk), .RN(i_rst_n), .Q(
        regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(i_data_Rd[31]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(i_data_Rd[30]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(i_data_Rd[29]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(i_data_Rd[28]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(i_data_Rd[27]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(i_data_Rd[26]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(i_data_Rd[25]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(i_data_Rd[24]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(i_data_Rd[23]), .E(n878), .C(i_clk), .RN(n861), 
        .Q(regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(i_data_Rd[22]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(i_data_Rd[21]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(i_data_Rd[20]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(i_data_Rd[19]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(i_data_Rd[18]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(i_data_Rd[17]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(i_data_Rd[16]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(i_data_Rd[15]), .E(n878), .C(i_clk), .RN(n869), 
        .Q(regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(i_data_Rd[14]), .E(n878), .C(i_clk), .RN(n868), 
        .Q(regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(i_data_Rd[13]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(i_data_Rd[12]), .E(n878), .C(i_clk), .RN(n868), 
        .Q(regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(i_data_Rd[11]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(i_data_Rd[10]), .E(n878), .C(i_clk), .RN(i_rst_n), .Q(regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(i_data_Rd[9]), .E(n878), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(i_data_Rd[8]), .E(n878), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(i_data_Rd[7]), .E(n878), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(i_data_Rd[6]), .E(n878), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(i_data_Rd[5]), .E(n878), .C(i_clk), .RN(n862), 
        .Q(regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(i_data_Rd[4]), .E(n878), .C(i_clk), .RN(n863), 
        .Q(regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(i_data_Rd[3]), .E(n878), .C(i_clk), .RN(n864), 
        .Q(regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(i_data_Rd[2]), .E(n878), .C(i_clk), .RN(n865), 
        .Q(regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(i_data_Rd[1]), .E(n878), .C(i_clk), .RN(n866), 
        .Q(regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(i_data_Rd[0]), .E(n878), .C(i_clk), .RN(n867), 
        .Q(regs[736]) );
  DFEC1 regs_reg_21__31_ ( .D(i_data_Rd[31]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(i_data_Rd[30]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(i_data_Rd[29]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(i_data_Rd[28]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(i_data_Rd[27]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(i_data_Rd[26]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(i_data_Rd[25]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(i_data_Rd[24]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(i_data_Rd[23]), .E(n880), .C(i_clk), .RN(n861), 
        .Q(regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(i_data_Rd[22]), .E(n880), .C(i_clk), .RN(n869), 
        .Q(regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(i_data_Rd[21]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(i_data_Rd[20]), .E(n880), .C(i_clk), .RN(n861), 
        .Q(regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(i_data_Rd[19]), .E(n880), .C(i_clk), .RN(n862), 
        .Q(regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(i_data_Rd[18]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(i_data_Rd[17]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(i_data_Rd[16]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(i_data_Rd[15]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(i_data_Rd[14]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(i_data_Rd[13]), .E(n880), .C(i_clk), .RN(n866), 
        .Q(regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(i_data_Rd[12]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(i_data_Rd[11]), .E(n880), .C(i_clk), .RN(n868), 
        .Q(regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(i_data_Rd[10]), .E(n880), .C(i_clk), .RN(i_rst_n), .Q(regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(i_data_Rd[9]), .E(n880), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(i_data_Rd[8]), .E(n880), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(i_data_Rd[7]), .E(n880), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(i_data_Rd[6]), .E(n880), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(i_data_Rd[5]), .E(n880), .C(i_clk), .RN(n864), 
        .Q(regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(i_data_Rd[4]), .E(n880), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(i_data_Rd[3]), .E(n880), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(i_data_Rd[2]), .E(n880), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(i_data_Rd[1]), .E(n880), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(i_data_Rd[0]), .E(n880), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[672]) );
  DFEC1 regs_reg_20__31_ ( .D(i_data_Rd[31]), .E(n881), .C(i_clk), .RN(n862), 
        .Q(regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(i_data_Rd[30]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(i_data_Rd[29]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(i_data_Rd[28]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(i_data_Rd[27]), .E(n881), .C(i_clk), .RN(n868), 
        .Q(regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(i_data_Rd[26]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(i_data_Rd[25]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(i_data_Rd[24]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(i_data_Rd[23]), .E(n881), .C(i_clk), .RN(n861), 
        .Q(regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(i_data_Rd[22]), .E(n881), .C(i_clk), .RN(n867), 
        .Q(regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(i_data_Rd[21]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(i_data_Rd[20]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(i_data_Rd[19]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(i_data_Rd[18]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(i_data_Rd[17]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(i_data_Rd[16]), .E(n881), .C(i_clk), .RN(n869), 
        .Q(regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(i_data_Rd[15]), .E(n881), .C(i_clk), .RN(n868), 
        .Q(regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(i_data_Rd[14]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(i_data_Rd[13]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(i_data_Rd[12]), .E(n881), .C(i_clk), .RN(n863), 
        .Q(regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(i_data_Rd[11]), .E(n881), .C(i_clk), .RN(n861), 
        .Q(regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(i_data_Rd[10]), .E(n881), .C(i_clk), .RN(i_rst_n), .Q(regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(i_data_Rd[9]), .E(n881), .C(i_clk), .RN(n868), 
        .Q(regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(i_data_Rd[8]), .E(n881), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(i_data_Rd[7]), .E(n881), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(i_data_Rd[6]), .E(n881), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(i_data_Rd[5]), .E(n881), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(i_data_Rd[4]), .E(n881), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(i_data_Rd[3]), .E(n881), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(i_data_Rd[2]), .E(n881), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(i_data_Rd[1]), .E(n881), .C(i_clk), .RN(n867), 
        .Q(regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(i_data_Rd[0]), .E(n881), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(i_data_Rd[31]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(i_data_Rd[30]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(i_data_Rd[29]), .E(n882), .C(i_clk), .RN(n864), 
        .Q(regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(i_data_Rd[28]), .E(n882), .C(i_clk), .RN(n862), 
        .Q(regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(i_data_Rd[27]), .E(n882), .C(i_clk), .RN(n861), 
        .Q(regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(i_data_Rd[26]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(i_data_Rd[25]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(n856), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(
        regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(i_data_Rd[23]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(n852), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(
        regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(i_data_Rd[21]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(n848), .E(n882), .C(i_clk), .RN(n861), .Q(
        regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(i_data_Rd[19]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(n844), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(
        regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(i_data_Rd[17]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(n840), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(
        regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(i_data_Rd[15]), .E(n882), .C(i_clk), .RN(n869), 
        .Q(regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(n836), .E(n882), .C(i_clk), .RN(n868), .Q(
        regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(i_data_Rd[13]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(n832), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(
        regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(i_data_Rd[11]), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(n828), .E(n882), .C(i_clk), .RN(n864), .Q(
        regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(n826), .E(n882), .C(i_clk), .RN(n865), .Q(
        regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(n824), .E(n882), .C(i_clk), .RN(n866), .Q(
        regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(i_data_Rd[7]), .E(n882), .C(i_clk), .RN(n867), 
        .Q(regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(i_data_Rd[6]), .E(n882), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(n818), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(
        regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(n815), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(
        regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(i_data_Rd[3]), .E(n882), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(n811), .E(n882), .C(i_clk), .RN(i_rst_n), .Q(
        regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(i_data_Rd[1]), .E(n882), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(i_data_Rd[0]), .E(n882), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[608]) );
  DFEC1 regs_reg_17__31_ ( .D(i_data_Rd[31]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(i_data_Rd[30]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(i_data_Rd[29]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(i_data_Rd[28]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(i_data_Rd[27]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(i_data_Rd[26]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(i_data_Rd[25]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(i_data_Rd[24]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(i_data_Rd[23]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(i_data_Rd[22]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(i_data_Rd[21]), .E(n884), .C(i_clk), .RN(n869), 
        .Q(regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(i_data_Rd[20]), .E(n884), .C(i_clk), .RN(n861), 
        .Q(regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(i_data_Rd[19]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(i_data_Rd[18]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(i_data_Rd[17]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(i_data_Rd[16]), .E(n884), .C(i_clk), .RN(n866), 
        .Q(regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(i_data_Rd[15]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(i_data_Rd[14]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(i_data_Rd[13]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(i_data_Rd[12]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(i_data_Rd[11]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(i_data_Rd[10]), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(i_data_Rd[9]), .E(n884), .C(i_clk), .RN(n866), 
        .Q(regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(i_data_Rd[8]), .E(n884), .C(i_clk), .RN(n865), 
        .Q(regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(i_data_Rd[7]), .E(n884), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(i_data_Rd[6]), .E(n884), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(i_data_Rd[5]), .E(n884), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(n816), .E(n884), .C(i_clk), .RN(i_rst_n), .Q(
        regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(i_data_Rd[3]), .E(n884), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(i_data_Rd[2]), .E(n884), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(i_data_Rd[1]), .E(n884), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(i_data_Rd[0]), .E(n884), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(i_data_Rd[31]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(i_data_Rd[30]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(i_data_Rd[29]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(i_data_Rd[28]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(i_data_Rd[27]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(i_data_Rd[26]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(i_data_Rd[25]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(n855), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(i_data_Rd[23]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(n851), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(i_data_Rd[21]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(n847), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(i_data_Rd[19]), .E(n885), .C(i_clk), .RN(n869), 
        .Q(regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(n843), .E(n885), .C(i_clk), .RN(n868), .Q(
        regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(i_data_Rd[17]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(n839), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(i_data_Rd[15]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(n835), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(i_data_Rd[13]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(n831), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(i_data_Rd[11]), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(n827), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(n825), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(n823), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(i_data_Rd[7]), .E(n885), .C(i_clk), .RN(n865), 
        .Q(regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(i_data_Rd[6]), .E(n885), .C(i_clk), .RN(n866), 
        .Q(regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(n817), .E(n885), .C(i_clk), .RN(n867), .Q(
        regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(n814), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(i_data_Rd[3]), .E(n885), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(n810), .E(n885), .C(i_clk), .RN(i_rst_n), .Q(
        regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(i_data_Rd[1]), .E(n885), .C(i_clk), .RN(n868), 
        .Q(regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(i_data_Rd[0]), .E(n885), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[512]) );
  DFEC1 regs_reg_15__31_ ( .D(n860), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(i_data_Rd[30]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(i_data_Rd[29]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(i_data_Rd[28]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(i_data_Rd[27]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(i_data_Rd[26]), .E(n887), .C(i_clk), .RN(n862), 
        .Q(regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(n858), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(i_data_Rd[24]), .E(n887), .C(i_clk), .RN(n867), 
        .Q(regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(n854), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(i_data_Rd[22]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(n850), .E(n887), .C(i_clk), .RN(n866), .Q(
        regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(i_data_Rd[20]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(n846), .E(n887), .C(i_clk), .RN(n864), .Q(
        regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(i_data_Rd[18]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(n842), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(i_data_Rd[16]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(n838), .E(n887), .C(i_clk), .RN(n866), .Q(
        regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(n834), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(i_data_Rd[12]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(n830), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(i_data_Rd[9]), .E(n887), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(i_data_Rd[8]), .E(n887), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(n822), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(n820), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(i_data_Rd[5]), .E(n887), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(n815), .E(n887), .C(i_clk), .RN(n864), .Q(
        regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(n813), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(i_data_Rd[2]), .E(n887), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(n809), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(n807), .E(n887), .C(i_clk), .RN(i_rst_n), .Q(
        regs[480]) );
  DFEC1 regs_reg_13__31_ ( .D(n860), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(i_data_Rd[30]), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(i_data_Rd[29]), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(i_data_Rd[28]), .E(n889), .C(i_clk), .RN(n862), 
        .Q(regs[444]) );
  DFEC1 regs_reg_13__27_ ( .D(i_data_Rd[27]), .E(n889), .C(i_clk), .RN(n863), 
        .Q(regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(i_data_Rd[26]), .E(n889), .C(i_clk), .RN(n864), 
        .Q(regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(n858), .E(n889), .C(i_clk), .RN(n865), .Q(
        regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(i_data_Rd[24]), .E(n889), .C(i_clk), .RN(n866), 
        .Q(regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(n854), .E(n889), .C(i_clk), .RN(n867), .Q(
        regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(i_data_Rd[22]), .E(n889), .C(i_clk), .RN(n865), 
        .Q(regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(n850), .E(n889), .C(i_clk), .RN(n863), .Q(
        regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(i_data_Rd[20]), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(n846), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(i_data_Rd[18]), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(n842), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(i_data_Rd[16]), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(n838), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(n834), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(i_data_Rd[12]), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(n830), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(i_data_Rd[9]), .E(n889), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(i_data_Rd[8]), .E(n889), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(n822), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(n820), .E(n889), .C(i_clk), .RN(n868), .Q(
        regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(i_data_Rd[5]), .E(n889), .C(i_clk), .RN(n869), 
        .Q(regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(n815), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(n813), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(i_data_Rd[2]), .E(n889), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(n809), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(n807), .E(n889), .C(i_clk), .RN(i_rst_n), .Q(
        regs[416]) );
  DFEC1 regs_reg_12__31_ ( .D(n860), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(i_data_Rd[30]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(i_data_Rd[29]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(i_data_Rd[28]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(i_data_Rd[27]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(i_data_Rd[26]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(n858), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(i_data_Rd[24]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(n854), .E(n890), .C(i_clk), .RN(n867), .Q(
        regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(i_data_Rd[22]), .E(n890), .C(i_clk), .RN(n865), 
        .Q(regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(n850), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(i_data_Rd[20]), .E(n890), .C(i_clk), .RN(n864), 
        .Q(regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(n846), .E(n890), .C(i_clk), .RN(n865), .Q(
        regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(i_data_Rd[18]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(n842), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(i_data_Rd[16]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(n838), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(n834), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(i_data_Rd[12]), .E(n890), .C(i_clk), .RN(n868), 
        .Q(regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(n830), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(i_data_Rd[9]), .E(n890), .C(i_clk), .RN(n862), 
        .Q(regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(i_data_Rd[8]), .E(n890), .C(i_clk), .RN(n868), 
        .Q(regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(n822), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(n820), .E(n890), .C(i_clk), .RN(n865), .Q(
        regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(i_data_Rd[5]), .E(n890), .C(i_clk), .RN(n869), 
        .Q(regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(n815), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(n813), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(i_data_Rd[2]), .E(n890), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(n809), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(n807), .E(n890), .C(i_clk), .RN(i_rst_n), .Q(
        regs[384]) );
  DFEC1 regs_reg_11__31_ ( .D(n860), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(i_data_Rd[30]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(i_data_Rd[29]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(i_data_Rd[28]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(i_data_Rd[27]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(i_data_Rd[26]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(n858), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(i_data_Rd[24]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(n854), .E(n891), .C(i_clk), .RN(n867), .Q(
        regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(i_data_Rd[22]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(n850), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(i_data_Rd[20]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(n846), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(i_data_Rd[18]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(n842), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(i_data_Rd[16]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(n838), .E(n891), .C(i_clk), .RN(n861), .Q(
        regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(n834), .E(n891), .C(i_clk), .RN(n862), .Q(
        regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(i_data_Rd[12]), .E(n891), .C(i_clk), .RN(n869), 
        .Q(regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(n830), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(i_data_Rd[10]), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(i_data_Rd[9]), .E(n891), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(i_data_Rd[8]), .E(n891), .C(i_clk), .RN(n863), 
        .Q(regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(n822), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(n820), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(i_data_Rd[5]), .E(n891), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(n815), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(n813), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(i_data_Rd[2]), .E(n891), .C(i_clk), .RN(n866), 
        .Q(regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(n809), .E(n891), .C(i_clk), .RN(n864), .Q(
        regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(n807), .E(n891), .C(i_clk), .RN(i_rst_n), .Q(
        regs[352]) );
  DFEC1 regs_reg_9__31_ ( .D(n860), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(i_data_Rd[30]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(i_data_Rd[29]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(i_data_Rd[28]), .E(n893), .C(i_clk), .RN(n861), 
        .Q(regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(i_data_Rd[27]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(i_data_Rd[26]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(n858), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(i_data_Rd[24]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(n854), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(i_data_Rd[22]), .E(n893), .C(i_clk), .RN(n864), 
        .Q(regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(n850), .E(n893), .C(i_clk), .RN(n862), .Q(
        regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(i_data_Rd[20]), .E(n893), .C(i_clk), .RN(n863), 
        .Q(regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(n846), .E(n893), .C(i_clk), .RN(n861), .Q(
        regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(i_data_Rd[18]), .E(n893), .C(i_clk), .RN(n862), 
        .Q(regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(n842), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(i_data_Rd[16]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(n838), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(i_data_Rd[14]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(n834), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(i_data_Rd[12]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(n830), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(i_data_Rd[10]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(i_data_Rd[9]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(i_data_Rd[8]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(n822), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(n820), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(i_data_Rd[5]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(n815), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(n813), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(i_data_Rd[2]), .E(n893), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(n809), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(n807), .E(n893), .C(i_clk), .RN(i_rst_n), .Q(
        regs[288]) );
  DFEC1 regs_reg_8__31_ ( .D(n860), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(i_data_Rd[30]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(i_data_Rd[29]), .E(n894), .C(i_clk), .RN(n862), 
        .Q(regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(i_data_Rd[28]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(i_data_Rd[27]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(i_data_Rd[26]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(n858), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(i_data_Rd[24]), .E(n894), .C(i_clk), .RN(n866), 
        .Q(regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(n854), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(i_data_Rd[22]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(n850), .E(n894), .C(i_clk), .RN(n861), .Q(
        regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(i_data_Rd[20]), .E(n894), .C(i_clk), .RN(n861), 
        .Q(regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(n846), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(i_data_Rd[18]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(n842), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(i_data_Rd[16]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(n838), .E(n894), .C(i_clk), .RN(n861), .Q(
        regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(i_data_Rd[14]), .E(n894), .C(i_clk), .RN(n863), 
        .Q(regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(n834), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(i_data_Rd[12]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(n830), .E(n894), .C(i_clk), .RN(n869), .Q(
        regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(i_data_Rd[10]), .E(n894), .C(i_clk), .RN(n866), 
        .Q(regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(i_data_Rd[9]), .E(n894), .C(i_clk), .RN(n861), .Q(
        regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(i_data_Rd[8]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(n822), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(n820), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(i_data_Rd[5]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(n815), .E(n894), .C(i_clk), .RN(n862), .Q(
        regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(n813), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(i_data_Rd[2]), .E(n894), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(n809), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(n807), .E(n894), .C(i_clk), .RN(i_rst_n), .Q(
        regs[256]) );
  DFEC1 regs_reg_7__31_ ( .D(n859), .E(n895), .C(i_clk), .RN(n864), .Q(
        regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(i_data_Rd[30]), .E(n895), .C(i_clk), .RN(n868), 
        .Q(regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(i_data_Rd[29]), .E(n895), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(i_data_Rd[28]), .E(n895), .C(i_clk), .RN(n868), 
        .Q(regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(i_data_Rd[27]), .E(n895), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(i_data_Rd[26]), .E(n895), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(n857), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(n855), .E(n895), .C(i_clk), .RN(n869), .Q(
        regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(n853), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(n851), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(n849), .E(n895), .C(i_clk), .RN(n867), .Q(
        regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(n847), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(n845), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(n843), .E(n895), .C(i_clk), .RN(n869), .Q(
        regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(n841), .E(n895), .C(i_clk), .RN(n868), .Q(
        regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(n839), .E(n895), .C(i_clk), .RN(n862), .Q(
        regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(n837), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(n835), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(n833), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(n831), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(n829), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(n827), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(n825), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(n823), .E(n895), .C(i_clk), .RN(n865), .Q(
        regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(n821), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(n819), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(n817), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(n814), .E(n895), .C(i_clk), .RN(n868), .Q(
        regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(n812), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(n810), .E(n895), .C(i_clk), .RN(i_rst_n), .Q(
        regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(n808), .E(n895), .C(i_clk), .RN(n865), .Q(
        regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(n806), .E(n895), .C(i_clk), .RN(n869), .Q(
        regs[224]) );
  DFEC1 regs_reg_5__31_ ( .D(n859), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(i_data_Rd[30]), .E(n897), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(i_data_Rd[29]), .E(n897), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(i_data_Rd[28]), .E(n897), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[188]) );
  DFEC1 regs_reg_5__27_ ( .D(i_data_Rd[27]), .E(n897), .C(i_clk), .RN(n865), 
        .Q(regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(i_data_Rd[26]), .E(n897), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(n857), .E(n897), .C(i_clk), .RN(n869), .Q(
        regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(n855), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(n853), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(n851), .E(n897), .C(i_clk), .RN(n863), .Q(
        regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(n849), .E(n897), .C(i_clk), .RN(n869), .Q(
        regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(n847), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(n845), .E(n897), .C(i_clk), .RN(n869), .Q(
        regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(n843), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(n841), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(n839), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(n837), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(n835), .E(n897), .C(i_clk), .RN(n863), .Q(
        regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(n833), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(n831), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(n829), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(n827), .E(n897), .C(i_clk), .RN(n864), .Q(
        regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(n825), .E(n897), .C(i_clk), .RN(n861), .Q(
        regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(n823), .E(n897), .C(i_clk), .RN(n865), .Q(
        regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(n821), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(n819), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(n817), .E(n897), .C(i_clk), .RN(n868), .Q(
        regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(n814), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(n812), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(n810), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(n808), .E(n897), .C(i_clk), .RN(i_rst_n), .Q(
        regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(n806), .E(n897), .C(i_clk), .RN(n867), .Q(
        regs[160]) );
  DFEC1 regs_reg_4__31_ ( .D(n859), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(i_data_Rd[30]), .E(n898), .C(i_clk), .RN(n867), 
        .Q(regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(i_data_Rd[29]), .E(n898), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(i_data_Rd[28]), .E(n898), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(i_data_Rd[27]), .E(n898), .C(i_clk), .RN(n865), 
        .Q(regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(i_data_Rd[26]), .E(n898), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(n857), .E(n898), .C(i_clk), .RN(n861), .Q(
        regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(n855), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(n853), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(n851), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(n849), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(n847), .E(n898), .C(i_clk), .RN(n866), .Q(
        regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(n845), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(n843), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(n841), .E(n898), .C(i_clk), .RN(n863), .Q(
        regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(n839), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(n837), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(n835), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(n833), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(n831), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(n829), .E(n898), .C(i_clk), .RN(n869), .Q(
        regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(n827), .E(n898), .C(i_clk), .RN(n868), .Q(
        regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(n825), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(n823), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(n821), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(n819), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(n817), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(n814), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(n812), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(n810), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(n808), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(n806), .E(n898), .C(i_clk), .RN(i_rst_n), .Q(
        regs[128]) );
  DFEC1 regs_reg_3__31_ ( .D(n859), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(i_data_Rd[30]), .E(n899), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(i_data_Rd[29]), .E(n899), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(i_data_Rd[28]), .E(n899), .C(i_clk), .RN(n862), 
        .Q(regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(i_data_Rd[27]), .E(n899), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(i_data_Rd[26]), .E(n899), .C(i_clk), .RN(n863), 
        .Q(regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(n857), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(n855), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(n853), .E(n899), .C(i_clk), .RN(n864), .Q(
        regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(n851), .E(n899), .C(i_clk), .RN(n862), .Q(
        regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(n849), .E(n899), .C(i_clk), .RN(n866), .Q(
        regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(n847), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(n845), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(n843), .E(n899), .C(i_clk), .RN(n868), .Q(
        regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(n841), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(n839), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(n837), .E(n899), .C(i_clk), .RN(n861), .Q(
        regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(n835), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(n833), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(n831), .E(n899), .C(i_clk), .RN(n868), .Q(
        regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(n829), .E(n899), .C(i_clk), .RN(n866), .Q(
        regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(n827), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(n825), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(n823), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(n821), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(n819), .E(n899), .C(i_clk), .RN(n862), .Q(
        regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(n817), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(n814), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(n812), .E(n899), .C(i_clk), .RN(n864), .Q(regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(n810), .E(n899), .C(i_clk), .RN(n869), .Q(regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(n808), .E(n899), .C(i_clk), .RN(i_rst_n), .Q(
        regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(n806), .E(n899), .C(i_clk), .RN(n861), .Q(regs[96]) );
  DFEC1 regs_reg_1__31_ ( .D(n859), .E(n901), .C(i_clk), .RN(n868), .Q(
        regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(i_data_Rd[30]), .E(n901), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(i_data_Rd[29]), .E(n901), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(i_data_Rd[28]), .E(n901), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(i_data_Rd[27]), .E(n901), .C(i_clk), .RN(n866), 
        .Q(regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(i_data_Rd[26]), .E(n901), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(n857), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(n855), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(n853), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(n851), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(n849), .E(n901), .C(i_clk), .RN(n868), .Q(
        regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(n847), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(n845), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(n843), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(n841), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(n839), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(n837), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(n835), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(n833), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(n831), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(n829), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(n827), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(n825), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(n823), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(n821), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(n819), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(n817), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(n814), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(n812), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(n810), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(n808), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(n806), .E(n901), .C(i_clk), .RN(i_rst_n), .Q(
        regs[32]) );
  DFEC1 regs_reg_0__31_ ( .D(n859), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(i_data_Rd[30]), .E(n902), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(i_data_Rd[29]), .E(n902), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(i_data_Rd[28]), .E(n902), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(i_data_Rd[27]), .E(n902), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(i_data_Rd[26]), .E(n902), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(n857), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(n855), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(n853), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(n851), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(n849), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(n847), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(n845), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(n843), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(n841), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(n839), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(n837), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(n835), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(n833), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(n831), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(n829), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(n827), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(n825), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(n823), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(n821), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(n819), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(n817), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(n814), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(n812), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(n810), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(n808), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(n806), .E(n902), .C(i_clk), .RN(i_rst_n), .Q(
        regs[0]) );
  IMUX41 U2 ( .A(n620), .B(n621), .C(n622), .D(n623), .S0(n749), .S1(n753), 
        .Q(n619) );
  IMUX41 U3 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n786), .S1(n776), .Q(n560) );
  IMUX41 U4 ( .A(n685), .B(n686), .C(n687), .D(n688), .S0(n746), .S1(n754), 
        .Q(n684) );
  CLKBU4 U5 ( .A(n783), .Q(n757) );
  BUF2 U6 ( .A(i_addr_Rs[0]), .Q(n805) );
  CLKBU4 U7 ( .A(n805), .Q(n800) );
  BUF6 U8 ( .A(n804), .Q(n798) );
  MUX22 U9 ( .A(n489), .B(n484), .S(n745), .Q(o_data_Rs[6]) );
  IMUX40 U10 ( .A(n485), .B(n486), .C(n487), .D(n488), .S0(n747), .S1(
        i_addr_Rs[2]), .Q(n484) );
  MUX22 U11 ( .A(n619), .B(n614), .S(i_addr_Rs[4]), .Q(o_data_Rs[19]) );
  IMUX40 U12 ( .A(n615), .B(n616), .C(n617), .D(n618), .S0(n749), .S1(n753), 
        .Q(n614) );
  MUX22 U13 ( .A(n459), .B(n454), .S(n744), .Q(o_data_Rs[3]) );
  IMUX40 U14 ( .A(n455), .B(n456), .C(n457), .D(n458), .S0(n747), .S1(n751), 
        .Q(n454) );
  IMUX40 U15 ( .A(n555), .B(n556), .C(n557), .D(n558), .S0(n748), .S1(n755), 
        .Q(n554) );
  BUF6 U16 ( .A(i_addr_Rs[0]), .Q(n803) );
  BUF6 U17 ( .A(n805), .Q(n786) );
  CLKBU4 U18 ( .A(n802), .Q(n796) );
  CLKBU4 U19 ( .A(n805), .Q(n791) );
  CLKBU4 U20 ( .A(n805), .Q(n788) );
  CLKBU4 U21 ( .A(n805), .Q(n787) );
  CLKBU4 U22 ( .A(n802), .Q(n790) );
  CLKBU4 U23 ( .A(n805), .Q(n801) );
  CLKBU4 U24 ( .A(n804), .Q(n799) );
  BUF2 U25 ( .A(i_addr_Rs[4]), .Q(n745) );
  BUF2 U26 ( .A(i_addr_Rt[4]), .Q(n366) );
  BUF2 U27 ( .A(n868), .Q(n867) );
  BUF2 U28 ( .A(n868), .Q(n866) );
  BUF2 U29 ( .A(n868), .Q(n865) );
  BUF2 U30 ( .A(n869), .Q(n864) );
  BUF2 U31 ( .A(n869), .Q(n863) );
  BUF2 U32 ( .A(n869), .Q(n862) );
  BUF2 U33 ( .A(n861), .Q(n868) );
  BUF2 U34 ( .A(n861), .Q(n869) );
  BUF2 U35 ( .A(n803), .Q(n789) );
  BUF2 U36 ( .A(n803), .Q(n792) );
  BUF2 U37 ( .A(n803), .Q(n793) );
  BUF2 U38 ( .A(n803), .Q(n794) );
  BUF2 U39 ( .A(n804), .Q(n795) );
  BUF2 U40 ( .A(n804), .Q(n797) );
  BUF2 U41 ( .A(n783), .Q(n762) );
  BUF2 U42 ( .A(n782), .Q(n763) );
  BUF2 U43 ( .A(n782), .Q(n764) );
  BUF2 U44 ( .A(n761), .Q(n765) );
  BUF2 U45 ( .A(n761), .Q(n766) );
  BUF2 U46 ( .A(n761), .Q(n767) );
  BUF2 U47 ( .A(n760), .Q(n768) );
  BUF2 U48 ( .A(n759), .Q(n769) );
  BUF2 U49 ( .A(n759), .Q(n770) );
  BUF2 U50 ( .A(n759), .Q(n771) );
  BUF2 U51 ( .A(n758), .Q(n772) );
  BUF2 U52 ( .A(n759), .Q(n773) );
  BUF2 U53 ( .A(n758), .Q(n774) );
  BUF2 U54 ( .A(n758), .Q(n775) );
  BUF2 U55 ( .A(n758), .Q(n776) );
  BUF2 U56 ( .A(n758), .Q(n777) );
  BUF2 U57 ( .A(n417), .Q(n396) );
  BUF2 U58 ( .A(n417), .Q(n397) );
  BUF2 U59 ( .A(n417), .Q(n398) );
  BUF2 U60 ( .A(n418), .Q(n399) );
  BUF2 U61 ( .A(n418), .Q(n400) );
  BUF2 U62 ( .A(n418), .Q(n401) );
  BUF2 U63 ( .A(n419), .Q(n402) );
  BUF2 U64 ( .A(n419), .Q(n403) );
  BUF2 U65 ( .A(n419), .Q(n404) );
  BUF2 U66 ( .A(n420), .Q(n405) );
  BUF2 U67 ( .A(n420), .Q(n406) );
  BUF2 U68 ( .A(n420), .Q(n407) );
  BUF2 U69 ( .A(n421), .Q(n408) );
  BUF2 U70 ( .A(n421), .Q(n409) );
  BUF2 U71 ( .A(n421), .Q(n410) );
  BUF2 U72 ( .A(n422), .Q(n411) );
  BUF2 U73 ( .A(n422), .Q(n412) );
  BUF2 U74 ( .A(n422), .Q(n413) );
  BUF2 U75 ( .A(n423), .Q(n414) );
  BUF2 U76 ( .A(n423), .Q(n415) );
  BUF2 U77 ( .A(n423), .Q(n416) );
  INV3 U78 ( .A(n55), .Q(n870) );
  NAND22 U79 ( .A(n41), .B(n56), .Q(n55) );
  BUF2 U80 ( .A(i_addr_Rt[1]), .Q(n382) );
  BUF2 U81 ( .A(n395), .Q(n383) );
  BUF2 U82 ( .A(n395), .Q(n384) );
  BUF2 U83 ( .A(n381), .Q(n385) );
  BUF2 U84 ( .A(n381), .Q(n386) );
  BUF2 U85 ( .A(n381), .Q(n387) );
  BUF2 U86 ( .A(n380), .Q(n388) );
  BUF2 U87 ( .A(n380), .Q(n389) );
  BUF2 U88 ( .A(n379), .Q(n390) );
  BUF2 U89 ( .A(n379), .Q(n391) );
  BUF2 U90 ( .A(n379), .Q(n392) );
  BUF2 U91 ( .A(n757), .Q(n778) );
  BUF2 U92 ( .A(n757), .Q(n779) );
  BUF2 U93 ( .A(i_rst_n), .Q(n861) );
  BUF2 U94 ( .A(i_addr_Rs[0]), .Q(n804) );
  BUF2 U95 ( .A(n784), .Q(n761) );
  BUF2 U96 ( .A(n784), .Q(n760) );
  BUF2 U97 ( .A(n784), .Q(n759) );
  BUF2 U98 ( .A(n783), .Q(n758) );
  NOR31 U99 ( .A(n907), .B(n886), .C(n903), .Q(n41) );
  NOR31 U100 ( .A(n905), .B(n906), .C(n904), .Q(n56) );
  INV3 U101 ( .A(n39), .Q(n878) );
  NAND22 U102 ( .A(n76), .B(n56), .Q(n39) );
  INV3 U103 ( .A(n40), .Q(n877) );
  NAND22 U104 ( .A(n41), .B(n42), .Q(n40) );
  INV3 U105 ( .A(n75), .Q(n885) );
  NAND22 U106 ( .A(n42), .B(n76), .Q(n75) );
  INV3 U107 ( .A(n77), .Q(n884) );
  NAND22 U108 ( .A(n44), .B(n76), .Q(n77) );
  INV3 U109 ( .A(n78), .Q(n883) );
  NAND22 U110 ( .A(n46), .B(n76), .Q(n78) );
  INV3 U111 ( .A(n79), .Q(n882) );
  NAND22 U112 ( .A(n48), .B(n76), .Q(n79) );
  INV3 U113 ( .A(n80), .Q(n881) );
  NAND22 U114 ( .A(n50), .B(n76), .Q(n80) );
  INV3 U115 ( .A(n81), .Q(n880) );
  NAND22 U116 ( .A(n52), .B(n76), .Q(n81) );
  INV3 U117 ( .A(n82), .Q(n879) );
  NAND22 U118 ( .A(n54), .B(n76), .Q(n82) );
  INV3 U119 ( .A(n43), .Q(n876) );
  NAND22 U120 ( .A(n44), .B(n41), .Q(n43) );
  INV3 U121 ( .A(n45), .Q(n875) );
  NAND22 U122 ( .A(n46), .B(n41), .Q(n45) );
  INV3 U123 ( .A(n47), .Q(n874) );
  NAND22 U124 ( .A(n48), .B(n41), .Q(n47) );
  INV3 U125 ( .A(n49), .Q(n873) );
  NAND22 U126 ( .A(n50), .B(n41), .Q(n49) );
  INV3 U127 ( .A(n51), .Q(n872) );
  NAND22 U128 ( .A(n52), .B(n41), .Q(n51) );
  INV3 U129 ( .A(n53), .Q(n871) );
  NAND22 U130 ( .A(n54), .B(n41), .Q(n53) );
  INV3 U131 ( .A(n57), .Q(n902) );
  NAND22 U132 ( .A(n58), .B(n42), .Q(n57) );
  INV3 U133 ( .A(n59), .Q(n901) );
  NAND22 U134 ( .A(n58), .B(n44), .Q(n59) );
  INV3 U135 ( .A(n60), .Q(n900) );
  NAND22 U136 ( .A(n58), .B(n46), .Q(n60) );
  INV3 U137 ( .A(n61), .Q(n899) );
  NAND22 U138 ( .A(n58), .B(n48), .Q(n61) );
  INV3 U139 ( .A(n62), .Q(n898) );
  NAND22 U140 ( .A(n58), .B(n50), .Q(n62) );
  INV3 U141 ( .A(n63), .Q(n897) );
  NAND22 U142 ( .A(n58), .B(n52), .Q(n63) );
  INV3 U143 ( .A(n64), .Q(n896) );
  NAND22 U144 ( .A(n58), .B(n54), .Q(n64) );
  INV3 U145 ( .A(n65), .Q(n895) );
  NAND22 U146 ( .A(n58), .B(n56), .Q(n65) );
  INV3 U147 ( .A(n66), .Q(n894) );
  NAND22 U148 ( .A(n67), .B(n42), .Q(n66) );
  INV3 U149 ( .A(n68), .Q(n893) );
  NAND22 U150 ( .A(n67), .B(n44), .Q(n68) );
  INV3 U151 ( .A(n69), .Q(n892) );
  NAND22 U152 ( .A(n67), .B(n46), .Q(n69) );
  INV3 U153 ( .A(n70), .Q(n891) );
  NAND22 U154 ( .A(n67), .B(n48), .Q(n70) );
  INV3 U155 ( .A(n71), .Q(n890) );
  NAND22 U156 ( .A(n67), .B(n50), .Q(n71) );
  INV3 U157 ( .A(n72), .Q(n889) );
  NAND22 U158 ( .A(n67), .B(n52), .Q(n72) );
  INV3 U159 ( .A(n73), .Q(n888) );
  NAND22 U160 ( .A(n67), .B(n54), .Q(n73) );
  INV3 U161 ( .A(n74), .Q(n887) );
  NAND22 U162 ( .A(n67), .B(n56), .Q(n74) );
  BUF2 U163 ( .A(n395), .Q(n393) );
  BUF2 U164 ( .A(n395), .Q(n394) );
  BUF2 U165 ( .A(n756), .Q(n780) );
  BUF2 U166 ( .A(n756), .Q(n781) );
  BUF2 U167 ( .A(n802), .Q(n785) );
  BUF2 U168 ( .A(i_addr_Rs[0]), .Q(n802) );
  BUF2 U169 ( .A(i_data_Rd[0]), .Q(n806) );
  BUF2 U170 ( .A(i_data_Rd[1]), .Q(n808) );
  BUF2 U171 ( .A(i_data_Rd[2]), .Q(n810) );
  BUF2 U172 ( .A(i_data_Rd[3]), .Q(n812) );
  BUF2 U173 ( .A(i_data_Rd[5]), .Q(n817) );
  BUF2 U174 ( .A(i_data_Rd[6]), .Q(n819) );
  BUF2 U175 ( .A(i_data_Rd[7]), .Q(n821) );
  BUF2 U176 ( .A(i_data_Rd[8]), .Q(n823) );
  BUF2 U177 ( .A(i_data_Rd[9]), .Q(n825) );
  BUF2 U178 ( .A(i_data_Rd[10]), .Q(n827) );
  BUF2 U179 ( .A(i_data_Rd[11]), .Q(n829) );
  BUF2 U180 ( .A(i_data_Rd[12]), .Q(n831) );
  BUF2 U181 ( .A(i_data_Rd[13]), .Q(n833) );
  BUF2 U182 ( .A(i_data_Rd[14]), .Q(n835) );
  BUF2 U183 ( .A(i_data_Rd[15]), .Q(n837) );
  BUF2 U184 ( .A(i_data_Rd[16]), .Q(n839) );
  BUF2 U185 ( .A(i_data_Rd[17]), .Q(n841) );
  BUF2 U186 ( .A(i_data_Rd[18]), .Q(n843) );
  BUF2 U187 ( .A(i_data_Rd[19]), .Q(n845) );
  BUF2 U188 ( .A(i_data_Rd[22]), .Q(n851) );
  BUF2 U189 ( .A(i_data_Rd[23]), .Q(n853) );
  BUF2 U190 ( .A(i_data_Rd[24]), .Q(n855) );
  BUF2 U191 ( .A(i_data_Rd[25]), .Q(n857) );
  BUF2 U192 ( .A(i_data_Rd[31]), .Q(n859) );
  BUF2 U193 ( .A(i_data_Rd[0]), .Q(n807) );
  BUF2 U194 ( .A(i_data_Rd[1]), .Q(n809) );
  BUF2 U195 ( .A(i_data_Rd[3]), .Q(n813) );
  BUF2 U196 ( .A(i_data_Rd[6]), .Q(n820) );
  BUF2 U197 ( .A(i_data_Rd[7]), .Q(n822) );
  BUF2 U198 ( .A(i_data_Rd[11]), .Q(n830) );
  BUF2 U199 ( .A(i_data_Rd[13]), .Q(n834) );
  BUF2 U200 ( .A(i_data_Rd[15]), .Q(n838) );
  BUF2 U201 ( .A(i_data_Rd[17]), .Q(n842) );
  BUF2 U202 ( .A(i_data_Rd[19]), .Q(n846) );
  BUF2 U203 ( .A(i_data_Rd[23]), .Q(n854) );
  BUF2 U204 ( .A(i_data_Rd[25]), .Q(n858) );
  BUF2 U205 ( .A(i_data_Rd[31]), .Q(n860) );
  BUF2 U206 ( .A(i_data_Rd[4]), .Q(n815) );
  BUF2 U207 ( .A(i_data_Rd[2]), .Q(n811) );
  BUF2 U208 ( .A(i_data_Rd[4]), .Q(n816) );
  BUF2 U209 ( .A(i_data_Rd[5]), .Q(n818) );
  BUF2 U210 ( .A(i_data_Rd[8]), .Q(n824) );
  BUF2 U211 ( .A(i_data_Rd[9]), .Q(n826) );
  BUF2 U212 ( .A(i_data_Rd[12]), .Q(n832) );
  BUF2 U213 ( .A(i_data_Rd[14]), .Q(n836) );
  BUF2 U214 ( .A(i_data_Rd[16]), .Q(n840) );
  BUF2 U215 ( .A(i_data_Rd[18]), .Q(n844) );
  BUF2 U216 ( .A(i_data_Rd[22]), .Q(n852) );
  BUF2 U217 ( .A(i_data_Rd[4]), .Q(n814) );
  BUF2 U218 ( .A(i_data_Rd[20]), .Q(n847) );
  BUF2 U219 ( .A(i_data_Rd[21]), .Q(n849) );
  BUF2 U220 ( .A(i_data_Rd[21]), .Q(n850) );
  BUF2 U221 ( .A(i_data_Rd[10]), .Q(n828) );
  BUF2 U222 ( .A(i_data_Rd[20]), .Q(n848) );
  BUF2 U223 ( .A(i_data_Rd[24]), .Q(n856) );
  BUF2 U224 ( .A(i_addr_Rt[0]), .Q(n417) );
  BUF2 U225 ( .A(i_addr_Rt[0]), .Q(n418) );
  BUF2 U226 ( .A(i_addr_Rt[0]), .Q(n419) );
  BUF2 U227 ( .A(i_addr_Rt[0]), .Q(n420) );
  BUF2 U228 ( .A(i_addr_Rt[0]), .Q(n421) );
  BUF2 U229 ( .A(i_addr_Rt[0]), .Q(n422) );
  BUF2 U230 ( .A(i_addr_Rt[0]), .Q(n423) );
  BUF2 U231 ( .A(i_addr_Rt[1]), .Q(n381) );
  BUF2 U232 ( .A(i_addr_Rt[1]), .Q(n380) );
  BUF2 U233 ( .A(i_addr_Rt[1]), .Q(n379) );
  IMUX40 U234 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n786), .S1(n761), .Q(n433) );
  IMUX40 U235 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n786), .S1(n760), .Q(n431) );
  IMUX40 U236 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n786), .S1(n784), .Q(n430) );
  IMUX40 U237 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(n785), .S1(n760), .Q(n428) );
  IMUX40 U238 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(n785), .S1(n762), .Q(n426) );
  IMUX40 U239 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n786), .S1(n756), .Q(n438) );
  IMUX40 U240 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n786), .S1(n757), .Q(n436) );
  IMUX40 U241 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n786), .S1(n759), .Q(n435) );
  IMUX40 U242 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n786), .S1(n759), .Q(n443) );
  IMUX40 U243 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n786), .S1(n766), .Q(n441) );
  IMUX40 U244 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n787), .S1(n763), .Q(n448) );
  IMUX40 U245 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n787), .S1(n758), .Q(n446) );
  IMUX40 U246 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n787), .S1(n764), .Q(n445) );
  IMUX40 U247 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n787), .S1(n782), .Q(n453) );
  IMUX40 U248 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n787), .S1(n762), .Q(n458) );
  IMUX40 U249 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n787), .S1(n759), .Q(n456) );
  IMUX40 U250 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n787), .S1(n767), .Q(n455) );
  IMUX40 U251 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n788), .S1(n757), .Q(n463) );
  IMUX40 U252 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n788), .S1(n760), .Q(n468) );
  IMUX40 U253 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n788), .S1(n758), .Q(n466) );
  IMUX40 U254 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n788), .S1(n759), .Q(n465) );
  IMUX40 U255 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n788), .S1(n783), .Q(n473) );
  IMUX40 U256 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n790), .S1(n782), .Q(n478) );
  IMUX40 U257 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n798), .S1(n764), .Q(n476) );
  IMUX40 U258 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n799), .S1(n783), .Q(n475) );
  IMUX40 U259 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n790), .S1(n782), .Q(n483) );
  IMUX40 U260 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n798), .S1(n759), .Q(n488) );
  IMUX40 U261 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n796), .S1(n762), .Q(n486) );
  IMUX40 U262 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n800), .S1(n762), .Q(n485) );
  IMUX40 U263 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n789), .S1(n762), .Q(n493) );
  IMUX40 U264 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n789), .S1(n762), .Q(n498) );
  IMUX40 U265 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n789), .S1(n762), .Q(n496) );
  IMUX40 U266 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n789), .S1(n763), .Q(n495) );
  IMUX40 U267 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n789), .S1(n763), .Q(n503) );
  IMUX40 U268 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n790), .S1(n763), .Q(n508) );
  IMUX40 U269 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n790), .S1(n763), .Q(n506) );
  IMUX40 U270 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n790), .S1(n764), .Q(n505) );
  IMUX40 U271 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n790), .S1(n764), .Q(n513) );
  IMUX40 U272 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n790), .S1(n764), .Q(n518) );
  IMUX40 U273 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n790), .S1(n764), .Q(n516) );
  IMUX40 U274 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n790), .S1(n764), .Q(n515) );
  IMUX40 U275 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n786), .S1(n765), .Q(n523) );
  IMUX40 U276 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n786), .S1(n765), .Q(n528) );
  IMUX40 U277 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n799), .S1(n765), .Q(n526) );
  IMUX40 U278 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n791), .S1(n765), .Q(n525) );
  IMUX40 U279 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n786), .S1(n765), .Q(n533) );
  IMUX40 U280 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n801), .S1(n766), .Q(n531) );
  IMUX40 U281 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n791), .S1(n766), .Q(n538) );
  IMUX40 U282 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n791), .S1(n766), .Q(n536) );
  IMUX40 U283 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n791), .S1(n766), .Q(n535) );
  IMUX40 U284 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n791), .S1(n766), .Q(n543) );
  IMUX40 U285 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n791), .S1(n766), .Q(n541) );
  IMUX40 U286 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n791), .S1(n767), .Q(n548) );
  IMUX40 U287 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n791), .S1(n767), .Q(n546) );
  IMUX40 U288 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n791), .S1(n767), .Q(n545) );
  IMUX40 U289 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n786), .S1(n767), .Q(n553) );
  IMUX40 U290 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n791), .S1(n767), .Q(n551) );
  IMUX40 U291 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n788), .S1(n762), .Q(n558) );
  IMUX40 U292 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n785), .S1(n760), .Q(n556) );
  IMUX40 U293 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n799), .S1(n775), .Q(n555) );
  IMUX40 U294 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n785), .S1(n764), .Q(n563) );
  IMUX40 U295 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n799), .S1(n762), .Q(n561) );
  IMUX40 U296 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n792), .S1(n768), .Q(n568) );
  IMUX40 U297 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n792), .S1(n768), .Q(n566) );
  IMUX40 U298 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n792), .S1(n768), .Q(n565) );
  IMUX40 U299 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n792), .S1(n768), .Q(n573) );
  IMUX40 U300 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n792), .S1(n768), .Q(n571) );
  IMUX40 U301 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n792), .S1(n768), .Q(n578) );
  IMUX40 U302 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n792), .S1(n778), .Q(n576) );
  IMUX40 U303 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n792), .S1(n763), .Q(n575) );
  IMUX40 U304 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n793), .S1(n781), .Q(n583) );
  IMUX40 U305 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n793), .S1(n772), .Q(n581) );
  IMUX40 U306 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n793), .S1(n760), .Q(n588) );
  IMUX40 U307 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n793), .S1(n767), .Q(n586) );
  IMUX40 U308 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n793), .S1(n769), .Q(n585) );
  IMUX40 U309 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n793), .S1(n769), .Q(n593) );
  IMUX40 U310 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n793), .S1(n769), .Q(n591) );
  IMUX40 U311 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n794), .S1(n769), .Q(n598) );
  IMUX40 U312 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n794), .S1(n769), .Q(n596) );
  IMUX40 U313 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n794), .S1(n770), .Q(n595) );
  IMUX40 U314 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n794), .S1(n770), .Q(n603) );
  IMUX40 U315 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n794), .S1(n770), .Q(n601) );
  IMUX40 U316 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n794), .S1(n770), .Q(n608) );
  IMUX40 U317 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n794), .S1(n770), .Q(n606) );
  IMUX40 U318 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n794), .S1(n770), .Q(n605) );
  IMUX40 U319 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n787), .S1(n771), .Q(n613) );
  IMUX40 U320 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n786), .S1(n771), .Q(n611) );
  IMUX40 U321 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n796), .S1(n771), .Q(n618) );
  IMUX40 U322 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n798), .S1(n771), .Q(n616) );
  IMUX40 U323 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n788), .S1(n771), .Q(n615) );
  IMUX40 U324 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n785), .S1(n771), .Q(n623) );
  IMUX40 U325 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n791), .S1(n772), .Q(n621) );
  IMUX40 U326 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n795), .S1(n772), .Q(n628) );
  IMUX40 U327 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n795), .S1(n772), .Q(n626) );
  IMUX40 U328 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n795), .S1(n772), .Q(n625) );
  IMUX40 U329 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n795), .S1(n772), .Q(n633) );
  IMUX40 U330 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n795), .S1(n772), .Q(n631) );
  IMUX40 U331 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n795), .S1(n773), .Q(n638) );
  IMUX40 U332 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n795), .S1(n773), .Q(n636) );
  IMUX40 U333 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n795), .S1(n773), .Q(n635) );
  IMUX40 U334 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n796), .S1(n773), .Q(n643) );
  IMUX40 U335 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n796), .S1(n773), .Q(n641) );
  IMUX40 U336 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n796), .S1(n774), .Q(n648) );
  IMUX40 U337 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n796), .S1(n774), .Q(n646) );
  IMUX40 U338 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n796), .S1(n774), .Q(n645) );
  IMUX40 U339 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n796), .S1(n774), .Q(n653) );
  IMUX40 U340 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n796), .S1(n774), .Q(n651) );
  IMUX40 U341 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n797), .S1(n775), .Q(n658) );
  IMUX40 U342 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n797), .S1(n775), .Q(n656) );
  IMUX40 U343 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n797), .S1(n775), .Q(n655) );
  IMUX40 U344 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n797), .S1(n775), .Q(n663) );
  IMUX40 U345 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n797), .S1(n775), .Q(n661) );
  IMUX40 U346 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n797), .S1(n775), .Q(n668) );
  IMUX40 U347 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n797), .S1(n776), .Q(n666) );
  IMUX40 U348 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n797), .S1(n776), .Q(n665) );
  IMUX40 U349 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n798), .S1(n776), .Q(n673) );
  IMUX40 U350 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n798), .S1(n776), .Q(n671) );
  IMUX40 U351 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n798), .S1(n776), .Q(n678) );
  IMUX40 U352 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n798), .S1(n776), .Q(n676) );
  IMUX40 U353 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n798), .S1(n777), .Q(n675) );
  IMUX40 U354 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n798), .S1(n777), .Q(n683) );
  IMUX40 U355 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n798), .S1(n777), .Q(n681) );
  IMUX40 U356 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n786), .S1(n765), .Q(n432) );
  IMUX40 U357 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n786), .S1(n763), .Q(n437) );
  IMUX40 U358 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n786), .S1(n767), .Q(n442) );
  IMUX40 U359 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n787), .S1(n757), .Q(n447) );
  IMUX40 U360 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n787), .S1(n763), .Q(n457) );
  IMUX40 U361 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n788), .S1(n757), .Q(n467) );
  IMUX40 U362 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n799), .S1(n756), .Q(n477) );
  IMUX40 U363 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n791), .S1(n762), .Q(n487) );
  IMUX40 U364 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n803), .S1(n763), .Q(n497) );
  IMUX40 U365 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n790), .S1(n763), .Q(n507) );
  IMUX40 U366 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n790), .S1(n764), .Q(n517) );
  IMUX40 U367 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n801), .S1(n765), .Q(n527) );
  IMUX40 U368 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n796), .S1(n766), .Q(n532) );
  IMUX40 U369 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n791), .S1(n766), .Q(n537) );
  IMUX40 U370 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n791), .S1(n767), .Q(n542) );
  IMUX40 U371 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n791), .S1(n767), .Q(n547) );
  IMUX40 U372 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n796), .S1(n767), .Q(n552) );
  IMUX40 U373 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n786), .S1(n762), .Q(n557) );
  IMUX40 U374 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n796), .S1(n780), .Q(n562) );
  IMUX40 U375 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n792), .S1(n768), .Q(n567) );
  IMUX40 U376 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n792), .S1(n768), .Q(n572) );
  IMUX40 U377 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n792), .S1(n779), .Q(n577) );
  IMUX40 U378 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n793), .S1(n766), .Q(n582) );
  IMUX40 U379 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n793), .S1(n769), .Q(n587) );
  IMUX40 U380 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n793), .S1(n769), .Q(n592) );
  IMUX40 U381 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n794), .S1(n769), .Q(n597) );
  IMUX40 U382 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n794), .S1(n770), .Q(n602) );
  IMUX40 U383 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n794), .S1(n770), .Q(n607) );
  IMUX40 U384 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n798), .S1(n771), .Q(n612) );
  IMUX40 U385 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n801), .S1(n771), .Q(n617) );
  IMUX40 U386 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n801), .S1(n772), .Q(n622) );
  IMUX40 U387 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n805), .S1(n772), .Q(n627) );
  IMUX40 U388 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n795), .S1(n773), .Q(n632) );
  IMUX40 U389 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n795), .S1(n773), .Q(n637) );
  IMUX40 U390 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n796), .S1(n773), .Q(n642) );
  IMUX40 U391 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n796), .S1(n774), .Q(n647) );
  IMUX40 U392 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n796), .S1(n774), .Q(n652) );
  IMUX40 U393 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(i_addr_Rs[0]), .S1(n775), .Q(n657) );
  IMUX40 U394 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n797), .S1(n775), .Q(n662) );
  IMUX40 U395 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n797), .S1(n776), .Q(n667) );
  IMUX40 U396 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n798), .S1(n776), .Q(n672) );
  IMUX40 U397 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n798), .S1(n777), .Q(n677) );
  IMUX40 U398 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n798), .S1(n777), .Q(n682) );
  MUX22 U399 ( .A(n429), .B(n424), .S(n744), .Q(o_data_Rs[0]) );
  IMUX40 U400 ( .A(n425), .B(n426), .C(n427), .D(n428), .S0(n746), .S1(n752), 
        .Q(n424) );
  IMUX40 U401 ( .A(n430), .B(n431), .C(n432), .D(n433), .S0(n746), .S1(n751), 
        .Q(n429) );
  MUX22 U402 ( .A(n439), .B(n434), .S(n744), .Q(o_data_Rs[1]) );
  IMUX40 U403 ( .A(n440), .B(n441), .C(n442), .D(n443), .S0(n746), .S1(n751), 
        .Q(n439) );
  IMUX40 U404 ( .A(n435), .B(n436), .C(n437), .D(n438), .S0(n746), .S1(n751), 
        .Q(n434) );
  IMUX40 U405 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n786), .S1(n762), .Q(n440) );
  MUX22 U406 ( .A(n449), .B(n444), .S(n744), .Q(o_data_Rs[2]) );
  IMUX40 U407 ( .A(n450), .B(n451), .C(n452), .D(n453), .S0(n747), .S1(n751), 
        .Q(n449) );
  IMUX40 U408 ( .A(n445), .B(n446), .C(n447), .D(n448), .S0(n747), .S1(n751), 
        .Q(n444) );
  IMUX40 U409 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n787), .S1(n782), .Q(n452) );
  IMUX40 U410 ( .A(n460), .B(n461), .C(n462), .D(n463), .S0(n747), .S1(n751), 
        .Q(n459) );
  IMUX40 U411 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n788), .S1(n760), .Q(n460) );
  MUX22 U412 ( .A(n469), .B(n464), .S(n744), .Q(o_data_Rs[4]) );
  IMUX40 U413 ( .A(n470), .B(n471), .C(n472), .D(n473), .S0(n747), .S1(n751), 
        .Q(n469) );
  IMUX40 U414 ( .A(n465), .B(n466), .C(n467), .D(n468), .S0(n747), .S1(n751), 
        .Q(n464) );
  IMUX40 U415 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n788), .S1(n760), .Q(n470) );
  MUX22 U416 ( .A(n479), .B(n474), .S(n744), .Q(o_data_Rs[5]) );
  IMUX40 U417 ( .A(n480), .B(n481), .C(n482), .D(n483), .S0(n747), .S1(
        i_addr_Rs[2]), .Q(n479) );
  IMUX40 U418 ( .A(n475), .B(n476), .C(n477), .D(n478), .S0(n747), .S1(n751), 
        .Q(n474) );
  IMUX40 U419 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n790), .S1(n767), .Q(n480) );
  IMUX40 U420 ( .A(n490), .B(n491), .C(n492), .D(n493), .S0(n747), .S1(
        i_addr_Rs[2]), .Q(n489) );
  IMUX40 U421 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n789), .S1(n762), .Q(n490) );
  MUX22 U422 ( .A(n499), .B(n494), .S(n745), .Q(o_data_Rs[7]) );
  IMUX40 U423 ( .A(n500), .B(n501), .C(n502), .D(n503), .S0(n747), .S1(
        i_addr_Rs[2]), .Q(n499) );
  IMUX40 U424 ( .A(n495), .B(n496), .C(n497), .D(n498), .S0(n747), .S1(n752), 
        .Q(n494) );
  IMUX40 U425 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n789), .S1(n763), .Q(n500) );
  MUX22 U426 ( .A(n509), .B(n504), .S(n745), .Q(o_data_Rs[8]) );
  IMUX40 U427 ( .A(n510), .B(n511), .C(n512), .D(n513), .S0(n748), .S1(n753), 
        .Q(n509) );
  IMUX40 U428 ( .A(n505), .B(n506), .C(n507), .D(n508), .S0(n748), .S1(n751), 
        .Q(n504) );
  IMUX40 U429 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n790), .S1(n764), .Q(n510) );
  MUX22 U430 ( .A(n519), .B(n514), .S(n745), .Q(o_data_Rs[9]) );
  IMUX40 U431 ( .A(n520), .B(n521), .C(n522), .D(n523), .S0(n748), .S1(n753), 
        .Q(n519) );
  IMUX40 U432 ( .A(n515), .B(n516), .C(n517), .D(n518), .S0(n748), .S1(n752), 
        .Q(n514) );
  IMUX40 U433 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n785), .S1(n765), .Q(n520) );
  BUF2 U434 ( .A(i_addr_Rs[1]), .Q(n784) );
  BUF2 U435 ( .A(i_addr_Rs[1]), .Q(n783) );
  MUX22 U436 ( .A(n529), .B(n524), .S(n745), .Q(o_data_Rs[10]) );
  IMUX40 U437 ( .A(n530), .B(n531), .C(n532), .D(n533), .S0(n748), .S1(n755), 
        .Q(n529) );
  IMUX40 U438 ( .A(n525), .B(n526), .C(n527), .D(n528), .S0(n748), .S1(n755), 
        .Q(n524) );
  IMUX40 U439 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n786), .S1(n766), .Q(n530) );
  MUX22 U440 ( .A(n539), .B(n534), .S(n745), .Q(o_data_Rs[11]) );
  IMUX40 U441 ( .A(n540), .B(n541), .C(n542), .D(n543), .S0(n748), .S1(n754), 
        .Q(n539) );
  IMUX40 U442 ( .A(n535), .B(n536), .C(n537), .D(n538), .S0(n748), .S1(n754), 
        .Q(n534) );
  IMUX40 U443 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n791), .S1(n767), .Q(n540) );
  MUX22 U444 ( .A(n549), .B(n544), .S(n745), .Q(o_data_Rs[12]) );
  IMUX40 U445 ( .A(n550), .B(n551), .C(n552), .D(n553), .S0(n748), .S1(n754), 
        .Q(n549) );
  IMUX40 U446 ( .A(n545), .B(n546), .C(n547), .D(n548), .S0(n748), .S1(n754), 
        .Q(n544) );
  IMUX40 U447 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n786), .S1(n760), .Q(n550) );
  MUX22 U448 ( .A(n559), .B(n554), .S(n745), .Q(o_data_Rs[13]) );
  IMUX40 U449 ( .A(n560), .B(n561), .C(n562), .D(n563), .S0(n748), .S1(n755), 
        .Q(n559) );
  MUX22 U450 ( .A(n569), .B(n564), .S(n745), .Q(o_data_Rs[14]) );
  IMUX40 U451 ( .A(n570), .B(n571), .C(n572), .D(n573), .S0(n749), .S1(n752), 
        .Q(n569) );
  IMUX40 U452 ( .A(n565), .B(n566), .C(n567), .D(n568), .S0(n749), .S1(n752), 
        .Q(n564) );
  IMUX40 U453 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n792), .S1(n768), .Q(n570) );
  MUX22 U454 ( .A(n579), .B(n574), .S(n745), .Q(o_data_Rs[15]) );
  IMUX40 U455 ( .A(n580), .B(n581), .C(n582), .D(n583), .S0(n749), .S1(n752), 
        .Q(n579) );
  IMUX40 U456 ( .A(n575), .B(n576), .C(n577), .D(n578), .S0(n749), .S1(n752), 
        .Q(n574) );
  IMUX40 U457 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n793), .S1(n765), .Q(n580) );
  MUX22 U458 ( .A(n589), .B(n584), .S(n745), .Q(o_data_Rs[16]) );
  IMUX40 U459 ( .A(n590), .B(n591), .C(n592), .D(n593), .S0(n749), .S1(n752), 
        .Q(n589) );
  IMUX40 U460 ( .A(n585), .B(n586), .C(n587), .D(n588), .S0(n749), .S1(n752), 
        .Q(n584) );
  IMUX40 U461 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n793), .S1(n769), .Q(n590) );
  MUX22 U462 ( .A(n599), .B(n594), .S(n745), .Q(o_data_Rs[17]) );
  IMUX40 U463 ( .A(n600), .B(n601), .C(n602), .D(n603), .S0(n749), .S1(n752), 
        .Q(n599) );
  IMUX40 U464 ( .A(n595), .B(n596), .C(n597), .D(n598), .S0(n749), .S1(n752), 
        .Q(n594) );
  IMUX40 U465 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n794), .S1(n770), .Q(n600) );
  MUX22 U466 ( .A(n609), .B(n604), .S(n745), .Q(o_data_Rs[18]) );
  IMUX40 U467 ( .A(n610), .B(n611), .C(n612), .D(n613), .S0(n749), .S1(n753), 
        .Q(n609) );
  IMUX40 U468 ( .A(n605), .B(n606), .C(n607), .D(n608), .S0(n749), .S1(n752), 
        .Q(n604) );
  IMUX40 U469 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n796), .S1(n771), .Q(n610) );
  IMUX40 U470 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n802), .S1(n772), .Q(n620) );
  MUX22 U471 ( .A(n629), .B(n624), .S(n744), .Q(o_data_Rs[20]) );
  IMUX40 U472 ( .A(n630), .B(n631), .C(n632), .D(n633), .S0(n750), .S1(n753), 
        .Q(n629) );
  IMUX40 U473 ( .A(n625), .B(n626), .C(n627), .D(n628), .S0(n750), .S1(n753), 
        .Q(n624) );
  IMUX40 U474 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n795), .S1(n773), .Q(n630) );
  MUX22 U475 ( .A(n639), .B(n634), .S(n744), .Q(o_data_Rs[21]) );
  IMUX40 U476 ( .A(n640), .B(n641), .C(n642), .D(n643), .S0(n750), .S1(n753), 
        .Q(n639) );
  IMUX40 U477 ( .A(n635), .B(n636), .C(n637), .D(n638), .S0(n750), .S1(n753), 
        .Q(n634) );
  IMUX40 U478 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n796), .S1(n774), .Q(n640) );
  MUX22 U479 ( .A(n649), .B(n644), .S(n744), .Q(o_data_Rs[22]) );
  IMUX40 U480 ( .A(n650), .B(n651), .C(n652), .D(n653), .S0(n750), .S1(n753), 
        .Q(n649) );
  IMUX40 U481 ( .A(n645), .B(n646), .C(n647), .D(n648), .S0(n750), .S1(n753), 
        .Q(n644) );
  IMUX40 U482 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n796), .S1(n774), .Q(n650) );
  MUX22 U483 ( .A(n659), .B(n654), .S(n744), .Q(o_data_Rs[23]) );
  IMUX40 U484 ( .A(n660), .B(n661), .C(n662), .D(n663), .S0(n750), .S1(n754), 
        .Q(n659) );
  IMUX40 U485 ( .A(n655), .B(n656), .C(n657), .D(n658), .S0(n750), .S1(n754), 
        .Q(n654) );
  IMUX40 U486 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n797), .S1(n775), .Q(n660) );
  MUX22 U487 ( .A(n669), .B(n664), .S(n744), .Q(o_data_Rs[24]) );
  IMUX40 U488 ( .A(n670), .B(n671), .C(n672), .D(n673), .S0(n750), .S1(n754), 
        .Q(n669) );
  IMUX40 U489 ( .A(n665), .B(n666), .C(n667), .D(n668), .S0(n750), .S1(n754), 
        .Q(n664) );
  IMUX40 U490 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n798), .S1(n776), .Q(n670) );
  MUX22 U491 ( .A(n679), .B(n674), .S(n744), .Q(o_data_Rs[25]) );
  IMUX40 U492 ( .A(n680), .B(n681), .C(n682), .D(n683), .S0(n750), .S1(n754), 
        .Q(n679) );
  IMUX40 U493 ( .A(n675), .B(n676), .C(n677), .D(n678), .S0(n750), .S1(n754), 
        .Q(n674) );
  IMUX40 U494 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n798), .S1(n777), .Q(n680) );
  NOR31 U495 ( .A(n886), .B(i_addr_Rd[3]), .C(n907), .Q(n76) );
  NOR31 U496 ( .A(i_addr_Rd[3]), .B(i_addr_Rd[4]), .C(n907), .Q(n58) );
  NOR31 U497 ( .A(n907), .B(i_addr_Rd[4]), .C(n903), .Q(n67) );
  NOR31 U498 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(i_addr_Rd[0]), .Q(n42)
         );
  NOR31 U499 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n904), .Q(n50) );
  NOR31 U500 ( .A(n906), .B(i_addr_Rd[1]), .C(n904), .Q(n52) );
  NOR31 U501 ( .A(n905), .B(i_addr_Rd[0]), .C(n904), .Q(n54) );
  NOR31 U502 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(n906), .Q(n44) );
  NOR31 U503 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[2]), .C(n905), .Q(n46) );
  NOR31 U504 ( .A(n906), .B(i_addr_Rd[2]), .C(n905), .Q(n48) );
  IMUX40 U505 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n396), .S1(n381), .Q(n10) );
  IMUX40 U506 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n396), .S1(i_addr_Rt[1]), .Q(n8) );
  IMUX40 U507 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n396), .S1(i_addr_Rt[1]), .Q(n7) );
  IMUX40 U508 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(i_addr_Rt[0]), .S1(n395), .Q(n5) );
  IMUX40 U509 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(i_addr_Rt[0]), .S1(n383), .Q(n3) );
  IMUX40 U510 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(i_addr_Rt[0]), .S1(n386), .Q(n2) );
  IMUX40 U511 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n396), .S1(n387), .Q(n15) );
  IMUX40 U512 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n396), .S1(i_addr_Rt[1]), .Q(n13) );
  IMUX40 U513 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n396), .S1(i_addr_Rt[1]), .Q(n12) );
  IMUX40 U514 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n396), .S1(n395), .Q(n20) );
  IMUX40 U515 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n396), .S1(i_addr_Rt[1]), .Q(n18) );
  IMUX40 U516 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n397), .S1(n383), .Q(n25) );
  IMUX40 U517 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n397), .S1(n380), .Q(n23) );
  IMUX40 U518 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n397), .S1(n380), .Q(n22) );
  IMUX40 U519 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n397), .S1(n382), .Q(n30) );
  IMUX40 U520 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n397), .S1(n383), .Q(n28) );
  IMUX40 U521 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n397), .S1(n393), .Q(n35) );
  IMUX40 U522 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n397), .S1(i_addr_Rt[1]), .Q(n33) );
  IMUX40 U523 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n397), .S1(i_addr_Rt[1]), .Q(n32) );
  IMUX40 U524 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n398), .S1(n384), .Q(n84) );
  IMUX40 U525 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n398), .S1(i_addr_Rt[1]), .Q(n38) );
  IMUX40 U526 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n398), .S1(n382), .Q(n89) );
  IMUX40 U527 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n398), .S1(n379), .Q(n87) );
  IMUX40 U528 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n398), .S1(n380), .Q(n86) );
  IMUX40 U529 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n398), .S1(n384), .Q(n94) );
  IMUX40 U530 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n398), .S1(n383), .Q(n92) );
  IMUX40 U531 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n399), .S1(n380), .Q(n99) );
  IMUX40 U532 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n399), .S1(n394), .Q(n97) );
  IMUX40 U533 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n399), .S1(n385), .Q(n96) );
  IMUX40 U534 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n399), .S1(n395), .Q(n104) );
  IMUX40 U535 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n399), .S1(n380), .Q(n102) );
  IMUX40 U536 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n399), .S1(n393), .Q(n109) );
  IMUX40 U537 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n399), .S1(n382), .Q(n107) );
  IMUX40 U538 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n399), .S1(n382), .Q(n106) );
  IMUX40 U539 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n400), .S1(n382), .Q(n114) );
  IMUX40 U540 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n400), .S1(n382), .Q(n112) );
  IMUX40 U541 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n400), .S1(n382), .Q(n119) );
  IMUX40 U542 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n400), .S1(n382), .Q(n117) );
  IMUX40 U543 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n400), .S1(n381), .Q(n116) );
  IMUX40 U544 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n400), .S1(n379), .Q(n124) );
  IMUX40 U545 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n400), .S1(n379), .Q(n122) );
  IMUX40 U546 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n401), .S1(n382), .Q(n129) );
  IMUX40 U547 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n401), .S1(n382), .Q(n127) );
  IMUX40 U548 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n401), .S1(n383), .Q(n126) );
  IMUX40 U549 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n401), .S1(n381), .Q(n134) );
  IMUX40 U550 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n401), .S1(n381), .Q(n132) );
  IMUX40 U551 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n401), .S1(n382), .Q(n139) );
  IMUX40 U552 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n401), .S1(n382), .Q(n137) );
  IMUX40 U553 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n401), .S1(n383), .Q(n136) );
  IMUX40 U554 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n402), .S1(n383), .Q(n144) );
  IMUX40 U555 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n402), .S1(n383), .Q(n142) );
  IMUX40 U556 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n402), .S1(n383), .Q(n149) );
  IMUX40 U557 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n402), .S1(n383), .Q(n147) );
  IMUX40 U558 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n402), .S1(n383), .Q(n146) );
  IMUX40 U559 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n402), .S1(n383), .Q(n154) );
  IMUX40 U560 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n402), .S1(n395), .Q(n152) );
  IMUX40 U561 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n403), .S1(n385), .Q(n159) );
  IMUX40 U562 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n403), .S1(n395), .Q(n157) );
  IMUX40 U563 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n403), .S1(n379), .Q(n156) );
  IMUX40 U564 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n403), .S1(n381), .Q(n164) );
  IMUX40 U565 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n403), .S1(n381), .Q(n162) );
  IMUX40 U566 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n403), .S1(n379), .Q(n169) );
  IMUX40 U567 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n403), .S1(n379), .Q(n167) );
  IMUX40 U568 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n403), .S1(n384), .Q(n166) );
  IMUX40 U569 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n404), .S1(n380), .Q(n174) );
  IMUX40 U570 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n404), .S1(n379), .Q(n172) );
  IMUX40 U571 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n404), .S1(n394), .Q(n179) );
  IMUX40 U572 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n404), .S1(n384), .Q(n177) );
  IMUX40 U573 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n404), .S1(n383), .Q(n176) );
  IMUX40 U574 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n404), .S1(n381), .Q(n184) );
  IMUX40 U575 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n404), .S1(n395), .Q(n182) );
  IMUX40 U576 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n405), .S1(n384), .Q(n189) );
  IMUX40 U577 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n405), .S1(n384), .Q(n187) );
  IMUX40 U578 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n405), .S1(n384), .Q(n186) );
  IMUX40 U579 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n405), .S1(n384), .Q(n194) );
  IMUX40 U580 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n405), .S1(n384), .Q(n192) );
  IMUX40 U581 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n405), .S1(n384), .Q(n199) );
  IMUX40 U582 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n405), .S1(n380), .Q(n197) );
  IMUX40 U583 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n405), .S1(n379), .Q(n196) );
  IMUX40 U584 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n406), .S1(n380), .Q(n204) );
  IMUX40 U585 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n406), .S1(n379), .Q(n202) );
  IMUX40 U586 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n406), .S1(n380), .Q(n209) );
  IMUX40 U587 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n406), .S1(n379), .Q(n207) );
  IMUX40 U588 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n406), .S1(n385), .Q(n206) );
  IMUX40 U589 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n406), .S1(n385), .Q(n214) );
  IMUX40 U590 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n406), .S1(n385), .Q(n212) );
  IMUX40 U591 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n407), .S1(n385), .Q(n219) );
  IMUX40 U592 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n407), .S1(n385), .Q(n217) );
  IMUX40 U593 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n407), .S1(n386), .Q(n216) );
  IMUX40 U594 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n407), .S1(n386), .Q(n224) );
  IMUX40 U595 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n407), .S1(n386), .Q(n222) );
  IMUX40 U596 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n407), .S1(n386), .Q(n229) );
  IMUX40 U597 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n407), .S1(n386), .Q(n227) );
  IMUX40 U598 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n407), .S1(n386), .Q(n226) );
  IMUX40 U599 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n408), .S1(n379), .Q(n234) );
  IMUX40 U600 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n408), .S1(n386), .Q(n232) );
  IMUX40 U601 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n408), .S1(n379), .Q(n239) );
  IMUX40 U602 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n408), .S1(n380), .Q(n237) );
  IMUX40 U603 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n408), .S1(n382), .Q(n236) );
  IMUX40 U604 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n408), .S1(n385), .Q(n244) );
  IMUX40 U605 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n408), .S1(n383), .Q(n242) );
  IMUX40 U606 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n409), .S1(n386), .Q(n249) );
  IMUX40 U607 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n409), .S1(n379), .Q(n247) );
  IMUX40 U608 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n409), .S1(n382), .Q(n246) );
  IMUX40 U609 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n409), .S1(n381), .Q(n254) );
  IMUX40 U610 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n409), .S1(n381), .Q(n252) );
  IMUX40 U611 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n409), .S1(n380), .Q(n259) );
  IMUX40 U612 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n409), .S1(n382), .Q(n257) );
  IMUX40 U613 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n409), .S1(n382), .Q(n256) );
  IMUX40 U614 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n410), .S1(n380), .Q(n264) );
  IMUX40 U615 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n410), .S1(n381), .Q(n262) );
  IMUX40 U616 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n410), .S1(n387), .Q(n269) );
  IMUX40 U617 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n410), .S1(n387), .Q(n267) );
  IMUX40 U618 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n410), .S1(n387), .Q(n266) );
  IMUX40 U619 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n410), .S1(n387), .Q(n274) );
  IMUX40 U620 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n410), .S1(n387), .Q(n272) );
  IMUX40 U621 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n411), .S1(n388), .Q(n279) );
  IMUX40 U622 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n411), .S1(n388), .Q(n277) );
  IMUX40 U623 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n411), .S1(n388), .Q(n276) );
  IMUX40 U624 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n411), .S1(n388), .Q(n284) );
  IMUX40 U625 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n411), .S1(n388), .Q(n282) );
  IMUX40 U626 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n411), .S1(n388), .Q(n289) );
  IMUX40 U627 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n411), .S1(n389), .Q(n287) );
  IMUX40 U628 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n411), .S1(n389), .Q(n286) );
  IMUX40 U629 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n412), .S1(n389), .Q(n294) );
  IMUX40 U630 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n412), .S1(n389), .Q(n292) );
  IMUX40 U631 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n412), .S1(n389), .Q(n299) );
  IMUX40 U632 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n412), .S1(n389), .Q(n297) );
  IMUX40 U633 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n412), .S1(n394), .Q(n296) );
  IMUX40 U634 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n412), .S1(n394), .Q(n304) );
  IMUX40 U635 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n412), .S1(n393), .Q(n302) );
  IMUX40 U636 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n413), .S1(n393), .Q(n309) );
  IMUX40 U637 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n413), .S1(n394), .Q(n307) );
  IMUX40 U638 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n413), .S1(n390), .Q(n306) );
  IMUX40 U639 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n413), .S1(n390), .Q(n314) );
  IMUX40 U640 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n413), .S1(n390), .Q(n312) );
  IMUX40 U641 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n413), .S1(n390), .Q(n319) );
  IMUX40 U642 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n413), .S1(n390), .Q(n317) );
  IMUX40 U643 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n413), .S1(n390), .Q(n316) );
  IMUX40 U644 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n414), .S1(n391), .Q(n324) );
  IMUX40 U645 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n414), .S1(n391), .Q(n322) );
  IMUX40 U646 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n414), .S1(n391), .Q(n329) );
  IMUX40 U647 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n414), .S1(n391), .Q(n327) );
  IMUX40 U648 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n414), .S1(n391), .Q(n326) );
  IMUX40 U649 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n414), .S1(n391), .Q(n334) );
  IMUX40 U650 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n414), .S1(n392), .Q(n332) );
  IMUX40 U651 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n415), .S1(n392), .Q(n339) );
  IMUX40 U652 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n415), .S1(n392), .Q(n337) );
  IMUX40 U653 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n415), .S1(n392), .Q(n336) );
  IMUX40 U654 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n415), .S1(n392), .Q(n344) );
  IMUX40 U655 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n415), .S1(n392), .Q(n342) );
  IMUX40 U656 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n415), .S1(n393), .Q(n349) );
  IMUX40 U657 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n415), .S1(n393), .Q(n347) );
  IMUX40 U658 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n415), .S1(n393), .Q(n346) );
  IMUX40 U659 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n416), .S1(n393), .Q(n354) );
  IMUX40 U660 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n416), .S1(n393), .Q(n352) );
  IMUX40 U661 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n416), .S1(n394), .Q(n359) );
  IMUX40 U662 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n416), .S1(n394), .Q(n357) );
  IMUX40 U663 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n416), .S1(n394), .Q(n356) );
  IMUX40 U664 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n416), .S1(n394), .Q(n364) );
  IMUX40 U665 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n416), .S1(n394), .Q(n362) );
  IMUX40 U666 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(n785), .S1(n760), .Q(n425) );
  IMUX40 U667 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n787), .S1(n764), .Q(n451) );
  IMUX40 U668 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n787), .S1(n783), .Q(n450) );
  IMUX40 U669 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n788), .S1(n766), .Q(n461) );
  IMUX40 U670 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n788), .S1(n759), .Q(n471) );
  IMUX40 U671 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n798), .S1(n760), .Q(n481) );
  IMUX40 U672 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n789), .S1(n762), .Q(n491) );
  IMUX40 U673 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n789), .S1(n763), .Q(n501) );
  IMUX40 U674 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n790), .S1(n764), .Q(n511) );
  IMUX40 U675 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n786), .S1(n765), .Q(n521) );
  IMUX40 U676 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n799), .S1(n777), .Q(n688) );
  IMUX40 U677 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n799), .S1(n777), .Q(n686) );
  IMUX40 U678 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n799), .S1(n774), .Q(n685) );
  IMUX40 U679 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n799), .S1(n757), .Q(n693) );
  IMUX40 U680 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n799), .S1(n780), .Q(n691) );
  IMUX40 U681 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n799), .S1(n766), .Q(n698) );
  IMUX40 U682 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n799), .S1(n776), .Q(n696) );
  IMUX40 U683 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n799), .S1(n777), .Q(n695) );
  IMUX40 U684 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n798), .S1(n778), .Q(n703) );
  IMUX40 U685 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n798), .S1(n778), .Q(n701) );
  IMUX40 U686 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n798), .S1(n778), .Q(n708) );
  IMUX40 U687 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n798), .S1(n778), .Q(n706) );
  IMUX40 U688 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n798), .S1(n778), .Q(n705) );
  IMUX40 U689 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n798), .S1(n778), .Q(n713) );
  IMUX40 U690 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n798), .S1(n779), .Q(n711) );
  IMUX40 U691 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n800), .S1(n779), .Q(n718) );
  IMUX40 U692 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n800), .S1(n779), .Q(n716) );
  IMUX40 U693 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n800), .S1(n779), .Q(n715) );
  IMUX40 U694 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n800), .S1(n779), .Q(n723) );
  IMUX40 U695 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n800), .S1(n779), .Q(n721) );
  IMUX40 U696 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n800), .S1(n780), .Q(n720) );
  IMUX40 U697 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n800), .S1(n780), .Q(n728) );
  IMUX40 U698 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n800), .S1(n780), .Q(n726) );
  IMUX40 U699 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n800), .S1(n780), .Q(n725) );
  IMUX40 U700 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n801), .S1(n780), .Q(n733) );
  IMUX40 U701 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n801), .S1(n781), .Q(n730) );
  IMUX40 U702 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n801), .S1(n780), .Q(n731) );
  IMUX40 U703 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n801), .S1(n781), .Q(n738) );
  IMUX40 U704 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n801), .S1(n781), .Q(n736) );
  IMUX40 U705 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n801), .S1(n781), .Q(n735) );
  IMUX40 U706 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n801), .S1(n781), .Q(n743) );
  IMUX40 U707 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n801), .S1(n781), .Q(n740) );
  IMUX40 U708 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n801), .S1(n781), .Q(n741) );
  IMUX40 U709 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n396), .S1(n382), .Q(n9) );
  IMUX40 U710 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(i_addr_Rt[0]), .S1(n382), .Q(n4) );
  IMUX40 U711 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n396), .S1(n395), .Q(n14) );
  IMUX40 U712 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n396), .S1(n386), .Q(n19) );
  IMUX40 U713 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n397), .S1(n387), .Q(n24) );
  IMUX40 U714 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n397), .S1(n380), .Q(n29) );
  IMUX40 U715 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n397), .S1(n382), .Q(n34) );
  IMUX40 U716 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n398), .S1(n381), .Q(n83) );
  IMUX40 U717 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n398), .S1(n382), .Q(n88) );
  IMUX40 U718 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n398), .S1(n385), .Q(n93) );
  IMUX40 U719 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n399), .S1(n382), .Q(n98) );
  IMUX40 U720 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n399), .S1(n387), .Q(n103) );
  IMUX40 U721 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n399), .S1(n382), .Q(n108) );
  IMUX40 U722 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n400), .S1(n382), .Q(n113) );
  IMUX40 U723 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n400), .S1(n387), .Q(n118) );
  IMUX40 U724 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n400), .S1(n395), .Q(n123) );
  IMUX40 U725 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n401), .S1(n381), .Q(n128) );
  IMUX40 U726 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n401), .S1(n382), .Q(n133) );
  IMUX40 U727 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n401), .S1(n382), .Q(n138) );
  IMUX40 U728 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n402), .S1(n383), .Q(n143) );
  IMUX40 U729 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n402), .S1(n383), .Q(n148) );
  IMUX40 U730 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n402), .S1(n386), .Q(n153) );
  IMUX40 U731 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n403), .S1(n384), .Q(n158) );
  IMUX40 U732 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n403), .S1(n379), .Q(n163) );
  IMUX40 U733 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n403), .S1(n380), .Q(n168) );
  IMUX40 U734 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n404), .S1(n380), .Q(n173) );
  IMUX40 U735 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n404), .S1(n394), .Q(n178) );
  IMUX40 U736 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n404), .S1(n387), .Q(n183) );
  IMUX40 U737 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n405), .S1(n384), .Q(n188) );
  IMUX40 U738 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n405), .S1(n384), .Q(n193) );
  IMUX40 U739 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n405), .S1(n379), .Q(n198) );
  IMUX40 U740 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n406), .S1(n379), .Q(n203) );
  IMUX40 U741 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n406), .S1(n385), .Q(n208) );
  IMUX40 U742 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n406), .S1(n385), .Q(n213) );
  IMUX40 U743 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n407), .S1(n385), .Q(n218) );
  IMUX40 U744 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n407), .S1(n386), .Q(n223) );
  IMUX40 U745 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n407), .S1(n386), .Q(n228) );
  IMUX40 U746 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n408), .S1(n380), .Q(n233) );
  IMUX40 U747 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n408), .S1(n380), .Q(n238) );
  IMUX40 U748 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n408), .S1(n381), .Q(n243) );
  IMUX40 U749 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n409), .S1(n385), .Q(n248) );
  IMUX40 U750 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n409), .S1(n380), .Q(n253) );
  IMUX40 U751 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n409), .S1(n382), .Q(n258) );
  IMUX40 U752 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n410), .S1(n382), .Q(n263) );
  IMUX40 U753 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n410), .S1(n387), .Q(n268) );
  IMUX40 U754 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n410), .S1(n387), .Q(n273) );
  IMUX40 U755 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n411), .S1(n388), .Q(n278) );
  IMUX40 U756 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n411), .S1(n388), .Q(n283) );
  IMUX40 U757 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n411), .S1(n389), .Q(n288) );
  IMUX40 U758 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n412), .S1(n389), .Q(n293) );
  IMUX40 U759 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n412), .S1(n394), .Q(n298) );
  IMUX40 U760 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n412), .S1(n393), .Q(n303) );
  IMUX40 U761 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n413), .S1(n394), .Q(n308) );
  IMUX40 U762 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n413), .S1(n390), .Q(n313) );
  IMUX40 U763 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n413), .S1(n390), .Q(n318) );
  IMUX40 U764 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n414), .S1(n391), .Q(n323) );
  IMUX40 U765 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n414), .S1(n391), .Q(n328) );
  IMUX40 U766 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n414), .S1(n392), .Q(n333) );
  IMUX40 U767 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n415), .S1(n392), .Q(n338) );
  IMUX40 U768 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n415), .S1(n393), .Q(n343) );
  IMUX40 U769 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n415), .S1(n393), .Q(n348) );
  IMUX40 U770 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n416), .S1(n393), .Q(n353) );
  IMUX40 U771 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n416), .S1(n394), .Q(n358) );
  IMUX40 U772 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n416), .S1(n394), .Q(n363) );
  IMUX40 U773 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(n785), .S1(n758), .Q(n427) );
  IMUX40 U774 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n788), .S1(n782), .Q(n462) );
  IMUX40 U775 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n788), .S1(n762), .Q(n472) );
  IMUX40 U776 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n799), .S1(n759), .Q(n482) );
  IMUX40 U777 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n789), .S1(n762), .Q(n492) );
  IMUX40 U778 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n789), .S1(n763), .Q(n502) );
  IMUX40 U779 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n790), .S1(n764), .Q(n512) );
  IMUX40 U780 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n798), .S1(n765), .Q(n522) );
  IMUX40 U781 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n799), .S1(n777), .Q(n687) );
  IMUX40 U782 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n799), .S1(n757), .Q(n692) );
  IMUX40 U783 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n799), .S1(n772), .Q(n697) );
  IMUX40 U784 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n798), .S1(n778), .Q(n702) );
  IMUX40 U785 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n798), .S1(n778), .Q(n707) );
  IMUX40 U786 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n800), .S1(n779), .Q(n712) );
  IMUX40 U787 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n800), .S1(n779), .Q(n717) );
  IMUX40 U788 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n800), .S1(n780), .Q(n727) );
  IMUX40 U789 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n801), .S1(n781), .Q(n737) );
  BUF2 U790 ( .A(i_addr_Rt[3]), .Q(n368) );
  BUF2 U791 ( .A(i_addr_Rt[3]), .Q(n369) );
  BUF2 U792 ( .A(i_addr_Rt[3]), .Q(n370) );
  BUF2 U793 ( .A(i_addr_Rt[3]), .Q(n371) );
  BUF2 U794 ( .A(i_addr_Rs[3]), .Q(n747) );
  BUF2 U795 ( .A(i_addr_Rs[3]), .Q(n748) );
  BUF2 U796 ( .A(i_addr_Rs[3]), .Q(n749) );
  BUF2 U797 ( .A(i_addr_Rs[3]), .Q(n750) );
  INV3 U798 ( .A(i_addr_Rd[0]), .Q(n906) );
  INV3 U799 ( .A(i_addr_Rd[1]), .Q(n905) );
  INV3 U800 ( .A(i_addr_Rd[2]), .Q(n904) );
  INV3 U801 ( .A(i_con_RegWr), .Q(n907) );
  BUF2 U802 ( .A(i_addr_Rs[4]), .Q(n744) );
  BUF2 U803 ( .A(i_addr_Rs[2]), .Q(n751) );
  BUF2 U804 ( .A(i_addr_Rs[2]), .Q(n752) );
  BUF2 U805 ( .A(i_addr_Rs[2]), .Q(n753) );
  BUF2 U806 ( .A(i_addr_Rs[2]), .Q(n754) );
  BUF2 U807 ( .A(i_addr_Rs[2]), .Q(n755) );
  INV3 U808 ( .A(i_addr_Rd[4]), .Q(n886) );
  INV3 U809 ( .A(i_addr_Rd[3]), .Q(n903) );
  BUF2 U810 ( .A(i_addr_Rs[3]), .Q(n746) );
  MUX22 U811 ( .A(n689), .B(n684), .S(n744), .Q(o_data_Rs[26]) );
  IMUX40 U812 ( .A(n690), .B(n691), .C(n692), .D(n693), .S0(n746), .S1(n754), 
        .Q(n689) );
  IMUX40 U813 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n799), .S1(n759), .Q(n690) );
  MUX22 U814 ( .A(n699), .B(n694), .S(n744), .Q(o_data_Rs[27]) );
  IMUX40 U815 ( .A(n700), .B(n701), .C(n702), .D(n703), .S0(n750), .S1(n755), 
        .Q(n699) );
  IMUX40 U816 ( .A(n695), .B(n696), .C(n697), .D(n698), .S0(n746), .S1(n754), 
        .Q(n694) );
  IMUX40 U817 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n800), .S1(n778), .Q(n700) );
  MUX22 U818 ( .A(n709), .B(n704), .S(n744), .Q(o_data_Rs[28]) );
  IMUX40 U819 ( .A(n710), .B(n711), .C(n712), .D(n713), .S0(n749), .S1(n755), 
        .Q(n709) );
  IMUX40 U820 ( .A(n705), .B(n706), .C(n707), .D(n708), .S0(n746), .S1(n755), 
        .Q(n704) );
  IMUX40 U821 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n800), .S1(n779), .Q(n710) );
  MUX22 U822 ( .A(n719), .B(n714), .S(n744), .Q(o_data_Rs[29]) );
  IMUX40 U823 ( .A(n720), .B(n721), .C(n722), .D(n723), .S0(n746), .S1(n755), 
        .Q(n719) );
  IMUX40 U824 ( .A(n715), .B(n716), .C(n717), .D(n718), .S0(n746), .S1(n755), 
        .Q(n714) );
  IMUX40 U825 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n800), .S1(n780), .Q(n722) );
  MUX22 U826 ( .A(n729), .B(n724), .S(i_addr_Rs[4]), .Q(o_data_Rs[30]) );
  IMUX40 U827 ( .A(n730), .B(n731), .C(n732), .D(n733), .S0(n750), .S1(n755), 
        .Q(n729) );
  IMUX40 U828 ( .A(n725), .B(n726), .C(n727), .D(n728), .S0(n746), .S1(n755), 
        .Q(n724) );
  IMUX40 U829 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n801), .S1(n780), .Q(n732) );
  MUX22 U830 ( .A(n739), .B(n734), .S(n744), .Q(o_data_Rs[31]) );
  IMUX40 U831 ( .A(n740), .B(n741), .C(n742), .D(n743), .S0(n746), .S1(n755), 
        .Q(n739) );
  IMUX40 U832 ( .A(n735), .B(n736), .C(n737), .D(n738), .S0(n746), .S1(n755), 
        .Q(n734) );
  IMUX40 U833 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n801), .S1(n781), .Q(n742) );
  BUF2 U834 ( .A(i_addr_Rt[1]), .Q(n395) );
  BUF2 U835 ( .A(n782), .Q(n756) );
  BUF2 U836 ( .A(i_addr_Rs[1]), .Q(n782) );
  MUX22 U837 ( .A(n6), .B(n1), .S(n365), .Q(o_data_Rt[0]) );
  IMUX40 U838 ( .A(n2), .B(n3), .C(n4), .D(n5), .S0(n367), .S1(i_addr_Rt[2]), 
        .Q(n1) );
  IMUX40 U839 ( .A(n7), .B(n8), .C(n9), .D(n10), .S0(n367), .S1(n372), .Q(n6)
         );
  MUX22 U840 ( .A(n16), .B(n11), .S(n365), .Q(o_data_Rt[1]) );
  IMUX40 U841 ( .A(n17), .B(n18), .C(n19), .D(n20), .S0(n367), .S1(n372), .Q(
        n16) );
  IMUX40 U842 ( .A(n12), .B(n13), .C(n14), .D(n15), .S0(n367), .S1(n372), .Q(
        n11) );
  IMUX40 U843 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n396), .S1(n379), .Q(n17) );
  MUX22 U844 ( .A(n26), .B(n21), .S(n365), .Q(o_data_Rt[2]) );
  IMUX40 U845 ( .A(n27), .B(n28), .C(n29), .D(n30), .S0(n368), .S1(n372), .Q(
        n26) );
  IMUX40 U846 ( .A(n22), .B(n23), .C(n24), .D(n25), .S0(n368), .S1(n372), .Q(
        n21) );
  IMUX40 U847 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n397), .S1(i_addr_Rt[1]), .Q(n27) );
  MUX22 U848 ( .A(n36), .B(n31), .S(n365), .Q(o_data_Rt[3]) );
  IMUX40 U849 ( .A(n37), .B(n38), .C(n83), .D(n84), .S0(n368), .S1(n372), .Q(
        n36) );
  IMUX40 U850 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(n368), .S1(n372), .Q(
        n31) );
  IMUX40 U851 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n398), .S1(n384), .Q(n37) );
  MUX22 U852 ( .A(n90), .B(n85), .S(n365), .Q(o_data_Rt[4]) );
  IMUX40 U853 ( .A(n91), .B(n92), .C(n93), .D(n94), .S0(n368), .S1(n372), .Q(
        n90) );
  IMUX40 U854 ( .A(n86), .B(n87), .C(n88), .D(n89), .S0(n368), .S1(n372), .Q(
        n85) );
  IMUX40 U855 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n398), .S1(n381), .Q(n91) );
  MUX22 U856 ( .A(n100), .B(n95), .S(n365), .Q(o_data_Rt[5]) );
  IMUX40 U857 ( .A(n101), .B(n102), .C(n103), .D(n104), .S0(n368), .S1(n373), 
        .Q(n100) );
  IMUX40 U858 ( .A(n96), .B(n97), .C(n98), .D(n99), .S0(n368), .S1(n373), .Q(
        n95) );
  IMUX40 U859 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n399), .S1(n395), .Q(n101) );
  MUX22 U860 ( .A(n110), .B(n105), .S(n366), .Q(o_data_Rt[6]) );
  IMUX40 U861 ( .A(n111), .B(n112), .C(n113), .D(n114), .S0(n368), .S1(n373), 
        .Q(n110) );
  IMUX40 U862 ( .A(n106), .B(n107), .C(n108), .D(n109), .S0(n368), .S1(n373), 
        .Q(n105) );
  IMUX40 U863 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n400), .S1(n382), .Q(n111) );
  MUX22 U864 ( .A(n120), .B(n115), .S(n366), .Q(o_data_Rt[7]) );
  IMUX40 U865 ( .A(n121), .B(n122), .C(n123), .D(n124), .S0(n368), .S1(n373), 
        .Q(n120) );
  IMUX40 U866 ( .A(n116), .B(n117), .C(n118), .D(n119), .S0(n368), .S1(n373), 
        .Q(n115) );
  IMUX40 U867 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n400), .S1(n379), .Q(n121) );
  MUX22 U868 ( .A(n130), .B(n125), .S(n366), .Q(o_data_Rt[8]) );
  IMUX40 U869 ( .A(n131), .B(n132), .C(n133), .D(n134), .S0(n369), .S1(n373), 
        .Q(n130) );
  IMUX40 U870 ( .A(n126), .B(n127), .C(n128), .D(n129), .S0(n369), .S1(n373), 
        .Q(n125) );
  IMUX40 U871 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n401), .S1(n393), .Q(n131) );
  MUX22 U872 ( .A(n140), .B(n135), .S(n366), .Q(o_data_Rt[9]) );
  IMUX40 U873 ( .A(n141), .B(n142), .C(n143), .D(n144), .S0(n369), .S1(n374), 
        .Q(n140) );
  IMUX40 U874 ( .A(n136), .B(n137), .C(n138), .D(n139), .S0(n369), .S1(n373), 
        .Q(n135) );
  IMUX40 U875 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n402), .S1(n383), .Q(n141) );
  MUX22 U876 ( .A(n150), .B(n145), .S(n366), .Q(o_data_Rt[10]) );
  IMUX40 U877 ( .A(n151), .B(n152), .C(n153), .D(n154), .S0(n369), .S1(n374), 
        .Q(n150) );
  IMUX40 U878 ( .A(n146), .B(n147), .C(n148), .D(n149), .S0(n369), .S1(n374), 
        .Q(n145) );
  IMUX40 U879 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n402), .S1(n382), .Q(n151) );
  MUX22 U880 ( .A(n160), .B(n155), .S(n366), .Q(o_data_Rt[11]) );
  IMUX40 U881 ( .A(n161), .B(n162), .C(n163), .D(n164), .S0(n369), .S1(n374), 
        .Q(n160) );
  IMUX40 U882 ( .A(n156), .B(n157), .C(n158), .D(n159), .S0(n369), .S1(n374), 
        .Q(n155) );
  IMUX40 U883 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n403), .S1(n380), .Q(n161) );
  MUX22 U884 ( .A(n170), .B(n165), .S(n366), .Q(o_data_Rt[12]) );
  IMUX40 U885 ( .A(n171), .B(n172), .C(n173), .D(n174), .S0(n369), .S1(n374), 
        .Q(n170) );
  IMUX40 U886 ( .A(n166), .B(n167), .C(n168), .D(n169), .S0(n369), .S1(n374), 
        .Q(n165) );
  IMUX40 U887 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n404), .S1(n384), .Q(n171) );
  MUX22 U888 ( .A(n180), .B(n175), .S(n366), .Q(o_data_Rt[13]) );
  IMUX40 U889 ( .A(n181), .B(n182), .C(n183), .D(n184), .S0(n369), .S1(n374), 
        .Q(n180) );
  IMUX40 U890 ( .A(n176), .B(n177), .C(n178), .D(n179), .S0(n369), .S1(n374), 
        .Q(n175) );
  IMUX40 U891 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n404), .S1(n384), .Q(n181) );
  MUX22 U892 ( .A(n190), .B(n185), .S(n366), .Q(o_data_Rt[14]) );
  IMUX40 U893 ( .A(n191), .B(n192), .C(n193), .D(n194), .S0(n370), .S1(n375), 
        .Q(n190) );
  IMUX40 U894 ( .A(n186), .B(n187), .C(n188), .D(n189), .S0(n370), .S1(n375), 
        .Q(n185) );
  IMUX40 U895 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n405), .S1(n384), .Q(n191) );
  MUX22 U896 ( .A(n200), .B(n195), .S(n366), .Q(o_data_Rt[15]) );
  IMUX40 U897 ( .A(n201), .B(n202), .C(n203), .D(n204), .S0(n370), .S1(n375), 
        .Q(n200) );
  IMUX40 U898 ( .A(n196), .B(n197), .C(n198), .D(n199), .S0(n370), .S1(n375), 
        .Q(n195) );
  IMUX40 U899 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n406), .S1(n379), .Q(n201) );
  MUX22 U900 ( .A(n210), .B(n205), .S(n366), .Q(o_data_Rt[16]) );
  IMUX40 U901 ( .A(n211), .B(n212), .C(n213), .D(n214), .S0(n370), .S1(n375), 
        .Q(n210) );
  IMUX40 U902 ( .A(n206), .B(n207), .C(n208), .D(n209), .S0(n370), .S1(n375), 
        .Q(n205) );
  IMUX40 U903 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n406), .S1(n385), .Q(n211) );
  MUX22 U904 ( .A(n220), .B(n215), .S(n366), .Q(o_data_Rt[17]) );
  IMUX40 U905 ( .A(n221), .B(n222), .C(n223), .D(n224), .S0(n370), .S1(n375), 
        .Q(n220) );
  IMUX40 U906 ( .A(n216), .B(n217), .C(n218), .D(n219), .S0(n370), .S1(n375), 
        .Q(n215) );
  IMUX40 U907 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n407), .S1(n386), .Q(n221) );
  MUX22 U908 ( .A(n230), .B(n225), .S(n366), .Q(o_data_Rt[18]) );
  IMUX40 U909 ( .A(n231), .B(n232), .C(n233), .D(n234), .S0(n370), .S1(n376), 
        .Q(n230) );
  IMUX40 U910 ( .A(n226), .B(n227), .C(n228), .D(n229), .S0(n370), .S1(n375), 
        .Q(n225) );
  IMUX40 U911 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n408), .S1(n393), .Q(n231) );
  MUX22 U912 ( .A(n240), .B(n235), .S(n365), .Q(o_data_Rt[19]) );
  IMUX40 U913 ( .A(n241), .B(n242), .C(n243), .D(n244), .S0(n370), .S1(n376), 
        .Q(n240) );
  IMUX40 U914 ( .A(n236), .B(n237), .C(n238), .D(n239), .S0(n370), .S1(n376), 
        .Q(n235) );
  IMUX40 U915 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n408), .S1(n380), .Q(n241) );
  MUX22 U916 ( .A(n250), .B(n245), .S(n365), .Q(o_data_Rt[20]) );
  IMUX40 U917 ( .A(n251), .B(n252), .C(n253), .D(n254), .S0(n371), .S1(n376), 
        .Q(n250) );
  IMUX40 U918 ( .A(n246), .B(n247), .C(n248), .D(n249), .S0(n371), .S1(n376), 
        .Q(n245) );
  IMUX40 U919 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n409), .S1(n379), .Q(n251) );
  MUX22 U920 ( .A(n260), .B(n255), .S(n365), .Q(o_data_Rt[21]) );
  IMUX40 U921 ( .A(n261), .B(n262), .C(n263), .D(n264), .S0(n371), .S1(n376), 
        .Q(n260) );
  IMUX40 U922 ( .A(n256), .B(n257), .C(n258), .D(n259), .S0(n371), .S1(n376), 
        .Q(n255) );
  IMUX40 U923 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n410), .S1(n387), .Q(n261) );
  MUX22 U924 ( .A(n270), .B(n265), .S(n365), .Q(o_data_Rt[22]) );
  IMUX40 U925 ( .A(n271), .B(n272), .C(n273), .D(n274), .S0(n371), .S1(n376), 
        .Q(n270) );
  IMUX40 U926 ( .A(n266), .B(n267), .C(n268), .D(n269), .S0(n371), .S1(n376), 
        .Q(n265) );
  IMUX40 U927 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n410), .S1(n387), .Q(n271) );
  MUX22 U928 ( .A(n280), .B(n275), .S(n365), .Q(o_data_Rt[23]) );
  IMUX40 U929 ( .A(n281), .B(n282), .C(n283), .D(n284), .S0(n371), .S1(n377), 
        .Q(n280) );
  IMUX40 U930 ( .A(n276), .B(n277), .C(n278), .D(n279), .S0(n371), .S1(n377), 
        .Q(n275) );
  IMUX40 U931 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n411), .S1(n388), .Q(n281) );
  MUX22 U932 ( .A(n290), .B(n285), .S(n365), .Q(o_data_Rt[24]) );
  IMUX40 U933 ( .A(n291), .B(n292), .C(n293), .D(n294), .S0(n371), .S1(n377), 
        .Q(n290) );
  IMUX40 U934 ( .A(n286), .B(n287), .C(n288), .D(n289), .S0(n371), .S1(n377), 
        .Q(n285) );
  IMUX40 U935 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n412), .S1(n389), .Q(n291) );
  MUX22 U936 ( .A(n300), .B(n295), .S(n365), .Q(o_data_Rt[25]) );
  IMUX40 U937 ( .A(n301), .B(n302), .C(n303), .D(n304), .S0(n371), .S1(n377), 
        .Q(n300) );
  IMUX40 U938 ( .A(n296), .B(n297), .C(n298), .D(n299), .S0(n371), .S1(n377), 
        .Q(n295) );
  IMUX40 U939 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n412), .S1(n393), .Q(n301) );
  MUX22 U940 ( .A(n310), .B(n305), .S(i_addr_Rt[4]), .Q(o_data_Rt[26]) );
  IMUX40 U941 ( .A(n311), .B(n312), .C(n313), .D(n314), .S0(n367), .S1(n377), 
        .Q(n310) );
  IMUX40 U942 ( .A(n306), .B(n307), .C(n308), .D(n309), .S0(n367), .S1(n377), 
        .Q(n305) );
  IMUX40 U943 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n413), .S1(n390), .Q(n311) );
  MUX22 U944 ( .A(n320), .B(n315), .S(i_addr_Rt[4]), .Q(o_data_Rt[27]) );
  IMUX40 U945 ( .A(n321), .B(n322), .C(n323), .D(n324), .S0(n367), .S1(n378), 
        .Q(n320) );
  IMUX40 U946 ( .A(n316), .B(n317), .C(n318), .D(n319), .S0(n367), .S1(n377), 
        .Q(n315) );
  IMUX40 U947 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n414), .S1(n391), .Q(n321) );
  MUX22 U948 ( .A(n330), .B(n325), .S(i_addr_Rt[4]), .Q(o_data_Rt[28]) );
  IMUX40 U949 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(i_addr_Rt[3]), 
        .S1(n378), .Q(n330) );
  IMUX40 U950 ( .A(n326), .B(n327), .C(n328), .D(n329), .S0(n367), .S1(n378), 
        .Q(n325) );
  IMUX40 U951 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n414), .S1(n392), .Q(n331) );
  MUX22 U952 ( .A(n340), .B(n335), .S(i_addr_Rt[4]), .Q(o_data_Rt[29]) );
  IMUX40 U953 ( .A(n341), .B(n342), .C(n343), .D(n344), .S0(i_addr_Rt[3]), 
        .S1(n378), .Q(n340) );
  IMUX40 U954 ( .A(n336), .B(n337), .C(n338), .D(n339), .S0(n367), .S1(n378), 
        .Q(n335) );
  IMUX40 U955 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n415), .S1(n393), .Q(n341) );
  MUX22 U956 ( .A(n350), .B(n345), .S(i_addr_Rt[4]), .Q(o_data_Rt[30]) );
  IMUX40 U957 ( .A(n351), .B(n352), .C(n353), .D(n354), .S0(i_addr_Rt[3]), 
        .S1(n378), .Q(n350) );
  IMUX40 U958 ( .A(n346), .B(n347), .C(n348), .D(n349), .S0(n367), .S1(n378), 
        .Q(n345) );
  IMUX40 U959 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n416), .S1(n394), .Q(n351) );
  MUX22 U960 ( .A(n360), .B(n355), .S(i_addr_Rt[4]), .Q(o_data_Rt[31]) );
  IMUX40 U961 ( .A(n361), .B(n362), .C(n363), .D(n364), .S0(i_addr_Rt[3]), 
        .S1(n378), .Q(n360) );
  IMUX40 U962 ( .A(n356), .B(n357), .C(n358), .D(n359), .S0(n367), .S1(n378), 
        .Q(n355) );
  IMUX40 U963 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n416), .S1(n394), .Q(n361) );
  BUF2 U964 ( .A(i_addr_Rt[4]), .Q(n365) );
  BUF2 U965 ( .A(i_addr_Rt[2]), .Q(n372) );
  BUF2 U966 ( .A(i_addr_Rt[2]), .Q(n373) );
  BUF2 U967 ( .A(i_addr_Rt[2]), .Q(n374) );
  BUF2 U968 ( .A(i_addr_Rt[2]), .Q(n375) );
  BUF2 U969 ( .A(i_addr_Rt[2]), .Q(n376) );
  BUF2 U970 ( .A(i_addr_Rt[2]), .Q(n377) );
  BUF2 U971 ( .A(i_addr_Rt[2]), .Q(n378) );
  BUF2 U972 ( .A(i_addr_Rt[3]), .Q(n367) );
endmodule


module D_shiftleft ( i_data_immE, o_data_immshiftl );
  input [15:0] i_data_immE;
  output [31:0] o_data_immshiftl;
  wire   n1;
  assign o_data_immshiftl[0] = o_data_immshiftl[1];
  assign o_data_immshiftl[27] = o_data_immshiftl[23];
  assign o_data_immshiftl[19] = o_data_immshiftl[23];
  assign o_data_immshiftl[24] = o_data_immshiftl[23];
  assign o_data_immshiftl[20] = o_data_immshiftl[23];
  assign o_data_immshiftl[29] = o_data_immshiftl[31];
  assign o_data_immshiftl[26] = o_data_immshiftl[31];
  assign o_data_immshiftl[25] = o_data_immshiftl[31];
  assign o_data_immshiftl[21] = o_data_immshiftl[31];
  assign o_data_immshiftl[30] = o_data_immshiftl[31];
  assign o_data_immshiftl[28] = i_data_immE[15];
  assign o_data_immshiftl[17] = i_data_immE[15];
  assign o_data_immshiftl[18] = i_data_immE[15];
  assign o_data_immshiftl[22] = i_data_immE[15];
  assign o_data_immshiftl[16] = i_data_immE[14];
  assign o_data_immshiftl[15] = i_data_immE[13];
  assign o_data_immshiftl[14] = i_data_immE[12];
  assign o_data_immshiftl[13] = i_data_immE[11];
  assign o_data_immshiftl[12] = i_data_immE[10];
  assign o_data_immshiftl[11] = i_data_immE[9];
  assign o_data_immshiftl[10] = i_data_immE[8];
  assign o_data_immshiftl[9] = i_data_immE[7];
  assign o_data_immshiftl[8] = i_data_immE[6];
  assign o_data_immshiftl[7] = i_data_immE[5];
  assign o_data_immshiftl[6] = i_data_immE[4];
  assign o_data_immshiftl[5] = i_data_immE[3];
  assign o_data_immshiftl[4] = i_data_immE[2];
  assign o_data_immshiftl[3] = i_data_immE[1];
  assign o_data_immshiftl[2] = i_data_immE[0];

  INV3 U2 ( .A(i_data_immE[15]), .Q(n1) );
  INV3 U3 ( .A(n1), .Q(o_data_immshiftl[23]) );
  INV3 U4 ( .A(n1), .Q(o_data_immshiftl[31]) );
  LOGIC0 U5 ( .Q(o_data_immshiftl[1]) );
endmodule


module D_sign_extend ( i_data_immD, i_con_signext, o_data_immD );
  input [15:0] i_data_immD;
  output [31:0] o_data_immD;
  input i_con_signext;
  wire   n2;
  assign o_data_immD[15] = i_data_immD[15];
  assign o_data_immD[14] = i_data_immD[14];
  assign o_data_immD[13] = i_data_immD[13];
  assign o_data_immD[12] = i_data_immD[12];
  assign o_data_immD[11] = i_data_immD[11];
  assign o_data_immD[10] = i_data_immD[10];
  assign o_data_immD[9] = i_data_immD[9];
  assign o_data_immD[8] = i_data_immD[8];
  assign o_data_immD[7] = i_data_immD[7];
  assign o_data_immD[6] = i_data_immD[6];
  assign o_data_immD[5] = i_data_immD[5];
  assign o_data_immD[4] = i_data_immD[4];
  assign o_data_immD[3] = i_data_immD[3];
  assign o_data_immD[2] = i_data_immD[2];
  assign o_data_immD[1] = i_data_immD[1];
  assign o_data_immD[0] = i_data_immD[0];
  assign o_data_immD[16] = o_data_immD[31];
  assign o_data_immD[17] = o_data_immD[31];
  assign o_data_immD[18] = o_data_immD[31];
  assign o_data_immD[19] = o_data_immD[31];
  assign o_data_immD[20] = o_data_immD[31];
  assign o_data_immD[21] = o_data_immD[31];
  assign o_data_immD[22] = o_data_immD[31];
  assign o_data_immD[23] = o_data_immD[31];
  assign o_data_immD[24] = o_data_immD[31];
  assign o_data_immD[25] = o_data_immD[31];
  assign o_data_immD[26] = o_data_immD[31];
  assign o_data_immD[27] = o_data_immD[31];
  assign o_data_immD[28] = o_data_immD[31];
  assign o_data_immD[29] = o_data_immD[31];
  assign o_data_immD[30] = o_data_immD[31];

  NAND20 U2 ( .A(i_con_signext), .B(i_data_immD[15]), .Q(n2) );
  INV3 U3 ( .A(n2), .Q(o_data_immD[31]) );
endmodule


module D_jump_ext ( i_addr_j, i_PC4_j, o_addr_j );
  input [25:0] i_addr_j;
  input [3:0] i_PC4_j;
  output [31:0] o_addr_j;

  assign o_addr_j[0] = o_addr_j[1];
  assign o_addr_j[31] = i_PC4_j[3];
  assign o_addr_j[30] = i_PC4_j[2];
  assign o_addr_j[29] = i_PC4_j[1];
  assign o_addr_j[28] = i_PC4_j[0];
  assign o_addr_j[27] = i_addr_j[25];
  assign o_addr_j[26] = i_addr_j[24];
  assign o_addr_j[25] = i_addr_j[23];
  assign o_addr_j[24] = i_addr_j[22];
  assign o_addr_j[23] = i_addr_j[21];
  assign o_addr_j[22] = i_addr_j[20];
  assign o_addr_j[21] = i_addr_j[19];
  assign o_addr_j[20] = i_addr_j[18];
  assign o_addr_j[19] = i_addr_j[17];
  assign o_addr_j[18] = i_addr_j[16];
  assign o_addr_j[17] = i_addr_j[15];
  assign o_addr_j[16] = i_addr_j[14];
  assign o_addr_j[15] = i_addr_j[13];
  assign o_addr_j[14] = i_addr_j[12];
  assign o_addr_j[13] = i_addr_j[11];
  assign o_addr_j[12] = i_addr_j[10];
  assign o_addr_j[11] = i_addr_j[9];
  assign o_addr_j[10] = i_addr_j[8];
  assign o_addr_j[9] = i_addr_j[7];
  assign o_addr_j[8] = i_addr_j[6];
  assign o_addr_j[7] = i_addr_j[5];
  assign o_addr_j[6] = i_addr_j[4];
  assign o_addr_j[5] = i_addr_j[3];
  assign o_addr_j[4] = i_addr_j[2];
  assign o_addr_j[3] = i_addr_j[1];
  assign o_addr_j[2] = i_addr_j[0];

  LOGIC0 U2 ( .Q(o_addr_j[1]) );
endmodule


module D_forward ( i_addr_rs, i_addr_rt, i_addr_rdE, i_addr_rdM, i_addr_rtM, 
        i_addr_rtW, i_con_regwriteE, i_con_regwriteM, i_con_memreadM, 
        i_con_memreadW, o_con_fa, o_con_fb );
  input [4:0] i_addr_rs;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rdE;
  input [4:0] i_addr_rdM;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  output [2:0] o_con_fa;
  output [2:0] o_con_fb;
  input i_con_regwriteE, i_con_regwriteM, i_con_memreadM, i_con_memreadW;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;

  NOR40 U1 ( .A(o_con_fa[2]), .B(n52), .C(n53), .D(n54), .Q(n51) );
  NAND41 U2 ( .A(n39), .B(n40), .C(n41), .D(n42), .Q(n3) );
  NOR21 U3 ( .A(n43), .B(n44), .Q(n41) );
  NOR31 U4 ( .A(i_addr_rs[2]), .B(i_addr_rs[4]), .C(i_addr_rs[3]), .Q(n85) );
  NAND22 U5 ( .A(n63), .B(n48), .Q(o_con_fa[2]) );
  NAND42 U6 ( .A(n55), .B(i_con_regwriteE), .C(n56), .D(n57), .Q(n46) );
  OAI211 U7 ( .A(n47), .B(n48), .C(n49), .Q(o_con_fa[0]) );
  NAND21 U8 ( .A(n4), .B(n10), .Q(o_con_fb[0]) );
  OAI310 U9 ( .A(n1), .B(n2), .C(n3), .D(n4), .Q(o_con_fb[2]) );
  NOR40 U10 ( .A(n5), .B(n6), .C(n7), .D(n8), .Q(o_con_fb[1]) );
  CLKIN0 U11 ( .A(n9), .Q(n6) );
  NAND40 U12 ( .A(n11), .B(i_con_regwriteM), .C(n12), .D(n13), .Q(n10) );
  NOR40 U13 ( .A(n14), .B(n15), .C(n16), .D(n17), .Q(n13) );
  XOR20 U14 ( .A(i_addr_rdM[4]), .B(i_addr_rt[4]), .Q(n17) );
  XNR20 U15 ( .A(n18), .B(i_addr_rt[2]), .Q(n16) );
  XNR20 U16 ( .A(n19), .B(i_addr_rt[1]), .Q(n15) );
  XNR20 U17 ( .A(n20), .B(i_addr_rt[0]), .Q(n14) );
  CLKIN0 U18 ( .A(n21), .Q(n12) );
  OAI210 U19 ( .A(n8), .B(n7), .C(n9), .Q(n21) );
  NAND40 U20 ( .A(n22), .B(n23), .C(n24), .D(n25), .Q(n7) );
  XNR20 U21 ( .A(i_addr_rt[0]), .B(i_addr_rdE[0]), .Q(n25) );
  NOR20 U22 ( .A(n26), .B(n27), .Q(n24) );
  XNR20 U23 ( .A(n28), .B(i_addr_rt[3]), .Q(n27) );
  XOR20 U24 ( .A(i_addr_rdE[1]), .B(i_addr_rt[1]), .Q(n26) );
  XNR20 U25 ( .A(i_addr_rt[2]), .B(i_addr_rdE[2]), .Q(n23) );
  XNR20 U26 ( .A(i_addr_rt[4]), .B(i_addr_rdE[4]), .Q(n22) );
  CLKIN0 U27 ( .A(i_con_regwriteE), .Q(n8) );
  XNR20 U28 ( .A(i_addr_rt[3]), .B(i_addr_rdM[3]), .Q(n11) );
  NAND20 U29 ( .A(n9), .B(n5), .Q(n4) );
  CLKIN0 U30 ( .A(n29), .Q(n5) );
  NAND40 U31 ( .A(n30), .B(i_con_memreadW), .C(n31), .D(n32), .Q(n29) );
  NOR30 U32 ( .A(n33), .B(n34), .C(n35), .Q(n32) );
  XOR20 U33 ( .A(i_addr_rtW[2]), .B(i_addr_rt[2]), .Q(n35) );
  XOR20 U34 ( .A(i_addr_rtW[4]), .B(i_addr_rt[4]), .Q(n34) );
  XOR20 U35 ( .A(i_addr_rtW[3]), .B(i_addr_rt[3]), .Q(n33) );
  XNR20 U36 ( .A(i_addr_rt[0]), .B(i_addr_rtW[0]), .Q(n31) );
  XNR20 U37 ( .A(i_addr_rt[1]), .B(i_addr_rtW[1]), .Q(n30) );
  AOI210 U38 ( .A(n36), .B(i_con_memreadM), .C(n2), .Q(n9) );
  NOR30 U39 ( .A(i_addr_rt[0]), .B(i_addr_rt[1]), .C(n37), .Q(n2) );
  CLKIN0 U40 ( .A(n38), .Q(n37) );
  NOR30 U41 ( .A(i_addr_rt[2]), .B(i_addr_rt[4]), .C(i_addr_rt[3]), .Q(n38) );
  CLKIN0 U42 ( .A(n3), .Q(n36) );
  XNR20 U43 ( .A(i_addr_rt[0]), .B(i_addr_rtM[0]), .Q(n42) );
  XOR20 U44 ( .A(i_addr_rtM[3]), .B(i_addr_rt[3]), .Q(n44) );
  XNR20 U45 ( .A(n45), .B(i_addr_rt[1]), .Q(n43) );
  XNR20 U46 ( .A(i_addr_rt[2]), .B(i_addr_rtM[2]), .Q(n40) );
  XNR20 U47 ( .A(i_addr_rt[4]), .B(i_addr_rtM[4]), .Q(n39) );
  NOR20 U48 ( .A(o_con_fa[2]), .B(n46), .Q(o_con_fa[1]) );
  NAND20 U49 ( .A(n50), .B(n51), .Q(n49) );
  XNR20 U50 ( .A(n20), .B(i_addr_rs[0]), .Q(n54) );
  CLKIN0 U51 ( .A(i_addr_rdM[0]), .Q(n20) );
  CLKIN0 U52 ( .A(i_con_regwriteM), .Q(n53) );
  CLKIN0 U53 ( .A(n46), .Q(n52) );
  NOR30 U54 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  XNR20 U55 ( .A(n28), .B(i_addr_rs[3]), .Q(n60) );
  CLKIN0 U56 ( .A(i_addr_rdE[3]), .Q(n28) );
  XOR20 U57 ( .A(i_addr_rdE[2]), .B(i_addr_rs[2]), .Q(n59) );
  IMUX20 U58 ( .A(n61), .B(i_addr_rs[4]), .S(i_addr_rdE[4]), .Q(n58) );
  NOR20 U59 ( .A(n62), .B(i_addr_rs[4]), .Q(n61) );
  NOR40 U60 ( .A(i_addr_rdE[3]), .B(i_addr_rdE[2]), .C(i_addr_rdE[1]), .D(
        i_addr_rdE[0]), .Q(n62) );
  XNR20 U61 ( .A(i_addr_rs[0]), .B(i_addr_rdE[0]), .Q(n56) );
  XNR20 U62 ( .A(i_addr_rs[1]), .B(i_addr_rdE[1]), .Q(n55) );
  NOR40 U63 ( .A(n64), .B(n65), .C(n66), .D(n67), .Q(n50) );
  IMUX20 U64 ( .A(n68), .B(i_addr_rs[4]), .S(i_addr_rdM[4]), .Q(n67) );
  NOR20 U65 ( .A(n69), .B(i_addr_rs[4]), .Q(n68) );
  NOR40 U66 ( .A(i_addr_rdM[3]), .B(i_addr_rdM[2]), .C(i_addr_rdM[1]), .D(
        i_addr_rdM[0]), .Q(n69) );
  XOR20 U67 ( .A(i_addr_rdM[3]), .B(i_addr_rs[3]), .Q(n66) );
  XNR20 U68 ( .A(n18), .B(i_addr_rs[2]), .Q(n65) );
  CLKIN0 U69 ( .A(i_addr_rdM[2]), .Q(n18) );
  XNR20 U70 ( .A(n19), .B(i_addr_rs[1]), .Q(n64) );
  CLKIN0 U71 ( .A(i_addr_rdM[1]), .Q(n19) );
  NAND40 U72 ( .A(n70), .B(n71), .C(n72), .D(n73), .Q(n48) );
  NOR40 U73 ( .A(n74), .B(n75), .C(n76), .D(n77), .Q(n73) );
  XOR20 U74 ( .A(i_addr_rtW[1]), .B(i_addr_rs[1]), .Q(n77) );
  XOR20 U75 ( .A(i_addr_rtW[0]), .B(i_addr_rs[0]), .Q(n76) );
  CLKIN0 U76 ( .A(i_con_memreadW), .Q(n75) );
  XNR20 U77 ( .A(i_addr_rtW[3]), .B(i_addr_rs[3]), .Q(n72) );
  XNR20 U78 ( .A(i_addr_rtW[4]), .B(i_addr_rs[4]), .Q(n71) );
  XNR20 U79 ( .A(i_addr_rtW[2]), .B(i_addr_rs[2]), .Q(n70) );
  CLKIN0 U80 ( .A(n63), .Q(n47) );
  NAND40 U81 ( .A(n78), .B(n79), .C(n80), .D(n81), .Q(n63) );
  NOR40 U82 ( .A(n74), .B(n1), .C(n82), .D(n83), .Q(n81) );
  XNR20 U83 ( .A(n45), .B(i_addr_rs[1]), .Q(n83) );
  CLKIN0 U84 ( .A(i_addr_rtM[1]), .Q(n45) );
  XOR20 U85 ( .A(i_addr_rtM[0]), .B(i_addr_rs[0]), .Q(n82) );
  CLKIN0 U86 ( .A(i_con_memreadM), .Q(n1) );
  NOR30 U87 ( .A(i_addr_rs[0]), .B(i_addr_rs[1]), .C(n84), .Q(n74) );
  CLKIN0 U88 ( .A(n85), .Q(n84) );
  XNR20 U89 ( .A(i_addr_rtM[3]), .B(i_addr_rs[3]), .Q(n80) );
  XNR20 U90 ( .A(i_addr_rtM[4]), .B(i_addr_rs[4]), .Q(n79) );
  XNR20 U91 ( .A(i_addr_rtM[2]), .B(i_addr_rs[2]), .Q(n78) );
endmodule


module decode ( i_clk, i_nrst, i_addr_pc4, i_data_instr, i_con_Wregwrite, 
        i_data_Wregwrite, i_addr_Wregwrite, i_addr_Erd, i_addr_Mrd, 
        i_con_Eregwrite, i_con_Mregwrite, i_addr_rtM, i_addr_rtW, 
        i_con_memreadM, i_con_memreadW, i_data_Wmemout, o_data_rs, o_data_rt, 
        o_addr_rd, o_addr_rt, o_data_jr, o_con_jump, o_addr_pc4, o_addr_branch, 
        o_addr_jump, o_con_Ealuop, o_con_Ealusrc, o_con_Eregdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_con_ifstall, o_con_Ebop, o_data_signext, 
        o_con_Efamux, o_con_Efbmux, o_data_Fmemout );
  input [31:0] i_addr_pc4;
  input [31:0] i_data_instr;
  input [31:0] i_data_Wregwrite;
  input [4:0] i_addr_Wregwrite;
  input [4:0] i_addr_Erd;
  input [4:0] i_addr_Mrd;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  input [31:0] i_data_Wmemout;
  output [31:0] o_data_rs;
  output [31:0] o_data_rt;
  output [4:0] o_addr_rd;
  output [4:0] o_addr_rt;
  output [31:0] o_data_jr;
  output [1:0] o_con_jump;
  output [31:0] o_addr_pc4;
  output [31:0] o_addr_branch;
  output [31:0] o_addr_jump;
  output [5:0] o_con_Ealuop;
  output [2:0] o_con_Ebop;
  output [31:0] o_data_signext;
  output [2:0] o_con_Efamux;
  output [2:0] o_con_Efbmux;
  output [31:0] o_data_Fmemout;
  input i_clk, i_nrst, i_con_Wregwrite, i_con_Eregwrite, i_con_Mregwrite,
         i_con_memreadM, i_con_memreadW;
  output o_con_Ealusrc, o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite,
         o_con_Malupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall;
  wire   n5, control_o_con_alusrc, control_o_con_regdst, jbcon_o_con_aluPC4,
         control_o_con_memread, control_o_con_memwrite, control_o_con_memtoreg,
         control_o_con_regwrite, signext_i_con_signext, n2, n4,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4;
  wire   [31:0] regbank_o_data_Rt;
  wire   [5:0] control_o_con_aluop;
  wire   [31:0] signext_o_data_immD;
  wire   [2:0] for_o_con_fa;
  wire   [2:0] for_o_con_fb;
  wire   [31:0] pcadd_o_addr_pcbranchE;
  wire   [2:0] jbcon_o_con_bop;
  wire   [31:2] pcadd_i_data_immshiftl;
  assign o_addr_jump[1] = o_addr_jump[0];

  DFC3 pipe_bop_reg_2_ ( .D(jbcon_o_con_bop[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[2]) );
  DFC3 pipe_bop_reg_1_ ( .D(jbcon_o_con_bop[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[1]) );
  DFC3 pipe_bop_reg_0_ ( .D(jbcon_o_con_bop[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[0]) );
  DFC3 pipe_data_rs_reg_13_ ( .D(o_data_jr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[13]) );
  DFC3 pipe_data_rt_reg_31_ ( .D(regbank_o_data_Rt[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[31]) );
  DFC3 pipe_data_rt_reg_29_ ( .D(regbank_o_data_Rt[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[29]) );
  DFC3 pipe_data_rt_reg_28_ ( .D(regbank_o_data_Rt[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28]) );
  DFC3 pipe_data_rt_reg_27_ ( .D(regbank_o_data_Rt[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27]) );
  DFC3 pipe_data_rt_reg_26_ ( .D(regbank_o_data_Rt[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26]) );
  DFC3 pipe_data_rt_reg_25_ ( .D(regbank_o_data_Rt[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25]) );
  DFC3 pipe_data_rt_reg_24_ ( .D(regbank_o_data_Rt[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24]) );
  DFC3 pipe_data_rt_reg_23_ ( .D(regbank_o_data_Rt[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23]) );
  DFC3 pipe_data_rt_reg_22_ ( .D(regbank_o_data_Rt[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC3 pipe_data_rt_reg_21_ ( .D(regbank_o_data_Rt[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21]) );
  DFC3 pipe_data_rt_reg_20_ ( .D(regbank_o_data_Rt[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20]) );
  DFC3 pipe_data_rt_reg_19_ ( .D(regbank_o_data_Rt[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19]) );
  DFC3 pipe_data_rt_reg_18_ ( .D(regbank_o_data_Rt[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18]) );
  DFC3 pipe_data_rt_reg_17_ ( .D(regbank_o_data_Rt[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17]) );
  DFC3 pipe_data_rt_reg_16_ ( .D(regbank_o_data_Rt[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC3 pipe_data_rt_reg_15_ ( .D(regbank_o_data_Rt[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15]) );
  DFC3 pipe_data_rt_reg_14_ ( .D(regbank_o_data_Rt[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14]) );
  DFC3 pipe_data_rt_reg_13_ ( .D(regbank_o_data_Rt[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC3 pipe_data_rt_reg_12_ ( .D(regbank_o_data_Rt[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12]) );
  DFC3 pipe_data_rt_reg_11_ ( .D(regbank_o_data_Rt[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11]) );
  DFC3 pipe_data_rt_reg_10_ ( .D(regbank_o_data_Rt[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC3 pipe_data_rt_reg_9_ ( .D(regbank_o_data_Rt[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[9]) );
  DFC3 pipe_data_rt_reg_8_ ( .D(regbank_o_data_Rt[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[8]) );
  DFC3 pipe_data_rt_reg_7_ ( .D(regbank_o_data_Rt[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[7]) );
  DFC3 pipe_data_rt_reg_6_ ( .D(regbank_o_data_Rt[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[6]) );
  DFC3 pipe_data_rt_reg_5_ ( .D(regbank_o_data_Rt[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[5]) );
  DFC3 pipe_data_rt_reg_4_ ( .D(regbank_o_data_Rt[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[4]) );
  DFC3 pipe_data_rt_reg_3_ ( .D(regbank_o_data_Rt[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[3]) );
  DFC3 pipe_data_rt_reg_2_ ( .D(regbank_o_data_Rt[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[2]) );
  DFC3 pipe_data_rt_reg_1_ ( .D(regbank_o_data_Rt[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[1]) );
  DFC3 pipe_data_rt_reg_0_ ( .D(regbank_o_data_Rt[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[0]) );
  DFC3 pipe_addr_rd_reg_3_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[3]) );
  DFC3 pipe_addr_rd_reg_2_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[2]) );
  DFC3 pipe_addr_rd_reg_1_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[1]) );
  DFC3 pipe_addr_rd_reg_0_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[0]) );
  DFC3 pipe_addr_rt_reg_4_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[0]) );
  DFC3 pipe_addr_pc4_reg_31_ ( .D(i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_addr_pc4_reg_30_ ( .D(i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_addr_pc4_reg_29_ ( .D(i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_addr_pc4_reg_28_ ( .D(i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_addr_pc4_reg_27_ ( .D(i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_addr_pc4_reg_26_ ( .D(i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_addr_pc4_reg_25_ ( .D(i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_addr_pc4_reg_24_ ( .D(i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_addr_pc4_reg_23_ ( .D(i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_addr_pc4_reg_22_ ( .D(i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_addr_pc4_reg_21_ ( .D(i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_addr_pc4_reg_20_ ( .D(i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_addr_pc4_reg_19_ ( .D(i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_addr_pc4_reg_18_ ( .D(i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_addr_pc4_reg_17_ ( .D(i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_addr_pc4_reg_16_ ( .D(i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_addr_pc4_reg_15_ ( .D(i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_addr_pc4_reg_14_ ( .D(i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_addr_pc4_reg_13_ ( .D(i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_addr_pc4_reg_12_ ( .D(i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_addr_pc4_reg_11_ ( .D(i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_addr_pc4_reg_10_ ( .D(i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_addr_pc4_reg_9_ ( .D(i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_addr_pc4_reg_8_ ( .D(i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_addr_pc4_reg_7_ ( .D(i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_addr_pc4_reg_6_ ( .D(i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_addr_pc4_reg_5_ ( .D(i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_addr_pc4_reg_4_ ( .D(i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_addr_pc4_reg_3_ ( .D(i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_addr_pc4_reg_1_ ( .D(i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_addr_pc4_reg_0_ ( .D(i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  DFC3 pipe_con_Ealuop_reg_5_ ( .D(control_o_con_aluop[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[5]) );
  DFC3 pipe_con_Ealuop_reg_4_ ( .D(control_o_con_aluop[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[4]) );
  DFC3 pipe_con_Ealuop_reg_3_ ( .D(control_o_con_aluop[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[3]) );
  DFC3 pipe_con_Ealuop_reg_2_ ( .D(control_o_con_aluop[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[2]) );
  DFC3 pipe_con_Ealuop_reg_1_ ( .D(control_o_con_aluop[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[1]) );
  DFC3 pipe_con_Ealuop_reg_0_ ( .D(control_o_con_aluop[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[0]) );
  DFC3 pipe_con_Ealusrc_reg ( .D(control_o_con_alusrc), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Ealusrc) );
  DFC3 pipe_con_Eregdst_reg ( .D(control_o_con_regdst), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Eregdst) );
  DFC3 pipe_con_MaluPC4_reg ( .D(jbcon_o_con_aluPC4), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Malupc8) );
  DFC3 pipe_con_Mmemread_reg ( .D(control_o_con_memread), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(control_o_con_memwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(control_o_con_memtoreg), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(control_o_con_regwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wregwrite) );
  DFC3 pipe_signext_o_data_immD_reg_27_ ( .D(signext_o_data_immD[27]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[27]) );
  DFC3 pipe_signext_o_data_immD_reg_26_ ( .D(signext_o_data_immD[26]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[26]) );
  DFC3 pipe_signext_o_data_immD_reg_25_ ( .D(signext_o_data_immD[25]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[25]) );
  DFC3 pipe_signext_o_data_immD_reg_24_ ( .D(signext_o_data_immD[24]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[24]) );
  DFC3 pipe_signext_o_data_immD_reg_23_ ( .D(signext_o_data_immD[23]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[23]) );
  DFC3 pipe_signext_o_data_immD_reg_22_ ( .D(signext_o_data_immD[22]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[22]) );
  DFC3 pipe_signext_o_data_immD_reg_21_ ( .D(signext_o_data_immD[21]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[21]) );
  DFC3 pipe_signext_o_data_immD_reg_20_ ( .D(signext_o_data_immD[20]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[20]) );
  DFC3 pipe_signext_o_data_immD_reg_19_ ( .D(signext_o_data_immD[19]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[19]) );
  DFC3 pipe_signext_o_data_immD_reg_18_ ( .D(signext_o_data_immD[18]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[18]) );
  DFC3 pipe_signext_o_data_immD_reg_17_ ( .D(signext_o_data_immD[17]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[17]) );
  DFC3 pipe_signext_o_data_immD_reg_16_ ( .D(signext_o_data_immD[16]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[16]) );
  DFC3 pipe_signext_o_data_immD_reg_14_ ( .D(signext_o_data_immD[14]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[14]) );
  DFC3 pipe_signext_o_data_immD_reg_13_ ( .D(signext_o_data_immD[13]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[13]) );
  DFC3 pipe_signext_o_data_immD_reg_12_ ( .D(signext_o_data_immD[12]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[12]) );
  DFC3 pipe_signext_o_data_immD_reg_11_ ( .D(signext_o_data_immD[11]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[11]) );
  DFC3 pipe_signext_o_data_immD_reg_10_ ( .D(signext_o_data_immD[10]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[10]) );
  DFC3 pipe_signext_o_data_immD_reg_9_ ( .D(signext_o_data_immD[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[9]) );
  DFC3 pipe_signext_o_data_immD_reg_8_ ( .D(signext_o_data_immD[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[8]) );
  DFC3 pipe_signext_o_data_immD_reg_7_ ( .D(signext_o_data_immD[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[7]) );
  DFC3 pipe_signext_o_data_immD_reg_6_ ( .D(signext_o_data_immD[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[6]) );
  DFC3 pipe_signext_o_data_immD_reg_5_ ( .D(signext_o_data_immD[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[5]) );
  DFC3 pipe_signext_o_data_immD_reg_4_ ( .D(signext_o_data_immD[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[4]) );
  DFC3 pipe_signext_o_data_immD_reg_3_ ( .D(signext_o_data_immD[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[3]) );
  DFC3 pipe_signext_o_data_immD_reg_2_ ( .D(signext_o_data_immD[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[2]) );
  DFC3 pipe_signext_o_data_immD_reg_1_ ( .D(signext_o_data_immD[1]), .C(i_clk), 
        .RN(i_nrst), .Q(n5) );
  DFC3 pipe_signext_o_data_immD_reg_0_ ( .D(signext_o_data_immD[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[0]) );
  DFC3 pipe_con_Efamux_reg_2_ ( .D(for_o_con_fa[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[2]) );
  DFC3 pipe_con_Efamux_reg_1_ ( .D(for_o_con_fa[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[1]) );
  DFC3 pipe_con_Efamux_reg_0_ ( .D(for_o_con_fa[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[0]) );
  DFC3 pipe_con_Efbmux_reg_2_ ( .D(for_o_con_fb[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[2]) );
  DFC3 pipe_con_Efbmux_reg_1_ ( .D(for_o_con_fb[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[1]) );
  DFC3 pipe_con_Efbmux_reg_0_ ( .D(for_o_con_fb[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[0]) );
  DFC3 pipe_FWmemout_reg_21_ ( .D(i_data_Wmemout[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[21]) );
  DFC3 pipe_FWmemout_reg_15_ ( .D(i_data_Wmemout[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[15]) );
  DFC3 pipe_FWmemout_reg_10_ ( .D(i_data_Wmemout[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[10]) );
  DFC3 pipe_FWmemout_reg_9_ ( .D(i_data_Wmemout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[9]) );
  DFC3 pipe_FWmemout_reg_6_ ( .D(i_data_Wmemout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[6]) );
  DFC3 pipe_addr_branch_reg_31_ ( .D(pcadd_o_addr_pcbranchE[31]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[31]) );
  DFC3 pipe_addr_branch_reg_30_ ( .D(pcadd_o_addr_pcbranchE[30]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[30]) );
  DFC3 pipe_addr_branch_reg_29_ ( .D(pcadd_o_addr_pcbranchE[29]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[29]) );
  DFC3 pipe_addr_branch_reg_24_ ( .D(pcadd_o_addr_pcbranchE[24]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[24]) );
  DFC3 pipe_addr_branch_reg_23_ ( .D(pcadd_o_addr_pcbranchE[23]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[23]) );
  DFC3 pipe_addr_branch_reg_22_ ( .D(pcadd_o_addr_pcbranchE[22]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[22]) );
  DFC3 pipe_addr_branch_reg_21_ ( .D(pcadd_o_addr_pcbranchE[21]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[21]) );
  DFC3 pipe_addr_branch_reg_20_ ( .D(pcadd_o_addr_pcbranchE[20]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[20]) );
  DFC3 pipe_addr_branch_reg_18_ ( .D(pcadd_o_addr_pcbranchE[18]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[18]) );
  DFC3 pipe_addr_branch_reg_17_ ( .D(pcadd_o_addr_pcbranchE[17]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[17]) );
  DFC3 pipe_addr_branch_reg_16_ ( .D(pcadd_o_addr_pcbranchE[16]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[16]) );
  DFC3 pipe_addr_branch_reg_13_ ( .D(pcadd_o_addr_pcbranchE[13]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[13]) );
  DFC3 pipe_addr_branch_reg_12_ ( .D(pcadd_o_addr_pcbranchE[12]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[12]) );
  DFC3 pipe_addr_branch_reg_10_ ( .D(pcadd_o_addr_pcbranchE[10]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[10]) );
  DFC3 pipe_addr_branch_reg_9_ ( .D(pcadd_o_addr_pcbranchE[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[9]) );
  DFC3 pipe_addr_branch_reg_8_ ( .D(pcadd_o_addr_pcbranchE[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[8]) );
  DFC3 pipe_addr_branch_reg_7_ ( .D(pcadd_o_addr_pcbranchE[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[7]) );
  DFC3 pipe_addr_branch_reg_6_ ( .D(pcadd_o_addr_pcbranchE[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[6]) );
  DFC3 pipe_addr_branch_reg_5_ ( .D(pcadd_o_addr_pcbranchE[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[5]) );
  DFC3 pipe_addr_branch_reg_4_ ( .D(pcadd_o_addr_pcbranchE[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[4]) );
  DFC3 pipe_addr_branch_reg_3_ ( .D(pcadd_o_addr_pcbranchE[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[3]) );
  DFC3 pipe_addr_branch_reg_2_ ( .D(pcadd_o_addr_pcbranchE[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[2]) );
  DFC3 pipe_addr_branch_reg_1_ ( .D(pcadd_o_addr_pcbranchE[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[1]) );
  DFC3 pipe_addr_branch_reg_0_ ( .D(pcadd_o_addr_pcbranchE[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[0]) );
  D_control u_control ( .o_con_regdst(control_o_con_regdst), .o_con_memread(
        control_o_con_memread), .o_con_memtoreg(control_o_con_memtoreg), 
        .o_con_memwrite(control_o_con_memwrite), .o_con_alusrc(
        control_o_con_alusrc), .o_con_regwrite(control_o_con_regwrite), 
        .o_con_ifsign(signext_i_con_signext), .o_con_aluop(control_o_con_aluop), .i_con_instru(i_data_instr[31:26]) );
  D_jb_control u_jb_control ( .o_con_jump(o_con_jump), .o_con_bop(
        jbcon_o_con_bop), .o_con_aluPC4(jbcon_o_con_aluPC4), .o_con_ifstall(
        o_con_ifstall), .i_con_instru(i_data_instr[31:26]), .i_con_func(
        i_data_instr[5:0]), .i_con_rt(i_data_instr[16]) );
  D_pcadd u_pcadd ( .i_addr_pcadd4E(i_addr_pc4), .i_data_immshiftl({
        pcadd_i_data_immshiftl, o_addr_jump[0], o_addr_jump[0]}), 
        .o_addr_pcbranchE(pcadd_o_addr_pcbranchE) );
  D_register_bank u_regbank ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_addr_Rs({
        i_data_instr[25:22], n4}), .i_addr_Rt(i_data_instr[20:16]), 
        .i_con_RegWr(i_con_Wregwrite), .i_addr_Rd(i_addr_Wregwrite), 
        .i_data_Rd(i_data_Wregwrite), .o_data_Rs(o_data_jr), .o_data_Rt(
        regbank_o_data_Rt) );
  D_shiftleft u_sl ( .i_data_immE(i_data_instr[15:0]), .o_data_immshiftl({
        pcadd_i_data_immshiftl, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}) );
  D_sign_extend u_signext ( .i_data_immD(i_data_instr[15:0]), .i_con_signext(
        signext_i_con_signext), .o_data_immD(signext_o_data_immD) );
  D_jump_ext u_jump_ext ( .i_addr_j({i_data_instr[25:22], n4, 
        i_data_instr[20:0]}), .i_PC4_j(i_addr_pc4[31:28]), .o_addr_j({
        o_addr_jump[31:2], SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4}) );
  D_forward u_forward ( .i_addr_rs({i_data_instr[25:22], n4}), .i_addr_rt(
        i_data_instr[20:16]), .i_addr_rdE(i_addr_Erd), .i_addr_rdM(i_addr_Mrd), 
        .i_addr_rtM(i_addr_rtM), .i_addr_rtW(i_addr_rtW), .i_con_regwriteE(
        i_con_Eregwrite), .i_con_regwriteM(i_con_Mregwrite), .i_con_memreadM(
        i_con_memreadM), .i_con_memreadW(i_con_memreadW), .o_con_fa(
        for_o_con_fa), .o_con_fb(for_o_con_fb) );
  DFC1 pipe_data_rs_reg_31_ ( .D(o_data_jr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[31]) );
  DFC1 pipe_data_rt_reg_30_ ( .D(regbank_o_data_Rt[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC1 pipe_data_rs_reg_7_ ( .D(o_data_jr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[7]) );
  DFC1 pipe_data_rs_reg_20_ ( .D(o_data_jr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[20]) );
  DFC1 pipe_data_rs_reg_28_ ( .D(o_data_jr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[28]) );
  DFC1 pipe_data_rs_reg_3_ ( .D(o_data_jr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[3]) );
  DFC1 pipe_data_rs_reg_1_ ( .D(o_data_jr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[1]) );
  DFC1 pipe_data_rs_reg_2_ ( .D(o_data_jr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[2]) );
  DFC1 pipe_data_rs_reg_11_ ( .D(o_data_jr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[11]) );
  DFC1 pipe_data_rs_reg_30_ ( .D(o_data_jr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[30]) );
  DFC1 pipe_data_rs_reg_29_ ( .D(o_data_jr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[29]) );
  DFC1 pipe_data_rs_reg_5_ ( .D(o_data_jr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[5]) );
  DFC1 pipe_data_rs_reg_8_ ( .D(o_data_jr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[8]) );
  DFC1 pipe_data_rs_reg_26_ ( .D(o_data_jr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[26]) );
  DFC1 pipe_data_rs_reg_12_ ( .D(o_data_jr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[12]) );
  DFC1 pipe_data_rs_reg_24_ ( .D(o_data_jr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[24]) );
  DFC1 pipe_data_rs_reg_14_ ( .D(o_data_jr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[14]) );
  DFC1 pipe_data_rs_reg_4_ ( .D(o_data_jr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[4]) );
  DFC1 pipe_data_rs_reg_19_ ( .D(o_data_jr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[19]) );
  DFC1 pipe_data_rs_reg_9_ ( .D(o_data_jr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[9]) );
  DFC1 pipe_data_rs_reg_16_ ( .D(o_data_jr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[16]) );
  DFC1 pipe_data_rs_reg_10_ ( .D(o_data_jr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[10]) );
  DFC1 pipe_data_rs_reg_21_ ( .D(o_data_jr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[21]) );
  DFC1 pipe_data_rs_reg_25_ ( .D(o_data_jr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[25]) );
  DFC1 pipe_data_rs_reg_18_ ( .D(o_data_jr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[18]) );
  DFC1 pipe_data_rs_reg_6_ ( .D(o_data_jr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[6]) );
  DFC1 pipe_data_rs_reg_22_ ( .D(o_data_jr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[22]) );
  DFC1 pipe_data_rs_reg_27_ ( .D(o_data_jr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[27]) );
  DFC1 pipe_data_rs_reg_23_ ( .D(o_data_jr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[23]) );
  DFC1 pipe_data_rs_reg_15_ ( .D(o_data_jr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[15]) );
  DFC1 pipe_data_rs_reg_17_ ( .D(o_data_jr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[17]) );
  DFC1 pipe_FWmemout_reg_7_ ( .D(i_data_Wmemout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[7]) );
  DFC1 pipe_FWmemout_reg_29_ ( .D(i_data_Wmemout[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[29]) );
  DFC1 pipe_FWmemout_reg_28_ ( .D(i_data_Wmemout[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[28]) );
  DFC1 pipe_FWmemout_reg_0_ ( .D(i_data_Wmemout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[0]) );
  DFC1 pipe_FWmemout_reg_3_ ( .D(i_data_Wmemout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[3]) );
  DFC1 pipe_FWmemout_reg_30_ ( .D(i_data_Wmemout[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[30]) );
  DFC1 pipe_FWmemout_reg_5_ ( .D(i_data_Wmemout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[5]) );
  DFC1 pipe_FWmemout_reg_8_ ( .D(i_data_Wmemout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[8]) );
  DFC1 pipe_FWmemout_reg_25_ ( .D(i_data_Wmemout[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[25]) );
  DFC1 pipe_FWmemout_reg_22_ ( .D(i_data_Wmemout[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[22]) );
  DFC1 pipe_FWmemout_reg_4_ ( .D(i_data_Wmemout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[4]) );
  DFC1 pipe_FWmemout_reg_14_ ( .D(i_data_Wmemout[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[14]) );
  DFC1 pipe_FWmemout_reg_2_ ( .D(i_data_Wmemout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[2]) );
  DFC1 pipe_FWmemout_reg_24_ ( .D(i_data_Wmemout[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[24]) );
  DFC1 pipe_FWmemout_reg_26_ ( .D(i_data_Wmemout[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[26]) );
  DFC1 pipe_FWmemout_reg_11_ ( .D(i_data_Wmemout[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[11]) );
  DFC1 pipe_FWmemout_reg_16_ ( .D(i_data_Wmemout[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[16]) );
  DFC1 pipe_FWmemout_reg_12_ ( .D(i_data_Wmemout[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[12]) );
  DFC1 pipe_FWmemout_reg_20_ ( .D(i_data_Wmemout[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[20]) );
  DFC1 pipe_FWmemout_reg_19_ ( .D(i_data_Wmemout[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[19]) );
  DFC1 pipe_FWmemout_reg_1_ ( .D(i_data_Wmemout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[1]) );
  DFC1 pipe_FWmemout_reg_17_ ( .D(i_data_Wmemout[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[17]) );
  DFC1 pipe_FWmemout_reg_18_ ( .D(i_data_Wmemout[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[18]) );
  DFC1 pipe_addr_branch_reg_28_ ( .D(pcadd_o_addr_pcbranchE[28]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[28]) );
  DFC1 pipe_addr_branch_reg_27_ ( .D(pcadd_o_addr_pcbranchE[27]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[27]) );
  DFC1 pipe_addr_branch_reg_26_ ( .D(pcadd_o_addr_pcbranchE[26]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[26]) );
  DFC1 pipe_addr_branch_reg_25_ ( .D(pcadd_o_addr_pcbranchE[25]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[25]) );
  DFC1 pipe_signext_o_data_immD_reg_29_ ( .D(signext_o_data_immD[29]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[29]) );
  DFC1 pipe_signext_o_data_immD_reg_30_ ( .D(signext_o_data_immD[30]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[30]) );
  DFC1 pipe_signext_o_data_immD_reg_31_ ( .D(signext_o_data_immD[31]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[31]) );
  DFC1 pipe_data_rs_reg_0_ ( .D(o_data_jr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[0]) );
  DFC1 pipe_signext_o_data_immD_reg_28_ ( .D(signext_o_data_immD[28]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[28]) );
  DFC1 pipe_addr_branch_reg_19_ ( .D(pcadd_o_addr_pcbranchE[19]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[19]) );
  DFC1 pipe_addr_branch_reg_15_ ( .D(pcadd_o_addr_pcbranchE[15]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[15]) );
  DFC1 pipe_addr_branch_reg_14_ ( .D(pcadd_o_addr_pcbranchE[14]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[14]) );
  DFC1 pipe_signext_o_data_immD_reg_15_ ( .D(signext_o_data_immD[15]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[15]) );
  DFC1 pipe_FWmemout_reg_27_ ( .D(i_data_Wmemout[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[27]) );
  DFC1 pipe_addr_branch_reg_11_ ( .D(pcadd_o_addr_pcbranchE[11]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[11]) );
  DFC1 pipe_addr_pc4_reg_2_ ( .D(i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC1 pipe_addr_rd_reg_4_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[4]) );
  DFC3 pipe_FWmemout_reg_13_ ( .D(i_data_Wmemout[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[13]) );
  DFC1 pipe_FWmemout_reg_23_ ( .D(i_data_Wmemout[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[23]) );
  DFC1 pipe_FWmemout_reg_31_ ( .D(i_data_Wmemout[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[31]) );
  LOGIC0 U3 ( .Q(o_addr_jump[0]) );
  BUF15 U4 ( .A(i_data_instr[21]), .Q(n4) );
  CLKIN6 U5 ( .A(n5), .Q(n2) );
  INV12 U6 ( .A(n2), .Q(o_data_signext[1]) );
endmodule


module E_alu_DW01_add_12 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;

  NOR23 U2 ( .A(n24), .B(n52), .Q(n28) );
  NOR22 U3 ( .A(n24), .B(n53), .Q(n21) );
  NOR24 U4 ( .A(B[2]), .B(A[2]), .Q(n53) );
  NAND21 U5 ( .A(n70), .B(n52), .Q(SUM[0]) );
  XNR20 U6 ( .A(n4), .B(A[4]), .Q(n40) );
  NAND24 U7 ( .A(n41), .B(n42), .Q(n32) );
  NAND22 U8 ( .A(B[0]), .B(A[0]), .Q(n52) );
  INV3 U9 ( .A(n24), .Q(n65) );
  NOR22 U10 ( .A(A[3]), .B(B[3]), .Q(n47) );
  NOR21 U11 ( .A(n25), .B(n26), .Q(n50) );
  XOR21 U12 ( .A(n56), .B(n59), .Q(SUM[2]) );
  NOR21 U13 ( .A(n33), .B(n34), .Q(n14) );
  NOR21 U14 ( .A(n35), .B(n33), .Q(n8) );
  NOR23 U15 ( .A(n44), .B(n43), .Q(n42) );
  INV2 U16 ( .A(n26), .Q(n19) );
  INV3 U17 ( .A(n1), .Q(n35) );
  NAND22 U18 ( .A(n39), .B(n5), .Q(n1) );
  CLKIN1 U19 ( .A(n58), .Q(n57) );
  NOR22 U20 ( .A(A[5]), .B(B[5]), .Q(n33) );
  NOR21 U21 ( .A(A[0]), .B(B[0]), .Q(n64) );
  CLKIN0 U22 ( .A(B[0]), .Q(n71) );
  INV0 U23 ( .A(A[4]), .Q(n39) );
  INV6 U24 ( .A(B[4]), .Q(n5) );
  NOR22 U25 ( .A(n47), .B(n53), .Q(n46) );
  NOR23 U26 ( .A(A[1]), .B(B[1]), .Q(n24) );
  NAND21 U27 ( .A(B[1]), .B(A[1]), .Q(n69) );
  INV1 U28 ( .A(B[1]), .Q(n49) );
  NAND21 U29 ( .A(B[3]), .B(A[3]), .Q(n23) );
  NOR21 U30 ( .A(B[3]), .B(A[3]), .Q(n25) );
  NOR21 U31 ( .A(B[0]), .B(A[0]), .Q(n26) );
  NAND42 U32 ( .A(n15), .B(n16), .C(n17), .D(n18), .Q(n10) );
  AOI221 U33 ( .A(B[5]), .B(A[5]), .C(n4), .D(A[4]), .Q(n34) );
  AOI212 U34 ( .A(n55), .B(n56), .C(n57), .Q(n54) );
  AOI222 U35 ( .A(n50), .B(n21), .C(n51), .D(n28), .Q(n41) );
  NOR20 U36 ( .A(n53), .B(n47), .Q(n51) );
  NAND24 U37 ( .A(n45), .B(n46), .Q(n16) );
  OAI2111 U38 ( .A(A[3]), .B(B[3]), .C(A[2]), .D(B[2]), .Q(n15) );
  XOR22 U39 ( .A(n36), .B(n37), .Q(SUM[5]) );
  XOR22 U40 ( .A(n30), .B(n31), .Q(SUM[6]) );
  AOI312 U41 ( .A(n19), .B(n20), .C(n21), .D(n22), .Q(n18) );
  OAI210 U42 ( .A(B[2]), .B(A[2]), .C(n58), .Q(n60) );
  INV6 U43 ( .A(n5), .Q(n4) );
  NOR20 U44 ( .A(n39), .B(n5), .Q(n38) );
  XOR22 U45 ( .A(n6), .B(n7), .Q(SUM[7]) );
  INV3 U46 ( .A(n29), .Q(n9) );
  XNR21 U47 ( .A(n2), .B(n54), .Q(SUM[3]) );
  XOR20 U48 ( .A(B[3]), .B(A[3]), .Q(n2) );
  NAND21 U49 ( .A(n64), .B(n52), .Q(n67) );
  NOR20 U50 ( .A(n66), .B(n24), .Q(n68) );
  CLKIN3 U51 ( .A(n60), .Q(n59) );
  CLKIN2 U52 ( .A(n64), .Q(n63) );
  NAND22 U53 ( .A(n27), .B(n28), .Q(n17) );
  NAND22 U54 ( .A(n15), .B(n23), .Q(n44) );
  INV3 U55 ( .A(n25), .Q(n20) );
  INV3 U56 ( .A(n53), .Q(n55) );
  XOR21 U57 ( .A(n67), .B(n68), .Q(SUM[1]) );
  NAND22 U58 ( .A(n61), .B(n62), .Q(n56) );
  NAND22 U59 ( .A(n63), .B(n65), .Q(n62) );
  AOI310 U60 ( .A(A[0]), .B(B[0]), .C(n65), .D(n66), .Q(n61) );
  NOR21 U61 ( .A(n48), .B(n49), .Q(n45) );
  XNR21 U62 ( .A(B[7]), .B(A[7]), .Q(n6) );
  NAND22 U63 ( .A(n12), .B(n13), .Q(n11) );
  NAND20 U64 ( .A(B[2]), .B(A[2]), .Q(n58) );
  NAND22 U65 ( .A(n14), .B(n9), .Q(n12) );
  NAND22 U66 ( .A(n3), .B(n71), .Q(n70) );
  INV0 U67 ( .A(A[0]), .Q(n3) );
  NOR21 U68 ( .A(n53), .B(n47), .Q(n27) );
  XNR21 U69 ( .A(n32), .B(n40), .Q(SUM[4]) );
  NAND20 U70 ( .A(B[6]), .B(A[6]), .Q(n13) );
  CLKIN0 U71 ( .A(A[1]), .Q(n48) );
  NOR21 U72 ( .A(A[6]), .B(B[6]), .Q(n29) );
  XNR20 U73 ( .A(B[6]), .B(A[6]), .Q(n30) );
  XNR20 U74 ( .A(B[5]), .B(A[5]), .Q(n36) );
  AOI312 U75 ( .A(n8), .B(n9), .C(n10), .D(n11), .Q(n7) );
  CLKIN3 U76 ( .A(n23), .Q(n22) );
  AOI212 U77 ( .A(n8), .B(n32), .C(n14), .Q(n31) );
  AOI212 U78 ( .A(n1), .B(n32), .C(n38), .Q(n37) );
  CLKIN3 U79 ( .A(n16), .Q(n43) );
  CLKIN3 U80 ( .A(n69), .Q(n66) );
endmodule


module E_alu_DW01_add_13 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55;

  NOR23 U2 ( .A(B[2]), .B(A[2]), .Q(n43) );
  NOR21 U3 ( .A(A[4]), .B(n3), .Q(n27) );
  CLKIN0 U4 ( .A(A[4]), .Q(n32) );
  XNR20 U5 ( .A(n3), .B(A[4]), .Q(n33) );
  NOR22 U6 ( .A(A[3]), .B(B[3]), .Q(n20) );
  NOR22 U7 ( .A(A[1]), .B(B[1]), .Q(n17) );
  NAND22 U8 ( .A(B[0]), .B(A[0]), .Q(n42) );
  NOR21 U9 ( .A(n25), .B(n26), .Q(n13) );
  NOR21 U10 ( .A(n27), .B(n25), .Q(n7) );
  CLKIN1 U11 ( .A(B[1]), .Q(n41) );
  NOR21 U12 ( .A(n52), .B(n17), .Q(n53) );
  XOR22 U13 ( .A(n22), .B(n23), .Q(SUM[6]) );
  XOR22 U14 ( .A(n5), .B(n6), .Q(SUM[7]) );
  NOR22 U15 ( .A(n20), .B(n43), .Q(n39) );
  NAND21 U16 ( .A(B[1]), .B(A[1]), .Q(n54) );
  AOI311 U17 ( .A(A[0]), .B(B[0]), .C(n51), .D(n52), .Q(n50) );
  NAND21 U18 ( .A(B[3]), .B(A[3]), .Q(n16) );
  AOI221 U19 ( .A(B[5]), .B(A[5]), .C(n3), .D(A[4]), .Q(n26) );
  NOR21 U20 ( .A(A[5]), .B(B[5]), .Q(n25) );
  OAI2111 U21 ( .A(A[3]), .B(B[3]), .C(A[2]), .D(B[2]), .Q(n14) );
  NAND24 U22 ( .A(n38), .B(n39), .Q(n15) );
  XOR22 U23 ( .A(n28), .B(n29), .Q(SUM[5]) );
  XNR20 U24 ( .A(B[5]), .B(A[5]), .Q(n28) );
  OAI210 U25 ( .A(B[2]), .B(A[2]), .C(n48), .Q(n49) );
  NAND26 U26 ( .A(n34), .B(n35), .Q(n24) );
  NOR24 U27 ( .A(n36), .B(n37), .Q(n35) );
  INV3 U28 ( .A(n54), .Q(n52) );
  XNR21 U29 ( .A(n46), .B(n49), .Q(SUM[2]) );
  CLKIN3 U30 ( .A(B[4]), .Q(n4) );
  INV3 U31 ( .A(n21), .Q(n8) );
  INV2 U32 ( .A(n48), .Q(n47) );
  MUX21 U33 ( .A(B[0]), .B(n55), .S(A[0]), .Q(SUM[0]) );
  XNR21 U34 ( .A(n2), .B(n44), .Q(SUM[3]) );
  XOR20 U35 ( .A(B[3]), .B(A[3]), .Q(n2) );
  INV2 U36 ( .A(n50), .Q(n46) );
  CLKIN0 U37 ( .A(B[0]), .Q(n55) );
  NAND22 U38 ( .A(n18), .B(n19), .Q(n34) );
  NAND22 U39 ( .A(n14), .B(n16), .Q(n37) );
  XNR21 U40 ( .A(B[7]), .B(A[7]), .Q(n5) );
  NAND41 U41 ( .A(n14), .B(n15), .C(n34), .D(n16), .Q(n9) );
  AOI211 U42 ( .A(n45), .B(n46), .C(n47), .Q(n44) );
  INV3 U43 ( .A(n43), .Q(n45) );
  XNR21 U44 ( .A(n42), .B(n53), .Q(SUM[1]) );
  NOR21 U45 ( .A(n40), .B(n41), .Q(n38) );
  NAND20 U46 ( .A(B[2]), .B(A[2]), .Q(n48) );
  NOR21 U47 ( .A(n43), .B(n20), .Q(n18) );
  NOR21 U48 ( .A(n17), .B(n42), .Q(n19) );
  INV3 U49 ( .A(n17), .Q(n51) );
  INV3 U50 ( .A(n27), .Q(n30) );
  INV3 U51 ( .A(n4), .Q(n3) );
  NOR21 U52 ( .A(n32), .B(n4), .Q(n31) );
  XNR20 U53 ( .A(B[6]), .B(A[6]), .Q(n22) );
  XNR21 U54 ( .A(n24), .B(n33), .Q(SUM[4]) );
  NAND22 U55 ( .A(n11), .B(n12), .Q(n10) );
  NAND20 U56 ( .A(B[6]), .B(A[6]), .Q(n12) );
  NAND22 U57 ( .A(n13), .B(n8), .Q(n11) );
  CLKIN0 U58 ( .A(A[1]), .Q(n40) );
  NOR21 U59 ( .A(A[6]), .B(B[6]), .Q(n21) );
  AOI312 U60 ( .A(n7), .B(n8), .C(n9), .D(n10), .Q(n6) );
  AOI212 U61 ( .A(n7), .B(n24), .C(n13), .Q(n23) );
  AOI212 U62 ( .A(n30), .B(n24), .C(n31), .Q(n29) );
  CLKIN3 U63 ( .A(n15), .Q(n36) );
endmodule


module E_alu_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   ML_int_1__31_, ML_int_1__30_, ML_int_1__29_, ML_int_1__28_,
         ML_int_1__27_, ML_int_1__26_, ML_int_1__25_, ML_int_1__24_,
         ML_int_1__23_, ML_int_1__22_, ML_int_1__21_, ML_int_1__20_,
         ML_int_1__19_, ML_int_1__18_, ML_int_1__17_, ML_int_1__16_,
         ML_int_1__15_, ML_int_1__14_, ML_int_1__13_, ML_int_1__12_,
         ML_int_1__11_, ML_int_1__10_, ML_int_1__9_, ML_int_1__8_,
         ML_int_1__7_, ML_int_1__6_, ML_int_1__5_, ML_int_1__4_, ML_int_1__3_,
         ML_int_1__2_, ML_int_1__1_, ML_int_1__0_, ML_int_2__31_,
         ML_int_2__30_, ML_int_2__29_, ML_int_2__28_, ML_int_2__27_,
         ML_int_2__26_, ML_int_2__25_, ML_int_2__24_, ML_int_2__23_,
         ML_int_2__22_, ML_int_2__21_, ML_int_2__20_, ML_int_2__19_,
         ML_int_2__18_, ML_int_2__17_, ML_int_2__16_, ML_int_2__15_,
         ML_int_2__14_, ML_int_2__13_, ML_int_2__12_, ML_int_2__11_,
         ML_int_2__10_, ML_int_2__9_, ML_int_2__8_, ML_int_2__7_, ML_int_2__6_,
         ML_int_2__5_, ML_int_2__4_, ML_int_2__3_, ML_int_2__2_, ML_int_2__1_,
         ML_int_2__0_, ML_int_3__31_, ML_int_3__30_, ML_int_3__29_,
         ML_int_3__28_, ML_int_3__27_, ML_int_3__26_, ML_int_3__25_,
         ML_int_3__24_, ML_int_3__23_, ML_int_3__22_, ML_int_3__21_,
         ML_int_3__20_, ML_int_3__19_, ML_int_3__18_, ML_int_3__17_,
         ML_int_3__16_, ML_int_3__15_, ML_int_3__14_, ML_int_3__13_,
         ML_int_3__12_, ML_int_3__11_, ML_int_3__10_, ML_int_3__9_,
         ML_int_3__8_, ML_int_3__7_, ML_int_3__6_, ML_int_3__5_, ML_int_3__4_,
         ML_int_3__3_, ML_int_3__2_, ML_int_3__1_, ML_int_3__0_, ML_int_4__31_,
         ML_int_4__30_, ML_int_4__29_, ML_int_4__28_, ML_int_4__27_,
         ML_int_4__26_, ML_int_4__25_, ML_int_4__24_, ML_int_4__23_,
         ML_int_4__22_, ML_int_4__21_, ML_int_4__20_, ML_int_4__19_,
         ML_int_4__18_, ML_int_4__17_, ML_int_4__15_, ML_int_4__14_,
         ML_int_4__13_, ML_int_4__12_, ML_int_4__11_, ML_int_4__10_,
         ML_int_4__9_, ML_int_4__8_, ML_int_4__7_, ML_int_4__6_, ML_int_4__5_,
         ML_int_4__4_, ML_int_4__3_, ML_int_4__2_, ML_int_4__1_, ML_int_4__0_,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;

  MUX21 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n41), .Q(ML_int_1__3_) );
  MUX22 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n41), .Q(ML_int_1__8_) );
  MUX22 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n43), .Q(ML_int_1__29_) );
  MUX22 M1_2_24 ( .A(ML_int_2__24_), .B(ML_int_2__20_), .S(n52), .Q(
        ML_int_3__24_) );
  MUX22 M1_3_24 ( .A(ML_int_3__24_), .B(ML_int_3__16_), .S(n58), .Q(
        ML_int_4__24_) );
  MUX22 M1_4_24 ( .A(ML_int_4__24_), .B(ML_int_4__8_), .S(SH[4]), .Q(B[24]) );
  MUX22 M1_2_28 ( .A(ML_int_2__28_), .B(ML_int_2__24_), .S(n53), .Q(
        ML_int_3__28_) );
  MUX22 M1_3_28 ( .A(ML_int_3__28_), .B(ML_int_3__20_), .S(n59), .Q(
        ML_int_4__28_) );
  MUX22 M1_2_26 ( .A(ML_int_2__26_), .B(ML_int_2__22_), .S(n53), .Q(
        ML_int_3__26_) );
  MUX22 M1_3_26 ( .A(ML_int_3__26_), .B(ML_int_3__18_), .S(n59), .Q(
        ML_int_4__26_) );
  MUX22 M1_4_26 ( .A(ML_int_4__26_), .B(ML_int_4__10_), .S(n61), .Q(B[26]) );
  MUX22 M1_4_27 ( .A(ML_int_4__27_), .B(ML_int_4__11_), .S(n61), .Q(B[27]) );
  MUX22 M1_4_23 ( .A(ML_int_4__23_), .B(ML_int_4__7_), .S(n61), .Q(B[23]) );
  MUX22 M1_2_25 ( .A(ML_int_2__25_), .B(ML_int_2__21_), .S(n53), .Q(
        ML_int_3__25_) );
  MUX22 M1_3_25 ( .A(ML_int_3__25_), .B(ML_int_3__17_), .S(n59), .Q(
        ML_int_4__25_) );
  MUX22 M1_4_25 ( .A(ML_int_4__25_), .B(ML_int_4__9_), .S(n61), .Q(B[25]) );
  MUX22 M1_1_30 ( .A(ML_int_1__30_), .B(ML_int_1__28_), .S(n46), .Q(
        ML_int_2__30_) );
  MUX22 M1_3_30 ( .A(ML_int_3__30_), .B(ML_int_3__22_), .S(n54), .Q(
        ML_int_4__30_) );
  MUX22 M1_1_31 ( .A(ML_int_1__31_), .B(ML_int_1__29_), .S(SH[1]), .Q(
        ML_int_2__31_) );
  MUX22 M1_2_31 ( .A(ML_int_2__31_), .B(ML_int_2__27_), .S(n53), .Q(
        ML_int_3__31_) );
  MUX22 M1_2_29 ( .A(ML_int_2__29_), .B(ML_int_2__25_), .S(n53), .Q(
        ML_int_3__29_) );
  MUX22 M1_3_14 ( .A(ML_int_3__14_), .B(ML_int_3__6_), .S(n56), .Q(
        ML_int_4__14_) );
  MUX22 M1_3_13 ( .A(ML_int_3__13_), .B(ML_int_3__5_), .S(n56), .Q(
        ML_int_4__13_) );
  MUX22 M1_2_7 ( .A(ML_int_2__7_), .B(ML_int_2__3_), .S(n49), .Q(ML_int_3__7_)
         );
  MUX22 M1_3_11 ( .A(ML_int_3__11_), .B(ML_int_3__3_), .S(n56), .Q(
        ML_int_4__11_) );
  MUX22 M1_3_9 ( .A(ML_int_3__9_), .B(ML_int_3__1_), .S(n55), .Q(ML_int_4__9_)
         );
  MUX22 M1_2_22 ( .A(ML_int_2__22_), .B(ML_int_2__18_), .S(n52), .Q(
        ML_int_3__22_) );
  MUX22 M1_1_23 ( .A(ML_int_1__23_), .B(ML_int_1__21_), .S(n47), .Q(
        ML_int_2__23_) );
  MUX21 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n43), .Q(ML_int_1__27_) );
  MUX22 M1_1_19 ( .A(ML_int_1__19_), .B(ML_int_1__17_), .S(n46), .Q(
        ML_int_2__19_) );
  MUX22 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n41), .Q(ML_int_1__6_) );
  MUX22 M1_1_5 ( .A(ML_int_1__5_), .B(ML_int_1__3_), .S(n46), .Q(ML_int_2__5_)
         );
  MUX22 M1_1_12 ( .A(ML_int_1__12_), .B(ML_int_1__10_), .S(n45), .Q(
        ML_int_2__12_) );
  MUX21 M1_1_29 ( .A(ML_int_1__29_), .B(ML_int_1__27_), .S(SH[1]), .Q(
        ML_int_2__29_) );
  MUX22 M1_4_19 ( .A(ML_int_4__19_), .B(ML_int_4__3_), .S(n61), .Q(B[19]) );
  MUX22 M1_2_9 ( .A(ML_int_2__9_), .B(ML_int_2__5_), .S(n49), .Q(ML_int_3__9_)
         );
  MUX22 M1_1_11 ( .A(ML_int_1__11_), .B(ML_int_1__9_), .S(n45), .Q(
        ML_int_2__11_) );
  MUX22 M1_1_28 ( .A(ML_int_1__28_), .B(ML_int_1__26_), .S(SH[1]), .Q(
        ML_int_2__28_) );
  MUX21 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n43), .Q(ML_int_1__31_) );
  MUX22 M1_1_17 ( .A(ML_int_1__17_), .B(ML_int_1__15_), .S(n46), .Q(
        ML_int_2__17_) );
  MUX22 M1_1_24 ( .A(ML_int_1__24_), .B(ML_int_1__22_), .S(n47), .Q(
        ML_int_2__24_) );
  MUX22 M1_2_5 ( .A(ML_int_2__5_), .B(ML_int_2__1_), .S(n49), .Q(ML_int_3__5_)
         );
  MUX22 M1_1_3 ( .A(ML_int_1__3_), .B(ML_int_1__1_), .S(n44), .Q(ML_int_2__3_)
         );
  MUX22 M1_3_10 ( .A(ML_int_3__10_), .B(ML_int_3__2_), .S(n56), .Q(
        ML_int_4__10_) );
  MUX22 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n41), .Q(ML_int_1__25_) );
  MUX22 M1_1_27 ( .A(ML_int_1__27_), .B(ML_int_1__25_), .S(n47), .Q(
        ML_int_2__27_) );
  MUX26 M1_2_6 ( .A(ML_int_2__6_), .B(ML_int_2__2_), .S(n49), .Q(ML_int_3__6_)
         );
  MUX24 M1_4_22 ( .A(ML_int_4__22_), .B(ML_int_4__6_), .S(n61), .Q(B[22]) );
  MUX22 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n41), .Q(ML_int_1__9_) );
  MUX24 M1_2_16 ( .A(ML_int_2__16_), .B(ML_int_2__12_), .S(n51), .Q(
        ML_int_3__16_) );
  MUX24 M1_2_19 ( .A(ML_int_2__19_), .B(ML_int_2__15_), .S(n51), .Q(
        ML_int_3__19_) );
  MUX22 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n41), .Q(ML_int_1__19_) );
  MUX22 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n41), .Q(ML_int_1__5_) );
  MUX22 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n42), .Q(ML_int_1__12_) );
  MUX24 M1_4_31 ( .A(ML_int_4__31_), .B(ML_int_4__15_), .S(SH[4]), .Q(B[31])
         );
  MUX22 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n42), .Q(ML_int_1__13_) );
  MUX26 M1_3_15 ( .A(ML_int_3__15_), .B(ML_int_3__7_), .S(n57), .Q(
        ML_int_4__15_) );
  MUX24 M1_2_10 ( .A(ML_int_2__10_), .B(ML_int_2__6_), .S(n50), .Q(
        ML_int_3__10_) );
  MUX22 M1_4_28 ( .A(ML_int_4__28_), .B(ML_int_4__12_), .S(SH[4]), .Q(B[28])
         );
  MUX22 M1_3_22 ( .A(ML_int_3__22_), .B(ML_int_3__14_), .S(n58), .Q(
        ML_int_4__22_) );
  MUX24 M1_4_18 ( .A(ML_int_4__18_), .B(ML_int_4__2_), .S(n60), .Q(B[18]) );
  MUX24 M1_2_27 ( .A(ML_int_2__27_), .B(ML_int_2__23_), .S(n53), .Q(
        ML_int_3__27_) );
  MUX22 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n42), .Q(ML_int_1__14_) );
  MUX22 M1_1_9 ( .A(ML_int_1__9_), .B(ML_int_1__7_), .S(n45), .Q(ML_int_2__9_)
         );
  MUX24 M1_4_20 ( .A(ML_int_4__20_), .B(ML_int_4__4_), .S(SH[4]), .Q(B[20]) );
  MUX22 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n42), .Q(ML_int_1__18_) );
  MUX26 M1_3_18 ( .A(ML_int_3__18_), .B(ML_int_3__10_), .S(n57), .Q(
        ML_int_4__18_) );
  MUX24 M1_2_23 ( .A(ML_int_2__23_), .B(ML_int_2__19_), .S(n52), .Q(
        ML_int_3__23_) );
  MUX24 M1_3_31 ( .A(ML_int_3__31_), .B(ML_int_3__23_), .S(n54), .Q(
        ML_int_4__31_) );
  MUX22 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n43), .Q(ML_int_1__4_) );
  MUX24 M1_1_8 ( .A(ML_int_1__8_), .B(ML_int_1__6_), .S(n44), .Q(ML_int_2__8_)
         );
  MUX26 M1_2_8 ( .A(ML_int_2__8_), .B(ML_int_2__4_), .S(n49), .Q(ML_int_3__8_)
         );
  MUX26 M1_3_19 ( .A(ML_int_3__19_), .B(ML_int_3__11_), .S(n57), .Q(
        ML_int_4__19_) );
  MUX22 M1_3_17 ( .A(ML_int_3__17_), .B(ML_int_3__9_), .S(n57), .Q(
        ML_int_4__17_) );
  MUX22 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n43), .Q(ML_int_1__23_) );
  MUX24 M1_3_21 ( .A(ML_int_3__21_), .B(ML_int_3__13_), .S(n58), .Q(
        ML_int_4__21_) );
  MUX26 M1_3_20 ( .A(ML_int_3__20_), .B(ML_int_3__12_), .S(n58), .Q(
        ML_int_4__20_) );
  MUX22 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n41), .Q(ML_int_1__17_) );
  MUX22 M1_1_4 ( .A(ML_int_1__4_), .B(ML_int_1__2_), .S(n44), .Q(ML_int_2__4_)
         );
  NOR24 U3 ( .A(n60), .B(n15), .Q(B[10]) );
  INV6 U4 ( .A(ML_int_4__10_), .Q(n15) );
  INV3 U5 ( .A(ML_int_3__1_), .Q(n32) );
  MUX22 U6 ( .A(ML_int_1__13_), .B(ML_int_1__11_), .S(n45), .Q(ML_int_2__13_)
         );
  NOR24 U7 ( .A(n60), .B(n11), .Q(B[14]) );
  NOR24 U8 ( .A(n60), .B(n13), .Q(B[12]) );
  IMUX21 U9 ( .A(n25), .B(n4), .S(n3), .Q(B[16]) );
  INV3 U10 ( .A(n50), .Q(n1) );
  NOR22 U11 ( .A(n48), .B(n39), .Q(ML_int_3__3_) );
  NAND22 U12 ( .A(n5), .B(n6), .Q(ML_int_3__4_) );
  MUX22 U13 ( .A(ML_int_2__12_), .B(ML_int_2__8_), .S(n50), .Q(ML_int_3__12_)
         );
  MUX22 U14 ( .A(ML_int_1__18_), .B(ML_int_1__16_), .S(n46), .Q(ML_int_2__18_)
         );
  MUX22 U15 ( .A(ML_int_2__20_), .B(ML_int_2__16_), .S(n52), .Q(ML_int_3__20_)
         );
  MUX22 U16 ( .A(ML_int_1__25_), .B(ML_int_1__23_), .S(SH[1]), .Q(
        ML_int_2__25_) );
  NOR22 U17 ( .A(n54), .B(n31), .Q(ML_int_4__2_) );
  MUX22 U18 ( .A(ML_int_3__12_), .B(ML_int_3__4_), .S(n56), .Q(ML_int_4__12_)
         );
  MUX22 U19 ( .A(ML_int_1__26_), .B(ML_int_1__24_), .S(SH[1]), .Q(
        ML_int_2__26_) );
  NOR22 U20 ( .A(n60), .B(n14), .Q(B[11]) );
  MUX22 U21 ( .A(ML_int_2__9_), .B(ML_int_2__13_), .S(n1), .Q(ML_int_3__13_)
         );
  MUX26 U22 ( .A(ML_int_4__17_), .B(ML_int_4__1_), .S(n60), .Q(B[17]) );
  INV3 U23 ( .A(ML_int_4__7_), .Q(n18) );
  CLKIN3 U24 ( .A(ML_int_4__13_), .Q(n12) );
  MUX26 U25 ( .A(ML_int_4__29_), .B(ML_int_4__13_), .S(SH[4]), .Q(B[29]) );
  NOR22 U26 ( .A(n60), .B(n16), .Q(B[9]) );
  MUX22 U27 ( .A(A[7]), .B(A[6]), .S(n41), .Q(ML_int_1__7_) );
  MUX22 U28 ( .A(A[26]), .B(A[25]), .S(n43), .Q(ML_int_1__26_) );
  BUF2 U29 ( .A(SH[2]), .Q(n51) );
  NOR23 U30 ( .A(n44), .B(n35), .Q(ML_int_2__0_) );
  MUX22 U31 ( .A(ML_int_2__11_), .B(ML_int_2__7_), .S(n50), .Q(ML_int_3__11_)
         );
  NOR22 U32 ( .A(n55), .B(n27), .Q(ML_int_4__6_) );
  INV3 U33 ( .A(ML_int_3__6_), .Q(n27) );
  INV3 U34 ( .A(n60), .Q(n3) );
  MUX22 U35 ( .A(A[30]), .B(A[29]), .S(n42), .Q(ML_int_1__30_) );
  NOR22 U36 ( .A(n55), .B(n28), .Q(ML_int_4__5_) );
  NAND22 U37 ( .A(n8), .B(n9), .Q(ML_int_3__15_) );
  INV3 U38 ( .A(ML_int_3__7_), .Q(n26) );
  NOR22 U39 ( .A(n54), .B(n29), .Q(ML_int_4__4_) );
  NOR22 U40 ( .A(n61), .B(n25), .Q(B[0]) );
  INV3 U41 ( .A(ML_int_4__2_), .Q(n23) );
  INV3 U42 ( .A(ML_int_4__12_), .Q(n13) );
  INV3 U43 ( .A(SH[0]), .Q(n2) );
  MUX22 U44 ( .A(ML_int_1__2_), .B(ML_int_1__0_), .S(n44), .Q(ML_int_2__2_) );
  NOR22 U45 ( .A(n48), .B(n38), .Q(ML_int_3__1_) );
  NOR22 U46 ( .A(n48), .B(n34), .Q(ML_int_3__0_) );
  INV3 U47 ( .A(ML_int_2__0_), .Q(n34) );
  MUX22 U48 ( .A(ML_int_1__14_), .B(ML_int_1__12_), .S(n45), .Q(ML_int_2__14_)
         );
  NOR22 U49 ( .A(n54), .B(n30), .Q(ML_int_4__3_) );
  MUX22 U50 ( .A(ML_int_3__8_), .B(ML_int_3__0_), .S(n55), .Q(ML_int_4__8_) );
  MUX22 U51 ( .A(ML_int_2__30_), .B(ML_int_2__26_), .S(n53), .Q(ML_int_3__30_)
         );
  NOR22 U52 ( .A(n60), .B(n18), .Q(B[7]) );
  INV3 U53 ( .A(ML_int_4__5_), .Q(n20) );
  MUX22 U54 ( .A(ML_int_3__27_), .B(ML_int_3__19_), .S(n59), .Q(ML_int_4__27_)
         );
  MUX22 U55 ( .A(ML_int_3__23_), .B(ML_int_3__15_), .S(n58), .Q(ML_int_4__23_)
         );
  MUX24 U56 ( .A(ML_int_1__22_), .B(ML_int_1__20_), .S(n47), .Q(ML_int_2__22_)
         );
  MUX22 U57 ( .A(A[10]), .B(A[9]), .S(n42), .Q(ML_int_1__10_) );
  NOR22 U58 ( .A(SH[0]), .B(n36), .Q(ML_int_1__0_) );
  INV2 U59 ( .A(A[0]), .Q(n36) );
  BUF2 U60 ( .A(SH[2]), .Q(n48) );
  CLKIN6 U61 ( .A(ML_int_2__2_), .Q(n37) );
  NOR22 U62 ( .A(n44), .B(n40), .Q(ML_int_2__1_) );
  MUX22 U63 ( .A(ML_int_1__6_), .B(ML_int_1__4_), .S(n47), .Q(ML_int_2__6_) );
  MUX22 U64 ( .A(ML_int_1__15_), .B(ML_int_1__13_), .S(n46), .Q(ML_int_2__15_)
         );
  MUX22 U65 ( .A(ML_int_1__16_), .B(ML_int_1__14_), .S(n46), .Q(ML_int_2__16_)
         );
  MUX24 U66 ( .A(ML_int_3__29_), .B(ML_int_3__21_), .S(n59), .Q(ML_int_4__29_)
         );
  MUX24 U67 ( .A(ML_int_2__21_), .B(ML_int_2__17_), .S(n52), .Q(ML_int_3__21_)
         );
  MUX22 U68 ( .A(ML_int_2__18_), .B(ML_int_2__14_), .S(n51), .Q(ML_int_3__18_)
         );
  MUX24 U69 ( .A(ML_int_2__17_), .B(ML_int_2__13_), .S(n51), .Q(ML_int_3__17_)
         );
  MUX22 U70 ( .A(A[20]), .B(A[19]), .S(n43), .Q(ML_int_1__20_) );
  MUX22 U71 ( .A(A[1]), .B(A[0]), .S(n42), .Q(ML_int_1__1_) );
  CLKIN3 U72 ( .A(ML_int_2__1_), .Q(n38) );
  MUX22 U73 ( .A(ML_int_1__7_), .B(ML_int_1__5_), .S(n45), .Q(ML_int_2__7_) );
  CLKIN2 U74 ( .A(ML_int_2__3_), .Q(n39) );
  MUX22 U75 ( .A(A[15]), .B(A[14]), .S(n42), .Q(ML_int_1__15_) );
  MUX22 U76 ( .A(A[10]), .B(A[11]), .S(n2), .Q(ML_int_1__11_) );
  MUX22 U77 ( .A(A[21]), .B(A[20]), .S(n43), .Q(ML_int_1__21_) );
  MUX22 U78 ( .A(A[16]), .B(A[15]), .S(n42), .Q(ML_int_1__16_) );
  MUX24 U79 ( .A(ML_int_1__10_), .B(ML_int_1__8_), .S(n45), .Q(ML_int_2__10_)
         );
  MUX22 U80 ( .A(A[24]), .B(A[23]), .S(n43), .Q(ML_int_1__24_) );
  MUX24 U81 ( .A(ML_int_4__30_), .B(ML_int_4__14_), .S(SH[4]), .Q(B[30]) );
  MUX22 U82 ( .A(A[22]), .B(A[21]), .S(n43), .Q(ML_int_1__22_) );
  MUX21 U83 ( .A(A[28]), .B(A[27]), .S(n43), .Q(ML_int_1__28_) );
  MUX26 U84 ( .A(ML_int_4__21_), .B(ML_int_4__5_), .S(SH[4]), .Q(B[21]) );
  INV2 U85 ( .A(ML_int_1__1_), .Q(n40) );
  MUX26 U86 ( .A(ML_int_2__14_), .B(ML_int_2__10_), .S(n50), .Q(ML_int_3__14_)
         );
  MUX22 U87 ( .A(ML_int_1__21_), .B(ML_int_1__19_), .S(n47), .Q(ML_int_2__21_)
         );
  MUX22 U88 ( .A(ML_int_1__20_), .B(ML_int_1__18_), .S(n47), .Q(ML_int_2__20_)
         );
  MUX22 U89 ( .A(A[1]), .B(A[2]), .S(n2), .Q(ML_int_1__2_) );
  CLKIN2 U90 ( .A(ML_int_4__3_), .Q(n22) );
  NOR22 U91 ( .A(n60), .B(n12), .Q(B[13]) );
  IMUX21 U92 ( .A(ML_int_3__16_), .B(ML_int_3__8_), .S(n57), .Q(n4) );
  NOR23 U93 ( .A(n54), .B(n33), .Q(ML_int_4__0_) );
  CLKIN4 U94 ( .A(ML_int_4__0_), .Q(n25) );
  NOR22 U95 ( .A(n54), .B(n32), .Q(ML_int_4__1_) );
  CLKIN3 U96 ( .A(ML_int_4__4_), .Q(n21) );
  NOR24 U97 ( .A(n55), .B(n26), .Q(ML_int_4__7_) );
  NOR24 U98 ( .A(n48), .B(n37), .Q(ML_int_3__2_) );
  CLKIN6 U99 ( .A(ML_int_4__15_), .Q(n10) );
  NAND21 U100 ( .A(ML_int_2__4_), .B(n7), .Q(n5) );
  NAND22 U101 ( .A(ML_int_2__0_), .B(n48), .Q(n6) );
  CLKIN2 U102 ( .A(ML_int_3__4_), .Q(n29) );
  NAND22 U103 ( .A(ML_int_2__15_), .B(n7), .Q(n8) );
  NAND22 U104 ( .A(ML_int_2__11_), .B(n51), .Q(n9) );
  INV3 U105 ( .A(n51), .Q(n7) );
  INV2 U106 ( .A(ML_int_3__2_), .Q(n31) );
  INV3 U107 ( .A(ML_int_1__0_), .Q(n35) );
  CLKIN3 U108 ( .A(ML_int_4__6_), .Q(n19) );
  INV2 U109 ( .A(ML_int_4__1_), .Q(n24) );
  INV2 U110 ( .A(ML_int_3__0_), .Q(n33) );
  INV3 U111 ( .A(ML_int_4__9_), .Q(n16) );
  INV3 U112 ( .A(ML_int_4__14_), .Q(n11) );
  INV3 U113 ( .A(ML_int_3__5_), .Q(n28) );
  INV3 U114 ( .A(ML_int_3__3_), .Q(n30) );
  INV3 U115 ( .A(ML_int_4__11_), .Q(n14) );
  NOR21 U116 ( .A(n60), .B(n19), .Q(B[6]) );
  NOR21 U117 ( .A(n60), .B(n17), .Q(B[8]) );
  INV3 U118 ( .A(ML_int_4__8_), .Q(n17) );
  NOR21 U119 ( .A(n60), .B(n10), .Q(B[15]) );
  NOR21 U120 ( .A(n61), .B(n22), .Q(B[3]) );
  NOR21 U121 ( .A(n61), .B(n20), .Q(B[5]) );
  NOR21 U122 ( .A(n61), .B(n24), .Q(B[1]) );
  NOR21 U123 ( .A(n61), .B(n21), .Q(B[4]) );
  NOR21 U124 ( .A(n61), .B(n23), .Q(B[2]) );
  BUF2 U125 ( .A(SH[0]), .Q(n41) );
  BUF2 U126 ( .A(SH[0]), .Q(n42) );
  BUF2 U127 ( .A(SH[4]), .Q(n60) );
  BUF2 U128 ( .A(SH[0]), .Q(n43) );
  BUF2 U129 ( .A(SH[2]), .Q(n49) );
  BUF2 U130 ( .A(SH[2]), .Q(n50) );
  BUF2 U131 ( .A(SH[1]), .Q(n47) );
  BUF2 U132 ( .A(SH[1]), .Q(n46) );
  BUF2 U133 ( .A(SH[2]), .Q(n53) );
  BUF2 U134 ( .A(SH[2]), .Q(n52) );
  BUF2 U135 ( .A(SH[3]), .Q(n56) );
  BUF2 U136 ( .A(SH[3]), .Q(n57) );
  BUF2 U137 ( .A(SH[3]), .Q(n58) );
  BUF2 U138 ( .A(SH[3]), .Q(n59) );
  BUF2 U139 ( .A(SH[1]), .Q(n44) );
  BUF2 U140 ( .A(SH[1]), .Q(n45) );
  BUF2 U141 ( .A(SH[3]), .Q(n55) );
  BUF2 U142 ( .A(SH[3]), .Q(n54) );
  BUF2 U143 ( .A(SH[4]), .Q(n61) );
endmodule


module E_alu_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187;

  CLKIN2 U3 ( .A(n50), .Q(n45) );
  OAI2112 U4 ( .A(n166), .B(n160), .C(n46), .D(n43), .Q(n165) );
  INV2 U5 ( .A(n159), .Q(n166) );
  INV10 U6 ( .A(B[11]), .Q(n37) );
  NOR24 U7 ( .A(A[4]), .B(n33), .Q(n184) );
  NAND28 U8 ( .A(n18), .B(n139), .Q(n137) );
  NAND24 U9 ( .A(n47), .B(n1), .Q(n18) );
  NAND24 U10 ( .A(n165), .B(n47), .Q(n163) );
  NOR24 U11 ( .A(n115), .B(n116), .Q(n114) );
  INV2 U12 ( .A(B[8]), .Q(n35) );
  NOR21 U13 ( .A(n16), .B(A[10]), .Q(n161) );
  CLKIN4 U14 ( .A(n61), .Q(n55) );
  INV4 U15 ( .A(A[2]), .Q(n182) );
  CLKIN12 U16 ( .A(A[1]), .Q(n180) );
  NAND26 U17 ( .A(n114), .B(n15), .Q(n111) );
  INV6 U18 ( .A(n12), .Q(n116) );
  CLKIN12 U19 ( .A(n32), .Q(n31) );
  INV6 U20 ( .A(B[0]), .Q(n32) );
  NAND23 U21 ( .A(A[7]), .B(n34), .Q(n122) );
  NOR23 U22 ( .A(n148), .B(n149), .Q(n144) );
  NAND22 U23 ( .A(n35), .B(A[8]), .Q(n1) );
  INV3 U24 ( .A(n13), .Q(n14) );
  NAND22 U25 ( .A(n57), .B(n126), .Q(n13) );
  INV6 U26 ( .A(B[9]), .Q(n141) );
  NAND23 U27 ( .A(n3), .B(n178), .Q(n113) );
  NAND24 U28 ( .A(n36), .B(A[10]), .Q(n156) );
  NAND23 U29 ( .A(n22), .B(n4), .Q(n25) );
  INV3 U30 ( .A(A[10]), .Q(n40) );
  INV6 U31 ( .A(B[7]), .Q(n34) );
  NOR24 U32 ( .A(A[9]), .B(n141), .Q(n148) );
  BUF2 U33 ( .A(B[8]), .Q(n28) );
  CLKIN6 U34 ( .A(n160), .Q(n158) );
  INV4 U35 ( .A(n174), .Q(n15) );
  NAND28 U36 ( .A(n10), .B(n57), .Q(n9) );
  INV8 U37 ( .A(n186), .Q(n10) );
  NAND28 U38 ( .A(n7), .B(n54), .Q(n131) );
  INV6 U39 ( .A(n10), .Q(n7) );
  CLKIN4 U40 ( .A(B[6]), .Q(n172) );
  INV10 U41 ( .A(B[10]), .Q(n36) );
  NAND23 U42 ( .A(n143), .B(n122), .Q(n20) );
  NAND26 U43 ( .A(n172), .B(A[6]), .Q(n54) );
  NAND28 U44 ( .A(n144), .B(n145), .Q(n129) );
  INV12 U45 ( .A(n129), .Q(n110) );
  NAND22 U46 ( .A(n136), .B(n137), .Q(n6) );
  NAND24 U47 ( .A(n136), .B(n137), .Q(n119) );
  CLKIN6 U48 ( .A(B[4]), .Q(n33) );
  NAND24 U49 ( .A(A[4]), .B(n33), .Q(n59) );
  INV6 U50 ( .A(n173), .Q(n67) );
  INV3 U51 ( .A(n115), .Q(n176) );
  NOR21 U52 ( .A(n31), .B(n38), .Q(n85) );
  NOR22 U53 ( .A(n182), .B(B[2]), .Q(n3) );
  NAND24 U54 ( .A(n159), .B(n21), .Q(n44) );
  NOR23 U55 ( .A(n121), .B(n122), .Q(n120) );
  XOR21 U56 ( .A(n133), .B(n132), .Q(DIFF[12]) );
  XOR21 U57 ( .A(n62), .B(n63), .Q(DIFF[6]) );
  INV3 U58 ( .A(n3), .Q(n82) );
  INV6 U59 ( .A(B[5]), .Q(n170) );
  NOR23 U60 ( .A(A[7]), .B(n34), .Q(n185) );
  NAND43 U61 ( .A(A[0]), .B(n77), .C(n178), .D(n179), .Q(n117) );
  NAND28 U62 ( .A(n112), .B(n113), .Q(n174) );
  NAND26 U63 ( .A(B[2]), .B(n182), .Q(n77) );
  NOR32 U64 ( .A(n9), .B(n184), .C(n185), .Q(n5) );
  NOR32 U65 ( .A(n9), .B(n184), .C(n185), .Q(n109) );
  NAND43 U66 ( .A(A[0]), .B(n77), .C(n178), .D(n179), .Q(n12) );
  INV3 U67 ( .A(A[8]), .Q(n39) );
  IMUX20 U68 ( .A(n31), .B(n32), .S(A[0]), .Q(DIFF[0]) );
  INV3 U69 ( .A(A[0]), .Q(n38) );
  INV3 U70 ( .A(n47), .Q(n138) );
  NAND23 U71 ( .A(A[9]), .B(n141), .Q(n47) );
  NOR20 U72 ( .A(A[13]), .B(n102), .Q(n101) );
  NAND20 U73 ( .A(n58), .B(n60), .Q(n68) );
  NAND21 U74 ( .A(B[5]), .B(n71), .Q(n58) );
  NAND23 U75 ( .A(n53), .B(n54), .Q(n51) );
  INV3 U76 ( .A(A[3]), .Q(n177) );
  OAI211 U77 ( .A(n80), .B(n84), .C(n81), .Q(n76) );
  INV3 U78 ( .A(n23), .Q(n4) );
  CLKIN3 U79 ( .A(B[1]), .Q(n183) );
  INV2 U80 ( .A(n164), .Q(n23) );
  CLKIN4 U81 ( .A(n163), .Q(n22) );
  NAND26 U82 ( .A(B[1]), .B(n180), .Q(n86) );
  NAND22 U83 ( .A(n61), .B(n59), .Q(n64) );
  NOR24 U84 ( .A(n130), .B(n129), .Q(n128) );
  NAND21 U85 ( .A(n28), .B(n39), .Q(n43) );
  NAND42 U86 ( .A(n108), .B(n5), .C(n110), .D(n111), .Q(n8) );
  NAND26 U87 ( .A(B[12]), .B(n125), .Q(n108) );
  NAND26 U88 ( .A(B[6]), .B(n187), .Q(n57) );
  NAND24 U89 ( .A(n131), .B(n108), .Q(n130) );
  INV0 U90 ( .A(A[5]), .Q(n71) );
  NAND24 U91 ( .A(A[1]), .B(n183), .Q(n81) );
  NOR24 U92 ( .A(n123), .B(n121), .Q(n118) );
  CLKIN2 U93 ( .A(A[6]), .Q(n187) );
  INV2 U94 ( .A(A[12]), .Q(n125) );
  INV0 U95 ( .A(n60), .Q(n65) );
  NAND20 U96 ( .A(n59), .B(n60), .Q(n56) );
  NAND34 U97 ( .A(n59), .B(n54), .C(n60), .Q(n127) );
  CLKIN2 U98 ( .A(n57), .Q(n168) );
  AOI222 U99 ( .A(n118), .B(n6), .C(n120), .D(n110), .Q(n11) );
  NOR22 U100 ( .A(B[3]), .B(n177), .Q(n115) );
  INV6 U101 ( .A(n86), .Q(n80) );
  NAND24 U102 ( .A(n117), .B(n176), .Q(n175) );
  NAND22 U103 ( .A(n163), .B(n23), .Q(n24) );
  NOR24 U104 ( .A(A[5]), .B(n170), .Q(n186) );
  XOR22 U105 ( .A(n51), .B(n52), .Q(DIFF[7]) );
  NOR24 U106 ( .A(n31), .B(n80), .Q(n179) );
  INV2 U107 ( .A(n6), .Q(n135) );
  IMUX21 U108 ( .A(n48), .B(n49), .S(n44), .Q(DIFF[8]) );
  NOR24 U109 ( .A(n146), .B(n147), .Q(n145) );
  NOR24 U110 ( .A(A[11]), .B(n37), .Q(n146) );
  NAND22 U111 ( .A(n159), .B(n158), .Q(n153) );
  INV6 U112 ( .A(n81), .Q(n181) );
  NAND43 U113 ( .A(n105), .B(n104), .C(n106), .D(n107), .Q(n91) );
  NAND34 U114 ( .A(n128), .B(n127), .C(n14), .Q(n104) );
  INV3 U115 ( .A(n108), .Q(n121) );
  NAND20 U116 ( .A(n77), .B(n82), .Q(n78) );
  INV1 U117 ( .A(B[13]), .Q(n102) );
  AOI210 U118 ( .A(n76), .B(n77), .C(n3), .Q(n75) );
  NAND24 U119 ( .A(n25), .B(n24), .Q(DIFF[10]) );
  CLKIN0 U120 ( .A(n140), .Q(n157) );
  CLKIN6 U121 ( .A(n156), .Q(n142) );
  BUF2 U122 ( .A(n36), .Q(n16) );
  INV1 U123 ( .A(n16), .Q(n19) );
  NAND42 U124 ( .A(n126), .B(n131), .C(n57), .D(n127), .Q(n143) );
  NOR24 U125 ( .A(A[10]), .B(n36), .Q(n149) );
  NOR24 U126 ( .A(A[10]), .B(n36), .Q(n140) );
  CLKIN6 U127 ( .A(n20), .Q(n21) );
  CLKIN3 U128 ( .A(n41), .Q(n17) );
  NAND28 U129 ( .A(n77), .B(n178), .Q(n26) );
  INV12 U130 ( .A(n26), .Q(n27) );
  INV3 U131 ( .A(n29), .Q(n103) );
  NAND33 U132 ( .A(n131), .B(n126), .C(n127), .Q(n169) );
  XNR22 U133 ( .A(n42), .B(n17), .Q(DIFF[9]) );
  XNR22 U134 ( .A(n103), .B(n30), .Q(DIFF[13]) );
  XNR22 U135 ( .A(n98), .B(n99), .Q(DIFF[14]) );
  AOI212 U136 ( .A(n64), .B(n58), .C(n65), .Q(n63) );
  NAND20 U137 ( .A(n57), .B(n54), .Q(n62) );
  NOR24 U138 ( .A(n148), .B(n140), .Q(n139) );
  AOI212 U139 ( .A(A[11]), .B(n37), .C(n142), .Q(n136) );
  INV1 U140 ( .A(A[7]), .Q(n171) );
  OAI2112 U141 ( .A(n55), .B(n56), .C(n57), .D(n58), .Q(n53) );
  NOR22 U142 ( .A(A[8]), .B(n35), .Q(n147) );
  NAND22 U143 ( .A(A[5]), .B(n170), .Q(n60) );
  NAND43 U144 ( .A(n108), .B(n109), .C(n110), .D(n111), .Q(n107) );
  CLKIN0 U145 ( .A(A[13]), .Q(n100) );
  NAND28 U146 ( .A(n181), .B(n27), .Q(n112) );
  XOR22 U147 ( .A(n151), .B(n150), .Q(DIFF[11]) );
  AOI212 U148 ( .A(n110), .B(n44), .C(n134), .Q(n132) );
  AOI312 U149 ( .A(n43), .B(n152), .C(n153), .D(n154), .Q(n150) );
  NAND24 U150 ( .A(n5), .B(n67), .Q(n159) );
  XNR22 U151 ( .A(n87), .B(n88), .Q(DIFF[15]) );
  NOR24 U152 ( .A(n174), .B(n175), .Q(n173) );
  NAND28 U153 ( .A(B[3]), .B(n177), .Q(n178) );
  NAND20 U154 ( .A(n86), .B(n81), .Q(n83) );
  NAND42 U155 ( .A(n105), .B(n104), .C(n8), .D(n11), .Q(n29) );
  NAND23 U156 ( .A(B[7]), .B(n171), .Q(n126) );
  OAI2112 U157 ( .A(n168), .B(n169), .C(n122), .D(n50), .Q(n160) );
  NOR20 U158 ( .A(B[12]), .B(n125), .Q(n124) );
  NOR22 U159 ( .A(A[11]), .B(n37), .Q(n123) );
  INV2 U160 ( .A(n184), .Q(n66) );
  INV3 U161 ( .A(n124), .Q(n105) );
  NAND20 U162 ( .A(n138), .B(n157), .Q(n155) );
  INV2 U163 ( .A(n85), .Q(n84) );
  AOI210 U164 ( .A(n28), .B(n39), .C(n45), .Q(n49) );
  XOR20 U165 ( .A(n28), .B(A[8]), .Q(n48) );
  NAND20 U166 ( .A(n155), .B(n156), .Q(n154) );
  NAND20 U167 ( .A(A[8]), .B(n35), .Q(n50) );
  NAND20 U168 ( .A(n46), .B(n47), .Q(n41) );
  NOR20 U169 ( .A(n184), .B(n70), .Q(n73) );
  INV2 U170 ( .A(n46), .Q(n162) );
  CLKIN3 U171 ( .A(n101), .Q(n89) );
  NAND22 U172 ( .A(n67), .B(n66), .Q(n61) );
  NOR21 U173 ( .A(n161), .B(n162), .Q(n152) );
  NOR21 U174 ( .A(n135), .B(n123), .Q(n134) );
  XOR20 U175 ( .A(n83), .B(n84), .Q(DIFF[1]) );
  XOR20 U176 ( .A(B[11]), .B(A[11]), .Q(n151) );
  XNR21 U177 ( .A(B[15]), .B(A[15]), .Q(n87) );
  XOR21 U178 ( .A(n68), .B(n69), .Q(DIFF[5]) );
  AOI210 U179 ( .A(n66), .B(n67), .C(n70), .Q(n69) );
  XOR21 U180 ( .A(n78), .B(n79), .Q(DIFF[2]) );
  IMUX20 U181 ( .A(n72), .B(n73), .S(n67), .Q(DIFF[4]) );
  XOR20 U182 ( .A(B[4]), .B(A[4]), .Q(n72) );
  AOI210 U183 ( .A(n19), .B(n40), .C(n142), .Q(n164) );
  INV3 U184 ( .A(n96), .Q(n94) );
  CLKIN0 U185 ( .A(B[14]), .Q(n97) );
  INV3 U186 ( .A(n93), .Q(n90) );
  INV0 U187 ( .A(A[14]), .Q(n95) );
  NAND20 U188 ( .A(B[9]), .B(n167), .Q(n46) );
  XNR20 U189 ( .A(B[13]), .B(A[13]), .Q(n30) );
  NOR21 U190 ( .A(B[13]), .B(n100), .Q(n96) );
  XNR20 U191 ( .A(B[14]), .B(A[14]), .Q(n98) );
  XNR21 U192 ( .A(n74), .B(n75), .Q(DIFF[3]) );
  XNR20 U193 ( .A(B[7]), .B(A[7]), .Q(n52) );
  NOR21 U194 ( .A(A[14]), .B(n97), .Q(n93) );
  XNR20 U195 ( .A(B[3]), .B(A[3]), .Q(n74) );
  INV0 U196 ( .A(A[9]), .Q(n167) );
  XOR20 U197 ( .A(B[12]), .B(A[12]), .Q(n133) );
  AOI212 U198 ( .A(n44), .B(n43), .C(n45), .Q(n42) );
  CLKIN3 U199 ( .A(n59), .Q(n70) );
  CLKIN3 U200 ( .A(n76), .Q(n79) );
  AOI312 U201 ( .A(n89), .B(n90), .C(n91), .D(n92), .Q(n88) );
  OAI222 U202 ( .A(n93), .B(n94), .C(B[14]), .D(n95), .Q(n92) );
  AOI212 U203 ( .A(n89), .B(n29), .C(n96), .Q(n99) );
  AOI222 U204 ( .A(n119), .B(n118), .C(n120), .D(n110), .Q(n106) );
endmodule


module E_alu_DW_rash_3 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324;

  AOI221 U3 ( .A(A[25]), .B(n219), .C(A[26]), .D(n220), .Q(n259) );
  NAND26 U4 ( .A(n293), .B(n294), .Q(n123) );
  NAND26 U5 ( .A(n302), .B(n303), .Q(n137) );
  NAND26 U6 ( .A(n285), .B(n284), .Q(n126) );
  AOI222 U7 ( .A(A[18]), .B(n12), .C(A[19]), .D(n218), .Q(n282) );
  NAND24 U8 ( .A(n216), .B(n217), .Q(n42) );
  NAND23 U9 ( .A(n312), .B(n313), .Q(n296) );
  AOI222 U10 ( .A(n116), .B(n55), .C(n30), .D(n54), .Q(n312) );
  AOI221 U11 ( .A(A[21]), .B(n13), .C(A[22]), .D(n218), .Q(n217) );
  BUF6 U12 ( .A(n51), .Q(n1) );
  INV3 U13 ( .A(n258), .Q(n2) );
  AOI222 U14 ( .A(A[27]), .B(n12), .C(A[28]), .D(n218), .Q(n258) );
  NAND23 U15 ( .A(n304), .B(n305), .Q(n52) );
  AOI222 U16 ( .A(n219), .B(A[18]), .C(A[19]), .D(n220), .Q(n304) );
  NAND22 U17 ( .A(n263), .B(n264), .Q(n70) );
  AOI221 U18 ( .A(n219), .B(A[17]), .C(A[18]), .D(n220), .Q(n263) );
  NAND28 U19 ( .A(n230), .B(n231), .Q(n31) );
  CLKIN3 U20 ( .A(n162), .Q(B[21]) );
  NOR24 U21 ( .A(n21), .B(n193), .Q(B[16]) );
  NAND26 U22 ( .A(n310), .B(n311), .Q(n152) );
  NOR22 U23 ( .A(n21), .B(n153), .Q(B[23]) );
  NOR22 U24 ( .A(n58), .B(n154), .Q(n153) );
  NOR23 U25 ( .A(n21), .B(n158), .Q(B[22]) );
  NOR20 U26 ( .A(n21), .B(n125), .Q(B[30]) );
  NOR23 U27 ( .A(n21), .B(n143), .Q(B[26]) );
  NOR22 U28 ( .A(n147), .B(n21), .Q(B[25]) );
  NOR23 U29 ( .A(n21), .B(n189), .Q(B[17]) );
  INV6 U30 ( .A(n2), .Q(n3) );
  NAND26 U31 ( .A(n281), .B(n282), .Q(n80) );
  NOR22 U32 ( .A(SH[4]), .B(n138), .Q(B[27]) );
  NOR20 U33 ( .A(n29), .B(n15), .Q(n229) );
  INV6 U34 ( .A(n15), .Q(n14) );
  NOR20 U35 ( .A(n29), .B(n15), .Q(n205) );
  AOI222 U36 ( .A(A[25]), .B(n10), .C(A[26]), .D(n218), .Q(n223) );
  NAND23 U37 ( .A(n116), .B(n122), .Q(n157) );
  NAND26 U38 ( .A(n259), .B(n260), .Q(n122) );
  NAND24 U39 ( .A(n166), .B(n167), .Q(n94) );
  NAND23 U40 ( .A(n116), .B(n42), .Q(n167) );
  NAND23 U41 ( .A(n276), .B(n277), .Q(n79) );
  AOI221 U42 ( .A(A[14]), .B(n10), .C(A[15]), .D(n218), .Q(n277) );
  NOR24 U43 ( .A(n21), .B(n149), .Q(B[24]) );
  NAND22 U44 ( .A(A[31]), .B(n219), .Q(n230) );
  NOR24 U45 ( .A(n168), .B(n21), .Q(B[20]) );
  NAND24 U46 ( .A(n14), .B(n135), .Q(n28) );
  NOR23 U47 ( .A(n306), .B(n307), .Q(n298) );
  NAND22 U48 ( .A(n30), .B(n152), .Q(n48) );
  NAND22 U49 ( .A(n59), .B(n152), .Q(n101) );
  NOR22 U50 ( .A(n21), .B(n185), .Q(B[18]) );
  NOR22 U51 ( .A(n186), .B(n187), .Q(n185) );
  NAND22 U52 ( .A(n130), .B(n188), .Q(n186) );
  INV3 U53 ( .A(n207), .Q(n206) );
  NAND23 U54 ( .A(n156), .B(n157), .Q(n58) );
  MUX22 U55 ( .A(n127), .B(n128), .S(n21), .Q(B[2]) );
  NAND41 U56 ( .A(n188), .B(n129), .C(n130), .D(n131), .Q(n128) );
  NAND21 U57 ( .A(n116), .B(n152), .Q(n136) );
  NAND22 U58 ( .A(n59), .B(n123), .Q(n188) );
  AOI220 U59 ( .A(A[14]), .B(n219), .C(A[15]), .D(n220), .Q(n314) );
  CLKIN6 U60 ( .A(n115), .Q(n111) );
  AOI222 U61 ( .A(n59), .B(n50), .C(n120), .D(n51), .Q(n313) );
  CLKIN6 U62 ( .A(n197), .Q(n306) );
  NAND28 U63 ( .A(n308), .B(n309), .Q(n53) );
  AOI222 U64 ( .A(A[22]), .B(n219), .C(A[23]), .D(n220), .Q(n308) );
  NAND24 U65 ( .A(n99), .B(n101), .Q(n169) );
  NAND24 U66 ( .A(n222), .B(n223), .Q(n135) );
  INV3 U67 ( .A(n195), .Q(n299) );
  NAND22 U68 ( .A(n129), .B(n131), .Q(n187) );
  INV3 U69 ( .A(n196), .Q(n307) );
  NAND24 U70 ( .A(n300), .B(n301), .Q(n195) );
  NAND22 U71 ( .A(n59), .B(n137), .Q(n301) );
  INV3 U72 ( .A(n215), .Q(n214) );
  INV3 U73 ( .A(n100), .Q(n170) );
  AOI211 U74 ( .A(n14), .B(n71), .C(n111), .Q(n183) );
  NAND33 U75 ( .A(n66), .B(n67), .C(n68), .Q(n61) );
  INV3 U76 ( .A(n113), .Q(n60) );
  AOI211 U77 ( .A(n27), .B(n28), .C(n29), .Q(n26) );
  NAND22 U78 ( .A(n233), .B(n234), .Q(n38) );
  NAND31 U79 ( .A(n44), .B(n45), .C(n43), .Q(B[8]) );
  NAND21 U80 ( .A(n99), .B(n100), .Q(n98) );
  AOI222 U81 ( .A(A[27]), .B(n219), .C(A[28]), .D(n220), .Q(n222) );
  NAND20 U82 ( .A(n41), .B(n135), .Q(n221) );
  AOI221 U83 ( .A(n116), .B(n71), .C(n59), .D(n117), .Q(n109) );
  NAND24 U84 ( .A(n261), .B(n262), .Q(n71) );
  CLKIN6 U85 ( .A(n142), .Q(n139) );
  AOI222 U86 ( .A(A[20]), .B(n11), .C(A[21]), .D(n218), .Q(n309) );
  AOI222 U87 ( .A(A[26]), .B(n219), .C(A[27]), .D(n220), .Q(n302) );
  NOR24 U88 ( .A(n169), .B(n170), .Q(n168) );
  NAND21 U89 ( .A(n48), .B(n49), .Q(n47) );
  AOI221 U90 ( .A(A[4]), .B(n10), .C(A[5]), .D(n218), .Q(n320) );
  AOI222 U91 ( .A(A[24]), .B(n11), .C(A[25]), .D(n218), .Q(n303) );
  INV3 U92 ( .A(SH[4]), .Q(n22) );
  INV3 U93 ( .A(n116), .Q(n15) );
  NAND21 U94 ( .A(n35), .B(n36), .Q(n34) );
  NAND22 U95 ( .A(n116), .B(n117), .Q(n142) );
  NAND21 U96 ( .A(n39), .B(n51), .Q(n244) );
  NAND28 U97 ( .A(n257), .B(n3), .Q(n117) );
  AOI221 U98 ( .A(A[20]), .B(n219), .C(A[21]), .D(n220), .Q(n281) );
  NAND22 U99 ( .A(n30), .B(n123), .Q(n77) );
  CLKIN6 U100 ( .A(n146), .Q(n145) );
  NAND22 U101 ( .A(n225), .B(n226), .Q(n36) );
  NOR22 U102 ( .A(n150), .B(n151), .Q(n149) );
  AOI222 U103 ( .A(A[24]), .B(n219), .C(A[25]), .D(n220), .Q(n284) );
  NOR23 U104 ( .A(n190), .B(n191), .Q(n189) );
  AOI221 U105 ( .A(n37), .B(n71), .C(n41), .D(n122), .Q(n249) );
  AOI220 U106 ( .A(n59), .B(n83), .C(n120), .D(n79), .Q(n133) );
  CLKIN3 U107 ( .A(n77), .Q(n160) );
  NAND31 U108 ( .A(n76), .B(n77), .C(n78), .Q(n75) );
  NAND22 U109 ( .A(n208), .B(n209), .Q(n207) );
  AOI221 U110 ( .A(A[19]), .B(n219), .C(A[20]), .D(n220), .Q(n233) );
  AOI220 U111 ( .A(A[15]), .B(n10), .C(A[16]), .D(n218), .Q(n264) );
  NAND33 U112 ( .A(n249), .B(n250), .C(n248), .Q(B[11]) );
  MUX26 U113 ( .A(n296), .B(n297), .S(n21), .Q(B[0]) );
  AOI222 U114 ( .A(A[23]), .B(n219), .C(A[24]), .D(n220), .Q(n216) );
  NAND20 U115 ( .A(n41), .B(n117), .Q(n202) );
  CLKIN1 U116 ( .A(n101), .Q(n97) );
  NOR20 U117 ( .A(n136), .B(n29), .Q(n247) );
  AOI222 U118 ( .A(A[23]), .B(n11), .C(A[24]), .D(n218), .Q(n260) );
  NAND20 U119 ( .A(n41), .B(n38), .Q(n90) );
  AOI220 U120 ( .A(A[19]), .B(n10), .C(A[20]), .D(n218), .Q(n262) );
  NAND21 U121 ( .A(n30), .B(n117), .Q(n156) );
  NAND22 U122 ( .A(n39), .B(n70), .Q(n204) );
  AOI221 U123 ( .A(A[17]), .B(n12), .C(A[18]), .D(n218), .Q(n234) );
  AOI221 U124 ( .A(n39), .B(n64), .C(n35), .D(n70), .Q(n248) );
  AOI220 U125 ( .A(n59), .B(n64), .C(n120), .D(n70), .Q(n119) );
  NAND22 U126 ( .A(n265), .B(n266), .Q(n64) );
  OAI222 U127 ( .A(n30), .B(n148), .C(n31), .D(n148), .Q(n147) );
  CLKIN12 U128 ( .A(n28), .Q(n148) );
  AOI221 U129 ( .A(n59), .B(n117), .C(n120), .D(n60), .Q(n184) );
  NAND21 U130 ( .A(n37), .B(n42), .Q(n215) );
  NAND42 U131 ( .A(n84), .B(n85), .C(n86), .D(n87), .Q(B[5]) );
  AOI221 U132 ( .A(A[16]), .B(n12), .C(n218), .D(A[17]), .Q(n305) );
  INV6 U133 ( .A(n323), .Q(n218) );
  NAND21 U134 ( .A(n120), .B(n31), .Q(n192) );
  AOI222 U135 ( .A(n206), .B(n29), .C(n206), .D(n125), .Q(B[14]) );
  AOI222 U136 ( .A(A[28]), .B(n219), .C(A[29]), .D(n220), .Q(n293) );
  NAND22 U137 ( .A(n120), .B(n152), .Q(n197) );
  NOR24 U138 ( .A(n61), .B(n62), .Q(n56) );
  NAND22 U139 ( .A(n39), .B(n36), .Q(n224) );
  NAND24 U140 ( .A(n298), .B(n299), .Q(n297) );
  NOR22 U141 ( .A(n194), .B(n195), .Q(n193) );
  AOI220 U142 ( .A(n37), .B(n79), .C(n41), .D(n80), .Q(n73) );
  NAND21 U143 ( .A(n37), .B(n80), .Q(n280) );
  AOI221 U144 ( .A(A[22]), .B(n13), .C(A[23]), .D(n218), .Q(n285) );
  NAND22 U145 ( .A(n30), .B(n126), .Q(n129) );
  NAND42 U146 ( .A(n23), .B(n24), .C(n34), .D(n25), .Q(B[9]) );
  AOI220 U147 ( .A(A[5]), .B(n13), .C(A[6]), .D(n218), .Q(n238) );
  CLKIN6 U148 ( .A(n76), .Q(n161) );
  NAND22 U149 ( .A(n14), .B(n126), .Q(n76) );
  NAND22 U150 ( .A(n37), .B(n122), .Q(n203) );
  AOI221 U151 ( .A(n37), .B(n126), .C(n41), .D(n123), .Q(n209) );
  AOI222 U152 ( .A(A[28]), .B(n12), .C(A[29]), .D(n218), .Q(n311) );
  AOI222 U153 ( .A(A[26]), .B(n11), .C(A[27]), .D(n218), .Q(n294) );
  NAND21 U154 ( .A(n30), .B(n135), .Q(n166) );
  AOI222 U155 ( .A(A[30]), .B(n10), .C(A[31]), .D(n218), .Q(n295) );
  AOI220 U156 ( .A(A[15]), .B(n219), .C(A[16]), .D(n220), .Q(n225) );
  AOI220 U157 ( .A(A[11]), .B(n13), .C(A[12]), .D(n218), .Q(n266) );
  NAND22 U158 ( .A(n196), .B(n197), .Q(n194) );
  AOI222 U159 ( .A(A[29]), .B(n10), .C(A[30]), .D(n218), .Q(n231) );
  AOI212 U160 ( .A(n94), .B(n22), .C(n163), .Q(n162) );
  NOR22 U161 ( .A(n164), .B(n165), .Q(n163) );
  NAND22 U162 ( .A(n30), .B(n53), .Q(n196) );
  CLKIN1 U163 ( .A(n177), .Q(n176) );
  CLKIN1 U164 ( .A(n178), .Q(n175) );
  INV1 U165 ( .A(SH[2]), .Q(n19) );
  CLKIN2 U166 ( .A(n104), .Q(n103) );
  NAND22 U167 ( .A(n120), .B(n144), .Q(n131) );
  CLKIN3 U168 ( .A(n275), .Q(n39) );
  NAND20 U169 ( .A(n30), .B(n31), .Q(n27) );
  NOR20 U170 ( .A(n113), .B(n114), .Q(n112) );
  AOI210 U171 ( .A(n120), .B(n31), .C(n179), .Q(n173) );
  NAND22 U172 ( .A(n37), .B(n36), .Q(n89) );
  NAND22 U173 ( .A(n180), .B(n178), .Q(n190) );
  CLKIN2 U174 ( .A(n224), .Q(n212) );
  INV2 U175 ( .A(n204), .Q(n200) );
  INV3 U176 ( .A(n232), .Q(n220) );
  NAND20 U177 ( .A(SH[1]), .B(n16), .Q(n232) );
  NAND20 U178 ( .A(SH[3]), .B(SH[2]), .Q(n114) );
  NAND20 U179 ( .A(SH[3]), .B(n19), .Q(n318) );
  NAND20 U180 ( .A(n16), .B(n18), .Q(n323) );
  NAND20 U181 ( .A(SH[2]), .B(n20), .Q(n256) );
  INV3 U182 ( .A(n17), .Q(n16) );
  CLKIN3 U183 ( .A(n49), .Q(n151) );
  CLKIN3 U184 ( .A(n180), .Q(n179) );
  AOI210 U185 ( .A(n292), .B(n146), .C(n29), .Q(n287) );
  NAND20 U186 ( .A(n30), .B(n144), .Q(n292) );
  NOR20 U187 ( .A(n154), .B(n58), .Q(n57) );
  INV2 U188 ( .A(n26), .Q(n25) );
  NAND20 U189 ( .A(n39), .B(n32), .Q(n85) );
  NAND20 U190 ( .A(n35), .B(n40), .Q(n84) );
  MUX22 U191 ( .A(n171), .B(n172), .S(n21), .Q(B[1]) );
  MUX22 U192 ( .A(n107), .B(n108), .S(n21), .Q(B[3]) );
  NAND20 U193 ( .A(n37), .B(n38), .Q(n24) );
  AOI220 U194 ( .A(A[13]), .B(n13), .C(A[14]), .D(n218), .Q(n226) );
  AOI220 U195 ( .A(A[13]), .B(n219), .C(A[14]), .D(n220), .Q(n265) );
  CLKIN3 U196 ( .A(n155), .Q(n154) );
  NAND21 U197 ( .A(n59), .B(n60), .Q(n155) );
  NOR20 U198 ( .A(n113), .B(n256), .Q(n255) );
  NAND20 U199 ( .A(n14), .B(n60), .Q(n121) );
  NOR20 U200 ( .A(SH[1]), .B(n16), .Q(n8) );
  NAND20 U201 ( .A(n35), .B(n79), .Q(n271) );
  NAND20 U202 ( .A(n35), .B(n50), .Q(n104) );
  AOI220 U203 ( .A(A[7]), .B(n13), .C(A[8]), .D(n218), .Q(n254) );
  AOI220 U204 ( .A(A[5]), .B(n219), .C(A[6]), .D(n220), .Q(n251) );
  AOI220 U205 ( .A(n14), .B(n65), .C(n30), .D(n69), .Q(n118) );
  CLKIN3 U206 ( .A(SH[1]), .Q(n18) );
  CLKIN1 U207 ( .A(SH[3]), .Q(n20) );
  NAND22 U208 ( .A(n30), .B(n137), .Q(n100) );
  NAND22 U209 ( .A(n116), .B(n137), .Q(n49) );
  NAND22 U210 ( .A(n30), .B(n122), .Q(n115) );
  NAND21 U211 ( .A(n116), .B(n144), .Q(n125) );
  NAND22 U212 ( .A(n30), .B(n42), .Q(n180) );
  AOI221 U213 ( .A(n56), .B(n29), .C(n57), .D(n56), .Q(B[7]) );
  NAND22 U214 ( .A(n116), .B(n53), .Q(n99) );
  NAND22 U215 ( .A(n30), .B(n60), .Q(n141) );
  INV3 U216 ( .A(n9), .Q(n10) );
  NOR21 U217 ( .A(n111), .B(n112), .Q(n110) );
  NOR21 U218 ( .A(n175), .B(n176), .Q(n174) );
  INV3 U219 ( .A(n9), .Q(n12) );
  INV3 U220 ( .A(n9), .Q(n11) );
  NAND22 U221 ( .A(n239), .B(n240), .Q(B[12]) );
  INV3 U222 ( .A(n247), .Q(n239) );
  NOR21 U223 ( .A(n241), .B(n242), .Q(n240) );
  NAND22 U224 ( .A(n267), .B(n268), .Q(B[10]) );
  NOR21 U225 ( .A(n269), .B(n270), .Q(n268) );
  INV3 U226 ( .A(n287), .Q(n267) );
  NAND22 U227 ( .A(n271), .B(n272), .Q(n270) );
  INV3 U228 ( .A(n9), .Q(n13) );
  INV3 U229 ( .A(n114), .Q(n120) );
  NAND22 U230 ( .A(n273), .B(n274), .Q(n83) );
  AOI220 U231 ( .A(A[21]), .B(n219), .C(A[22]), .D(n220), .Q(n261) );
  NAND22 U232 ( .A(n315), .B(n314), .Q(n51) );
  AOI220 U233 ( .A(n39), .B(n40), .C(n41), .D(n42), .Q(n23) );
  AOI220 U234 ( .A(A[16]), .B(n219), .C(A[17]), .D(n220), .Q(n276) );
  INV3 U235 ( .A(n88), .Q(n87) );
  NAND22 U236 ( .A(A[31]), .B(n11), .Q(n113) );
  NAND22 U237 ( .A(n235), .B(n236), .Q(n40) );
  AOI221 U238 ( .A(n59), .B(n40), .C(n120), .D(n36), .Q(n182) );
  NAND22 U239 ( .A(n95), .B(n96), .Q(B[4]) );
  AOI2110 U240 ( .A(n37), .B(n1), .C(n102), .D(n103), .Q(n95) );
  NAND22 U241 ( .A(n105), .B(n106), .Q(n102) );
  NAND22 U242 ( .A(n37), .B(n70), .Q(n67) );
  NAND22 U243 ( .A(n39), .B(n69), .Q(n68) );
  NAND22 U244 ( .A(n41), .B(n71), .Q(n66) );
  AOI221 U245 ( .A(n39), .B(n79), .C(n35), .D(n80), .Q(n208) );
  NOR21 U246 ( .A(SH[3]), .B(SH[2]), .Q(n116) );
  AOI220 U247 ( .A(n39), .B(n50), .C(n35), .D(n1), .Q(n44) );
  AOI220 U248 ( .A(n37), .B(n52), .C(n53), .D(n41), .Q(n43) );
  NAND22 U249 ( .A(n46), .B(n47), .Q(n45) );
  NAND22 U250 ( .A(n59), .B(n135), .Q(n178) );
  NAND22 U251 ( .A(n14), .B(n38), .Q(n177) );
  NAND31 U252 ( .A(n73), .B(n74), .C(n72), .Q(B[6]) );
  AOI220 U253 ( .A(n39), .B(n82), .C(n35), .D(n83), .Q(n72) );
  NAND22 U254 ( .A(n46), .B(n75), .Q(n74) );
  NAND22 U255 ( .A(n14), .B(n123), .Q(n146) );
  NOR21 U256 ( .A(n21), .B(n136), .Q(B[28]) );
  NAND22 U257 ( .A(n59), .B(n144), .Q(n78) );
  NAND22 U258 ( .A(n116), .B(n52), .Q(n300) );
  NAND22 U259 ( .A(n116), .B(n80), .Q(n130) );
  INV3 U260 ( .A(n8), .Q(n9) );
  NAND21 U261 ( .A(n39), .B(n83), .Q(n272) );
  NAND22 U262 ( .A(n245), .B(n246), .Q(n241) );
  NAND20 U263 ( .A(n41), .B(n137), .Q(n245) );
  NAND20 U264 ( .A(n37), .B(n53), .Q(n246) );
  NAND22 U265 ( .A(n279), .B(n280), .Q(n269) );
  NAND20 U266 ( .A(n41), .B(n126), .Q(n279) );
  NAND22 U267 ( .A(n202), .B(n203), .Q(n201) );
  NAND22 U268 ( .A(n243), .B(n244), .Q(n242) );
  NAND20 U269 ( .A(n35), .B(n52), .Q(n243) );
  NAND22 U270 ( .A(n39), .B(n54), .Q(n106) );
  NAND22 U271 ( .A(n89), .B(n90), .Q(n88) );
  NAND20 U272 ( .A(n41), .B(n52), .Q(n105) );
  NOR31 U273 ( .A(n159), .B(n160), .C(n161), .Q(n158) );
  NAND22 U274 ( .A(n192), .B(n177), .Q(n191) );
  NOR21 U275 ( .A(n21), .B(n121), .Q(B[31]) );
  NAND22 U276 ( .A(n46), .B(n91), .Q(n86) );
  NAND22 U277 ( .A(n92), .B(n93), .Q(n91) );
  NAND21 U278 ( .A(n59), .B(n31), .Q(n93) );
  INV3 U279 ( .A(n94), .Q(n92) );
  NAND22 U280 ( .A(n198), .B(n199), .Q(B[15]) );
  AOI220 U281 ( .A(n35), .B(n71), .C(n205), .D(n60), .Q(n198) );
  NOR21 U282 ( .A(n200), .B(n201), .Q(n199) );
  NAND22 U283 ( .A(n210), .B(n211), .Q(B[13]) );
  AOI220 U284 ( .A(n35), .B(n38), .C(n229), .D(n31), .Q(n210) );
  NOR31 U285 ( .A(n212), .B(n213), .C(n214), .Q(n211) );
  NOR21 U286 ( .A(n21), .B(n134), .Q(B[29]) );
  NAND20 U287 ( .A(n14), .B(n31), .Q(n134) );
  NOR21 U288 ( .A(n139), .B(n140), .Q(n138) );
  INV3 U289 ( .A(n141), .Q(n140) );
  INV3 U290 ( .A(n221), .Q(n213) );
  CLKIN3 U291 ( .A(n63), .Q(n62) );
  NAND22 U292 ( .A(n35), .B(n64), .Q(n63) );
  NAND22 U293 ( .A(n132), .B(n133), .Q(n127) );
  NAND22 U294 ( .A(n181), .B(n182), .Q(n171) );
  NAND22 U295 ( .A(n173), .B(n174), .Q(n172) );
  NAND22 U296 ( .A(n118), .B(n119), .Q(n107) );
  NAND22 U297 ( .A(n109), .B(n110), .Q(n108) );
  INV3 U298 ( .A(n21), .Q(n29) );
  INV3 U299 ( .A(n256), .Q(n30) );
  NAND22 U300 ( .A(n237), .B(n238), .Q(n32) );
  INV3 U301 ( .A(n324), .Q(n219) );
  NAND22 U302 ( .A(SH[1]), .B(n17), .Q(n324) );
  NAND22 U303 ( .A(n316), .B(n317), .Q(n50) );
  NAND22 U304 ( .A(n319), .B(n320), .Q(n54) );
  AOI220 U305 ( .A(A[6]), .B(n219), .C(A[7]), .D(n220), .Q(n319) );
  NAND22 U306 ( .A(n116), .B(n22), .Q(n275) );
  AOI221 U307 ( .A(n116), .B(n33), .C(n30), .D(n32), .Q(n181) );
  NAND22 U308 ( .A(n227), .B(n228), .Q(n33) );
  NAND22 U309 ( .A(n251), .B(n252), .Q(n65) );
  AOI221 U310 ( .A(n14), .B(n81), .C(n30), .D(n82), .Q(n132) );
  NAND22 U311 ( .A(n288), .B(n289), .Q(n81) );
  AOI220 U312 ( .A(A[4]), .B(n219), .C(A[5]), .D(n220), .Q(n288) );
  NAND22 U313 ( .A(n321), .B(n322), .Q(n55) );
  NAND22 U314 ( .A(n253), .B(n254), .Q(n69) );
  NAND22 U315 ( .A(n290), .B(n291), .Q(n82) );
  AOI220 U316 ( .A(A[6]), .B(n12), .C(A[7]), .D(n218), .Q(n291) );
  NAND22 U317 ( .A(n59), .B(n22), .Q(n165) );
  INV3 U318 ( .A(n22), .Q(n21) );
  INV3 U319 ( .A(n318), .Q(n59) );
  INV3 U320 ( .A(n278), .Q(n35) );
  NAND22 U321 ( .A(n30), .B(n22), .Q(n278) );
  INV3 U322 ( .A(n283), .Q(n37) );
  NAND22 U323 ( .A(n59), .B(n22), .Q(n283) );
  INV3 U324 ( .A(n286), .Q(n41) );
  NAND22 U325 ( .A(n120), .B(n22), .Q(n286) );
  INV3 U326 ( .A(SH[0]), .Q(n17) );
  CLKIN6 U327 ( .A(n295), .Q(n144) );
  OAI222 U328 ( .A(n183), .B(n21), .C(n184), .D(n21), .Q(B[19]) );
  OAI222 U329 ( .A(n30), .B(n145), .C(n144), .D(n145), .Q(n143) );
  AOI220 U330 ( .A(A[7]), .B(n219), .C(A[8]), .D(n220), .Q(n237) );
  AOI220 U331 ( .A(A[8]), .B(n219), .C(A[9]), .D(n220), .Q(n290) );
  AOI220 U332 ( .A(A[8]), .B(n11), .C(A[9]), .D(n218), .Q(n317) );
  AOI220 U333 ( .A(A[1]), .B(n13), .C(A[2]), .D(n218), .Q(n228) );
  AOI220 U334 ( .A(A[9]), .B(n13), .C(A[10]), .D(n218), .Q(n236) );
  AOI220 U335 ( .A(A[10]), .B(n13), .C(A[11]), .D(n218), .Q(n274) );
  AOI220 U336 ( .A(A[10]), .B(n219), .C(A[11]), .D(n220), .Q(n316) );
  AOI220 U337 ( .A(A[9]), .B(n219), .C(A[10]), .D(n220), .Q(n253) );
  AOI220 U338 ( .A(n11), .B(A[0]), .C(A[1]), .D(n218), .Q(n322) );
  AOI220 U339 ( .A(A[11]), .B(n219), .C(A[12]), .D(n220), .Q(n235) );
  AOI220 U340 ( .A(A[12]), .B(n219), .C(A[13]), .D(n220), .Q(n273) );
  AOI220 U341 ( .A(A[12]), .B(n12), .C(A[13]), .D(n218), .Q(n315) );
  AOI220 U342 ( .A(A[2]), .B(n12), .C(A[3]), .D(n218), .Q(n289) );
  AOI220 U343 ( .A(A[3]), .B(n219), .C(A[4]), .D(n220), .Q(n227) );
  AOI220 U344 ( .A(A[2]), .B(n219), .C(A[3]), .D(n220), .Q(n321) );
  AOI220 U345 ( .A(A[3]), .B(n13), .C(A[4]), .D(n218), .Q(n252) );
  OAI212 U346 ( .A(n97), .B(n98), .C(n46), .Q(n96) );
  CLKIN3 U347 ( .A(n48), .Q(n150) );
  CLKIN3 U348 ( .A(n78), .Q(n159) );
  CLKIN3 U349 ( .A(n31), .Q(n164) );
  OAI212 U350 ( .A(n139), .B(n255), .C(n46), .Q(n250) );
  CLKIN3 U351 ( .A(n29), .Q(n46) );
  AOI222 U352 ( .A(A[29]), .B(n219), .C(A[30]), .D(n220), .Q(n257) );
  AOI222 U353 ( .A(A[30]), .B(n219), .C(A[31]), .D(n220), .Q(n310) );
endmodule


module E_alu_DW01_add_23 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111;

  NOR22 U2 ( .A(A[6]), .B(B[6]), .Q(n1) );
  NOR23 U3 ( .A(A[6]), .B(B[6]), .Q(n45) );
  CLKIN1 U4 ( .A(n38), .Q(n87) );
  INV2 U5 ( .A(n1), .Q(n61) );
  INV8 U6 ( .A(n13), .Q(n14) );
  INV6 U7 ( .A(n4), .Q(n96) );
  NAND28 U8 ( .A(n11), .B(n8), .Q(n4) );
  NAND24 U9 ( .A(n17), .B(A[0]), .Q(n104) );
  NOR24 U10 ( .A(A[1]), .B(B[1]), .Q(n56) );
  XOR22 U11 ( .A(n64), .B(n65), .Q(SUM[7]) );
  NOR22 U12 ( .A(n66), .B(n67), .Q(n65) );
  INV4 U13 ( .A(A[7]), .Q(n16) );
  NOR23 U14 ( .A(n29), .B(n28), .Q(n27) );
  CLKIN3 U15 ( .A(n61), .Q(n2) );
  INV6 U16 ( .A(n2), .Q(n3) );
  NAND42 U17 ( .A(n4), .B(n61), .C(n7), .D(n62), .Q(n24) );
  XOR22 U18 ( .A(n78), .B(n79), .Q(SUM[6]) );
  NOR20 U19 ( .A(n108), .B(n56), .Q(n109) );
  NAND20 U20 ( .A(A[4]), .B(n12), .Q(n81) );
  INV8 U21 ( .A(A[4]), .Q(n8) );
  NOR22 U22 ( .A(A[4]), .B(n12), .Q(n82) );
  INV10 U23 ( .A(n11), .Q(n12) );
  NOR22 U24 ( .A(n36), .B(n96), .Q(n51) );
  NAND22 U25 ( .A(n12), .B(A[4]), .Q(n97) );
  NAND22 U26 ( .A(B[1]), .B(A[1]), .Q(n63) );
  NOR21 U27 ( .A(A[5]), .B(B[5]), .Q(n38) );
  NOR22 U28 ( .A(n23), .B(n18), .Q(n91) );
  NAND21 U29 ( .A(n87), .B(n35), .Q(n83) );
  NOR23 U30 ( .A(n47), .B(n50), .Q(n49) );
  AOI2111 U31 ( .A(n60), .B(n20), .C(n47), .D(n63), .Q(n62) );
  INV6 U32 ( .A(n15), .Q(n47) );
  NAND23 U33 ( .A(n51), .B(n52), .Q(n39) );
  INV4 U34 ( .A(n37), .Q(n31) );
  CLKIN6 U35 ( .A(n22), .Q(n21) );
  INV3 U36 ( .A(n53), .Q(n94) );
  INV3 U37 ( .A(n94), .Q(n5) );
  NAND22 U38 ( .A(n95), .B(n19), .Q(n77) );
  INV10 U39 ( .A(B[4]), .Q(n11) );
  NAND22 U40 ( .A(n48), .B(n77), .Q(n6) );
  NOR21 U41 ( .A(n44), .B(n82), .Q(n74) );
  NOR22 U42 ( .A(n47), .B(n48), .Q(n46) );
  NOR22 U43 ( .A(A[7]), .B(n21), .Q(n30) );
  INV6 U44 ( .A(n20), .Q(n19) );
  INV6 U45 ( .A(n18), .Q(n17) );
  INV3 U46 ( .A(n6), .Q(n70) );
  AOI211 U47 ( .A(n74), .B(n80), .C(n69), .Q(n79) );
  NAND22 U48 ( .A(A[2]), .B(n19), .Q(n50) );
  INV3 U49 ( .A(A[0]), .Q(n23) );
  CLKIN3 U50 ( .A(B[0]), .Q(n18) );
  INV6 U51 ( .A(n9), .Q(n10) );
  INV3 U52 ( .A(n49), .Q(n40) );
  CLKIN3 U53 ( .A(B[7]), .Q(n22) );
  INV12 U54 ( .A(B[2]), .Q(n20) );
  NOR21 U55 ( .A(n19), .B(A[2]), .Q(n76) );
  INV2 U56 ( .A(n103), .Q(n102) );
  NOR24 U57 ( .A(n53), .B(n44), .Q(n9) );
  NAND20 U58 ( .A(n19), .B(A[2]), .Q(n103) );
  INV2 U59 ( .A(n10), .Q(n7) );
  NAND22 U60 ( .A(n46), .B(n4), .Q(n41) );
  NOR20 U61 ( .A(n96), .B(n86), .Q(n89) );
  NOR24 U62 ( .A(n10), .B(n56), .Q(n59) );
  NOR41 U63 ( .A(n104), .B(n76), .C(n56), .D(n5), .Q(n75) );
  NAND28 U64 ( .A(n27), .B(n14), .Q(SUM[8]) );
  AOI212 U65 ( .A(n60), .B(n20), .C(n47), .Q(n57) );
  NAND21 U66 ( .A(n60), .B(n20), .Q(n93) );
  NOR23 U67 ( .A(n36), .B(n96), .Q(n58) );
  NAND43 U68 ( .A(n91), .B(n57), .C(n59), .D(n58), .Q(n25) );
  NAND22 U69 ( .A(B[6]), .B(A[6]), .Q(n55) );
  AOI2111 U70 ( .A(n60), .B(n20), .C(n56), .D(n5), .Q(n92) );
  NAND34 U71 ( .A(n24), .B(n25), .C(n26), .Q(n13) );
  NOR22 U72 ( .A(B[6]), .B(A[6]), .Q(n36) );
  OAI312 U73 ( .A(n97), .B(n30), .C(n31), .D(n32), .Q(n29) );
  NOR21 U74 ( .A(n30), .B(n1), .Q(n33) );
  NOR24 U75 ( .A(A[5]), .B(B[5]), .Q(n44) );
  NOR22 U76 ( .A(n38), .B(n45), .Q(n37) );
  NAND21 U77 ( .A(n68), .B(n55), .Q(n67) );
  NAND43 U78 ( .A(n77), .B(n48), .C(n71), .D(n90), .Q(n80) );
  NOR22 U79 ( .A(n45), .B(n44), .Q(n43) );
  NAND21 U80 ( .A(B[5]), .B(A[5]), .Q(n35) );
  AOI312 U81 ( .A(n70), .B(n71), .C(n72), .D(n73), .Q(n66) );
  NAND22 U82 ( .A(B[3]), .B(A[3]), .Q(n48) );
  NAND22 U83 ( .A(n69), .B(n3), .Q(n68) );
  NAND21 U84 ( .A(n74), .B(n3), .Q(n73) );
  INV2 U85 ( .A(n75), .Q(n72) );
  NOR20 U86 ( .A(n104), .B(n56), .Q(n107) );
  NAND22 U87 ( .A(n63), .B(n104), .Q(n101) );
  NOR21 U88 ( .A(n53), .B(n44), .Q(n52) );
  NOR24 U89 ( .A(A[3]), .B(B[3]), .Q(n53) );
  NOR21 U90 ( .A(n53), .B(n60), .Q(n95) );
  AOI210 U91 ( .A(n60), .B(n20), .C(n56), .Q(n100) );
  INV2 U92 ( .A(A[2]), .Q(n60) );
  NAND42 U93 ( .A(A[1]), .B(B[1]), .C(n93), .D(n94), .Q(n71) );
  AOI212 U94 ( .A(n85), .B(n80), .C(n86), .Q(n84) );
  IMUX21 U95 ( .A(n88), .B(n89), .S(n80), .Q(SUM[4]) );
  OAI211 U96 ( .A(n44), .B(n81), .C(n35), .Q(n69) );
  NAND22 U97 ( .A(n22), .B(n16), .Q(n15) );
  INV1 U98 ( .A(n63), .Q(n108) );
  NOR20 U99 ( .A(n17), .B(n23), .Q(n111) );
  XNR21 U100 ( .A(n104), .B(n109), .Q(SUM[1]) );
  INV3 U101 ( .A(n111), .Q(n110) );
  INV3 U102 ( .A(n82), .Q(n85) );
  XOR21 U103 ( .A(n83), .B(n84), .Q(SUM[5]) );
  XOR21 U104 ( .A(n105), .B(n106), .Q(SUM[2]) );
  NOR21 U105 ( .A(n107), .B(n108), .Q(n106) );
  NAND22 U106 ( .A(n91), .B(n92), .Q(n90) );
  INV3 U107 ( .A(n54), .Q(n26) );
  XNR20 U108 ( .A(n12), .B(A[4]), .Q(n88) );
  AOI211 U109 ( .A(n100), .B(n101), .C(n102), .Q(n99) );
  NAND20 U110 ( .A(n3), .B(n55), .Q(n78) );
  NAND22 U111 ( .A(n33), .B(n34), .Q(n32) );
  INV3 U112 ( .A(n43), .Q(n42) );
  XOR21 U113 ( .A(n98), .B(n99), .Q(SUM[3]) );
  XNR20 U114 ( .A(B[3]), .B(A[3]), .Q(n98) );
  OAI210 U115 ( .A(n19), .B(A[2]), .C(n103), .Q(n105) );
  XNR20 U116 ( .A(n21), .B(A[7]), .Q(n64) );
  CLKIN3 U117 ( .A(n35), .Q(n34) );
  OAI222 U118 ( .A(n39), .B(n40), .C(n41), .D(n42), .Q(n28) );
  OAI222 U119 ( .A(n55), .B(n30), .C(n16), .D(n22), .Q(n54) );
  CLKIN3 U120 ( .A(n97), .Q(n86) );
  OAI212 U121 ( .A(A[0]), .B(n18), .C(n110), .Q(SUM[0]) );
endmodule


module E_alu_DW01_sub_10 ( A, B, CI, DIFF, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325;

  INV8 U3 ( .A(n110), .Q(n75) );
  CLKIN3 U4 ( .A(n321), .Q(n108) );
  INV8 U5 ( .A(B[11]), .Q(n59) );
  INV2 U6 ( .A(n303), .Q(n316) );
  NAND22 U7 ( .A(n177), .B(n176), .Q(n169) );
  INV10 U8 ( .A(n40), .Q(n41) );
  NAND33 U9 ( .A(n150), .B(n151), .C(n152), .Q(n48) );
  NOR22 U10 ( .A(n222), .B(n223), .Q(n212) );
  CLKIN6 U11 ( .A(B[3]), .Q(n309) );
  CLKIN1 U12 ( .A(n159), .Q(n175) );
  NAND20 U13 ( .A(n205), .B(n206), .Q(n282) );
  NAND23 U14 ( .A(n246), .B(n17), .Q(n56) );
  NAND24 U15 ( .A(B[13]), .B(n252), .Q(n163) );
  NOR24 U16 ( .A(A[3]), .B(n309), .Q(n215) );
  INV6 U17 ( .A(n215), .Q(n313) );
  INV2 U18 ( .A(n146), .Q(n1) );
  INV1 U19 ( .A(B[15]), .Q(n146) );
  INV12 U20 ( .A(n157), .Q(n153) );
  NAND20 U21 ( .A(n159), .B(n154), .Q(n189) );
  CLKIN12 U22 ( .A(B[8]), .Q(n58) );
  NAND20 U23 ( .A(n22), .B(n159), .Q(n158) );
  INV12 U24 ( .A(A[11]), .Q(n63) );
  NAND34 U25 ( .A(n20), .B(n164), .C(n163), .Q(n2) );
  NAND32 U26 ( .A(n20), .B(n164), .C(n163), .Q(n139) );
  NAND24 U27 ( .A(n73), .B(n41), .Q(n86) );
  NAND23 U28 ( .A(A[7]), .B(n304), .Q(n79) );
  AOI210 U29 ( .A(n76), .B(n77), .C(n78), .Q(n67) );
  INV10 U30 ( .A(B[6]), .Q(n298) );
  CLKIN3 U31 ( .A(B[10]), .Q(n322) );
  CLKIN3 U32 ( .A(A[14]), .Q(n226) );
  INV1 U33 ( .A(A[6]), .Q(n112) );
  NAND28 U34 ( .A(n145), .B(n76), .Q(n44) );
  NAND26 U35 ( .A(n242), .B(n243), .Q(n77) );
  CLKIN12 U36 ( .A(B[13]), .Q(n251) );
  NAND23 U37 ( .A(n322), .B(A[10]), .Q(n263) );
  NOR22 U38 ( .A(n178), .B(n179), .Q(n177) );
  INV6 U39 ( .A(A[10]), .Q(n323) );
  NAND22 U40 ( .A(n95), .B(n96), .Q(n38) );
  INV2 U41 ( .A(A[13]), .Q(n252) );
  NAND24 U42 ( .A(A[13]), .B(n251), .Q(n157) );
  CLKIN6 U43 ( .A(n57), .Q(n325) );
  NOR22 U44 ( .A(n103), .B(n100), .Q(n102) );
  INV3 U45 ( .A(n319), .Q(n107) );
  NOR23 U46 ( .A(n319), .B(n320), .Q(n318) );
  NOR22 U47 ( .A(A[4]), .B(n115), .Q(n319) );
  NAND24 U48 ( .A(n299), .B(n300), .Q(n244) );
  INV3 U49 ( .A(n301), .Q(n300) );
  NAND24 U50 ( .A(n141), .B(n142), .Q(n140) );
  INV3 U51 ( .A(n207), .Q(n171) );
  NOR21 U52 ( .A(n237), .B(n238), .Q(n236) );
  NOR22 U53 ( .A(n301), .B(n321), .Q(n317) );
  INV6 U54 ( .A(n22), .Q(n160) );
  NOR22 U55 ( .A(B[4]), .B(n119), .Q(n205) );
  INV12 U56 ( .A(B[0]), .Q(n57) );
  NAND26 U57 ( .A(n124), .B(n313), .Q(n110) );
  NOR23 U58 ( .A(n226), .B(B[14]), .Q(n55) );
  NOR23 U59 ( .A(A[5]), .B(n116), .Q(n321) );
  INV3 U60 ( .A(B[4]), .Q(n115) );
  NOR32 U61 ( .A(n161), .B(n162), .C(n24), .Q(n136) );
  NAND22 U62 ( .A(n107), .B(n108), .Q(n98) );
  NOR22 U63 ( .A(n171), .B(n195), .Q(n193) );
  NAND23 U64 ( .A(B[6]), .B(n112), .Q(n96) );
  INV2 U65 ( .A(B[9]), .Q(n6) );
  NOR22 U66 ( .A(A[0]), .B(n57), .Q(n237) );
  NOR22 U67 ( .A(n74), .B(n109), .Q(n105) );
  NOR22 U68 ( .A(n74), .B(n234), .Q(n268) );
  NAND24 U69 ( .A(n235), .B(n123), .Q(n222) );
  NOR21 U70 ( .A(n325), .B(n219), .Q(n135) );
  NAND20 U71 ( .A(A[4]), .B(n115), .Q(n99) );
  INV6 U72 ( .A(n36), .Q(n37) );
  INV6 U73 ( .A(A[8]), .Q(n66) );
  NOR23 U74 ( .A(n55), .B(n153), .Q(n151) );
  INV0 U75 ( .A(n16), .Q(n3) );
  INV6 U76 ( .A(B[8]), .Q(n16) );
  INV6 U77 ( .A(n79), .Q(n142) );
  NOR23 U78 ( .A(n203), .B(n204), .Q(n198) );
  INV3 U79 ( .A(n205), .Q(n204) );
  INV2 U80 ( .A(A[5]), .Q(n302) );
  NOR22 U81 ( .A(n201), .B(n202), .Q(n200) );
  CLKIN12 U82 ( .A(n244), .Q(n199) );
  NAND23 U83 ( .A(B[14]), .B(n226), .Q(n159) );
  CLKIN4 U84 ( .A(B[2]), .Q(n310) );
  NOR22 U85 ( .A(n13), .B(n303), .Q(n271) );
  NOR24 U86 ( .A(n229), .B(n230), .Q(n228) );
  OAI211 U87 ( .A(n179), .B(n196), .C(n5), .Q(n195) );
  NOR20 U88 ( .A(n179), .B(n201), .Q(n241) );
  CLKIN6 U89 ( .A(n46), .Q(n47) );
  INV6 U90 ( .A(A[1]), .Q(n133) );
  NOR24 U91 ( .A(A[1]), .B(n315), .Q(n218) );
  OAI212 U92 ( .A(A[3]), .B(n309), .C(A[1]), .Q(n312) );
  NAND23 U93 ( .A(n184), .B(n142), .Q(n207) );
  BUF2 U94 ( .A(n263), .Q(n10) );
  INV3 U95 ( .A(n32), .Q(n33) );
  XNR21 U96 ( .A(n125), .B(n122), .Q(DIFF[2]) );
  INV6 U97 ( .A(B[14]), .Q(n166) );
  INV6 U98 ( .A(A[15]), .Q(n23) );
  INV3 U99 ( .A(n26), .Q(n216) );
  INV3 U100 ( .A(n199), .Q(n27) );
  NAND22 U101 ( .A(n69), .B(n172), .Q(n178) );
  NAND22 U102 ( .A(A[3]), .B(n309), .Q(n71) );
  INV3 U103 ( .A(n243), .Q(n266) );
  INV8 U104 ( .A(n63), .Q(n62) );
  NAND31 U105 ( .A(n69), .B(n288), .C(n43), .Q(n287) );
  NOR22 U106 ( .A(n181), .B(n180), .Q(n168) );
  NOR21 U107 ( .A(n182), .B(n183), .Q(n181) );
  NAND24 U108 ( .A(n29), .B(n30), .Q(n28) );
  CLKIN6 U109 ( .A(n222), .Q(n29) );
  INV6 U110 ( .A(n156), .Q(n259) );
  CLKIN3 U111 ( .A(n145), .Q(n24) );
  NOR24 U112 ( .A(n264), .B(n13), .Q(n261) );
  NOR24 U113 ( .A(n50), .B(n63), .Q(n156) );
  NOR24 U114 ( .A(n62), .B(n59), .Q(n250) );
  INV3 U115 ( .A(n235), .Q(n126) );
  NAND24 U116 ( .A(B[1]), .B(n133), .Q(n235) );
  INV3 U117 ( .A(n99), .Q(n97) );
  XOR20 U118 ( .A(n1), .B(A[15]), .Q(n4) );
  INV12 U119 ( .A(n162), .Q(n141) );
  CLKIN3 U120 ( .A(n72), .Q(n11) );
  NOR21 U121 ( .A(n283), .B(n284), .Q(n280) );
  NOR23 U122 ( .A(n276), .B(n277), .Q(n275) );
  NAND26 U123 ( .A(n9), .B(n39), .Q(n94) );
  CLKIN8 U124 ( .A(n25), .Q(n60) );
  BUF6 U125 ( .A(B[11]), .Q(n50) );
  BUF2 U126 ( .A(n197), .Q(n5) );
  NAND22 U127 ( .A(A[12]), .B(n25), .Q(n197) );
  INV6 U128 ( .A(n11), .Q(n12) );
  INV2 U129 ( .A(A[0]), .Q(n219) );
  AOI310 U130 ( .A(n235), .B(n123), .C(n273), .D(n75), .Q(n269) );
  NOR24 U131 ( .A(A[6]), .B(n298), .Q(n301) );
  NAND26 U132 ( .A(n260), .B(n47), .Q(n152) );
  CLKIN2 U133 ( .A(n237), .Q(n224) );
  IMUX21 U134 ( .A(n117), .B(n118), .S(n9), .Q(DIFF[4]) );
  INV3 U135 ( .A(n245), .Q(n264) );
  NAND22 U136 ( .A(n6), .B(n7), .Q(n8) );
  NAND24 U137 ( .A(n8), .B(n263), .Q(n262) );
  INV2 U138 ( .A(n61), .Q(n7) );
  CLKIN3 U139 ( .A(A[12]), .Q(n249) );
  INV3 U140 ( .A(n210), .Q(n185) );
  CLKIN3 U141 ( .A(B[5]), .Q(n116) );
  NAND34 U142 ( .A(n77), .B(n141), .C(n45), .Q(n144) );
  BUF2 U143 ( .A(n217), .Q(n26) );
  NAND22 U144 ( .A(n69), .B(n70), .Q(n68) );
  NAND32 U145 ( .A(n73), .B(n28), .C(n33), .Q(n70) );
  NAND28 U146 ( .A(n73), .B(n41), .Q(n9) );
  NOR24 U147 ( .A(n311), .B(n312), .Q(n74) );
  NOR21 U148 ( .A(B[5]), .B(n302), .Q(n299) );
  NAND28 U149 ( .A(B[10]), .B(n323), .Q(n245) );
  INV12 U150 ( .A(B[12]), .Q(n25) );
  INV3 U151 ( .A(n18), .Q(n19) );
  NOR21 U152 ( .A(n97), .B(n11), .Q(n106) );
  AOI222 U153 ( .A(n209), .B(n208), .C(n14), .D(n187), .Q(n192) );
  NOR21 U154 ( .A(n179), .B(n161), .Q(n208) );
  NAND22 U155 ( .A(n211), .B(n105), .Q(n209) );
  NAND26 U156 ( .A(B[7]), .B(n297), .Q(n76) );
  NOR23 U157 ( .A(n265), .B(n266), .Q(n258) );
  NAND24 U158 ( .A(n267), .B(n27), .Q(n265) );
  NAND43 U159 ( .A(n110), .B(n233), .C(n268), .D(n12), .Q(n176) );
  NAND21 U160 ( .A(n77), .B(n76), .Q(n182) );
  NAND21 U161 ( .A(n16), .B(A[8]), .Q(n80) );
  NAND21 U162 ( .A(A[5]), .B(n116), .Q(n104) );
  NAND21 U163 ( .A(n172), .B(n187), .Q(n186) );
  NOR33 U164 ( .A(n214), .B(n215), .C(n216), .Q(n213) );
  NOR24 U165 ( .A(n62), .B(n59), .Q(n13) );
  AOI211 U166 ( .A(n107), .B(n9), .C(n97), .Q(n114) );
  INV6 U167 ( .A(n111), .Q(n53) );
  CLKIN6 U168 ( .A(n185), .Q(n14) );
  NAND33 U169 ( .A(n206), .B(n96), .C(n205), .Q(n243) );
  NAND21 U170 ( .A(n184), .B(n172), .Q(n183) );
  NAND30 U171 ( .A(n17), .B(n96), .C(n76), .Q(n283) );
  NOR20 U172 ( .A(n129), .B(n126), .Q(n132) );
  INV6 U173 ( .A(n56), .Q(n272) );
  NAND24 U174 ( .A(n314), .B(n217), .Q(n51) );
  INV2 U175 ( .A(n57), .Q(n15) );
  NAND22 U176 ( .A(B[12]), .B(n249), .Q(n20) );
  NOR21 U177 ( .A(n325), .B(n221), .Q(n220) );
  INV3 U178 ( .A(n306), .Q(n30) );
  NAND22 U179 ( .A(B[10]), .B(n323), .Q(n17) );
  CLKIN6 U180 ( .A(n188), .Q(n172) );
  NOR22 U181 ( .A(n185), .B(n186), .Q(n180) );
  NOR24 U182 ( .A(A[8]), .B(n16), .Q(n303) );
  INV6 U183 ( .A(B[1]), .Q(n315) );
  NOR24 U184 ( .A(n66), .B(n250), .Q(n260) );
  AOI312 U185 ( .A(n69), .B(n288), .C(n9), .D(n293), .Q(n292) );
  INV2 U186 ( .A(A[4]), .Q(n119) );
  NOR21 U187 ( .A(n54), .B(n133), .Q(n129) );
  INV2 U188 ( .A(n163), .Q(n194) );
  NAND21 U189 ( .A(n163), .B(n159), .Q(n188) );
  AOI312 U190 ( .A(n157), .B(n154), .C(n174), .D(n175), .Q(n173) );
  AOI222 U191 ( .A(n66), .B(n31), .C(n67), .D(n68), .Q(n65) );
  XNR22 U192 ( .A(n274), .B(n275), .Q(DIFF[11]) );
  AOI311 U193 ( .A(n268), .B(n12), .C(n286), .D(n287), .Q(n276) );
  OAI220 U194 ( .A(n235), .B(n75), .C(n289), .D(n75), .Q(n286) );
  XOR22 U195 ( .A(n90), .B(n91), .Q(DIFF[7]) );
  NAND34 U196 ( .A(n92), .B(n93), .C(n94), .Q(n91) );
  NAND23 U197 ( .A(B[3]), .B(n307), .Q(n225) );
  INV3 U198 ( .A(A[3]), .Q(n307) );
  NOR24 U199 ( .A(n142), .B(n53), .Q(n267) );
  OAI312 U200 ( .A(n198), .B(n53), .C(n199), .D(n200), .Q(n196) );
  INV6 U201 ( .A(A[9]), .Q(n61) );
  NAND21 U202 ( .A(A[9]), .B(n6), .Q(n305) );
  NAND22 U203 ( .A(n245), .B(n246), .Q(n18) );
  NAND34 U204 ( .A(n248), .B(n247), .C(n19), .Q(n179) );
  INV2 U205 ( .A(n13), .Q(n247) );
  XNR22 U206 ( .A(n167), .B(n4), .Q(DIFF[15]) );
  NOR24 U207 ( .A(n74), .B(n75), .Q(n73) );
  XOR22 U208 ( .A(n291), .B(n292), .Q(DIFF[10]) );
  NAND23 U209 ( .A(n316), .B(n246), .Q(n284) );
  AOI311 U210 ( .A(n105), .B(n28), .C(n106), .D(n98), .Q(n103) );
  INV0 U211 ( .A(n309), .Q(n21) );
  NAND28 U212 ( .A(n23), .B(B[15]), .Q(n22) );
  INV0 U213 ( .A(n315), .Q(n54) );
  NOR24 U214 ( .A(n325), .B(n221), .Q(n314) );
  NOR22 U215 ( .A(n24), .B(n140), .Q(n138) );
  NAND20 U216 ( .A(n17), .B(n225), .Q(n42) );
  INV6 U217 ( .A(n179), .Q(n184) );
  NAND24 U218 ( .A(n143), .B(n144), .Q(n137) );
  INV6 U219 ( .A(n2), .Q(n145) );
  NAND21 U220 ( .A(n69), .B(n141), .Q(n270) );
  OAI210 U221 ( .A(n81), .B(n285), .C(n17), .Q(n278) );
  NAND20 U222 ( .A(n17), .B(n10), .Q(n291) );
  AOI311 U223 ( .A(n268), .B(n12), .C(n269), .D(n270), .Q(n256) );
  NAND24 U224 ( .A(n170), .B(n169), .Q(n36) );
  INV3 U225 ( .A(n176), .Q(n231) );
  NAND21 U226 ( .A(n244), .B(n111), .Q(n296) );
  NOR24 U227 ( .A(A[14]), .B(n166), .Q(n165) );
  NOR23 U228 ( .A(A[7]), .B(n304), .Q(n320) );
  NAND28 U229 ( .A(n271), .B(n272), .Q(n162) );
  NAND20 U230 ( .A(n210), .B(n187), .Q(n239) );
  NAND22 U231 ( .A(n35), .B(n185), .Q(n257) );
  NOR24 U232 ( .A(n219), .B(n218), .Q(n217) );
  NAND21 U233 ( .A(n172), .B(n155), .Q(n174) );
  INV12 U234 ( .A(n161), .Q(n69) );
  NAND22 U235 ( .A(n110), .B(n71), .Q(n109) );
  NOR23 U236 ( .A(n212), .B(n213), .Q(n211) );
  NAND31 U237 ( .A(n152), .B(n150), .C(n259), .Q(n210) );
  NOR24 U238 ( .A(n153), .B(n191), .Q(n190) );
  INV6 U239 ( .A(n51), .Q(n52) );
  INV2 U240 ( .A(n206), .Q(n203) );
  INV3 U241 ( .A(n98), .Q(n95) );
  XOR22 U242 ( .A(n227), .B(n228), .Q(DIFF[13]) );
  INV6 U243 ( .A(B[7]), .Q(n304) );
  NOR23 U244 ( .A(A[2]), .B(n310), .Q(n221) );
  XOR22 U245 ( .A(n64), .B(n65), .Q(DIFF[9]) );
  NAND23 U246 ( .A(B[2]), .B(n308), .Q(n123) );
  NAND33 U247 ( .A(n239), .B(n5), .C(n240), .Q(n229) );
  BUF2 U248 ( .A(n3), .Q(n31) );
  AOI211 U249 ( .A(n122), .B(n123), .C(n124), .Q(n121) );
  INV3 U250 ( .A(n220), .Q(n214) );
  NAND28 U251 ( .A(n317), .B(n318), .Q(n161) );
  OAI2112 U252 ( .A(n266), .B(n296), .C(n288), .D(n76), .Q(n295) );
  INV4 U253 ( .A(n284), .Q(n288) );
  AOI212 U254 ( .A(n79), .B(n80), .C(n284), .Q(n285) );
  OAI212 U255 ( .A(A[2]), .B(n310), .C(n315), .Q(n311) );
  NAND31 U256 ( .A(n27), .B(n111), .C(n282), .Q(n281) );
  NAND34 U257 ( .A(n245), .B(n246), .C(n58), .Q(n46) );
  INV2 U258 ( .A(n55), .Q(n154) );
  NAND34 U259 ( .A(n72), .B(n28), .C(n71), .Q(n40) );
  NOR24 U260 ( .A(n160), .B(n165), .Q(n164) );
  NAND24 U261 ( .A(n262), .B(n261), .Q(n150) );
  INV6 U262 ( .A(n44), .Q(n45) );
  NOR24 U263 ( .A(n53), .B(n199), .Q(n242) );
  NAND28 U264 ( .A(n52), .B(n313), .Q(n72) );
  INV6 U265 ( .A(n48), .Q(n49) );
  INV2 U266 ( .A(A[2]), .Q(n308) );
  AOI212 U267 ( .A(n192), .B(n193), .C(n194), .Q(n191) );
  INV2 U268 ( .A(A[7]), .Q(n297) );
  AOI211 U269 ( .A(n69), .B(n9), .C(n87), .Q(n85) );
  INV2 U270 ( .A(n123), .Q(n290) );
  IMUX22 U271 ( .A(n253), .B(n254), .S(n255), .Q(DIFF[12]) );
  NAND22 U272 ( .A(n72), .B(n71), .Q(n32) );
  NAND33 U273 ( .A(n34), .B(n76), .C(n141), .Q(n35) );
  INV2 U274 ( .A(n258), .Q(n34) );
  INV3 U275 ( .A(n76), .Q(n201) );
  NOR23 U276 ( .A(n256), .B(n257), .Q(n255) );
  NAND24 U277 ( .A(n168), .B(n37), .Q(n167) );
  AOI212 U278 ( .A(n171), .B(n172), .C(n173), .Q(n170) );
  INV3 U279 ( .A(n38), .Q(n39) );
  XOR22 U280 ( .A(n189), .B(n190), .Q(DIFF[14]) );
  NAND22 U281 ( .A(n76), .B(n77), .Q(n88) );
  NOR22 U282 ( .A(n155), .B(n156), .Q(n149) );
  AOI222 U283 ( .A(A[15]), .B(n146), .C(n148), .D(n147), .Q(n143) );
  NAND24 U284 ( .A(n49), .B(n149), .Q(n148) );
  NAND21 U285 ( .A(n79), .B(n80), .Q(n78) );
  NAND21 U286 ( .A(n79), .B(n88), .Q(n87) );
  OAI212 U287 ( .A(n126), .B(n127), .C(n128), .Q(n122) );
  NAND28 U288 ( .A(B[9]), .B(n61), .Q(n246) );
  NAND22 U289 ( .A(A[6]), .B(n298), .Q(n111) );
  AOI212 U290 ( .A(n60), .B(n249), .C(n303), .Q(n248) );
  INV3 U291 ( .A(n42), .Q(n43) );
  NAND21 U292 ( .A(n60), .B(n249), .Q(n187) );
  NAND31 U293 ( .A(n123), .B(n236), .C(n235), .Q(n233) );
  NOR21 U294 ( .A(n81), .B(n285), .Q(n294) );
  NAND22 U295 ( .A(n280), .B(n281), .Q(n279) );
  NAND20 U296 ( .A(n108), .B(n104), .Q(n113) );
  XNR20 U297 ( .A(n50), .B(n62), .Q(n274) );
  NAND31 U298 ( .A(n278), .B(n10), .C(n279), .Q(n277) );
  NAND20 U299 ( .A(n96), .B(n111), .Q(n101) );
  NAND22 U300 ( .A(n224), .B(n225), .Q(n223) );
  INV3 U301 ( .A(n130), .Q(n127) );
  NAND31 U302 ( .A(n96), .B(n97), .C(n95), .Q(n93) );
  XOR20 U303 ( .A(n130), .B(n132), .Q(DIFF[1]) );
  AOI210 U304 ( .A(n15), .B(n219), .C(n290), .Q(n289) );
  AOI210 U305 ( .A(n100), .B(n96), .C(n53), .Q(n92) );
  INV2 U306 ( .A(n135), .Q(n134) );
  NAND22 U307 ( .A(n241), .B(n77), .Q(n240) );
  NAND21 U308 ( .A(n69), .B(n184), .Q(n232) );
  INV2 U309 ( .A(n129), .Q(n128) );
  NOR20 U310 ( .A(n81), .B(n82), .Q(n64) );
  INV0 U311 ( .A(n246), .Q(n82) );
  AOI210 U312 ( .A(n15), .B(n219), .C(n238), .Q(n273) );
  XOR21 U313 ( .A(n101), .B(n102), .Q(DIFF[6]) );
  NAND20 U314 ( .A(n163), .B(n157), .Q(n227) );
  INV3 U315 ( .A(n131), .Q(n124) );
  INV3 U316 ( .A(n197), .Q(n155) );
  IMUX21 U317 ( .A(n83), .B(n84), .S(n85), .Q(DIFF[8]) );
  AOI210 U318 ( .A(B[4]), .B(n119), .C(n97), .Q(n118) );
  AOI311 U319 ( .A(n157), .B(n154), .C(n139), .D(n158), .Q(n147) );
  XNR21 U320 ( .A(n120), .B(n121), .Q(DIFF[3]) );
  NAND22 U321 ( .A(B[5]), .B(n302), .Q(n206) );
  AOI210 U322 ( .A(n60), .B(n249), .C(n155), .Q(n253) );
  NAND22 U323 ( .A(n324), .B(n134), .Q(DIFF[0]) );
  NAND22 U324 ( .A(n134), .B(n237), .Q(n130) );
  NAND20 U325 ( .A(n219), .B(n15), .Q(n324) );
  NAND20 U326 ( .A(n123), .B(n131), .Q(n125) );
  NAND22 U327 ( .A(A[2]), .B(n310), .Q(n131) );
  AOI210 U328 ( .A(n31), .B(n66), .C(n89), .Q(n83) );
  XOR21 U329 ( .A(n113), .B(n114), .Q(DIFF[5]) );
  XNR20 U330 ( .A(B[7]), .B(A[7]), .Q(n90) );
  XOR20 U331 ( .A(B[4]), .B(A[4]), .Q(n117) );
  XOR20 U332 ( .A(n31), .B(A[8]), .Q(n84) );
  XOR20 U333 ( .A(n60), .B(A[12]), .Q(n254) );
  NAND22 U334 ( .A(n294), .B(n295), .Q(n293) );
  XNR20 U335 ( .A(n21), .B(A[3]), .Q(n120) );
  CLKIN3 U336 ( .A(n80), .Q(n89) );
  CLKIN3 U337 ( .A(n104), .Q(n100) );
  AOI2112 U338 ( .A(n136), .B(n86), .C(n138), .D(n137), .Q(DIFF[16]) );
  CLKIN3 U339 ( .A(n96), .Q(n202) );
  OAI212 U340 ( .A(n232), .B(n231), .C(n207), .Q(n230) );
  CLKIN3 U341 ( .A(n225), .Q(n238) );
  CLKIN3 U342 ( .A(n71), .Q(n234) );
  CLKIN3 U343 ( .A(n305), .Q(n81) );
  OAI212 U344 ( .A(A[0]), .B(n57), .C(n225), .Q(n306) );
endmodule


module E_alu_DW01_cmp2_4 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262;

  INV0 U1 ( .A(A[5]), .Q(n115) );
  NOR23 U2 ( .A(n59), .B(n60), .Q(n57) );
  NOR23 U3 ( .A(n197), .B(n198), .Q(n196) );
  INV3 U4 ( .A(B[20]), .Q(n14) );
  NAND22 U5 ( .A(n61), .B(B[7]), .Q(n60) );
  NAND24 U6 ( .A(A[15]), .B(n240), .Q(n135) );
  NAND22 U7 ( .A(n206), .B(n207), .Q(n205) );
  INV6 U8 ( .A(n166), .Q(n197) );
  NAND40 U9 ( .A(B[20]), .B(n165), .C(n166), .D(n167), .Q(n209) );
  AOI312 U10 ( .A(n175), .B(n174), .C(n49), .D(n176), .Q(n168) );
  CLKIN6 U11 ( .A(n44), .Q(n4) );
  NAND21 U12 ( .A(A[14]), .B(n183), .Q(n133) );
  INV4 U13 ( .A(n213), .Q(n204) );
  INV15 U14 ( .A(n2), .Q(n3) );
  NOR23 U15 ( .A(n190), .B(n191), .Q(n189) );
  INV4 U16 ( .A(B[22]), .Q(n262) );
  NAND22 U17 ( .A(A[20]), .B(n14), .Q(n206) );
  NAND23 U18 ( .A(n214), .B(n49), .Q(n188) );
  INV2 U19 ( .A(A[18]), .Q(n256) );
  NAND23 U20 ( .A(n202), .B(n203), .Q(n192) );
  NOR22 U21 ( .A(n204), .B(n205), .Q(n203) );
  INV1 U22 ( .A(A[13]), .Q(n134) );
  INV6 U23 ( .A(n51), .Q(n35) );
  NOR22 U24 ( .A(n32), .B(n51), .Q(n31) );
  NOR20 U25 ( .A(n51), .B(n33), .Q(n30) );
  NOR24 U26 ( .A(A[31]), .B(n52), .Q(n51) );
  NAND41 U27 ( .A(n1), .B(n62), .C(n150), .D(n151), .Q(n149) );
  INV2 U28 ( .A(B[21]), .Q(n255) );
  INV6 U29 ( .A(B[15]), .Q(n240) );
  NAND24 U30 ( .A(A[17]), .B(n249), .Q(n62) );
  NOR23 U31 ( .A(n208), .B(n209), .Q(n190) );
  INV3 U32 ( .A(n46), .Q(n5) );
  NAND42 U33 ( .A(n70), .B(n71), .C(n72), .D(n73), .Q(n46) );
  NOR21 U34 ( .A(n260), .B(n261), .Q(n245) );
  NAND22 U35 ( .A(n146), .B(n147), .Q(n145) );
  NOR23 U36 ( .A(n8), .B(B[23]), .Q(n7) );
  NOR22 U37 ( .A(n77), .B(n92), .Q(n129) );
  NOR32 U38 ( .A(n125), .B(A[8]), .C(n78), .Q(n124) );
  NOR22 U39 ( .A(n229), .B(n230), .Q(n228) );
  NAND24 U40 ( .A(A[25]), .B(n259), .Q(n167) );
  NAND21 U41 ( .A(n68), .B(n19), .Q(n141) );
  INV3 U42 ( .A(n68), .Q(n78) );
  INV2 U43 ( .A(B[9]), .Q(n10) );
  CLKIN10 U44 ( .A(n3), .Q(n61) );
  NOR23 U45 ( .A(n55), .B(n56), .Q(n48) );
  CLKIN12 U46 ( .A(n74), .Q(n58) );
  NAND24 U47 ( .A(n133), .B(n135), .Q(n238) );
  NOR21 U48 ( .A(B[13]), .B(n134), .Q(n239) );
  NAND28 U49 ( .A(n17), .B(A[27]), .Q(n165) );
  INV2 U50 ( .A(B[28]), .Q(n18) );
  NOR21 U51 ( .A(A[28]), .B(n18), .Q(n229) );
  NAND23 U52 ( .A(n50), .B(n35), .Q(n38) );
  INV6 U53 ( .A(n7), .Q(n2) );
  INV2 U54 ( .A(B[30]), .Q(n34) );
  NOR21 U55 ( .A(n92), .B(n93), .Q(n241) );
  NAND21 U56 ( .A(n167), .B(n22), .Q(n224) );
  NAND33 U57 ( .A(n116), .B(n117), .C(n118), .Q(n42) );
  NAND22 U58 ( .A(n119), .B(n49), .Q(n118) );
  NOR21 U59 ( .A(n36), .B(n37), .Q(n28) );
  NOR21 U60 ( .A(n38), .B(n40), .Q(n36) );
  INV3 U61 ( .A(B[24]), .Q(n15) );
  NAND21 U62 ( .A(n1), .B(n256), .Q(n261) );
  NOR22 U63 ( .A(n200), .B(n201), .Q(n199) );
  INV6 U64 ( .A(n62), .Q(n92) );
  NAND22 U65 ( .A(n123), .B(n124), .Q(n120) );
  INV2 U66 ( .A(B[8]), .Q(n9) );
  INV1 U67 ( .A(A[19]), .Q(n207) );
  NOR20 U68 ( .A(A[11]), .B(n77), .Q(n172) );
  NOR21 U69 ( .A(n7), .B(n12), .Q(n151) );
  INV1 U70 ( .A(B[6]), .Q(n84) );
  NAND21 U71 ( .A(B[18]), .B(n61), .Q(n260) );
  NAND20 U72 ( .A(n133), .B(n134), .Q(n132) );
  NAND20 U73 ( .A(A[7]), .B(n85), .Q(n82) );
  CLKIN0 U74 ( .A(A[7]), .Q(n69) );
  NOR21 U75 ( .A(n197), .B(n221), .Q(n218) );
  CLKIN0 U76 ( .A(n107), .Q(n106) );
  INV0 U77 ( .A(A[0]), .Q(n107) );
  CLKIN0 U78 ( .A(B[4]), .Q(n87) );
  NAND23 U79 ( .A(n168), .B(n169), .Q(n144) );
  OAI312 U80 ( .A(n90), .B(n89), .C(n88), .D(n91), .Q(n44) );
  NOR21 U81 ( .A(A[29]), .B(n41), .Q(n53) );
  INV2 U82 ( .A(B[29]), .Q(n41) );
  NAND22 U83 ( .A(n170), .B(n49), .Q(n169) );
  CLKIN3 U84 ( .A(n206), .Q(n254) );
  NOR21 U85 ( .A(n74), .B(n171), .Q(n170) );
  NAND42 U86 ( .A(B[19]), .B(n165), .C(n166), .D(n199), .Q(n193) );
  INV6 U87 ( .A(n237), .Q(n74) );
  NAND20 U88 ( .A(B[5]), .B(n115), .Q(n86) );
  NOR23 U89 ( .A(n144), .B(n145), .Q(n25) );
  NAND41 U90 ( .A(A[4]), .B(n80), .C(n86), .D(n87), .Q(n70) );
  CLKIN2 U91 ( .A(B[2]), .Q(n101) );
  NOR21 U92 ( .A(n38), .B(n39), .Q(n37) );
  NAND22 U93 ( .A(A[11]), .B(n11), .Q(n143) );
  INV2 U94 ( .A(B[12]), .Q(n12) );
  NAND33 U95 ( .A(n4), .B(n49), .C(n5), .Q(n6) );
  NOR22 U96 ( .A(n93), .B(n3), .Q(n202) );
  NOR20 U97 ( .A(n3), .B(n142), .Q(n236) );
  INV1 U98 ( .A(B[7]), .Q(n85) );
  NAND24 U99 ( .A(A[22]), .B(n262), .Q(n1) );
  INV2 U100 ( .A(B[1]), .Q(n104) );
  INV2 U101 ( .A(B[17]), .Q(n249) );
  NAND24 U102 ( .A(A[22]), .B(n262), .Q(n64) );
  NAND22 U103 ( .A(A[21]), .B(n255), .Q(n213) );
  NAND20 U104 ( .A(n1), .B(n62), .Q(n157) );
  NAND20 U105 ( .A(n1), .B(n217), .Q(n215) );
  NAND20 U106 ( .A(n1), .B(n162), .Q(n159) );
  NAND24 U107 ( .A(n250), .B(n251), .Q(n45) );
  NAND22 U108 ( .A(n58), .B(n122), .Q(n121) );
  NOR21 U109 ( .A(n66), .B(n141), .Q(n140) );
  NAND21 U110 ( .A(B[17]), .B(n61), .Q(n216) );
  INV3 U111 ( .A(B[26]), .Q(n16) );
  NAND21 U112 ( .A(B[6]), .B(n95), .Q(n80) );
  INV2 U113 ( .A(A[23]), .Q(n8) );
  INV0 U114 ( .A(A[24]), .Q(n22) );
  NAND24 U115 ( .A(A[24]), .B(n15), .Q(n161) );
  NOR20 U116 ( .A(B[0]), .B(n107), .Q(n105) );
  NAND24 U117 ( .A(n231), .B(n232), .Q(n184) );
  AOI222 U118 ( .A(n245), .B(n49), .C(n246), .D(n49), .Q(n231) );
  NOR22 U119 ( .A(n257), .B(n258), .Q(n250) );
  NAND22 U120 ( .A(n167), .B(n161), .Q(n257) );
  NAND21 U121 ( .A(B[24]), .B(n165), .Q(n225) );
  NOR21 U122 ( .A(n3), .B(n11), .Q(n173) );
  NAND21 U123 ( .A(A[1]), .B(n104), .Q(n103) );
  NOR21 U124 ( .A(A[27]), .B(n17), .Q(n230) );
  NOR23 U125 ( .A(n120), .B(n121), .Q(n119) );
  NAND42 U126 ( .A(n167), .B(n161), .C(n195), .D(n196), .Q(n194) );
  INV4 U127 ( .A(B[14]), .Q(n183) );
  INV0 U128 ( .A(A[9]), .Q(n19) );
  NOR24 U129 ( .A(n234), .B(n235), .Q(n233) );
  NOR21 U130 ( .A(A[22]), .B(n3), .Q(n195) );
  NAND21 U131 ( .A(n165), .B(B[22]), .Q(n198) );
  INV10 U132 ( .A(n63), .Q(n77) );
  NAND22 U133 ( .A(n161), .B(n61), .Q(n160) );
  NAND24 U134 ( .A(A[26]), .B(n16), .Q(n166) );
  INV1 U135 ( .A(B[3]), .Q(n112) );
  INV1 U136 ( .A(B[10]), .Q(n142) );
  CLKIN15 U137 ( .A(n45), .Q(n49) );
  NOR31 U138 ( .A(n247), .B(n93), .C(n248), .Q(n246) );
  NAND21 U139 ( .A(B[16]), .B(n61), .Q(n247) );
  NAND22 U140 ( .A(A[10]), .B(n142), .Q(n68) );
  NAND21 U141 ( .A(n68), .B(n69), .Q(n67) );
  NOR42 U142 ( .A(n252), .B(n253), .C(n254), .D(n204), .Q(n251) );
  NOR21 U143 ( .A(B[18]), .B(n256), .Q(n252) );
  NAND22 U144 ( .A(n58), .B(n139), .Q(n138) );
  NOR31 U145 ( .A(n3), .B(n93), .C(n10), .Q(n139) );
  NAND21 U146 ( .A(B[15]), .B(n61), .Q(n155) );
  NOR21 U147 ( .A(n74), .B(n149), .Q(n148) );
  NAND24 U148 ( .A(n6), .B(n47), .Q(n43) );
  AOI212 U149 ( .A(n48), .B(n49), .C(n38), .Q(n47) );
  NOR21 U150 ( .A(n3), .B(n200), .Q(n210) );
  NOR32 U151 ( .A(n224), .B(n197), .C(n225), .Q(n223) );
  NAND22 U152 ( .A(n75), .B(n76), .Q(n59) );
  NOR31 U153 ( .A(n3), .B(n93), .C(n9), .Q(n122) );
  NOR23 U154 ( .A(n222), .B(n223), .Q(n186) );
  NOR24 U155 ( .A(n43), .B(n42), .Q(n26) );
  CLKIN0 U156 ( .A(B[5]), .Q(n79) );
  NOR21 U157 ( .A(B[19]), .B(n207), .Q(n253) );
  NAND22 U158 ( .A(n167), .B(n8), .Q(n220) );
  NAND20 U159 ( .A(n166), .B(n167), .Q(n163) );
  INV3 U160 ( .A(n167), .Q(n201) );
  NOR24 U161 ( .A(n184), .B(n185), .Q(n24) );
  NAND43 U162 ( .A(n186), .B(n187), .C(n188), .D(n189), .Q(n185) );
  INV2 U163 ( .A(B[11]), .Q(n11) );
  NAND22 U164 ( .A(n148), .B(n49), .Q(n147) );
  AOI221 U165 ( .A(n152), .B(n153), .C(n154), .D(n49), .Q(n146) );
  NAND42 U166 ( .A(n1), .B(n62), .C(n172), .D(n173), .Q(n171) );
  NOR22 U167 ( .A(n59), .B(n74), .Q(n73) );
  NAND21 U168 ( .A(n126), .B(n49), .Q(n117) );
  AOI312 U169 ( .A(n24), .B(n25), .C(n26), .D(n27), .Q(LT_LE) );
  NAND22 U170 ( .A(n236), .B(n58), .Q(n235) );
  NAND21 U171 ( .A(n213), .B(n21), .Q(n212) );
  INV12 U172 ( .A(n64), .Q(n93) );
  NAND42 U173 ( .A(n62), .B(n63), .C(n1), .D(n65), .Q(n55) );
  AOI2112 U174 ( .A(A[12]), .B(n12), .C(n239), .D(n238), .Q(n237) );
  NAND24 U175 ( .A(A[16]), .B(n13), .Q(n63) );
  NAND22 U176 ( .A(A[9]), .B(n10), .Q(n75) );
  INV3 U177 ( .A(n135), .Q(n131) );
  NAND22 U178 ( .A(n135), .B(n182), .Q(n180) );
  CLKIN0 U179 ( .A(A[26]), .Q(n23) );
  NAND22 U180 ( .A(n136), .B(n49), .Q(n116) );
  NAND22 U181 ( .A(n233), .B(n49), .Q(n232) );
  NOR30 U182 ( .A(n3), .B(n93), .C(n183), .Q(n174) );
  CLKIN0 U183 ( .A(A[20]), .Q(n21) );
  NOR21 U184 ( .A(n127), .B(n128), .Q(n126) );
  NOR21 U185 ( .A(n93), .B(n212), .Q(n211) );
  XNR20 U186 ( .A(B[31]), .B(A[31]), .Q(n32) );
  NAND20 U187 ( .A(B[26]), .B(n23), .Q(n227) );
  NOR20 U188 ( .A(n200), .B(n220), .Q(n219) );
  NAND22 U189 ( .A(n111), .B(n96), .Q(n110) );
  NAND20 U190 ( .A(n143), .B(n244), .Q(n243) );
  NOR21 U191 ( .A(n159), .B(n160), .Q(n153) );
  NOR21 U192 ( .A(n177), .B(n178), .Q(n176) );
  NAND22 U193 ( .A(n218), .B(n219), .Q(n187) );
  INV3 U194 ( .A(B[16]), .Q(n13) );
  NAND41 U195 ( .A(n86), .B(n108), .C(n109), .D(n110), .Q(n88) );
  NOR21 U196 ( .A(n99), .B(n100), .Q(n89) );
  NOR30 U197 ( .A(n3), .B(n92), .C(n93), .Q(n91) );
  NAND31 U198 ( .A(n96), .B(B[0]), .C(n97), .Q(n100) );
  NAND22 U199 ( .A(n28), .B(n29), .Q(n27) );
  NAND22 U200 ( .A(n57), .B(n58), .Q(n56) );
  NOR31 U201 ( .A(n155), .B(n156), .C(n157), .Q(n154) );
  NAND20 U202 ( .A(n63), .B(n158), .Q(n156) );
  NAND20 U203 ( .A(n62), .B(n20), .Q(n248) );
  INV0 U204 ( .A(A[16]), .Q(n20) );
  INV3 U205 ( .A(n143), .Q(n66) );
  NAND22 U206 ( .A(n210), .B(n211), .Q(n208) );
  NAND31 U207 ( .A(B[13]), .B(n1), .C(n61), .Q(n128) );
  NAND22 U208 ( .A(n129), .B(n130), .Q(n127) );
  NOR21 U209 ( .A(n163), .B(n164), .Q(n152) );
  NAND20 U210 ( .A(B[21]), .B(n165), .Q(n164) );
  NOR21 U211 ( .A(n137), .B(n138), .Q(n136) );
  NAND22 U212 ( .A(n129), .B(n140), .Q(n137) );
  NOR21 U213 ( .A(n131), .B(n132), .Q(n130) );
  NOR21 U214 ( .A(n30), .B(n31), .Q(n29) );
  NOR21 U215 ( .A(n215), .B(n216), .Q(n214) );
  NAND22 U216 ( .A(n241), .B(n242), .Q(n234) );
  NAND20 U217 ( .A(n165), .B(B[23]), .Q(n221) );
  INV3 U218 ( .A(B[31]), .Q(n52) );
  INV3 U219 ( .A(B[27]), .Q(n17) );
  NAND22 U220 ( .A(n94), .B(n80), .Q(n90) );
  INV2 U221 ( .A(B[25]), .Q(n259) );
  NAND22 U222 ( .A(n82), .B(n83), .Q(n81) );
  NOR21 U223 ( .A(n53), .B(n54), .Q(n50) );
  NOR20 U224 ( .A(A[30]), .B(n34), .Q(n54) );
  NAND20 U225 ( .A(A[30]), .B(n34), .Q(n33) );
  NAND22 U226 ( .A(n102), .B(n103), .Q(n99) );
  NOR21 U227 ( .A(n105), .B(n106), .Q(n102) );
  NAND20 U228 ( .A(B[4]), .B(n114), .Q(n108) );
  NOR21 U229 ( .A(n66), .B(n67), .Q(n65) );
  NOR21 U230 ( .A(n180), .B(n181), .Q(n175) );
  NAND20 U231 ( .A(n62), .B(n63), .Q(n181) );
  INV0 U232 ( .A(A[21]), .Q(n162) );
  NAND20 U233 ( .A(B[25]), .B(n165), .Q(n178) );
  NAND20 U234 ( .A(n166), .B(n179), .Q(n177) );
  NAND22 U235 ( .A(n165), .B(n166), .Q(n258) );
  NOR31 U236 ( .A(n77), .B(n78), .C(n66), .Q(n72) );
  INV0 U237 ( .A(A[1]), .Q(n98) );
  NAND20 U238 ( .A(A[6]), .B(n84), .Q(n83) );
  CLKIN0 U239 ( .A(A[6]), .Q(n95) );
  CLKIN0 U240 ( .A(A[14]), .Q(n182) );
  NAND22 U241 ( .A(A[3]), .B(n112), .Q(n96) );
  NOR20 U242 ( .A(A[2]), .B(n101), .Q(n111) );
  NAND20 U243 ( .A(A[2]), .B(n101), .Q(n97) );
  INV0 U244 ( .A(A[4]), .Q(n114) );
  NAND40 U245 ( .A(B[1]), .B(n96), .C(n97), .D(n98), .Q(n94) );
  CLKIN0 U246 ( .A(A[17]), .Q(n217) );
  CLKIN0 U247 ( .A(A[15]), .Q(n158) );
  NOR21 U248 ( .A(n77), .B(n243), .Q(n242) );
  NOR31 U249 ( .A(n77), .B(n66), .C(n92), .Q(n123) );
  NAND20 U250 ( .A(A[8]), .B(n9), .Q(n76) );
  INV0 U251 ( .A(A[10]), .Q(n244) );
  NAND20 U252 ( .A(B[3]), .B(n113), .Q(n109) );
  AOI311 U253 ( .A(A[5]), .B(n79), .C(n80), .D(n81), .Q(n71) );
  INV1 U254 ( .A(A[3]), .Q(n113) );
  NAND20 U255 ( .A(A[29]), .B(n41), .Q(n40) );
  INV0 U256 ( .A(A[25]), .Q(n179) );
  NOR20 U257 ( .A(A[12]), .B(n77), .Q(n150) );
  NAND20 U258 ( .A(A[28]), .B(n18), .Q(n39) );
  CLKIN3 U259 ( .A(n75), .Q(n125) );
  OAI212 U260 ( .A(n193), .B(n192), .C(n194), .Q(n191) );
  CLKIN3 U261 ( .A(n161), .Q(n200) );
  OAI212 U262 ( .A(n226), .B(n227), .C(n228), .Q(n222) );
  CLKIN3 U263 ( .A(n165), .Q(n226) );
endmodule


module E_alu_DW01_sub_13 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202;

  NAND21 U3 ( .A(n72), .B(n63), .Q(n66) );
  NAND28 U4 ( .A(n87), .B(n185), .Q(n127) );
  BUF2 U5 ( .A(n51), .Q(n1) );
  NAND28 U6 ( .A(n35), .B(A[8]), .Q(n50) );
  INV6 U7 ( .A(B[11]), .Q(n37) );
  NOR24 U8 ( .A(n11), .B(B[4]), .Q(n9) );
  NAND26 U9 ( .A(n36), .B(A[10]), .Q(n13) );
  OAI312 U10 ( .A(n180), .B(n160), .C(n181), .D(n56), .Q(n177) );
  XOR22 U11 ( .A(n61), .B(n62), .Q(DIFF[7]) );
  INV6 U12 ( .A(A[5]), .Q(n79) );
  NOR24 U13 ( .A(n165), .B(n60), .Q(n164) );
  CLKIN6 U14 ( .A(n28), .Q(n165) );
  INV6 U15 ( .A(n93), .Q(n87) );
  NAND28 U16 ( .A(n188), .B(n18), .Q(n128) );
  CLKIN8 U17 ( .A(n144), .Q(n122) );
  NAND26 U18 ( .A(n67), .B(n198), .Q(n145) );
  NAND33 U19 ( .A(n146), .B(n145), .C(n194), .Q(n141) );
  INV12 U20 ( .A(B[9]), .Q(n200) );
  INV1 U21 ( .A(A[9]), .Q(n179) );
  NAND26 U22 ( .A(n50), .B(n52), .Q(n153) );
  CLKIN10 U23 ( .A(A[4]), .Q(n11) );
  NAND26 U24 ( .A(n133), .B(n134), .Q(n132) );
  AOI212 U25 ( .A(n56), .B(n47), .C(n57), .Q(n55) );
  NAND28 U26 ( .A(n158), .B(n159), .Q(n47) );
  NAND24 U27 ( .A(n13), .B(n155), .Q(n154) );
  INV4 U28 ( .A(A[2]), .Q(n192) );
  NAND28 U29 ( .A(n152), .B(n51), .Q(n19) );
  INV1 U30 ( .A(n152), .Q(n170) );
  INV12 U31 ( .A(A[1]), .Q(n193) );
  NAND31 U32 ( .A(n1), .B(n15), .C(n46), .Q(n172) );
  NAND22 U33 ( .A(B[8]), .B(n40), .Q(n46) );
  INV3 U34 ( .A(n185), .Q(n189) );
  NAND24 U35 ( .A(n179), .B(B[9]), .Q(n51) );
  AOI211 U36 ( .A(n171), .B(n177), .C(n178), .Q(n176) );
  NOR22 U37 ( .A(n156), .B(n157), .Q(n151) );
  INV3 U38 ( .A(B[1]), .Q(n187) );
  NAND22 U39 ( .A(A[2]), .B(n31), .Q(n93) );
  NAND23 U40 ( .A(n110), .B(n104), .Q(n108) );
  NAND23 U41 ( .A(n44), .B(n45), .Q(n43) );
  NOR22 U42 ( .A(n175), .B(n176), .Q(n174) );
  NOR23 U43 ( .A(A[7]), .B(n34), .Q(n27) );
  NOR21 U44 ( .A(A[4]), .B(n33), .Q(n82) );
  NAND22 U45 ( .A(n68), .B(n69), .Q(n72) );
  NOR24 U46 ( .A(A[5]), .B(n78), .Q(n198) );
  INV12 U47 ( .A(B[8]), .Q(n35) );
  NOR23 U48 ( .A(n49), .B(n57), .Q(n171) );
  NOR24 U49 ( .A(A[8]), .B(n35), .Q(n60) );
  NAND28 U50 ( .A(n127), .B(n124), .Q(n181) );
  NOR23 U51 ( .A(n197), .B(n9), .Q(n196) );
  CLKIN3 U52 ( .A(A[10]), .Q(n41) );
  NOR24 U53 ( .A(A[6]), .B(n199), .Q(n147) );
  INV12 U54 ( .A(B[3]), .Q(n32) );
  CLKIN3 U55 ( .A(n120), .Q(n131) );
  INV2 U56 ( .A(B[2]), .Q(n31) );
  NAND24 U57 ( .A(n47), .B(n26), .Q(n45) );
  INV3 U58 ( .A(n23), .Q(n24) );
  INV6 U59 ( .A(n128), .Q(n160) );
  INV2 U60 ( .A(A[12]), .Q(n136) );
  NAND33 U61 ( .A(n92), .B(n86), .C(n30), .Q(n17) );
  NAND24 U62 ( .A(n196), .B(n67), .Q(n146) );
  INV6 U63 ( .A(B[7]), .Q(n34) );
  NOR21 U64 ( .A(n27), .B(n122), .Q(n143) );
  NAND22 U65 ( .A(B[4]), .B(n11), .Q(n10) );
  BUF2 U66 ( .A(n67), .Q(n3) );
  NAND26 U67 ( .A(B[1]), .B(n193), .Q(n92) );
  XOR21 U68 ( .A(n149), .B(n148), .Q(DIFF[12]) );
  NOR22 U69 ( .A(n168), .B(n169), .Q(n167) );
  INV3 U70 ( .A(A[3]), .Q(n190) );
  NAND21 U71 ( .A(n56), .B(n46), .Q(n25) );
  NOR24 U72 ( .A(n38), .B(n30), .Q(n96) );
  NAND26 U73 ( .A(B[12]), .B(n136), .Q(n144) );
  NOR21 U74 ( .A(A[14]), .B(n107), .Q(n103) );
  INV3 U75 ( .A(B[14]), .Q(n107) );
  INV6 U76 ( .A(n39), .Q(n38) );
  INV4 U77 ( .A(A[0]), .Q(n39) );
  INV1 U78 ( .A(A[8]), .Q(n40) );
  INV3 U79 ( .A(n2), .Q(n49) );
  NOR21 U80 ( .A(B[13]), .B(n111), .Q(n106) );
  INV3 U81 ( .A(n106), .Q(n104) );
  INV3 U82 ( .A(n97), .Q(n202) );
  XNR21 U83 ( .A(B[15]), .B(A[15]), .Q(n16) );
  NOR20 U84 ( .A(A[13]), .B(n113), .Q(n112) );
  CLKIN0 U85 ( .A(A[13]), .Q(n111) );
  XOR21 U86 ( .A(n76), .B(n77), .Q(DIFF[5]) );
  OAI212 U87 ( .A(n125), .B(n90), .C(n91), .Q(n85) );
  NAND24 U88 ( .A(A[1]), .B(n187), .Q(n91) );
  INV3 U89 ( .A(n59), .Q(n157) );
  NAND24 U90 ( .A(B[6]), .B(n183), .Q(n63) );
  NOR23 U91 ( .A(n39), .B(n189), .Q(n188) );
  IMUX20 U92 ( .A(n80), .B(n81), .S(n47), .Q(DIFF[4]) );
  AOI211 U93 ( .A(n75), .B(n47), .C(n9), .Q(n77) );
  NAND20 U94 ( .A(n92), .B(n91), .Q(n94) );
  NAND20 U95 ( .A(A[8]), .B(n35), .Q(n2) );
  NOR23 U96 ( .A(n27), .B(n198), .Q(n182) );
  AOI211 U97 ( .A(n57), .B(n46), .C(n49), .Q(n44) );
  NOR23 U98 ( .A(A[11]), .B(n37), .Q(n140) );
  NAND26 U99 ( .A(n59), .B(n58), .Q(n57) );
  INV4 U100 ( .A(B[5]), .Q(n78) );
  NAND24 U101 ( .A(A[11]), .B(n37), .Q(n155) );
  NAND26 U102 ( .A(B[10]), .B(n41), .Q(n152) );
  NAND20 U103 ( .A(n1), .B(n46), .Q(n178) );
  INV6 U104 ( .A(B[0]), .Q(n30) );
  OAI210 U105 ( .A(n170), .B(n52), .C(n13), .Q(n169) );
  CLKIN1 U106 ( .A(A[6]), .Q(n183) );
  NAND28 U107 ( .A(A[9]), .B(n200), .Q(n52) );
  BUF6 U108 ( .A(n86), .Q(n4) );
  NOR22 U109 ( .A(B[5]), .B(n79), .Q(n197) );
  INV2 U110 ( .A(B[4]), .Q(n33) );
  INV4 U111 ( .A(B[10]), .Q(n36) );
  NAND21 U112 ( .A(B[5]), .B(n79), .Q(n73) );
  NAND22 U113 ( .A(n9), .B(n73), .Q(n68) );
  INV8 U114 ( .A(B[6]), .Q(n199) );
  NOR24 U115 ( .A(n8), .B(n120), .Q(n119) );
  NAND28 U116 ( .A(n164), .B(n20), .Q(n120) );
  NAND28 U117 ( .A(B[3]), .B(n190), .Q(n185) );
  INV0 U118 ( .A(n63), .Q(n5) );
  INV3 U119 ( .A(n5), .Q(n6) );
  AOI212 U120 ( .A(n64), .B(n47), .C(n72), .Q(n71) );
  NAND21 U121 ( .A(n66), .B(n3), .Q(n65) );
  NAND28 U122 ( .A(A[6]), .B(n199), .Q(n67) );
  NOR23 U123 ( .A(n122), .B(n121), .Q(n7) );
  CLKIN6 U124 ( .A(n7), .Q(n8) );
  CLKIN3 U125 ( .A(n103), .Q(n100) );
  NAND24 U126 ( .A(n115), .B(n116), .Q(n101) );
  XOR21 U127 ( .A(n70), .B(n71), .Q(DIFF[6]) );
  INV3 U128 ( .A(n96), .Q(n129) );
  INV0 U129 ( .A(n52), .Q(n175) );
  NAND26 U130 ( .A(n138), .B(n137), .Q(n133) );
  AOI211 U131 ( .A(n85), .B(n4), .C(n87), .Q(n84) );
  NOR21 U132 ( .A(B[0]), .B(n39), .Q(n97) );
  INV1 U133 ( .A(B[13]), .Q(n113) );
  INV1 U134 ( .A(n138), .Q(n14) );
  NAND21 U135 ( .A(A[5]), .B(n78), .Q(n69) );
  NOR22 U136 ( .A(n140), .B(n122), .Q(n137) );
  INV12 U137 ( .A(n21), .Q(n22) );
  NAND28 U138 ( .A(n10), .B(n63), .Q(n21) );
  INV2 U139 ( .A(n170), .Q(n15) );
  BUF2 U140 ( .A(n120), .Q(n12) );
  OAI222 U141 ( .A(n151), .B(n12), .C(n140), .D(n14), .Q(n150) );
  INV6 U142 ( .A(n147), .Q(n194) );
  XNR22 U143 ( .A(n42), .B(n43), .Q(DIFF[9]) );
  INV6 U144 ( .A(n139), .Q(n138) );
  NAND26 U145 ( .A(n184), .B(n185), .Q(n124) );
  XOR22 U146 ( .A(n173), .B(n174), .Q(DIFF[10]) );
  NAND22 U147 ( .A(n101), .B(n99), .Q(n110) );
  NOR24 U148 ( .A(n186), .B(n91), .Q(n184) );
  XNR22 U149 ( .A(n166), .B(n167), .Q(DIFF[11]) );
  INV12 U150 ( .A(n19), .Q(n20) );
  XNR22 U151 ( .A(n16), .B(n98), .Q(DIFF[15]) );
  NAND22 U152 ( .A(n123), .B(n124), .Q(n118) );
  AOI312 U153 ( .A(n56), .B(n131), .C(n47), .D(n150), .Q(n148) );
  AOI312 U154 ( .A(n6), .B(n64), .C(n47), .D(n65), .Q(n61) );
  OAI220 U155 ( .A(n103), .B(n104), .C(B[14]), .D(n105), .Q(n102) );
  NOR23 U156 ( .A(n96), .B(n121), .Q(n191) );
  NOR23 U157 ( .A(A[3]), .B(n32), .Q(n121) );
  OAI2112 U158 ( .A(n125), .B(n126), .C(n127), .D(n128), .Q(n117) );
  NAND22 U159 ( .A(B[11]), .B(n29), .Q(n28) );
  XNR20 U160 ( .A(B[13]), .B(A[13]), .Q(n114) );
  AOI212 U161 ( .A(n58), .B(n141), .C(n142), .Q(n130) );
  XOR22 U162 ( .A(n108), .B(n109), .Q(DIFF[14]) );
  NAND26 U163 ( .A(B[2]), .B(n192), .Q(n86) );
  NAND22 U164 ( .A(n92), .B(n86), .Q(n23) );
  CLKIN6 U165 ( .A(n86), .Q(n186) );
  NAND22 U166 ( .A(n129), .B(n4), .Q(n126) );
  INV6 U167 ( .A(n17), .Q(n18) );
  NAND28 U168 ( .A(n182), .B(n22), .Q(n48) );
  INV12 U169 ( .A(n48), .Q(n56) );
  NAND24 U170 ( .A(n191), .B(n24), .Q(n163) );
  INV3 U171 ( .A(n163), .Q(n162) );
  INV3 U172 ( .A(n25), .Q(n26) );
  NAND43 U173 ( .A(n195), .B(n145), .C(n194), .D(n146), .Q(n59) );
  IMUX21 U174 ( .A(n53), .B(n54), .S(n55), .Q(DIFF[8]) );
  AOI212 U175 ( .A(n130), .B(n131), .C(n132), .Q(n115) );
  NAND22 U176 ( .A(n163), .B(n123), .Q(n180) );
  OAI2112 U177 ( .A(n118), .B(n117), .C(n56), .D(n119), .Q(n116) );
  CLKIN2 U178 ( .A(A[11]), .Q(n29) );
  INV2 U179 ( .A(n92), .Q(n125) );
  NAND22 U180 ( .A(A[3]), .B(n32), .Q(n123) );
  INV2 U181 ( .A(n82), .Q(n75) );
  NAND22 U182 ( .A(n75), .B(n73), .Q(n74) );
  XOR20 U183 ( .A(n94), .B(n90), .Q(DIFF[1]) );
  NAND20 U184 ( .A(n73), .B(n69), .Q(n76) );
  NAND20 U185 ( .A(n51), .B(n52), .Q(n42) );
  CLKIN3 U186 ( .A(n143), .Q(n142) );
  CLKIN3 U187 ( .A(n135), .Q(n134) );
  CLKIN3 U188 ( .A(n112), .Q(n99) );
  NAND22 U189 ( .A(n202), .B(n96), .Q(n95) );
  NOR20 U190 ( .A(n82), .B(n9), .Q(n81) );
  INV3 U191 ( .A(n27), .Q(n195) );
  XNR20 U192 ( .A(B[11]), .B(A[11]), .Q(n166) );
  NOR20 U193 ( .A(n60), .B(n49), .Q(n53) );
  NAND20 U194 ( .A(n63), .B(n3), .Q(n70) );
  NOR23 U195 ( .A(n161), .B(n162), .Q(n158) );
  NAND20 U196 ( .A(n15), .B(n13), .Q(n173) );
  XOR21 U197 ( .A(n88), .B(n89), .Q(DIFF[2]) );
  NAND20 U198 ( .A(n4), .B(n93), .Q(n88) );
  NAND22 U199 ( .A(n201), .B(n202), .Q(DIFF[0]) );
  NAND20 U200 ( .A(n39), .B(B[0]), .Q(n201) );
  XNR21 U201 ( .A(n83), .B(n84), .Q(DIFF[3]) );
  INV0 U202 ( .A(A[14]), .Q(n105) );
  XOR20 U203 ( .A(n101), .B(n114), .Q(DIFF[13]) );
  NAND22 U204 ( .A(A[7]), .B(n34), .Q(n58) );
  XOR20 U205 ( .A(B[4]), .B(A[4]), .Q(n80) );
  XOR20 U206 ( .A(B[12]), .B(A[12]), .Q(n149) );
  NOR21 U207 ( .A(B[12]), .B(n136), .Q(n135) );
  XOR20 U208 ( .A(B[8]), .B(A[8]), .Q(n54) );
  XOR20 U209 ( .A(B[7]), .B(A[7]), .Q(n62) );
  XNR20 U210 ( .A(B[14]), .B(A[14]), .Q(n109) );
  XNR20 U211 ( .A(B[3]), .B(A[3]), .Q(n83) );
  CLKIN3 U212 ( .A(n74), .Q(n64) );
  CLKIN3 U213 ( .A(n85), .Q(n89) );
  CLKIN3 U214 ( .A(n95), .Q(n90) );
  AOI312 U215 ( .A(n99), .B(n100), .C(n101), .D(n102), .Q(n98) );
  AOI312 U216 ( .A(n51), .B(n153), .C(n152), .D(n154), .Q(n139) );
  CLKIN3 U217 ( .A(n58), .Q(n156) );
  NOR24 U218 ( .A(n160), .B(n181), .Q(n159) );
  CLKIN3 U219 ( .A(n123), .Q(n161) );
  AOI212 U220 ( .A(n171), .B(n177), .C(n172), .Q(n168) );
endmodule


module E_alu_DW01_add_27 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103;

  INV8 U2 ( .A(n24), .Q(n20) );
  NAND28 U3 ( .A(n71), .B(n72), .Q(n24) );
  NAND21 U4 ( .A(A[2]), .B(B[2]), .Q(n81) );
  NAND22 U5 ( .A(B[4]), .B(A[4]), .Q(n21) );
  INV6 U6 ( .A(n40), .Q(n44) );
  NOR23 U7 ( .A(A[2]), .B(B[2]), .Q(n40) );
  INV1 U8 ( .A(B[2]), .Q(n14) );
  CLKIN6 U9 ( .A(n4), .Q(n5) );
  NOR22 U10 ( .A(n38), .B(n45), .Q(n88) );
  INV2 U11 ( .A(A[6]), .Q(n72) );
  INV1 U12 ( .A(A[2]), .Q(n84) );
  NAND26 U13 ( .A(n62), .B(n46), .Q(n56) );
  NAND24 U14 ( .A(n87), .B(n88), .Q(n62) );
  NAND23 U15 ( .A(n55), .B(n21), .Q(n52) );
  INV2 U16 ( .A(A[1]), .Q(n85) );
  NAND24 U17 ( .A(n83), .B(n82), .Q(n47) );
  NOR23 U18 ( .A(n66), .B(n65), .Q(n64) );
  NOR23 U19 ( .A(n39), .B(n81), .Q(n48) );
  INV6 U20 ( .A(n48), .Q(n60) );
  XOR22 U21 ( .A(n90), .B(n91), .Q(SUM[3]) );
  CLKIN3 U22 ( .A(n13), .Q(n103) );
  NAND21 U23 ( .A(n13), .B(n15), .Q(n2) );
  NOR22 U24 ( .A(n13), .B(n15), .Q(n4) );
  NOR22 U25 ( .A(n38), .B(n39), .Q(n37) );
  INV3 U26 ( .A(n2), .Q(n89) );
  INV4 U27 ( .A(B[6]), .Q(n71) );
  NOR21 U28 ( .A(n20), .B(n32), .Q(n29) );
  AOI312 U29 ( .A(A[5]), .B(B[5]), .C(n24), .D(n25), .Q(n23) );
  INV3 U30 ( .A(A[0]), .Q(n15) );
  INV3 U31 ( .A(n38), .Q(n42) );
  INV3 U32 ( .A(n22), .Q(n51) );
  NOR24 U33 ( .A(n70), .B(n48), .Q(n69) );
  NAND23 U34 ( .A(n43), .B(n44), .Q(n33) );
  NAND33 U35 ( .A(n46), .B(n60), .C(n47), .Q(n27) );
  INV10 U36 ( .A(B[0]), .Q(n13) );
  INV2 U37 ( .A(n20), .Q(n3) );
  CLKIN2 U38 ( .A(n45), .Q(n43) );
  INV0 U39 ( .A(n42), .Q(n1) );
  NOR22 U40 ( .A(B[3]), .B(A[3]), .Q(n45) );
  NAND22 U41 ( .A(B[3]), .B(A[3]), .Q(n46) );
  NAND21 U42 ( .A(B[1]), .B(A[1]), .Q(n96) );
  CLKIN3 U43 ( .A(B[1]), .Q(n86) );
  NAND22 U44 ( .A(B[6]), .B(A[6]), .Q(n26) );
  NOR21 U45 ( .A(n5), .B(n40), .Q(n36) );
  NOR20 U46 ( .A(A[4]), .B(B[4]), .Q(n77) );
  INV3 U47 ( .A(n51), .Q(n6) );
  NAND23 U48 ( .A(n19), .B(n9), .Q(n17) );
  NOR21 U49 ( .A(n93), .B(n40), .Q(n95) );
  NOR22 U50 ( .A(n22), .B(n31), .Q(n30) );
  NAND22 U51 ( .A(n7), .B(n8), .Q(n9) );
  INV0 U52 ( .A(A[7]), .Q(n7) );
  INV0 U53 ( .A(B[7]), .Q(n8) );
  NAND24 U54 ( .A(n17), .B(n18), .Q(n11) );
  BUF2 U55 ( .A(n26), .Q(n10) );
  NAND26 U56 ( .A(n16), .B(n12), .Q(SUM[8]) );
  NAND21 U57 ( .A(n103), .B(A[0]), .Q(n101) );
  INV6 U58 ( .A(n11), .Q(n12) );
  NOR21 U59 ( .A(n31), .B(n76), .Q(n79) );
  CLKIN6 U60 ( .A(n47), .Q(n70) );
  INV3 U61 ( .A(n21), .Q(n76) );
  NOR22 U62 ( .A(n85), .B(n86), .Q(n82) );
  XOR22 U63 ( .A(n49), .B(n50), .Q(SUM[7]) );
  NAND34 U64 ( .A(n37), .B(n44), .C(n80), .Q(n61) );
  AOI212 U65 ( .A(n59), .B(n75), .C(n76), .Q(n74) );
  INV6 U66 ( .A(n61), .Q(n57) );
  NOR22 U67 ( .A(n40), .B(n89), .Q(n87) );
  OAI210 U68 ( .A(n20), .B(n54), .C(n10), .Q(n53) );
  OAI312 U69 ( .A(n20), .B(n21), .C(n22), .D(n23), .Q(n19) );
  OAI2112 U70 ( .A(n28), .B(n27), .C(n29), .D(n30), .Q(n16) );
  NAND21 U71 ( .A(n60), .B(n47), .Q(n58) );
  XOR22 U72 ( .A(n63), .B(n64), .Q(SUM[6]) );
  AOI212 U73 ( .A(n92), .B(n44), .C(n93), .Q(n91) );
  IMUX22 U74 ( .A(n78), .B(n79), .S(n75), .Q(SUM[4]) );
  NAND42 U75 ( .A(n46), .B(n62), .C(n69), .D(n61), .Q(n75) );
  AOI212 U76 ( .A(n21), .B(n67), .C(n6), .Q(n65) );
  NOR22 U77 ( .A(A[5]), .B(B[5]), .Q(n22) );
  XOR20 U78 ( .A(n98), .B(n99), .Q(SUM[1]) );
  OAI210 U79 ( .A(A[0]), .B(n103), .C(n101), .Q(SUM[0]) );
  NOR20 U80 ( .A(A[0]), .B(n103), .Q(n102) );
  NAND20 U81 ( .A(n15), .B(n13), .Q(n41) );
  INV2 U82 ( .A(n94), .Q(n93) );
  NAND20 U83 ( .A(n51), .B(n54), .Q(n73) );
  NAND22 U84 ( .A(n41), .B(n42), .Q(n34) );
  NAND22 U85 ( .A(n36), .B(n37), .Q(n35) );
  NAND22 U86 ( .A(n101), .B(n102), .Q(n98) );
  NAND22 U87 ( .A(n96), .B(n97), .Q(n92) );
  NAND22 U88 ( .A(n98), .B(n42), .Q(n97) );
  NOR20 U89 ( .A(n100), .B(n1), .Q(n99) );
  XOR21 U90 ( .A(n73), .B(n74), .Q(SUM[5]) );
  XOR21 U91 ( .A(n92), .B(n95), .Q(SUM[2]) );
  CLKIN3 U92 ( .A(n77), .Q(n59) );
  NOR22 U93 ( .A(n15), .B(n13), .Q(n80) );
  NAND20 U94 ( .A(n3), .B(n10), .Q(n63) );
  NAND22 U95 ( .A(n69), .B(n61), .Q(n68) );
  NAND20 U96 ( .A(B[5]), .B(A[5]), .Q(n54) );
  INV3 U97 ( .A(n26), .Q(n25) );
  XNR20 U98 ( .A(B[4]), .B(A[4]), .Q(n78) );
  NOR21 U99 ( .A(B[4]), .B(A[4]), .Q(n31) );
  NAND20 U100 ( .A(B[2]), .B(A[2]), .Q(n94) );
  NAND20 U101 ( .A(B[7]), .B(A[7]), .Q(n18) );
  NOR20 U102 ( .A(B[7]), .B(A[7]), .Q(n32) );
  AOI212 U103 ( .A(n14), .B(n84), .C(n39), .Q(n83) );
  NOR24 U104 ( .A(A[3]), .B(B[3]), .Q(n39) );
  XNR20 U105 ( .A(B[3]), .B(A[3]), .Q(n90) );
  XNR20 U106 ( .A(B[7]), .B(A[7]), .Q(n49) );
  OAI212 U107 ( .A(n33), .B(n34), .C(n35), .Q(n28) );
  AOI312 U108 ( .A(n3), .B(n51), .C(n52), .D(n53), .Q(n50) );
  OAI312 U109 ( .A(n56), .B(n57), .C(n58), .D(n59), .Q(n55) );
  CLKIN3 U110 ( .A(n54), .Q(n66) );
  OAI212 U111 ( .A(n68), .B(n56), .C(n59), .Q(n67) );
  NOR24 U112 ( .A(A[1]), .B(B[1]), .Q(n38) );
  CLKIN3 U113 ( .A(n96), .Q(n100) );
endmodule


module E_alu_DW01_add_24 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95;

  INV3 U2 ( .A(A[5]), .Q(n68) );
  NOR23 U3 ( .A(n23), .B(n24), .Q(n45) );
  BUF15 U4 ( .A(B[2]), .Q(n13) );
  INV1 U5 ( .A(n92), .Q(n1) );
  INV3 U6 ( .A(n30), .Q(n92) );
  INV2 U7 ( .A(n94), .Q(n2) );
  INV1 U8 ( .A(n89), .Q(n94) );
  NAND26 U9 ( .A(B[1]), .B(A[1]), .Q(n89) );
  CLKIN3 U10 ( .A(A[6]), .Q(n61) );
  INV3 U11 ( .A(n29), .Q(n20) );
  AOI212 U12 ( .A(n23), .B(n24), .C(n25), .Q(n22) );
  NAND26 U13 ( .A(n33), .B(n34), .Q(n19) );
  BUF2 U14 ( .A(n59), .Q(n3) );
  NAND23 U15 ( .A(n58), .B(n3), .Q(n53) );
  NAND23 U16 ( .A(B[0]), .B(A[0]), .Q(n79) );
  NOR22 U17 ( .A(n13), .B(n15), .Q(n80) );
  INV4 U18 ( .A(n44), .Q(n25) );
  NAND34 U19 ( .A(n43), .B(n44), .C(n45), .Q(n42) );
  NAND22 U20 ( .A(B[6]), .B(A[6]), .Q(n48) );
  NAND21 U21 ( .A(n2), .B(n90), .Q(n86) );
  NAND24 U22 ( .A(n41), .B(n42), .Q(n39) );
  NOR23 U23 ( .A(A[1]), .B(B[1]), .Q(n30) );
  XOR21 U24 ( .A(n81), .B(n82), .Q(SUM[3]) );
  BUF6 U25 ( .A(A[2]), .Q(n15) );
  CLKBU4 U26 ( .A(A[2]), .Q(n16) );
  INV12 U27 ( .A(B[4]), .Q(n24) );
  NAND28 U28 ( .A(n18), .B(n17), .Q(SUM[8]) );
  CLKIN6 U29 ( .A(n74), .Q(n6) );
  NAND26 U30 ( .A(B[5]), .B(A[5]), .Q(n55) );
  INV6 U31 ( .A(n64), .Q(n58) );
  INV6 U32 ( .A(B[6]), .Q(n60) );
  INV2 U33 ( .A(n24), .Q(n4) );
  NOR24 U34 ( .A(n13), .B(n15), .Q(n75) );
  CLKIN6 U35 ( .A(n9), .Q(n10) );
  BUF2 U36 ( .A(n48), .Q(n5) );
  INV6 U37 ( .A(n6), .Q(n7) );
  AOI212 U38 ( .A(n26), .B(n27), .C(n28), .Q(n21) );
  NOR24 U39 ( .A(n30), .B(n79), .Q(n77) );
  NAND20 U40 ( .A(n14), .B(n16), .Q(n83) );
  OAI210 U41 ( .A(n14), .B(n16), .C(n83), .Q(n88) );
  INV6 U42 ( .A(n55), .Q(n46) );
  IMUX21 U43 ( .A(n69), .B(n70), .S(n58), .Q(SUM[4]) );
  BUF2 U44 ( .A(B[3]), .Q(n8) );
  NOR24 U45 ( .A(n15), .B(n13), .Q(n32) );
  CLKIN2 U46 ( .A(n49), .Q(n38) );
  OAI210 U47 ( .A(n28), .B(n55), .C(n5), .Q(n54) );
  NAND28 U48 ( .A(n60), .B(n61), .Q(n43) );
  NAND20 U49 ( .A(B[4]), .B(A[4]), .Q(n59) );
  CLKIN6 U50 ( .A(n43), .Q(n28) );
  NOR22 U51 ( .A(n26), .B(n27), .Q(n40) );
  INV1 U52 ( .A(A[7]), .Q(n26) );
  AOI212 U53 ( .A(n76), .B(n77), .C(n36), .Q(n71) );
  NOR22 U54 ( .A(n32), .B(n7), .Q(n31) );
  AOI212 U55 ( .A(n46), .B(n43), .C(n47), .Q(n41) );
  CLKBU12 U56 ( .A(B[2]), .Q(n14) );
  NAND24 U57 ( .A(n31), .B(n77), .Q(n29) );
  CLKIN2 U58 ( .A(A[4]), .Q(n23) );
  NOR24 U59 ( .A(n74), .B(n89), .Q(n9) );
  INV2 U60 ( .A(n3), .Q(n65) );
  INV6 U61 ( .A(B[5]), .Q(n67) );
  XOR22 U62 ( .A(n12), .B(n50), .Q(SUM[7]) );
  INV3 U63 ( .A(B[7]), .Q(n27) );
  XOR22 U64 ( .A(n56), .B(n57), .Q(SUM[6]) );
  AOI312 U65 ( .A(n52), .B(n44), .C(n53), .D(n46), .Q(n57) );
  NOR24 U66 ( .A(n36), .B(n37), .Q(n33) );
  NOR21 U67 ( .A(n80), .B(n7), .Q(n76) );
  NOR24 U68 ( .A(n7), .B(n73), .Q(n35) );
  NAND24 U69 ( .A(n16), .B(n14), .Q(n73) );
  NAND28 U70 ( .A(n67), .B(n68), .Q(n44) );
  NAND20 U71 ( .A(n44), .B(n55), .Q(n62) );
  NOR21 U72 ( .A(n35), .B(n37), .Q(n72) );
  CLKIN6 U73 ( .A(n35), .Q(n34) );
  NOR24 U74 ( .A(A[3]), .B(B[3]), .Q(n74) );
  NOR24 U75 ( .A(n75), .B(n10), .Q(n37) );
  INV2 U76 ( .A(n87), .Q(n85) );
  AOI212 U77 ( .A(n38), .B(n39), .C(n40), .Q(n17) );
  XNR20 U78 ( .A(n86), .B(n88), .Q(SUM[2]) );
  NOR20 U79 ( .A(n94), .B(n1), .Q(n93) );
  XOR20 U80 ( .A(n91), .B(n93), .Q(SUM[1]) );
  NOR20 U81 ( .A(n13), .B(n15), .Q(n87) );
  MUX21 U82 ( .A(B[0]), .B(n95), .S(A[0]), .Q(SUM[0]) );
  INV2 U83 ( .A(n66), .Q(n52) );
  XNR20 U84 ( .A(B[7]), .B(A[7]), .Q(n12) );
  INV2 U85 ( .A(n79), .Q(n91) );
  NOR20 U86 ( .A(n25), .B(n28), .Q(n51) );
  NAND20 U87 ( .A(n43), .B(n5), .Q(n56) );
  NAND22 U88 ( .A(n91), .B(n92), .Q(n90) );
  XOR21 U89 ( .A(n62), .B(n63), .Q(SUM[5]) );
  AOI211 U90 ( .A(n52), .B(n64), .C(n65), .Q(n63) );
  NAND22 U91 ( .A(n71), .B(n72), .Q(n64) );
  INV0 U92 ( .A(B[0]), .Q(n95) );
  AOI210 U93 ( .A(n23), .B(n24), .C(n65), .Q(n69) );
  NAND22 U94 ( .A(n83), .B(n84), .Q(n81) );
  NAND22 U95 ( .A(n85), .B(n86), .Q(n84) );
  NOR20 U96 ( .A(A[4]), .B(n4), .Q(n66) );
  NAND21 U97 ( .A(B[3]), .B(A[3]), .Q(n78) );
  NOR21 U98 ( .A(A[7]), .B(B[7]), .Q(n49) );
  XNR20 U99 ( .A(n4), .B(A[4]), .Q(n70) );
  XOR20 U100 ( .A(n8), .B(A[3]), .Q(n82) );
  OAI2112 U101 ( .A(n19), .B(n20), .C(n22), .D(n21), .Q(n18) );
  CLKIN3 U102 ( .A(n48), .Q(n47) );
  AOI312 U103 ( .A(n51), .B(n52), .C(n53), .D(n54), .Q(n50) );
  CLKIN3 U104 ( .A(n78), .Q(n36) );
endmodule


module E_alu_DW01_add_25 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97;

  CLKIN3 U2 ( .A(n65), .Q(n59) );
  CLKIN10 U3 ( .A(n44), .Q(n43) );
  NAND23 U4 ( .A(n65), .B(n8), .Q(n9) );
  NAND33 U5 ( .A(n69), .B(n70), .C(n71), .Q(n65) );
  NAND23 U6 ( .A(n1), .B(n21), .Q(n47) );
  NAND24 U7 ( .A(n11), .B(n77), .Q(n46) );
  CLKIN6 U8 ( .A(n33), .Q(n32) );
  CLKIN3 U9 ( .A(n47), .Q(n74) );
  NOR20 U10 ( .A(A[4]), .B(B[4]), .Q(n60) );
  CLKIN15 U11 ( .A(n22), .Q(n21) );
  INV8 U12 ( .A(A[3]), .Q(n22) );
  XNR22 U13 ( .A(n57), .B(n7), .Q(SUM[6]) );
  NAND23 U14 ( .A(B[4]), .B(A[4]), .Q(n28) );
  NAND26 U15 ( .A(n9), .B(n28), .Q(n53) );
  INV3 U16 ( .A(n43), .Q(n3) );
  INV3 U17 ( .A(n12), .Q(n13) );
  NAND22 U18 ( .A(n77), .B(n79), .Q(n12) );
  NOR23 U19 ( .A(n15), .B(n19), .Q(n80) );
  NOR22 U20 ( .A(n29), .B(n38), .Q(n37) );
  NAND22 U21 ( .A(n78), .B(n13), .Q(n70) );
  NAND22 U22 ( .A(B[0]), .B(A[0]), .Q(n76) );
  XOR21 U23 ( .A(n50), .B(n51), .Q(SUM[7]) );
  NOR22 U24 ( .A(B[4]), .B(A[4]), .Q(n38) );
  XOR20 U25 ( .A(n1), .B(n22), .Q(n85) );
  INV6 U26 ( .A(B[6]), .Q(n61) );
  NAND24 U27 ( .A(n43), .B(n5), .Q(n42) );
  NOR22 U28 ( .A(n82), .B(n83), .Q(n69) );
  NOR22 U29 ( .A(n27), .B(n39), .Q(n36) );
  INV4 U30 ( .A(A[1]), .Q(n20) );
  INV12 U31 ( .A(B[1]), .Q(n16) );
  CLKIN4 U32 ( .A(n18), .Q(n1) );
  INV12 U33 ( .A(B[3]), .Q(n18) );
  NOR23 U34 ( .A(n75), .B(n76), .Q(n73) );
  INV6 U35 ( .A(n31), .Q(n27) );
  INV3 U36 ( .A(n56), .Q(n7) );
  INV6 U37 ( .A(n20), .Q(n19) );
  XOR22 U38 ( .A(n85), .B(n86), .Q(SUM[3]) );
  INV2 U39 ( .A(n81), .Q(n78) );
  INV1 U40 ( .A(n48), .Q(n83) );
  XOR21 U41 ( .A(n63), .B(n64), .Q(SUM[5]) );
  AOI212 U42 ( .A(n65), .B(n8), .C(n66), .Q(n64) );
  INV4 U43 ( .A(n17), .Q(n10) );
  INV2 U44 ( .A(A[6]), .Q(n62) );
  OAI210 U45 ( .A(n27), .B(n55), .C(n33), .Q(n54) );
  NOR24 U46 ( .A(n49), .B(n44), .Q(n77) );
  BUF2 U47 ( .A(n31), .Q(n2) );
  INV6 U48 ( .A(n80), .Q(n79) );
  NAND24 U49 ( .A(n10), .B(n22), .Q(n11) );
  CLKIN6 U50 ( .A(n4), .Q(n5) );
  NAND24 U51 ( .A(n15), .B(n19), .Q(n4) );
  AOI2112 U52 ( .A(n10), .B(n22), .C(n84), .D(n3), .Q(n82) );
  NAND22 U53 ( .A(n15), .B(n19), .Q(n84) );
  NAND22 U54 ( .A(n43), .B(n45), .Q(n41) );
  NOR23 U55 ( .A(B[0]), .B(A[0]), .Q(n49) );
  INV2 U56 ( .A(n88), .Q(n6) );
  CLKIN1 U57 ( .A(n44), .Q(n88) );
  NOR21 U58 ( .A(B[7]), .B(A[7]), .Q(n39) );
  NAND28 U59 ( .A(n61), .B(n62), .Q(n31) );
  NAND21 U60 ( .A(n2), .B(n33), .Q(n56) );
  NAND23 U61 ( .A(B[6]), .B(A[6]), .Q(n33) );
  CLKIN15 U62 ( .A(n16), .Q(n15) );
  NAND22 U63 ( .A(n20), .B(n16), .Q(n45) );
  NOR23 U64 ( .A(n21), .B(n17), .Q(n75) );
  NOR23 U65 ( .A(A[5]), .B(B[5]), .Q(n29) );
  OAI212 U66 ( .A(A[7]), .B(B[7]), .C(n26), .Q(n24) );
  OAI312 U67 ( .A(n27), .B(n28), .C(n29), .D(n30), .Q(n26) );
  OAI2111 U68 ( .A(n21), .B(n1), .C(B[0]), .D(A[0]), .Q(n40) );
  CLKIN15 U69 ( .A(n18), .Q(n17) );
  AOI311 U70 ( .A(A[5]), .B(B[5]), .C(n31), .D(n32), .Q(n30) );
  OAI211 U71 ( .A(n15), .B(n19), .C(n93), .Q(n92) );
  NOR20 U72 ( .A(n89), .B(n6), .Q(n90) );
  AOI211 U73 ( .A(n20), .B(n16), .C(n44), .Q(n72) );
  OAI210 U74 ( .A(n15), .B(n19), .C(n84), .Q(n94) );
  AOI212 U75 ( .A(n87), .B(n88), .C(n89), .Q(n86) );
  INV1 U76 ( .A(n60), .Q(n8) );
  AOI312 U77 ( .A(n2), .B(n52), .C(n53), .D(n54), .Q(n51) );
  AOI212 U78 ( .A(n53), .B(n52), .C(n58), .Q(n57) );
  OAI2112 U79 ( .A(n21), .B(n17), .C(B[2]), .D(A[2]), .Q(n48) );
  NAND34 U80 ( .A(n23), .B(n24), .C(n25), .Q(SUM[8]) );
  OAI2112 U81 ( .A(n35), .B(n34), .C(n36), .D(n37), .Q(n23) );
  OAI2112 U82 ( .A(n80), .B(n46), .C(n47), .D(n48), .Q(n34) );
  INV3 U83 ( .A(n29), .Q(n52) );
  NOR24 U84 ( .A(A[2]), .B(B[2]), .Q(n44) );
  NAND21 U85 ( .A(n52), .B(n55), .Q(n63) );
  XOR20 U86 ( .A(n87), .B(n90), .Q(SUM[2]) );
  XNR20 U87 ( .A(n93), .B(n94), .Q(SUM[1]) );
  NOR20 U88 ( .A(n17), .B(n21), .Q(n81) );
  NAND22 U89 ( .A(n84), .B(n92), .Q(n87) );
  NAND20 U90 ( .A(B[5]), .B(A[5]), .Q(n55) );
  NAND22 U91 ( .A(n95), .B(n76), .Q(n93) );
  NOR20 U92 ( .A(A[0]), .B(B[0]), .Q(n95) );
  IMUX20 U93 ( .A(n67), .B(n68), .S(n59), .Q(SUM[4]) );
  NOR20 U94 ( .A(n38), .B(n66), .Q(n67) );
  NAND22 U95 ( .A(n96), .B(n76), .Q(SUM[0]) );
  NAND22 U96 ( .A(n14), .B(n97), .Q(n96) );
  INV0 U97 ( .A(A[0]), .Q(n14) );
  INV0 U98 ( .A(B[0]), .Q(n97) );
  XNR20 U99 ( .A(B[7]), .B(A[7]), .Q(n50) );
  NAND20 U100 ( .A(B[7]), .B(A[7]), .Q(n25) );
  NAND20 U101 ( .A(B[2]), .B(A[2]), .Q(n91) );
  XNR20 U102 ( .A(B[4]), .B(A[4]), .Q(n68) );
  OAI222 U103 ( .A(n40), .B(n41), .C(n42), .D(n75), .Q(n35) );
  CLKIN3 U104 ( .A(n55), .Q(n58) );
  AOI212 U105 ( .A(n72), .B(n73), .C(n74), .Q(n71) );
  CLKIN3 U106 ( .A(n28), .Q(n66) );
  CLKIN3 U107 ( .A(n91), .Q(n89) );
endmodule


module E_alu_DW01_add_26 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82;

  CLKIN1 U2 ( .A(n24), .Q(n61) );
  NOR24 U3 ( .A(A[2]), .B(B[2]), .Q(n41) );
  OAI2112 U4 ( .A(n17), .B(B[3]), .C(B[2]), .D(A[2]), .Q(n44) );
  INV6 U5 ( .A(n18), .Q(n17) );
  CLKIN4 U6 ( .A(B[6]), .Q(n56) );
  IMUX21 U7 ( .A(n62), .B(n63), .S(n54), .Q(SUM[4]) );
  NAND22 U8 ( .A(B[4]), .B(A[4]), .Q(n24) );
  NAND26 U9 ( .A(n56), .B(n57), .Q(n27) );
  INV12 U10 ( .A(B[3]), .Q(n14) );
  NAND24 U11 ( .A(n22), .B(n3), .Q(n20) );
  INV2 U12 ( .A(A[6]), .Q(n57) );
  NOR22 U13 ( .A(n25), .B(n34), .Q(n33) );
  NAND24 U14 ( .A(n64), .B(n65), .Q(n60) );
  NAND23 U15 ( .A(n11), .B(n15), .Q(n77) );
  NAND22 U16 ( .A(B[0]), .B(A[0]), .Q(n81) );
  INV3 U17 ( .A(n7), .Q(n43) );
  INV6 U18 ( .A(n4), .Q(n73) );
  NAND22 U19 ( .A(n1), .B(n2), .Q(n3) );
  INV0 U20 ( .A(A[7]), .Q(n1) );
  INV1 U21 ( .A(B[7]), .Q(n2) );
  NOR23 U22 ( .A(A[2]), .B(B[2]), .Q(n4) );
  NAND33 U23 ( .A(n40), .B(n15), .C(n11), .Q(n39) );
  CLKIN6 U24 ( .A(B[1]), .Q(n12) );
  NAND23 U25 ( .A(n9), .B(n24), .Q(n48) );
  NAND23 U26 ( .A(n60), .B(n8), .Q(n9) );
  XOR21 U27 ( .A(n51), .B(n52), .Q(SUM[6]) );
  INV3 U28 ( .A(n60), .Q(n54) );
  NOR22 U29 ( .A(n23), .B(n35), .Q(n32) );
  NOR22 U30 ( .A(n68), .B(n69), .Q(n64) );
  XOR21 U31 ( .A(n45), .B(n46), .Q(SUM[7]) );
  NAND24 U32 ( .A(n42), .B(n73), .Q(n37) );
  NOR22 U33 ( .A(B[4]), .B(A[4]), .Q(n34) );
  CLKIN6 U34 ( .A(A[3]), .Q(n18) );
  INV2 U35 ( .A(n44), .Q(n69) );
  INV12 U36 ( .A(n14), .Q(n13) );
  INV3 U37 ( .A(n29), .Q(n28) );
  INV3 U38 ( .A(n25), .Q(n47) );
  BUF2 U39 ( .A(n29), .Q(n5) );
  INV0 U40 ( .A(n23), .Q(n6) );
  INV8 U41 ( .A(n27), .Q(n23) );
  INV2 U42 ( .A(n76), .Q(n74) );
  NOR24 U43 ( .A(n18), .B(n14), .Q(n7) );
  NOR23 U44 ( .A(A[5]), .B(B[5]), .Q(n25) );
  AOI210 U45 ( .A(n16), .B(n12), .C(n41), .Q(n66) );
  CLKIN6 U46 ( .A(n41), .Q(n40) );
  NAND22 U47 ( .A(n47), .B(n50), .Q(n58) );
  INV3 U48 ( .A(A[1]), .Q(n16) );
  AOI311 U49 ( .A(A[5]), .B(B[5]), .C(n27), .D(n28), .Q(n26) );
  NAND22 U50 ( .A(n44), .B(n43), .Q(n30) );
  NOR22 U51 ( .A(n38), .B(n81), .Q(n67) );
  OAI2111 U52 ( .A(B[3]), .B(n17), .C(B[0]), .D(A[0]), .Q(n36) );
  OAI210 U53 ( .A(n23), .B(n50), .C(n5), .Q(n49) );
  XOR21 U54 ( .A(n70), .B(n71), .Q(SUM[3]) );
  NAND21 U55 ( .A(B[7]), .B(A[7]), .Q(n21) );
  NOR20 U56 ( .A(A[4]), .B(B[4]), .Q(n55) );
  NOR22 U57 ( .A(B[7]), .B(A[7]), .Q(n35) );
  NOR24 U58 ( .A(n17), .B(n13), .Q(n38) );
  AOI212 U59 ( .A(n8), .B(n60), .C(n61), .Q(n59) );
  XOR22 U60 ( .A(n58), .B(n59), .Q(SUM[5]) );
  AOI2111 U61 ( .A(n14), .B(n18), .C(n77), .D(n41), .Q(n68) );
  OAI210 U62 ( .A(n11), .B(n15), .C(n77), .Q(n80) );
  NAND21 U63 ( .A(n12), .B(n16), .Q(n42) );
  INV2 U64 ( .A(n55), .Q(n8) );
  AOI312 U65 ( .A(n6), .B(n47), .C(n48), .D(n49), .Q(n46) );
  AOI212 U66 ( .A(n48), .B(n47), .C(n53), .Q(n52) );
  NAND34 U67 ( .A(n19), .B(n20), .C(n21), .Q(SUM[8]) );
  OAI2112 U68 ( .A(n30), .B(n31), .C(n32), .D(n33), .Q(n19) );
  CLKIN6 U69 ( .A(n12), .Q(n11) );
  NAND20 U70 ( .A(n27), .B(n5), .Q(n51) );
  XNR20 U71 ( .A(n13), .B(n17), .Q(n70) );
  AOI211 U72 ( .A(n72), .B(n73), .C(n74), .Q(n71) );
  XNR20 U73 ( .A(n79), .B(n80), .Q(SUM[1]) );
  INV3 U74 ( .A(n16), .Q(n15) );
  NAND22 U75 ( .A(n77), .B(n78), .Q(n72) );
  NOR20 U76 ( .A(n34), .B(n61), .Q(n62) );
  MUX21 U77 ( .A(B[0]), .B(n82), .S(A[0]), .Q(SUM[0]) );
  XOR21 U78 ( .A(n72), .B(n75), .Q(SUM[2]) );
  NAND20 U79 ( .A(B[5]), .B(A[5]), .Q(n50) );
  INV2 U80 ( .A(n81), .Q(n79) );
  INV0 U81 ( .A(B[0]), .Q(n82) );
  NAND22 U82 ( .A(B[6]), .B(A[6]), .Q(n29) );
  XNR20 U83 ( .A(B[7]), .B(A[7]), .Q(n45) );
  NOR20 U84 ( .A(n74), .B(n4), .Q(n75) );
  NAND20 U85 ( .A(B[2]), .B(A[2]), .Q(n76) );
  XNR20 U86 ( .A(B[4]), .B(A[4]), .Q(n63) );
  OAI312 U87 ( .A(n23), .B(n24), .C(n25), .D(n26), .Q(n22) );
  OAI222 U88 ( .A(n37), .B(n36), .C(n39), .D(n38), .Q(n31) );
  CLKIN3 U89 ( .A(n50), .Q(n53) );
  AOI212 U90 ( .A(n66), .B(n67), .C(n7), .Q(n65) );
  OAI212 U91 ( .A(n11), .B(n15), .C(n79), .Q(n78) );
endmodule


module E_alu ( o_data_AluRes, i_data_A, i_data_B, i_con_AluCtrl, i_data_shamt
 );
  output [31:0] o_data_AluRes;
  input [31:0] i_data_A;
  input [31:0] i_data_B;
  input [3:0] i_con_AluCtrl;
  input [4:0] i_data_shamt;
  wire   N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N306, n41, n42,
         n161, n169, n176, n183, n190, n198, n221, n333, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n162, n163, n164, n165, n166, n167, n168, n170, n171, n172, n173,
         n174, n175, n177, n178, n179, n180, n181, n182, n184, n185, n186,
         n187, n188, n189, n191, n192, n193, n194, n195, n196, n197, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536;
  wire   [8:0] sum_1;
  wire   [8:0] pre_sum_2a;
  wire   [8:0] pre_sum_2b;
  wire   [8:0] pre_sum_3a;
  wire   [8:0] pre_sum_3b;
  wire   [7:0] pre_sum_4a;
  wire   [7:0] pre_sum_4b;
  wire   [16:0] half_sub;
  wire   [15:0] pre_suba;
  wire   [15:0] pre_subb;

  E_alu_DW01_add_12 add_1_root_add_31_2 ( .A({n128, i_data_A[30:28], n166, 
        n164, i_data_A[25], n162}), .B({n126, n124, n123, n156, n7, n21, n120, 
        n100}), .CI(n41), .SUM(pre_sum_4b) );
  E_alu_DW01_add_13 add_30 ( .A({n128, i_data_A[30:28], n166, n164, 
        i_data_A[25], n162}), .B({n126, n124, n123, n156, n6, n21, n120, n101}), .CI(n42), .SUM(pre_sum_4a) );
  E_alu_DW01_ash_1 sll_56 ( .A({n125, n124, n122, n156, n7, n21, n120, n100, 
        n4, n118, n117, n97, n50, n22, n114, n153, n84, n111, n11, n151, n20, 
        n109, n147, n19, i_data_B[7:1], n143}), .DATA_TC(n42), .SH(
        i_data_shamt), .SH_TC(n42), .B({N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, 
        N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193}) );
  E_alu_DW01_sub_7 sub_1_root_sub_35_2 ( .A({n127, i_data_A[30:28], n166, n164, 
        i_data_A[25], n162, i_data_A[23:21], n159, i_data_A[19:17], n157}), 
        .B({n126, n124, n122, n156, n6, n103, n121, i_data_B[24], n99, n119, 
        n116, n96, n49, n154, n115, n153}), .CI(n41), .DIFF(pre_subb) );
  E_alu_DW_rash_3 r130 ( .A({n125, n124, n123, n156, n7, n103, n121, n101, n99, 
        n118, n117, n96, n49, n22, n85, n153, n113, n111, n11, n151, n20, n109, 
        n13, n19, i_data_B[7:6], n15, i_data_B[4], n34, n18, n36, n143}), 
        .DATA_TC(n42), .SH(i_data_shamt), .SH_TC(n42), .B({N256, N255, N254, 
        N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, 
        N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, 
        N229, N228, N227, N226, N225}) );
  E_alu_DW01_add_23 add_28 ( .A({n42, i_data_A[23:21], n159, i_data_A[19:17], 
        n157}), .B({n42, i_data_B[23], n118, n116, n96, n49, n22, n85, n153}), 
        .CI(n42), .SUM(pre_sum_3a) );
  E_alu_DW01_sub_10 sub_33 ( .A({n42, i_data_A[15:0]}), .B({n42, n113, n112, 
        n110, n151, n149, n108, n147, n145, i_data_B[7:1], n143}), .CI(n42), 
        .DIFF(half_sub) );
  E_alu_DW01_cmp2_4 r131 ( .A({n127, i_data_A[30:28], n166, n164, i_data_A[25], 
        n162, i_data_A[23:21], n159, i_data_A[19:17], n157, i_data_A[15:10], 
        n31, i_data_A[8:0]}), .B({n126, n124, n123, n156, n7, n103, n121, n102, 
        n99, n118, n117, n97, n50, n22, n114, n153, n84, n112, n110, n151, n20, 
        n109, n13, n19, i_data_B[7:4], n34, i_data_B[2], n36, n143}), .LEQ(n42), .TC(n42), .LT_LE(N306) );
  E_alu_DW01_sub_13 sub_34 ( .A({n127, i_data_A[30:28], n166, n164, 
        i_data_A[25], n162, i_data_A[23:21], n159, i_data_A[19:17], n157}), 
        .B({n126, n124, n122, n156, n6, n103, n121, n102, n155, n119, n116, 
        n96, n50, n154, n114, n153}), .CI(n42), .DIFF(pre_suba) );
  E_alu_DW01_add_27 add_1_root_add_29_2 ( .A({n42, i_data_A[23:21], n159, 
        i_data_A[19:17], n157}), .B({n42, n4, n119, n117, n96, n50, n154, n85, 
        n153}), .CI(n41), .SUM(pre_sum_3b) );
  E_alu_DW01_add_24 add_25 ( .A({n42, i_data_A[7:0]}), .B({n42, i_data_B[7:1], 
        n143}), .CI(n42), .SUM(sum_1) );
  E_alu_DW01_add_25 add_1_root_add_27_2 ( .A({n42, i_data_A[15:8]}), .B({n42, 
        n84, n111, n11, n151, n149, n108, n147, n145}), .CI(n41), .SUM(
        pre_sum_2b) );
  E_alu_DW01_add_26 add_26 ( .A({n42, i_data_A[15:8]}), .B({n42, n84, n112, 
        n11, n151, n20, n109, n147, n19}), .CI(n42), .SUM(pre_sum_2a) );
  INV4 U3 ( .A(n179), .Q(n24) );
  NAND43 U4 ( .A(n308), .B(n309), .C(n307), .D(n306), .Q(o_data_AluRes[15]) );
  OAI2110 U5 ( .A(i_data_A[5]), .B(n139), .C(n133), .D(n176), .Q(n220) );
  INV2 U6 ( .A(i_data_B[5]), .Q(n386) );
  AOI212 U7 ( .A(n136), .B(n393), .C(n129), .Q(n394) );
  CLKIN12 U8 ( .A(n320), .Q(n414) );
  INV12 U9 ( .A(n531), .Q(n39) );
  NAND24 U10 ( .A(n269), .B(n83), .Q(o_data_AluRes[11]) );
  CLKIN4 U11 ( .A(n180), .Q(n1) );
  INV10 U12 ( .A(i_con_AluCtrl[1]), .Q(n180) );
  CLKIN4 U13 ( .A(n320), .Q(n8) );
  BUF12 U14 ( .A(i_data_B[21]), .Q(n117) );
  INV15 U15 ( .A(n152), .Q(n151) );
  CLKBU15 U16 ( .A(i_data_B[17]), .Q(n85) );
  NAND22 U17 ( .A(n517), .B(n393), .Q(n395) );
  CLKIN12 U18 ( .A(n150), .Q(n20) );
  BUF2 U19 ( .A(i_data_B[7]), .Q(n2) );
  NAND24 U20 ( .A(n366), .B(n367), .Q(n71) );
  CLKIN0 U21 ( .A(n84), .Q(n521) );
  BUF8 U22 ( .A(i_data_B[26]), .Q(n21) );
  INV3 U23 ( .A(n139), .Q(n37) );
  CLKIN10 U24 ( .A(n155), .Q(n3) );
  INV12 U25 ( .A(n3), .Q(n4) );
  CLKIN6 U26 ( .A(n93), .Q(n94) );
  INV10 U27 ( .A(i_data_A[20]), .Q(n160) );
  NAND23 U28 ( .A(i_con_AluCtrl[0]), .B(n91), .Q(n77) );
  IMUX22 U29 ( .A(n334), .B(n332), .S(n85), .Q(n339) );
  AOI211 U30 ( .A(n136), .B(n344), .C(n129), .Q(n345) );
  INV10 U31 ( .A(i_data_B[11]), .Q(n150) );
  AOI2111 U32 ( .A(i_data_A[28]), .B(n486), .C(n484), .D(n485), .Q(n490) );
  NAND24 U33 ( .A(n270), .B(n268), .Q(n65) );
  OAI212 U34 ( .A(n107), .B(n51), .C(n465), .Q(n468) );
  AOI2112 U35 ( .A(N246), .B(n141), .C(n388), .D(n387), .Q(n392) );
  CLKIN10 U36 ( .A(n474), .Q(n55) );
  IMUX22 U37 ( .A(n383), .B(n382), .S(n117), .Q(n388) );
  NAND23 U38 ( .A(half_sub[15]), .B(n325), .Q(n307) );
  AOI211 U39 ( .A(n136), .B(n290), .C(n129), .Q(n288) );
  CLKIN15 U40 ( .A(n137), .Q(n136) );
  AOI222 U41 ( .A(N200), .B(n81), .C(sum_1[7]), .D(n471), .Q(n235) );
  BUF15 U42 ( .A(i_data_B[24]), .Q(n101) );
  INV6 U43 ( .A(n86), .Q(n87) );
  NAND22 U44 ( .A(n530), .B(pre_suba[9]), .Q(n446) );
  CLKIN4 U45 ( .A(half_sub[16]), .Q(n323) );
  INV15 U46 ( .A(n167), .Q(n166) );
  CLKIN6 U47 ( .A(i_data_A[27]), .Q(n167) );
  NAND23 U48 ( .A(half_sub[7]), .B(n325), .Q(n234) );
  NAND32 U49 ( .A(n180), .B(n313), .C(n179), .Q(n503) );
  BUF12 U50 ( .A(i_data_B[31]), .Q(n125) );
  NAND33 U51 ( .A(n314), .B(n91), .C(n45), .Q(n462) );
  BUF6 U52 ( .A(n527), .Q(n141) );
  INV12 U53 ( .A(n92), .Q(n325) );
  BUF6 U54 ( .A(n175), .Q(n92) );
  INV12 U55 ( .A(n165), .Q(n164) );
  INV6 U56 ( .A(i_con_AluCtrl[3]), .Q(n179) );
  CLKBU12 U57 ( .A(n503), .Q(n104) );
  INV3 U58 ( .A(i_data_A[24]), .Q(n163) );
  BUF6 U59 ( .A(i_data_B[31]), .Q(n126) );
  CLKIN8 U60 ( .A(n12), .Q(n13) );
  BUF6 U61 ( .A(n312), .Q(n45) );
  NAND23 U62 ( .A(n343), .B(n342), .Q(n67) );
  AOI221 U63 ( .A(N194), .B(n81), .C(N226), .D(n141), .Q(n204) );
  INV12 U64 ( .A(n163), .Q(n162) );
  INV3 U65 ( .A(n73), .Q(n74) );
  AOI221 U66 ( .A(pre_sum_2b[6]), .B(n305), .C(N207), .D(n81), .Q(n297) );
  CLKIN15 U67 ( .A(n144), .Q(n143) );
  CLKIN15 U68 ( .A(n90), .Q(n91) );
  CLKIN6 U69 ( .A(n326), .Q(n14) );
  INV12 U70 ( .A(n324), .Q(n530) );
  CLKIN12 U71 ( .A(n326), .Q(n531) );
  BUF8 U72 ( .A(i_data_B[17]), .Q(n114) );
  BUF6 U73 ( .A(i_data_B[17]), .Q(n115) );
  BUF8 U74 ( .A(i_data_B[24]), .Q(n100) );
  INV12 U75 ( .A(i_data_B[8]), .Q(n146) );
  NAND24 U76 ( .A(n377), .B(n376), .Q(n93) );
  INV12 U77 ( .A(n150), .Q(n149) );
  CLKIN15 U78 ( .A(n241), .Q(n305) );
  BUF12 U79 ( .A(i_data_B[10]), .Q(n109) );
  INV10 U80 ( .A(i_data_B[0]), .Q(n144) );
  CLKIN6 U81 ( .A(n433), .Q(n5) );
  NAND23 U82 ( .A(half_sub[14]), .B(n325), .Q(n296) );
  CLKIN4 U83 ( .A(sum_1[8]), .Q(n431) );
  NAND23 U84 ( .A(n430), .B(pre_sum_3b[8]), .Q(n470) );
  INV10 U85 ( .A(n433), .Q(n529) );
  AOI222 U86 ( .A(N202), .B(n81), .C(half_sub[9]), .D(n325), .Q(n253) );
  BUF12 U87 ( .A(i_data_B[13]), .Q(n110) );
  CLKBU4 U88 ( .A(i_data_B[2]), .Q(n18) );
  BUF6 U89 ( .A(i_data_B[1]), .Q(n36) );
  NAND32 U90 ( .A(n402), .B(n401), .C(n64), .Q(o_data_AluRes[22]) );
  OAI211 U91 ( .A(n129), .B(n384), .C(i_data_A[21]), .Q(n385) );
  OAI212 U92 ( .A(n106), .B(n349), .C(n348), .Q(n350) );
  OAI211 U93 ( .A(n129), .B(n335), .C(i_data_A[17]), .Q(n336) );
  AOI2112 U94 ( .A(N240), .B(n141), .C(n303), .D(n302), .Q(n309) );
  AOI211 U95 ( .A(n301), .B(n132), .C(n300), .Q(n302) );
  AOI221 U96 ( .A(n531), .B(pre_subb[8]), .C(pre_suba[8]), .D(n25), .Q(n434)
         );
  NAND21 U97 ( .A(pre_subb[9]), .B(n531), .Q(n447) );
  CLKBU4 U98 ( .A(n462), .Q(n26) );
  NAND24 U99 ( .A(half_sub[16]), .B(n325), .Q(n326) );
  AOI2112 U100 ( .A(N256), .B(n141), .C(n526), .D(n525), .Q(n535) );
  BUF12 U101 ( .A(i_data_B[13]), .Q(n11) );
  NAND24 U102 ( .A(n528), .B(pre_sum_4b[7]), .Q(n534) );
  CLKIN6 U103 ( .A(n474), .Q(n528) );
  NAND34 U104 ( .A(n532), .B(n534), .C(n535), .Q(n86) );
  XNR21 U105 ( .A(n126), .B(n128), .Q(n524) );
  INV3 U106 ( .A(n88), .Q(n79) );
  NAND24 U107 ( .A(n60), .B(n471), .Q(n241) );
  BUF12 U108 ( .A(n523), .Q(n137) );
  NAND22 U109 ( .A(N193), .B(n80), .Q(n186) );
  BUF12 U110 ( .A(i_data_B[3]), .Q(n34) );
  INV12 U111 ( .A(n137), .Q(n135) );
  INV12 U112 ( .A(n462), .Q(n517) );
  BUF6 U113 ( .A(n527), .Q(n142) );
  INV6 U114 ( .A(n174), .Q(n471) );
  INV6 U115 ( .A(n168), .Q(n314) );
  NAND22 U116 ( .A(i_con_AluCtrl[3]), .B(n180), .Q(n168) );
  NOR21 U117 ( .A(n126), .B(n128), .Q(n516) );
  BUF6 U118 ( .A(n503), .Q(n105) );
  BUF2 U119 ( .A(i_data_A[31]), .Q(n128) );
  INV6 U120 ( .A(i_data_A[26]), .Q(n165) );
  NAND23 U121 ( .A(n404), .B(n403), .Q(n63) );
  NAND24 U122 ( .A(N215), .B(n80), .Q(n403) );
  NAND22 U123 ( .A(N211), .B(n80), .Q(n354) );
  NAND23 U124 ( .A(n330), .B(n329), .Q(n73) );
  NAND22 U125 ( .A(N209), .B(n81), .Q(n329) );
  NAND23 U126 ( .A(N213), .B(n80), .Q(n375) );
  NOR22 U127 ( .A(n38), .B(n39), .Q(n40) );
  INV3 U128 ( .A(pre_subb[4]), .Q(n38) );
  NAND23 U129 ( .A(N306), .B(n196), .Q(n197) );
  AOI2111 U130 ( .A(N254), .B(n141), .C(n498), .D(n497), .Q(n502) );
  NAND22 U131 ( .A(pre_sum_2a[6]), .B(n304), .Q(n294) );
  NAND22 U132 ( .A(half_sub[2]), .B(n325), .Q(n208) );
  AOI221 U133 ( .A(N196), .B(n80), .C(N228), .D(n141), .Q(n214) );
  AOI221 U134 ( .A(pre_sum_2b[4]), .B(n305), .C(N237), .D(n141), .Q(n278) );
  NAND23 U135 ( .A(n1), .B(n179), .Q(n173) );
  OAI211 U136 ( .A(n130), .B(n315), .C(n157), .Q(n316) );
  AOI221 U137 ( .A(sum_1[3]), .B(n471), .C(i_data_A[3]), .D(n130), .Q(n212) );
  NAND22 U138 ( .A(n199), .B(n197), .Q(o_data_AluRes[0]) );
  BUF15 U139 ( .A(i_data_B[10]), .Q(n108) );
  AOI222 U140 ( .A(pre_suba[5]), .B(n25), .C(pre_subb[5]), .D(n14), .Q(n389)
         );
  BUF15 U141 ( .A(i_data_B[27]), .Q(n6) );
  BUF15 U142 ( .A(i_data_B[27]), .Q(n7) );
  OAI212 U143 ( .A(n107), .B(n152), .C(n480), .Q(n485) );
  BUF6 U144 ( .A(i_data_B[20]), .Q(n97) );
  INV12 U145 ( .A(n79), .Q(n80) );
  NAND26 U146 ( .A(n314), .B(n78), .Q(n523) );
  CLKBU12 U147 ( .A(i_data_B[29]), .Q(n122) );
  BUF12 U148 ( .A(i_data_B[14]), .Q(n111) );
  CLKIN6 U149 ( .A(n322), .Q(n413) );
  NAND20 U150 ( .A(n517), .B(n344), .Q(n346) );
  CLKIN0 U151 ( .A(i_data_A[19]), .Q(n356) );
  AOI221 U152 ( .A(n530), .B(pre_suba[3]), .C(pre_subb[3]), .D(n14), .Q(n364)
         );
  NAND32 U153 ( .A(n365), .B(n364), .C(n72), .Q(o_data_AluRes[19]) );
  AOI221 U154 ( .A(n8), .B(pre_sum_3b[3]), .C(pre_sum_3a[3]), .D(n53), .Q(n365) );
  CLKIN12 U155 ( .A(n428), .Q(n46) );
  NAND20 U156 ( .A(i_data_A[6]), .B(n536), .Q(n169) );
  INV0 U157 ( .A(n19), .Q(n9) );
  INV3 U158 ( .A(n9), .Q(n10) );
  INV12 U159 ( .A(n146), .Q(n19) );
  OAI210 U160 ( .A(i_data_A[11]), .B(n138), .C(n133), .Q(n266) );
  CLKIN15 U161 ( .A(n160), .Q(n159) );
  CLKBU8 U162 ( .A(n134), .Q(n133) );
  INV6 U163 ( .A(i_data_B[9]), .Q(n148) );
  CLKIN0 U164 ( .A(i_data_A[14]), .Q(n290) );
  NAND20 U165 ( .A(i_data_A[7]), .B(n536), .Q(n161) );
  OAI2110 U166 ( .A(i_data_A[7]), .B(n139), .C(n133), .D(n161), .Q(n233) );
  AOI220 U167 ( .A(sum_1[0]), .B(n471), .C(half_sub[0]), .D(n325), .Q(n177) );
  OAI211 U168 ( .A(n106), .B(n144), .C(n316), .Q(n317) );
  INV6 U169 ( .A(n147), .Q(n12) );
  INV12 U170 ( .A(pre_sum_2a[8]), .Q(n429) );
  OAI2111 U171 ( .A(i_data_A[3]), .B(n139), .C(n133), .D(n190), .Q(n210) );
  NAND20 U172 ( .A(i_data_A[3]), .B(n536), .Q(n190) );
  NAND20 U173 ( .A(n517), .B(n170), .Q(n172) );
  BUF15 U174 ( .A(i_data_B[15]), .Q(n113) );
  AOI221 U175 ( .A(N197), .B(n80), .C(N229), .D(n142), .Q(n219) );
  NAND22 U176 ( .A(n369), .B(n132), .Q(n373) );
  NAND22 U177 ( .A(n392), .B(n391), .Q(n75) );
  NAND23 U178 ( .A(N214), .B(n81), .Q(n391) );
  INV3 U179 ( .A(n75), .Q(n76) );
  IMUX21 U180 ( .A(n138), .B(n105), .S(n123), .Q(n491) );
  NAND23 U181 ( .A(N249), .B(n142), .Q(n420) );
  BUF15 U182 ( .A(i_data_B[22]), .Q(n118) );
  CLKIN6 U183 ( .A(n386), .Q(n15) );
  BUF2 U184 ( .A(n118), .Q(n16) );
  CLKIN0 U185 ( .A(i_data_A[30]), .Q(n507) );
  NAND32 U186 ( .A(n328), .B(n327), .C(n74), .Q(o_data_AluRes[16]) );
  AOI221 U187 ( .A(pre_sum_3b[0]), .B(n8), .C(pre_sum_3a[0]), .D(n53), .Q(n328) );
  BUF2 U188 ( .A(n13), .Q(n17) );
  IMUX30 U189 ( .A(n517), .B(n135), .C(n215), .S0(i_data_A[4]), .S1(n32), .Q(
        n216) );
  IMUX20 U190 ( .A(n135), .B(n536), .S(n100), .Q(n419) );
  CLKIN0 U191 ( .A(n18), .Q(n349) );
  IMUX21 U192 ( .A(n138), .B(n104), .S(n22), .Q(n347) );
  CLKIN0 U193 ( .A(n111), .Q(n506) );
  INV8 U194 ( .A(i_data_A[16]), .Q(n158) );
  CLKIN0 U195 ( .A(n153), .Q(n47) );
  NAND22 U196 ( .A(half_sub[4]), .B(n325), .Q(n218) );
  BUF15 U197 ( .A(i_data_B[19]), .Q(n50) );
  OAI212 U198 ( .A(n106), .B(n398), .C(n397), .Q(n399) );
  AOI2112 U199 ( .A(N241), .B(n141), .C(n318), .D(n317), .Q(n330) );
  AOI221 U200 ( .A(sum_1[5]), .B(n471), .C(i_data_A[5]), .D(n130), .Q(n223) );
  CLKIN0 U201 ( .A(n126), .Q(n520) );
  IMUX20 U202 ( .A(n464), .B(n463), .S(n7), .Q(n465) );
  NAND23 U203 ( .A(N221), .B(n80), .Q(n489) );
  NAND26 U204 ( .A(N225), .B(n142), .Q(n182) );
  BUF8 U205 ( .A(n523), .Q(n139) );
  NAND22 U206 ( .A(n517), .B(n160), .Q(n371) );
  NAND24 U207 ( .A(N210), .B(n81), .Q(n342) );
  CLKBU12 U208 ( .A(n523), .Q(n138) );
  INV12 U209 ( .A(n59), .Q(n60) );
  AOI222 U210 ( .A(N204), .B(n80), .C(half_sub[11]), .D(n325), .Q(n269) );
  CLKIN6 U211 ( .A(n91), .Q(n313) );
  NAND21 U212 ( .A(i_data_A[5]), .B(n536), .Q(n176) );
  INV12 U213 ( .A(n324), .Q(n25) );
  CLKIN0 U214 ( .A(n2), .Q(n407) );
  OAI211 U215 ( .A(n106), .B(n386), .C(n385), .Q(n387) );
  NAND20 U216 ( .A(n517), .B(n165), .Q(n454) );
  BUF15 U217 ( .A(i_data_B[18]), .Q(n22) );
  AOI222 U218 ( .A(n25), .B(pre_suba[0]), .C(pre_subb[0]), .D(n14), .Q(n327)
         );
  BUF6 U219 ( .A(i_data_B[25]), .Q(n120) );
  BUF2 U220 ( .A(n194), .Q(n23) );
  CLKIN4 U221 ( .A(n322), .Q(n53) );
  CLKIN4 U222 ( .A(n71), .Q(n72) );
  CLKIN15 U223 ( .A(n98), .Q(n99) );
  IMUX21 U224 ( .A(n138), .B(n105), .S(n50), .Q(n359) );
  NAND31 U225 ( .A(n91), .B(n185), .C(n45), .Q(n175) );
  NAND28 U226 ( .A(n323), .B(n325), .Q(n324) );
  IMUX20 U227 ( .A(n138), .B(n105), .S(n99), .Q(n405) );
  INV15 U228 ( .A(n39), .Q(n27) );
  INV6 U229 ( .A(n518), .Q(n134) );
  OAI2111 U230 ( .A(i_data_A[1]), .B(n139), .C(n133), .D(n333), .Q(n200) );
  INV12 U231 ( .A(n429), .Q(n48) );
  NAND22 U232 ( .A(n517), .B(n439), .Q(n441) );
  IMUX20 U233 ( .A(n136), .B(n536), .S(n156), .Q(n479) );
  IMUX22 U234 ( .A(n371), .B(n370), .S(n97), .Q(n372) );
  NAND21 U235 ( .A(n517), .B(n163), .Q(n422) );
  NAND22 U236 ( .A(N219), .B(n81), .Q(n460) );
  INV15 U237 ( .A(n148), .Q(n147) );
  CLKIN6 U238 ( .A(pre_sum_3a[8]), .Q(n28) );
  INV6 U239 ( .A(n28), .Q(n29) );
  CLKIN0 U240 ( .A(n11), .Q(n493) );
  IMUX21 U241 ( .A(n283), .B(n282), .S(n110), .Q(n284) );
  AOI211 U242 ( .A(n136), .B(n331), .C(n129), .Q(n332) );
  NAND34 U243 ( .A(n374), .B(n375), .C(n94), .Q(n378) );
  INV1 U244 ( .A(i_data_A[9]), .Q(n30) );
  INV3 U245 ( .A(n30), .Q(n31) );
  OAI2111 U246 ( .A(i_data_A[2]), .B(n140), .C(n133), .D(n221), .Q(n205) );
  IMUX20 U247 ( .A(n137), .B(n104), .S(n143), .Q(n178) );
  BUF2 U248 ( .A(i_data_B[4]), .Q(n32) );
  AOI221 U249 ( .A(n530), .B(pre_suba[7]), .C(pre_subb[7]), .D(n14), .Q(n415)
         );
  IMUX21 U250 ( .A(n129), .B(n517), .S(n516), .Q(n519) );
  IMUX23 U251 ( .A(n441), .B(n440), .S(n120), .Q(n442) );
  AOI2112 U252 ( .A(n141), .B(N247), .C(n400), .D(n399), .Q(n404) );
  AOI222 U253 ( .A(pre_sum_2b[7]), .B(n305), .C(pre_sum_2a[7]), .D(n304), .Q(
        n306) );
  BUF6 U254 ( .A(n522), .Q(n107) );
  BUF6 U255 ( .A(n522), .Q(n106) );
  INV6 U256 ( .A(n61), .Q(n62) );
  INV12 U257 ( .A(n155), .Q(n98) );
  NAND24 U258 ( .A(n432), .B(n29), .Q(n469) );
  IMUX21 U259 ( .A(n140), .B(n105), .S(n117), .Q(n384) );
  INV3 U260 ( .A(n45), .Q(n33) );
  BUF4 U261 ( .A(n134), .Q(n132) );
  BUF2 U262 ( .A(n20), .Q(n35) );
  IMUX20 U263 ( .A(n140), .B(n105), .S(n120), .Q(n438) );
  NAND33 U264 ( .A(n285), .B(n287), .C(n62), .Q(o_data_AluRes[13]) );
  AOI222 U265 ( .A(N206), .B(n80), .C(half_sub[13]), .D(n325), .Q(n285) );
  NOR24 U266 ( .A(n40), .B(n378), .Q(n380) );
  NAND21 U267 ( .A(n33), .B(n185), .Q(n193) );
  INV6 U268 ( .A(n173), .Q(n185) );
  OAI212 U269 ( .A(n106), .B(n361), .C(n360), .Q(n362) );
  INV4 U270 ( .A(n82), .Q(n83) );
  MUX21 U271 ( .A(n517), .B(n136), .S(i_data_A[6]), .Q(n43) );
  IMUX21 U272 ( .A(n43), .B(n226), .S(n44), .Q(n227) );
  AOI222 U273 ( .A(N203), .B(n81), .C(half_sub[10]), .D(n325), .Q(n261) );
  NAND21 U274 ( .A(n536), .B(n128), .Q(n198) );
  BUF2 U275 ( .A(i_data_B[6]), .Q(n44) );
  IMUX20 U276 ( .A(n135), .B(n536), .S(n52), .Q(n256) );
  AOI211 U277 ( .A(n136), .B(n158), .C(n129), .Q(n310) );
  AOI2112 U278 ( .A(N243), .B(n141), .C(n350), .D(n351), .Q(n355) );
  BUF15 U279 ( .A(i_data_B[20]), .Q(n96) );
  INV12 U280 ( .A(pre_sum_2b[8]), .Q(n428) );
  INV2 U281 ( .A(n181), .Q(n527) );
  INV6 U282 ( .A(i_con_AluCtrl[0]), .Q(n312) );
  IMUX21 U283 ( .A(n454), .B(n453), .S(n21), .Q(n455) );
  AOI211 U284 ( .A(n136), .B(n381), .C(n129), .Q(n382) );
  IMUX21 U285 ( .A(n136), .B(n536), .S(n97), .Q(n369) );
  AOI2112 U286 ( .A(N242), .B(n141), .C(n339), .D(n338), .Q(n343) );
  IMUX21 U287 ( .A(n310), .B(n311), .S(n47), .Q(n318) );
  AOI2112 U288 ( .A(N252), .B(n141), .C(n468), .D(n467), .Q(n478) );
  OAI210 U289 ( .A(i_data_A[13]), .B(n138), .C(n133), .Q(n282) );
  BUF15 U290 ( .A(i_data_B[19]), .Q(n49) );
  NAND32 U291 ( .A(n185), .B(n313), .C(n45), .Q(n174) );
  NAND31 U292 ( .A(n314), .B(n313), .C(n45), .Q(n522) );
  OAI220 U293 ( .A(n195), .B(n23), .C(n313), .D(n193), .Q(n196) );
  AOI222 U294 ( .A(n414), .B(pre_sum_3b[7]), .C(pre_sum_3a[7]), .D(n53), .Q(
        n416) );
  INV0 U295 ( .A(n35), .Q(n51) );
  CLKBU12 U296 ( .A(i_data_B[15]), .Q(n84) );
  IMUX22 U297 ( .A(n358), .B(n357), .S(n50), .Q(n363) );
  AOI211 U298 ( .A(n136), .B(n356), .C(n129), .Q(n357) );
  OAI210 U299 ( .A(n130), .B(n178), .C(i_data_A[0]), .Q(n184) );
  CLKBU15 U300 ( .A(n134), .Q(n131) );
  INV6 U301 ( .A(n65), .Q(n66) );
  AOI221 U302 ( .A(i_data_A[11]), .B(n265), .C(pre_sum_2a[3]), .D(n304), .Q(
        n271) );
  CLKIN12 U303 ( .A(n239), .Q(n304) );
  OAI312 U304 ( .A(n23), .B(n524), .C(n187), .D(n186), .Q(n188) );
  AOI221 U305 ( .A(n414), .B(pre_sum_3b[1]), .C(n413), .D(pre_sum_3a[1]), .Q(
        n341) );
  AOI221 U306 ( .A(pre_sum_3b[2]), .B(n8), .C(pre_sum_3a[2]), .D(n53), .Q(n353) );
  IMUX20 U307 ( .A(n135), .B(n536), .S(n10), .Q(n238) );
  NAND20 U308 ( .A(n248), .B(n133), .Q(n249) );
  BUF2 U309 ( .A(n109), .Q(n52) );
  AOI222 U310 ( .A(N205), .B(n80), .C(half_sub[12]), .D(n325), .Q(n277) );
  NAND22 U311 ( .A(n431), .B(n471), .Q(n239) );
  INV6 U312 ( .A(i_con_AluCtrl[2]), .Q(n90) );
  CLKIN15 U313 ( .A(sum_1[8]), .Q(n59) );
  INV0 U314 ( .A(n17), .Q(n54) );
  CLKIN0 U315 ( .A(i_data_A[21]), .Q(n381) );
  NAND42 U316 ( .A(n461), .B(n460), .C(n459), .D(n458), .Q(o_data_AluRes[26])
         );
  AOI2112 U317 ( .A(N239), .B(n141), .C(n293), .D(n292), .Q(n295) );
  AOI222 U318 ( .A(pre_sum_3b[6]), .B(n8), .C(pre_sum_3a[6]), .D(n53), .Q(n402) );
  NAND22 U319 ( .A(n56), .B(n57), .Q(n58) );
  NAND22 U320 ( .A(n58), .B(n227), .Q(n229) );
  INV0 U321 ( .A(n132), .Q(n56) );
  INV3 U322 ( .A(n228), .Q(n57) );
  AOI212 U323 ( .A(sum_1[6]), .B(n471), .C(n229), .Q(n230) );
  IMUX21 U324 ( .A(n289), .B(n288), .S(n111), .Q(n293) );
  NAND24 U325 ( .A(n355), .B(n354), .Q(n69) );
  AOI2112 U326 ( .A(n162), .B(n425), .C(n424), .D(n423), .Q(n437) );
  AOI221 U327 ( .A(n31), .B(n249), .C(pre_sum_2a[1]), .D(n304), .Q(n255) );
  AOI221 U328 ( .A(pre_sum_2b[0]), .B(n305), .C(N233), .D(n141), .Q(n246) );
  NAND26 U329 ( .A(n319), .B(n471), .Q(n320) );
  OAI210 U330 ( .A(n129), .B(n396), .C(i_data_A[22]), .Q(n397) );
  OAI210 U331 ( .A(n129), .B(n347), .C(i_data_A[18]), .Q(n348) );
  AOI212 U332 ( .A(n136), .B(n160), .C(n129), .Q(n370) );
  CLKIN6 U333 ( .A(n63), .Q(n64) );
  AOI222 U334 ( .A(N224), .B(n80), .C(n5), .D(pre_sum_4a[7]), .Q(n533) );
  AOI221 U335 ( .A(N232), .B(n142), .C(i_data_A[7]), .D(n130), .Q(n237) );
  NAND42 U336 ( .A(n490), .B(n489), .C(n488), .D(n487), .Q(o_data_AluRes[28])
         );
  AOI222 U337 ( .A(n529), .B(pre_sum_4a[1]), .C(pre_sum_4b[1]), .D(n55), .Q(
        n449) );
  AOI222 U338 ( .A(N223), .B(n80), .C(n529), .D(pre_sum_4a[6]), .Q(n513) );
  AOI222 U339 ( .A(pre_sum_4a[3]), .B(n529), .C(pre_sum_4b[3]), .D(n55), .Q(
        n476) );
  AOI222 U340 ( .A(N222), .B(n81), .C(n5), .D(pre_sum_4a[5]), .Q(n500) );
  CLKIN3 U341 ( .A(n131), .Q(n130) );
  NAND24 U342 ( .A(n321), .B(n471), .Q(n322) );
  NAND32 U343 ( .A(n389), .B(n390), .C(n76), .Q(o_data_AluRes[21]) );
  NAND23 U344 ( .A(n380), .B(n379), .Q(o_data_AluRes[20]) );
  IMUX20 U345 ( .A(n275), .B(n274), .S(n151), .Q(n276) );
  CLKIN0 U346 ( .A(n44), .Q(n398) );
  AOI220 U347 ( .A(i_data_A[13]), .B(n281), .C(pre_sum_2a[5]), .D(n304), .Q(
        n287) );
  AOI2112 U348 ( .A(N244), .B(n141), .C(n363), .D(n362), .Q(n367) );
  NAND23 U349 ( .A(n87), .B(n533), .Q(o_data_AluRes[31]) );
  IMUX20 U350 ( .A(n135), .B(n536), .S(n151), .Q(n272) );
  IMUX21 U351 ( .A(n267), .B(n266), .S(n35), .Q(n268) );
  CLKIN15 U352 ( .A(n131), .Q(n129) );
  IMUX21 U353 ( .A(n137), .B(n105), .S(n124), .Q(n504) );
  IMUX20 U354 ( .A(n140), .B(n105), .S(n16), .Q(n396) );
  AOI221 U355 ( .A(pre_subb[13]), .B(n531), .C(n25), .D(pre_suba[13]), .Q(n499) );
  NAND24 U356 ( .A(n286), .B(n284), .Q(n61) );
  AOI222 U357 ( .A(pre_sum_2b[5]), .B(n305), .C(N238), .D(n142), .Q(n286) );
  AOI221 U358 ( .A(N198), .B(n80), .C(N230), .D(n141), .Q(n225) );
  AOI2112 U359 ( .A(n164), .B(n457), .C(n456), .D(n455), .Q(n461) );
  AOI222 U360 ( .A(n59), .B(n429), .C(n60), .D(n428), .Q(n430) );
  AOI212 U361 ( .A(N250), .B(n142), .C(n442), .Q(n443) );
  BUF15 U362 ( .A(i_data_B[28]), .Q(n156) );
  AOI222 U363 ( .A(n32), .B(n368), .C(N245), .D(n142), .Q(n377) );
  NAND42 U364 ( .A(n295), .B(n294), .C(n297), .D(n296), .Q(o_data_AluRes[14])
         );
  AOI212 U365 ( .A(n159), .B(n373), .C(n372), .Q(n376) );
  AOI222 U366 ( .A(pre_sum_2b[3]), .B(n305), .C(N236), .D(n142), .Q(n270) );
  AOI222 U367 ( .A(n59), .B(n48), .C(n46), .D(n60), .Q(n432) );
  IMUX21 U368 ( .A(n395), .B(n394), .S(n16), .Q(n400) );
  OAI2111 U369 ( .A(i_data_A[6]), .B(n139), .C(n169), .D(n132), .Q(n226) );
  INV6 U370 ( .A(i_data_B[12]), .Q(n152) );
  NOR42 U371 ( .A(n192), .B(n191), .C(n189), .D(n188), .Q(n199) );
  NAND24 U372 ( .A(n184), .B(n182), .Q(n189) );
  AOI212 U373 ( .A(n48), .B(n59), .C(pre_sum_3a[8]), .Q(n426) );
  AOI221 U374 ( .A(n414), .B(pre_sum_3b[5]), .C(n413), .D(pre_sum_3a[5]), .Q(
        n390) );
  NAND34 U375 ( .A(n469), .B(n470), .C(n471), .Q(n433) );
  AOI222 U376 ( .A(pre_subb[10]), .B(n27), .C(n25), .D(pre_suba[10]), .Q(n458)
         );
  BUF15 U377 ( .A(i_data_B[30]), .Q(n124) );
  AOI222 U378 ( .A(pre_subb[14]), .B(n27), .C(pre_suba[14]), .D(n25), .Q(n512)
         );
  OAI2112 U379 ( .A(n107), .B(n54), .C(n444), .D(n443), .Q(n445) );
  NAND42 U380 ( .A(n255), .B(n254), .C(n253), .D(n252), .Q(o_data_AluRes[9])
         );
  BUF15 U381 ( .A(i_data_B[29]), .Q(n123) );
  AOI221 U382 ( .A(pre_sum_2b[8]), .B(sum_1[8]), .C(n48), .D(n59), .Q(n321) );
  AOI222 U383 ( .A(n25), .B(pre_suba[11]), .C(pre_subb[11]), .D(n27), .Q(n475)
         );
  BUF15 U384 ( .A(i_data_B[16]), .Q(n153) );
  NAND34 U385 ( .A(n473), .B(n472), .C(n471), .Q(n474) );
  NAND42 U386 ( .A(n279), .B(n278), .C(n277), .D(n276), .Q(o_data_AluRes[12])
         );
  IMUX22 U387 ( .A(n429), .B(n428), .S(sum_1[8]), .Q(n319) );
  INV15 U388 ( .A(n158), .Q(n157) );
  AOI221 U389 ( .A(n530), .B(pre_suba[6]), .C(pre_subb[6]), .D(n14), .Q(n401)
         );
  NAND24 U390 ( .A(n271), .B(n66), .Q(n82) );
  NAND32 U391 ( .A(n340), .B(n341), .C(n68), .Q(o_data_AluRes[17]) );
  CLKIN6 U392 ( .A(n67), .Q(n68) );
  NAND32 U393 ( .A(n353), .B(n352), .C(n70), .Q(o_data_AluRes[18]) );
  INV6 U394 ( .A(n69), .Q(n70) );
  CLKIN6 U395 ( .A(n77), .Q(n78) );
  BUF6 U396 ( .A(n523), .Q(n140) );
  AOI212 U397 ( .A(N218), .B(n80), .C(n445), .Q(n448) );
  AOI222 U398 ( .A(n25), .B(pre_suba[12]), .C(n27), .D(pre_subb[12]), .Q(n487)
         );
  AOI222 U399 ( .A(pre_sum_3b[4]), .B(n414), .C(pre_sum_3a[4]), .D(n413), .Q(
        n374) );
  INV6 U400 ( .A(n79), .Q(n81) );
  INV15 U401 ( .A(n104), .Q(n536) );
  BUF15 U402 ( .A(i_data_B[21]), .Q(n116) );
  BUF15 U403 ( .A(i_data_B[24]), .Q(n102) );
  BUF15 U404 ( .A(i_data_B[26]), .Q(n103) );
  BUF15 U405 ( .A(i_data_B[23]), .Q(n155) );
  AOI222 U406 ( .A(pre_subb[15]), .B(n531), .C(pre_suba[15]), .D(n530), .Q(
        n532) );
  CLKIN0 U407 ( .A(n313), .Q(n89) );
  IMUX30 U408 ( .A(n517), .B(n135), .C(n205), .S0(i_data_A[2]), .S1(n18), .Q(
        n206) );
  AOI221 U409 ( .A(N195), .B(n80), .C(N227), .D(n141), .Q(n209) );
  NAND41 U410 ( .A(n219), .B(n218), .C(n216), .D(n217), .Q(o_data_AluRes[4])
         );
  AOI221 U411 ( .A(N231), .B(n142), .C(N199), .D(n80), .Q(n232) );
  AOI221 U412 ( .A(pre_sum_2b[2]), .B(n305), .C(N235), .D(n141), .Q(n262) );
  OAI210 U413 ( .A(n130), .B(n504), .C(i_data_A[30]), .Q(n505) );
  AOI221 U414 ( .A(N201), .B(n80), .C(half_sub[8]), .D(n325), .Q(n245) );
  NAND22 U415 ( .A(half_sub[3]), .B(n325), .Q(n213) );
  IMUX20 U416 ( .A(n135), .B(n536), .S(n17), .Q(n248) );
  NAND22 U417 ( .A(half_sub[5]), .B(n325), .Q(n224) );
  AOI211 U418 ( .A(n466), .B(n132), .C(n167), .Q(n467) );
  AOI211 U419 ( .A(n291), .B(n132), .C(n290), .Q(n292) );
  NOR22 U420 ( .A(n193), .B(n89), .Q(n88) );
  INV2 U421 ( .A(n177), .Q(n191) );
  NAND41 U422 ( .A(n214), .B(n213), .C(n212), .D(n211), .Q(o_data_AluRes[3])
         );
  IMUX21 U423 ( .A(n496), .B(n495), .S(n123), .Q(n497) );
  NAND41 U424 ( .A(n204), .B(n203), .C(n202), .D(n201), .Q(o_data_AluRes[1])
         );
  IMUX20 U425 ( .A(n138), .B(n104), .S(n85), .Q(n335) );
  INV0 U426 ( .A(i_data_A[28]), .Q(n481) );
  INV0 U427 ( .A(i_data_A[0]), .Q(n170) );
  IMUX21 U428 ( .A(n299), .B(n298), .S(n84), .Q(n303) );
  AOI210 U429 ( .A(n136), .B(n300), .C(n129), .Q(n298) );
  IMUX20 U430 ( .A(n135), .B(n536), .S(n84), .Q(n301) );
  NAND41 U431 ( .A(n263), .B(n262), .C(n261), .D(n260), .Q(o_data_AluRes[10])
         );
  NAND31 U432 ( .A(n232), .B(n231), .C(n230), .Q(o_data_AluRes[6]) );
  IMUX20 U433 ( .A(n135), .B(n536), .S(n111), .Q(n291) );
  AOI210 U434 ( .A(n136), .B(n165), .C(n129), .Q(n453) );
  IMUX21 U435 ( .A(n422), .B(n421), .S(n101), .Q(n423) );
  AOI210 U436 ( .A(n136), .B(n163), .C(n129), .Q(n421) );
  IMUX20 U437 ( .A(n136), .B(n536), .S(n21), .Q(n450) );
  IMUX20 U438 ( .A(n135), .B(n536), .S(n11), .Q(n280) );
  IMUX20 U439 ( .A(n136), .B(n536), .S(n7), .Q(n466) );
  IMUX20 U440 ( .A(n251), .B(n250), .S(n17), .Q(n252) );
  NAND41 U441 ( .A(n245), .B(n246), .C(n247), .D(n244), .Q(o_data_AluRes[8])
         );
  NAND41 U442 ( .A(n237), .B(n236), .C(n235), .D(n234), .Q(o_data_AluRes[7])
         );
  NAND41 U443 ( .A(n209), .B(n208), .C(n207), .D(n206), .Q(o_data_AluRes[2])
         );
  NAND41 U444 ( .A(n225), .B(n224), .C(n223), .D(n222), .Q(o_data_AluRes[5])
         );
  NAND20 U445 ( .A(half_sub[1]), .B(n325), .Q(n203) );
  AOI210 U446 ( .A(n136), .B(n481), .C(n129), .Q(n482) );
  NOR20 U447 ( .A(n166), .B(n462), .Q(n464) );
  NOR20 U448 ( .A(i_data_A[13]), .B(n26), .Q(n283) );
  IMUX21 U449 ( .A(n410), .B(n409), .S(n99), .Q(n411) );
  AOI210 U450 ( .A(n136), .B(n408), .C(n129), .Q(n409) );
  AOI210 U451 ( .A(n136), .B(n494), .C(n129), .Q(n495) );
  AOI210 U452 ( .A(n136), .B(n170), .C(n129), .Q(n171) );
  IMUX21 U453 ( .A(n509), .B(n508), .S(n124), .Q(n510) );
  AOI210 U454 ( .A(n136), .B(n507), .C(n129), .Q(n508) );
  NOR20 U455 ( .A(i_data_A[11]), .B(n462), .Q(n267) );
  BUF2 U456 ( .A(i_data_A[31]), .Q(n127) );
  LOGIC0 U457 ( .Q(n42) );
  LOGIC1 U458 ( .Q(n41) );
  INV0 U459 ( .A(i_data_A[15]), .Q(n300) );
  IMUX20 U460 ( .A(n135), .B(n536), .S(n35), .Q(n264) );
  NAND30 U461 ( .A(n33), .B(n314), .C(n313), .Q(n194) );
  CLKIN0 U462 ( .A(i_data_A[25]), .Q(n439) );
  NAND20 U463 ( .A(i_data_A[1]), .B(n536), .Q(n333) );
  INV0 U464 ( .A(i_data_A[6]), .Q(n228) );
  NAND30 U465 ( .A(n91), .B(n180), .C(n179), .Q(n181) );
  NOR20 U466 ( .A(n31), .B(n26), .Q(n251) );
  OAI210 U467 ( .A(n31), .B(n139), .C(n133), .Q(n250) );
  AOI220 U468 ( .A(sum_1[2]), .B(n471), .C(i_data_A[2]), .D(n130), .Q(n207) );
  NAND20 U469 ( .A(i_data_A[2]), .B(n536), .Q(n221) );
  AOI220 U470 ( .A(sum_1[4]), .B(n471), .C(i_data_A[4]), .D(n130), .Q(n217) );
  NAND20 U471 ( .A(i_data_A[4]), .B(n536), .Q(n183) );
  IMUX21 U472 ( .A(n483), .B(n482), .S(n156), .Q(n484) );
  AOI212 U473 ( .A(n37), .B(n439), .C(n129), .Q(n440) );
  IMUX20 U474 ( .A(n243), .B(n242), .S(n10), .Q(n244) );
  CLKIN0 U475 ( .A(i_data_A[17]), .Q(n331) );
  INV15 U476 ( .A(n146), .Q(n145) );
  IMUX21 U477 ( .A(n346), .B(n345), .S(n22), .Q(n351) );
  IMUX21 U478 ( .A(n138), .B(n104), .S(n153), .Q(n315) );
  OAI210 U479 ( .A(n129), .B(n405), .C(i_data_A[23]), .Q(n406) );
  CLKIN0 U480 ( .A(i_data_A[18]), .Q(n344) );
  CLKIN0 U481 ( .A(n36), .Q(n337) );
  OAI210 U482 ( .A(i_data_A[8]), .B(n139), .C(n133), .Q(n242) );
  NOR20 U483 ( .A(i_data_A[8]), .B(n26), .Q(n243) );
  AOI220 U484 ( .A(i_data_A[8]), .B(n240), .C(pre_sum_2a[0]), .D(n304), .Q(
        n247) );
  INV0 U485 ( .A(n10), .Q(n95) );
  INV0 U486 ( .A(n34), .Q(n361) );
  IMUX21 U487 ( .A(n259), .B(n258), .S(n52), .Q(n260) );
  INV2 U488 ( .A(n52), .Q(n452) );
  AOI221 U489 ( .A(i_data_A[12]), .B(n273), .C(pre_sum_2a[4]), .D(n304), .Q(
        n279) );
  IMUX21 U490 ( .A(n172), .B(n171), .S(n143), .Q(n192) );
  IMUX30 U491 ( .A(n517), .B(n135), .C(n220), .S0(i_data_A[5]), .S1(n15), .Q(
        n222) );
  NOR20 U492 ( .A(i_data_A[10]), .B(n26), .Q(n259) );
  OAI210 U493 ( .A(n129), .B(n359), .C(i_data_A[19]), .Q(n360) );
  IMUX30 U494 ( .A(n517), .B(n135), .C(n233), .S0(i_data_A[7]), .S1(n2), .Q(
        n236) );
  AOI221 U495 ( .A(n530), .B(pre_suba[2]), .C(pre_subb[2]), .D(n14), .Q(n352)
         );
  AOI221 U496 ( .A(n25), .B(pre_suba[1]), .C(pre_subb[1]), .D(n14), .Q(n340)
         );
  CLKIN0 U497 ( .A(i_data_A[22]), .Q(n393) );
  NAND41 U498 ( .A(n449), .B(n448), .C(n447), .D(n446), .Q(o_data_AluRes[25])
         );
  AOI220 U499 ( .A(sum_1[1]), .B(n471), .C(i_data_A[1]), .D(n130), .Q(n202) );
  IMUX30 U500 ( .A(n517), .B(n135), .C(n200), .S0(i_data_A[1]), .S1(n36), .Q(
        n201) );
  CLKIN0 U501 ( .A(i_data_A[23]), .Q(n408) );
  OAI2110 U502 ( .A(i_data_A[4]), .B(n139), .C(n133), .D(n183), .Q(n215) );
  INV0 U503 ( .A(i_data_A[29]), .Q(n494) );
  OAI210 U504 ( .A(n129), .B(n491), .C(i_data_A[29]), .Q(n492) );
  OAI210 U505 ( .A(n130), .B(n438), .C(i_data_A[25]), .Q(n444) );
  NOR20 U506 ( .A(i_data_A[12]), .B(n26), .Q(n275) );
  OAI210 U507 ( .A(i_data_A[12]), .B(n138), .C(n133), .Q(n274) );
  NOR42 U508 ( .A(n312), .B(i_con_AluCtrl[1]), .C(n91), .D(n24), .Q(n518) );
  OAI210 U509 ( .A(i_data_A[10]), .B(n139), .C(n133), .Q(n258) );
  AOI220 U510 ( .A(i_data_A[10]), .B(n257), .C(pre_sum_2a[2]), .D(n304), .Q(
        n263) );
  NAND21 U511 ( .A(n530), .B(pre_suba[4]), .Q(n379) );
  IMUX30 U512 ( .A(n517), .B(n135), .C(n210), .S0(i_data_A[3]), .S1(n34), .Q(
        n211) );
  BUF15 U513 ( .A(i_data_B[14]), .Q(n112) );
  BUF15 U514 ( .A(i_data_B[22]), .Q(n119) );
  BUF15 U515 ( .A(i_data_B[25]), .Q(n121) );
  BUF15 U516 ( .A(i_data_B[18]), .Q(n154) );
  CLKIN3 U517 ( .A(n128), .Q(n187) );
  CLKIN3 U518 ( .A(n524), .Q(n195) );
  NAND22 U519 ( .A(half_sub[6]), .B(n325), .Q(n231) );
  NAND22 U520 ( .A(n238), .B(n133), .Q(n240) );
  AOI222 U521 ( .A(pre_sum_2b[1]), .B(n305), .C(N234), .D(n141), .Q(n254) );
  NAND22 U522 ( .A(n256), .B(n133), .Q(n257) );
  NAND22 U523 ( .A(n264), .B(n133), .Q(n265) );
  NAND22 U524 ( .A(n272), .B(n133), .Q(n273) );
  NAND22 U525 ( .A(n280), .B(n133), .Q(n281) );
  NAND22 U526 ( .A(n517), .B(n290), .Q(n289) );
  NAND22 U527 ( .A(n517), .B(n300), .Q(n299) );
  NAND22 U528 ( .A(N208), .B(n80), .Q(n308) );
  NAND22 U529 ( .A(n517), .B(n158), .Q(n311) );
  NAND22 U530 ( .A(n517), .B(n331), .Q(n334) );
  OAI212 U531 ( .A(n106), .B(n337), .C(n336), .Q(n338) );
  NAND22 U532 ( .A(n517), .B(n356), .Q(n358) );
  NAND22 U533 ( .A(N212), .B(n80), .Q(n366) );
  CLKIN3 U534 ( .A(n107), .Q(n368) );
  NAND22 U535 ( .A(n517), .B(n381), .Q(n383) );
  OAI212 U536 ( .A(n106), .B(n407), .C(n406), .Q(n412) );
  NAND22 U537 ( .A(n517), .B(n408), .Q(n410) );
  AOI2112 U538 ( .A(N248), .B(n141), .C(n412), .D(n411), .Q(n418) );
  NAND22 U539 ( .A(N216), .B(n80), .Q(n417) );
  NAND42 U540 ( .A(n418), .B(n417), .C(n416), .D(n415), .Q(o_data_AluRes[23])
         );
  NAND22 U541 ( .A(n419), .B(n132), .Q(n425) );
  OAI212 U542 ( .A(n107), .B(n95), .C(n420), .Q(n424) );
  NAND22 U543 ( .A(N217), .B(n80), .Q(n436) );
  OAI212 U544 ( .A(n431), .B(n428), .C(n426), .Q(n473) );
  AOI212 U545 ( .A(n59), .B(n429), .C(pre_sum_3b[8]), .Q(n427) );
  OAI212 U546 ( .A(n46), .B(n431), .C(n427), .Q(n472) );
  AOI222 U547 ( .A(n55), .B(pre_sum_4b[0]), .C(n5), .D(pre_sum_4a[0]), .Q(n435) );
  NAND42 U548 ( .A(n437), .B(n436), .C(n434), .D(n435), .Q(o_data_AluRes[24])
         );
  NAND22 U549 ( .A(n450), .B(n132), .Q(n457) );
  NAND22 U550 ( .A(N251), .B(n142), .Q(n451) );
  OAI212 U551 ( .A(n107), .B(n452), .C(n451), .Q(n456) );
  AOI222 U552 ( .A(n528), .B(pre_sum_4b[2]), .C(n5), .D(pre_sum_4a[2]), .Q(
        n459) );
  OAI212 U553 ( .A(n166), .B(n138), .C(n133), .Q(n463) );
  NAND22 U554 ( .A(N220), .B(n80), .Q(n477) );
  NAND42 U555 ( .A(n478), .B(n477), .C(n476), .D(n475), .Q(o_data_AluRes[27])
         );
  NAND22 U556 ( .A(n479), .B(n132), .Q(n486) );
  NAND22 U557 ( .A(N253), .B(n142), .Q(n480) );
  NAND22 U558 ( .A(n517), .B(n481), .Q(n483) );
  AOI222 U559 ( .A(pre_sum_4a[4]), .B(n529), .C(pre_sum_4b[4]), .D(n55), .Q(
        n488) );
  OAI212 U560 ( .A(n107), .B(n493), .C(n492), .Q(n498) );
  NAND22 U561 ( .A(n517), .B(n494), .Q(n496) );
  NAND22 U562 ( .A(n55), .B(pre_sum_4b[5]), .Q(n501) );
  NAND42 U563 ( .A(n502), .B(n501), .C(n500), .D(n499), .Q(o_data_AluRes[29])
         );
  OAI212 U564 ( .A(n107), .B(n506), .C(n505), .Q(n511) );
  NAND22 U565 ( .A(n517), .B(n507), .Q(n509) );
  AOI2112 U566 ( .A(N255), .B(n141), .C(n511), .D(n510), .Q(n515) );
  NAND22 U567 ( .A(n55), .B(pre_sum_4b[6]), .Q(n514) );
  NAND42 U568 ( .A(n515), .B(n514), .C(n513), .D(n512), .Q(o_data_AluRes[30])
         );
  OAI212 U569 ( .A(n198), .B(n520), .C(n519), .Q(n526) );
  OAI222 U570 ( .A(n524), .B(n140), .C(n106), .D(n521), .Q(n525) );
endmodule


module E_alu_control ( o_con_AluCtrl, i_con_AluOp, i_con_FuncCode );
  output [3:0] o_con_AluCtrl;
  input [5:0] i_con_AluOp;
  input [5:0] i_con_FuncCode;
  wire   n22, n24, n27, n28, n29, n30, n38, n43, n45, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n23, n25, n26, n31, n32, n33, n34, n35, n36, n37, n39, n40, n41,
         n42, n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;

  INV3 U3 ( .A(n6), .Q(n40) );
  NOR33 U4 ( .A(n36), .B(n5), .C(n68), .Q(n57) );
  INV6 U5 ( .A(n4), .Q(n5) );
  CLKIN8 U6 ( .A(i_con_FuncCode[2]), .Q(n11) );
  BUF12 U7 ( .A(n48), .Q(n10) );
  INV2 U8 ( .A(n68), .Q(n7) );
  NAND34 U9 ( .A(n41), .B(n40), .C(n39), .Q(o_con_AluCtrl[1]) );
  IMUX22 U10 ( .A(n35), .B(n34), .S(i_con_AluOp[0]), .Q(n41) );
  NOR22 U11 ( .A(n37), .B(n58), .Q(n39) );
  INV6 U12 ( .A(n60), .Q(n17) );
  INV6 U13 ( .A(i_con_FuncCode[5]), .Q(n14) );
  NAND43 U14 ( .A(n11), .B(i_con_FuncCode[1]), .C(i_con_FuncCode[5]), .D(
        i_con_FuncCode[3]), .Q(n1) );
  NOR32 U15 ( .A(n7), .B(n8), .C(n56), .Q(n9) );
  INV3 U16 ( .A(i_con_FuncCode[1]), .Q(n61) );
  NOR23 U17 ( .A(n2), .B(n57), .Q(n38) );
  NAND21 U18 ( .A(n36), .B(i_con_AluOp[0]), .Q(n29) );
  INV6 U19 ( .A(n1), .Q(n47) );
  INV3 U20 ( .A(n32), .Q(n33) );
  NAND26 U21 ( .A(n12), .B(n59), .Q(n42) );
  NAND32 U22 ( .A(i_con_FuncCode[5]), .B(n11), .C(n13), .Q(n59) );
  CLKIN6 U23 ( .A(i_con_FuncCode[3]), .Q(n13) );
  NAND22 U24 ( .A(n49), .B(i_con_FuncCode[1]), .Q(n51) );
  NOR24 U25 ( .A(n56), .B(i_con_AluOp[1]), .Q(n2) );
  NAND21 U26 ( .A(n17), .B(i_con_FuncCode[0]), .Q(n18) );
  NAND26 U27 ( .A(n47), .B(n15), .Q(n46) );
  OAI2112 U28 ( .A(n53), .B(n52), .C(n51), .D(n50), .Q(n3) );
  NAND24 U29 ( .A(n46), .B(n44), .Q(n53) );
  NOR23 U30 ( .A(n43), .B(n56), .Q(n4) );
  INV3 U31 ( .A(n22), .Q(n68) );
  INV6 U32 ( .A(i_con_AluOp[0]), .Q(n56) );
  NAND22 U33 ( .A(n59), .B(n33), .Q(n35) );
  INV1 U34 ( .A(n62), .Q(n64) );
  NAND31 U35 ( .A(i_con_FuncCode[2]), .B(i_con_FuncCode[5]), .C(n13), .Q(n48)
         );
  NAND22 U36 ( .A(n47), .B(i_con_FuncCode[0]), .Q(n62) );
  NOR40 U37 ( .A(n36), .B(n43), .C(n68), .D(n56), .Q(n6) );
  NOR22 U38 ( .A(i_con_AluOp[5]), .B(i_con_AluOp[4]), .Q(n43) );
  CLKIN6 U39 ( .A(n42), .Q(n44) );
  OAI211 U40 ( .A(n32), .B(n21), .C(n20), .Q(n31) );
  CLKIN2 U41 ( .A(n30), .Q(n67) );
  INV6 U42 ( .A(n46), .Q(n54) );
  INV6 U43 ( .A(n10), .Q(n49) );
  OAI212 U44 ( .A(n54), .B(n63), .C(n20), .Q(n55) );
  NAND26 U45 ( .A(n38), .B(n45), .Q(n30) );
  OAI2112 U46 ( .A(n27), .B(n28), .C(n29), .D(n67), .Q(o_con_AluCtrl[2]) );
  NOR42 U47 ( .A(i_con_AluOp[4]), .B(i_con_AluOp[3]), .C(n66), .D(n69), .Q(n36) );
  NAND41 U48 ( .A(n43), .B(i_con_AluOp[2]), .C(i_con_AluOp[3]), .D(
        i_con_AluOp[0]), .Q(n45) );
  NOR32 U49 ( .A(n65), .B(n64), .C(n3), .Q(n27) );
  NOR24 U50 ( .A(n9), .B(n30), .Q(n24) );
  INV0 U51 ( .A(n66), .Q(n8) );
  CLKIN6 U52 ( .A(n24), .Q(n23) );
  OAI220 U53 ( .A(n61), .B(n60), .C(n61), .D(n59), .Q(n65) );
  CLKIN0 U54 ( .A(n28), .Q(n20) );
  INV3 U55 ( .A(i_con_FuncCode[4]), .Q(n50) );
  NAND22 U56 ( .A(n10), .B(n62), .Q(n52) );
  AOI210 U57 ( .A(n17), .B(n61), .C(i_con_FuncCode[4]), .Q(n16) );
  NAND30 U58 ( .A(n43), .B(i_con_AluOp[0]), .C(i_con_AluOp[3]), .Q(n26) );
  OAI2110 U59 ( .A(n19), .B(n10), .C(n18), .D(n46), .Q(n21) );
  NOR20 U60 ( .A(i_con_AluOp[3]), .B(i_con_AluOp[2]), .Q(n34) );
  CLKIN6 U61 ( .A(i_con_AluOp[2]), .Q(n66) );
  NAND34 U62 ( .A(i_con_AluOp[3]), .B(i_con_AluOp[4]), .C(n69), .Q(n22) );
  CLKIN6 U63 ( .A(i_con_AluOp[5]), .Q(n69) );
  XNR20 U64 ( .A(i_con_FuncCode[1]), .B(i_con_FuncCode[0]), .Q(n19) );
  NAND34 U65 ( .A(n31), .B(n26), .C(n25), .Q(o_con_AluCtrl[0]) );
  NAND22 U66 ( .A(i_con_AluOp[1]), .B(n56), .Q(n28) );
  CLKIN3 U67 ( .A(i_con_FuncCode[0]), .Q(n15) );
  NAND33 U68 ( .A(n13), .B(n11), .C(n14), .Q(n60) );
  OAI212 U69 ( .A(i_con_FuncCode[1]), .B(n15), .C(n17), .Q(n12) );
  OAI312 U70 ( .A(n42), .B(n49), .C(n54), .D(n16), .Q(n32) );
  CLKIN3 U71 ( .A(n29), .Q(n37) );
  NOR24 U72 ( .A(n37), .B(n23), .Q(n25) );
  CLKIN3 U73 ( .A(i_con_AluOp[1]), .Q(n58) );
  OAI2112 U74 ( .A(n53), .B(n52), .C(n51), .D(n50), .Q(n63) );
  OAI2112 U75 ( .A(n22), .B(n56), .C(n24), .D(n55), .Q(o_con_AluCtrl[3]) );
endmodule


module E_famux5 ( i_data_rs, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fa, o_data_alusra );
  input [31:0] i_data_rs;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fa;
  output [31:0] o_data_alusra;
  wire   n164, n165, n166, n167, n168, n169, n170, n171, n1, n2, n3, n4, n5,
         n6, n7, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n35, n36,
         n38, n40, n42, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163;

  CLKIN6 U1 ( .A(n168), .Q(n36) );
  NAND26 U2 ( .A(n15), .B(n16), .Q(n77) );
  INV6 U3 ( .A(n158), .Q(n17) );
  AOI222 U4 ( .A(n160), .B(i_data_lwM[23]), .C(i_data_lwW[23]), .D(n29), .Q(
        n132) );
  NAND21 U5 ( .A(i_data_alures[29]), .B(n20), .Q(n153) );
  NAND23 U6 ( .A(i_data_alures[19]), .B(n20), .Q(n120) );
  NAND22 U7 ( .A(i_data_alures[2]), .B(n18), .Q(n63) );
  NAND34 U8 ( .A(n99), .B(n97), .C(n98), .Q(n167) );
  INV6 U9 ( .A(n171), .Q(n45) );
  AOI222 U10 ( .A(n160), .B(i_data_lwM[25]), .C(i_data_alures[25]), .D(n18), 
        .Q(n139) );
  NAND21 U11 ( .A(i_data_rs[9]), .B(n148), .Q(n84) );
  AOI221 U12 ( .A(i_data_rs[28]), .B(n148), .C(i_data_writeres[28]), .D(n44), 
        .Q(n151) );
  NAND22 U13 ( .A(i_data_alures[4]), .B(n19), .Q(n69) );
  INV15 U14 ( .A(n6), .Q(n19) );
  INV15 U15 ( .A(n77), .Q(n10) );
  INV10 U16 ( .A(n166), .Q(n38) );
  BUF15 U17 ( .A(n165), .Q(o_data_alusra[22]) );
  NAND33 U18 ( .A(n76), .B(n74), .C(n75), .Q(o_data_alusra[6]) );
  INV10 U19 ( .A(n167), .Q(n42) );
  NAND23 U20 ( .A(i_data_alures[12]), .B(n19), .Q(n95) );
  NAND34 U21 ( .A(n96), .B(n94), .C(n95), .Q(o_data_alusra[12]) );
  NAND34 U22 ( .A(n54), .B(n53), .C(n52), .Q(n171) );
  CLKIN15 U23 ( .A(n51), .Q(n29) );
  CLKBU15 U24 ( .A(n164), .Q(o_data_alusra[28]) );
  INV10 U25 ( .A(n58), .Q(n148) );
  NAND34 U26 ( .A(n124), .B(n123), .C(n122), .Q(o_data_alusra[20]) );
  NAND26 U27 ( .A(i_data_writeres[10]), .B(n44), .Q(n89) );
  INV12 U28 ( .A(n48), .Q(n44) );
  AOI221 U29 ( .A(i_data_lwM[20]), .B(n160), .C(i_data_lwW[20]), .D(n29), .Q(
        n122) );
  NAND26 U30 ( .A(n20), .B(i_data_alures[10]), .Q(n88) );
  AOI222 U31 ( .A(i_data_rs[3]), .B(n31), .C(i_data_writeres[3]), .D(n1), .Q(
        n67) );
  NAND34 U32 ( .A(n67), .B(n66), .C(n65), .Q(o_data_alusra[3]) );
  CLKIN4 U33 ( .A(i_con_fa[2]), .Q(n27) );
  CLKIN6 U34 ( .A(i_con_fa[2]), .Q(n56) );
  AOI222 U35 ( .A(n160), .B(i_data_lwM[19]), .C(i_data_lwW[19]), .D(n159), .Q(
        n119) );
  AOI222 U36 ( .A(n32), .B(i_data_lwM[3]), .C(i_data_lwW[3]), .D(n29), .Q(n65)
         );
  NAND22 U37 ( .A(n141), .B(i_data_rs[17]), .Q(n7) );
  NAND24 U38 ( .A(n111), .B(n110), .Q(n112) );
  NAND23 U39 ( .A(i_data_alures[17]), .B(n18), .Q(n110) );
  AOI221 U40 ( .A(i_data_lwM[1]), .B(n32), .C(i_data_lwW[1]), .D(n29), .Q(n59)
         );
  INV3 U41 ( .A(n7), .Q(n113) );
  NAND33 U42 ( .A(n134), .B(n132), .C(n133), .Q(o_data_alusra[23]) );
  INV8 U43 ( .A(n109), .Q(n141) );
  CLKIN6 U44 ( .A(n13), .Q(n14) );
  AOI222 U45 ( .A(i_data_rs[6]), .B(n148), .C(i_data_writeres[6]), .D(n1), .Q(
        n76) );
  AOI221 U46 ( .A(i_data_rs[29]), .B(n10), .C(i_data_writeres[29]), .D(n1), 
        .Q(n154) );
  NAND21 U47 ( .A(i_data_alures[1]), .B(n19), .Q(n60) );
  NAND21 U48 ( .A(i_data_alures[26]), .B(n19), .Q(n143) );
  AOI222 U49 ( .A(i_data_alures[18]), .B(n18), .C(i_data_writeres[18]), .D(n44), .Q(n118) );
  CLKIN15 U50 ( .A(n40), .Q(o_data_alusra[10]) );
  CLKIN15 U51 ( .A(n36), .Q(o_data_alusra[11]) );
  AOI222 U52 ( .A(i_data_rs[2]), .B(n31), .C(i_data_writeres[2]), .D(n1), .Q(
        n64) );
  AOI222 U53 ( .A(n10), .B(i_data_rs[13]), .C(i_data_writeres[13]), .D(n1), 
        .Q(n99) );
  AOI222 U54 ( .A(i_data_rs[23]), .B(n10), .C(i_data_writeres[23]), .D(n1), 
        .Q(n134) );
  NAND33 U55 ( .A(n131), .B(n130), .C(n129), .Q(n165) );
  AOI222 U56 ( .A(n32), .B(i_data_lwM[22]), .C(i_data_lwW[22]), .D(n159), .Q(
        n129) );
  AOI222 U57 ( .A(i_data_rs[19]), .B(n31), .C(i_data_writeres[19]), .D(n1), 
        .Q(n121) );
  AOI222 U58 ( .A(i_data_rs[22]), .B(n10), .C(i_data_writeres[22]), .D(n1), 
        .Q(n131) );
  CLKIN12 U59 ( .A(n35), .Q(n23) );
  NAND22 U60 ( .A(n141), .B(i_data_rs[18]), .Q(n116) );
  NAND33 U61 ( .A(n61), .B(n60), .C(n59), .Q(o_data_alusra[1]) );
  AOI221 U62 ( .A(i_data_rs[1]), .B(n148), .C(i_data_writeres[1]), .D(n1), .Q(
        n61) );
  NAND33 U63 ( .A(n118), .B(n117), .C(n116), .Q(o_data_alusra[18]) );
  INV6 U64 ( .A(n21), .Q(n22) );
  CLKIN6 U65 ( .A(n13), .Q(n2) );
  INV6 U66 ( .A(n169), .Q(n40) );
  CLKIN3 U67 ( .A(n47), .Q(n24) );
  NOR24 U68 ( .A(n113), .B(n112), .Q(n115) );
  INV15 U69 ( .A(n48), .Q(n1) );
  NAND28 U70 ( .A(n13), .B(n30), .Q(n11) );
  CLKIN15 U71 ( .A(n57), .Q(n30) );
  NAND22 U72 ( .A(n160), .B(i_data_lwM[17]), .Q(n111) );
  CLKIN15 U73 ( .A(n35), .Q(n50) );
  NAND26 U74 ( .A(n26), .B(n25), .Q(n31) );
  AOI221 U75 ( .A(i_data_lwM[31]), .B(n160), .C(i_data_lwW[31]), .D(n159), .Q(
        n161) );
  CLKIN15 U76 ( .A(n45), .Q(o_data_alusra[0]) );
  NAND21 U77 ( .A(n10), .B(i_data_rs[21]), .Q(n125) );
  NAND22 U78 ( .A(i_data_alures[3]), .B(n19), .Q(n66) );
  NAND34 U79 ( .A(n108), .B(n107), .C(n106), .Q(o_data_alusra[16]) );
  AOI222 U80 ( .A(i_data_writeres[16]), .B(n1), .C(i_data_lwW[16]), .D(n159), 
        .Q(n108) );
  NAND33 U81 ( .A(n157), .B(n156), .C(n155), .Q(o_data_alusra[30]) );
  NAND21 U82 ( .A(i_data_alures[30]), .B(n18), .Q(n156) );
  NAND20 U83 ( .A(i_data_alures[31]), .B(n19), .Q(n162) );
  NAND21 U84 ( .A(i_data_alures[15]), .B(n19), .Q(n104) );
  NAND21 U85 ( .A(i_data_alures[20]), .B(n20), .Q(n123) );
  NAND21 U86 ( .A(i_data_alures[24]), .B(n20), .Q(n136) );
  NAND21 U87 ( .A(i_data_alures[27]), .B(n20), .Q(n146) );
  AOI222 U88 ( .A(n160), .B(i_data_lwM[10]), .C(i_data_lwW[10]), .D(n159), .Q(
        n90) );
  INV8 U89 ( .A(n49), .Q(n160) );
  CLKIN15 U90 ( .A(n49), .Q(n32) );
  NAND21 U91 ( .A(i_data_alures[5]), .B(n20), .Q(n72) );
  NAND22 U92 ( .A(i_data_alures[21]), .B(n20), .Q(n126) );
  NAND21 U93 ( .A(i_data_alures[14]), .B(n20), .Q(n101) );
  NAND24 U94 ( .A(n11), .B(n12), .Q(n58) );
  NAND22 U95 ( .A(n47), .B(n13), .Q(n25) );
  INV10 U96 ( .A(n51), .Q(n159) );
  NAND33 U97 ( .A(n144), .B(n143), .C(n142), .Q(o_data_alusra[26]) );
  NAND32 U98 ( .A(n151), .B(n150), .C(n149), .Q(n164) );
  NAND33 U99 ( .A(n70), .B(n69), .C(n68), .Q(n170) );
  INV3 U100 ( .A(n47), .Q(n3) );
  NAND22 U101 ( .A(n2), .B(n47), .Q(n5) );
  AOI221 U102 ( .A(n141), .B(i_data_rs[8]), .C(i_data_writeres[8]), .D(n44), 
        .Q(n83) );
  NAND22 U103 ( .A(n13), .B(n3), .Q(n4) );
  NAND24 U104 ( .A(n4), .B(n5), .Q(n109) );
  NAND24 U105 ( .A(n115), .B(n114), .Q(o_data_alusra[17]) );
  NAND22 U106 ( .A(n50), .B(n24), .Q(n26) );
  INV15 U107 ( .A(n158), .Q(n6) );
  CLKIN15 U108 ( .A(n11), .Q(n158) );
  AOI221 U109 ( .A(i_data_rs[12]), .B(n31), .C(i_data_writeres[12]), .D(n44), 
        .Q(n96) );
  NAND22 U110 ( .A(i_data_alures[13]), .B(n19), .Q(n98) );
  NAND33 U111 ( .A(n105), .B(n104), .C(n103), .Q(o_data_alusra[15]) );
  CLKIN15 U112 ( .A(n17), .Q(n18) );
  BUF15 U113 ( .A(n170), .Q(o_data_alusra[4]) );
  AOI222 U114 ( .A(n32), .B(i_data_lwM[4]), .C(n29), .D(i_data_lwW[4]), .Q(n68) );
  NAND33 U115 ( .A(n147), .B(n146), .C(n145), .Q(o_data_alusra[27]) );
  NAND33 U116 ( .A(n64), .B(n63), .C(n62), .Q(o_data_alusra[2]) );
  AOI222 U117 ( .A(n32), .B(i_data_lwM[2]), .C(i_data_lwW[2]), .D(n29), .Q(n62) );
  AOI221 U118 ( .A(i_data_lwM[6]), .B(n160), .C(i_data_lwW[6]), .D(n159), .Q(
        n74) );
  AOI222 U119 ( .A(n32), .B(i_data_lwM[0]), .C(n159), .D(i_data_lwW[0]), .Q(
        n52) );
  NAND26 U120 ( .A(n56), .B(n55), .Q(n47) );
  AOI221 U121 ( .A(n141), .B(i_data_rs[20]), .C(i_data_writeres[20]), .D(n1), 
        .Q(n124) );
  NAND22 U122 ( .A(n141), .B(i_data_rs[16]), .Q(n106) );
  AOI221 U123 ( .A(i_data_lwM[16]), .B(n160), .C(i_data_alures[16]), .D(n18), 
        .Q(n107) );
  INV15 U124 ( .A(n38), .Q(o_data_alusra[19]) );
  AOI221 U125 ( .A(n10), .B(i_data_rs[15]), .C(i_data_writeres[15]), .D(n1), 
        .Q(n105) );
  NAND22 U126 ( .A(i_data_alures[22]), .B(n20), .Q(n130) );
  AOI221 U127 ( .A(i_data_lwM[15]), .B(n160), .C(i_data_lwW[15]), .D(n159), 
        .Q(n103) );
  NAND28 U128 ( .A(n50), .B(n22), .Q(n48) );
  NAND22 U129 ( .A(n57), .B(n2), .Q(n12) );
  INV6 U130 ( .A(n34), .Q(n13) );
  NAND43 U131 ( .A(n89), .B(n88), .C(n87), .D(n90), .Q(n169) );
  CLKIN15 U132 ( .A(n6), .Q(n20) );
  INV12 U133 ( .A(n34), .Q(n35) );
  CLKIN8 U134 ( .A(i_con_fa[1]), .Q(n34) );
  NAND22 U135 ( .A(n13), .B(n30), .Q(n15) );
  NAND22 U136 ( .A(n57), .B(n14), .Q(n16) );
  INV15 U137 ( .A(n42), .Q(o_data_alusra[13]) );
  NAND22 U138 ( .A(n31), .B(i_data_rs[10]), .Q(n87) );
  NAND34 U139 ( .A(n28), .B(i_con_fa[0]), .C(n50), .Q(n51) );
  AOI221 U140 ( .A(i_data_lwM[12]), .B(n160), .C(i_data_lwW[12]), .D(n159), 
        .Q(n94) );
  NAND22 U141 ( .A(i_con_fa[0]), .B(n56), .Q(n21) );
  NAND34 U142 ( .A(n119), .B(n121), .C(n120), .Q(n166) );
  NAND33 U143 ( .A(n137), .B(n136), .C(n135), .Q(o_data_alusra[24]) );
  AOI221 U144 ( .A(n10), .B(i_data_rs[30]), .C(i_data_writeres[30]), .D(n1), 
        .Q(n157) );
  NAND28 U145 ( .A(n55), .B(n56), .Q(n57) );
  AOI222 U146 ( .A(i_data_writeres[25]), .B(n44), .C(n159), .D(i_data_lwW[25]), 
        .Q(n140) );
  NAND21 U147 ( .A(i_data_alures[8]), .B(n20), .Q(n82) );
  NAND22 U148 ( .A(i_data_writeres[21]), .B(n44), .Q(n127) );
  NAND33 U149 ( .A(n73), .B(n72), .C(n71), .Q(o_data_alusra[5]) );
  AOI221 U150 ( .A(n32), .B(i_data_lwM[18]), .C(i_data_lwW[18]), .D(n159), .Q(
        n117) );
  NAND33 U151 ( .A(n83), .B(n82), .C(n81), .Q(o_data_alusra[8]) );
  AOI221 U152 ( .A(n32), .B(i_data_lwM[8]), .C(i_data_lwW[8]), .D(n29), .Q(n81) );
  AOI222 U153 ( .A(i_data_rs[0]), .B(n31), .C(i_data_writeres[0]), .D(n44), 
        .Q(n54) );
  AOI221 U154 ( .A(i_data_writeres[9]), .B(n1), .C(i_data_lwW[9]), .D(n159), 
        .Q(n86) );
  AOI222 U155 ( .A(n141), .B(i_data_rs[4]), .C(i_data_writeres[4]), .D(n44), 
        .Q(n70) );
  AOI221 U156 ( .A(n32), .B(i_data_lwM[30]), .C(i_data_lwW[30]), .D(n29), .Q(
        n155) );
  INV6 U157 ( .A(n27), .Q(n28) );
  NAND33 U158 ( .A(n80), .B(n78), .C(n79), .Q(o_data_alusra[7]) );
  AOI221 U159 ( .A(n160), .B(i_data_lwM[7]), .C(i_data_lwW[7]), .D(n159), .Q(
        n78) );
  AOI221 U160 ( .A(i_data_lwM[28]), .B(n32), .C(i_data_lwW[28]), .D(n29), .Q(
        n149) );
  AOI221 U161 ( .A(i_data_rs[7]), .B(n10), .C(i_data_writeres[7]), .D(n1), .Q(
        n80) );
  NAND34 U162 ( .A(n86), .B(n85), .C(n84), .Q(o_data_alusra[9]) );
  NAND33 U163 ( .A(n154), .B(n153), .C(n152), .Q(o_data_alusra[29]) );
  AOI221 U164 ( .A(n32), .B(i_data_lwM[29]), .C(i_data_lwW[29]), .D(n29), .Q(
        n152) );
  AOI221 U165 ( .A(i_data_lwM[5]), .B(n32), .C(i_data_lwW[5]), .D(n29), .Q(n71) );
  AOI221 U166 ( .A(n32), .B(i_data_lwM[11]), .C(i_data_lwW[11]), .D(n29), .Q(
        n91) );
  AOI221 U167 ( .A(n10), .B(i_data_rs[14]), .C(i_data_writeres[14]), .D(n1), 
        .Q(n102) );
  AOI221 U168 ( .A(i_data_rs[5]), .B(n148), .C(i_data_writeres[5]), .D(n1), 
        .Q(n73) );
  NAND33 U169 ( .A(n93), .B(n92), .C(n91), .Q(n168) );
  NAND21 U170 ( .A(i_data_alures[11]), .B(n20), .Q(n92) );
  NAND34 U171 ( .A(n28), .B(n55), .C(n23), .Q(n49) );
  AOI221 U172 ( .A(i_data_rs[11]), .B(n148), .C(i_data_writeres[11]), .D(n44), 
        .Q(n93) );
  AOI221 U173 ( .A(n160), .B(i_data_lwM[9]), .C(i_data_alures[9]), .D(n19), 
        .Q(n85) );
  NAND33 U174 ( .A(n140), .B(n139), .C(n138), .Q(o_data_alusra[25]) );
  AOI221 U175 ( .A(i_data_rs[27]), .B(n148), .C(i_data_writeres[27]), .D(n1), 
        .Q(n147) );
  AOI221 U176 ( .A(n141), .B(i_data_rs[24]), .C(i_data_writeres[24]), .D(n1), 
        .Q(n137) );
  AOI221 U177 ( .A(n32), .B(i_data_lwM[24]), .C(i_data_lwW[24]), .D(n29), .Q(
        n135) );
  AOI220 U178 ( .A(i_data_rs[31]), .B(n10), .C(i_data_writeres[31]), .D(n1), 
        .Q(n163) );
  AOI221 U179 ( .A(i_data_lwM[26]), .B(n32), .C(i_data_lwW[26]), .D(n29), .Q(
        n142) );
  AOI221 U180 ( .A(n141), .B(i_data_rs[26]), .C(i_data_writeres[26]), .D(n1), 
        .Q(n144) );
  AOI221 U181 ( .A(n32), .B(i_data_lwM[27]), .C(i_data_lwW[27]), .D(n29), .Q(
        n145) );
  AOI221 U182 ( .A(i_data_lwW[17]), .B(n159), .C(i_data_writeres[17]), .D(n44), 
        .Q(n114) );
  NAND33 U183 ( .A(n102), .B(n101), .C(n100), .Q(o_data_alusra[14]) );
  AOI221 U184 ( .A(n32), .B(i_data_lwM[14]), .C(i_data_lwW[14]), .D(n29), .Q(
        n100) );
  AOI221 U185 ( .A(i_data_lwM[13]), .B(n160), .C(i_data_lwW[13]), .D(n159), 
        .Q(n97) );
  CLKIN12 U186 ( .A(i_con_fa[0]), .Q(n55) );
  NAND43 U187 ( .A(n128), .B(n127), .C(n126), .D(n125), .Q(o_data_alusra[21])
         );
  NAND22 U188 ( .A(i_data_alures[0]), .B(n19), .Q(n53) );
  NAND22 U189 ( .A(i_data_alures[6]), .B(n19), .Q(n75) );
  NAND22 U190 ( .A(i_data_alures[7]), .B(n19), .Q(n79) );
  AOI222 U191 ( .A(i_data_lwM[21]), .B(n32), .C(i_data_lwW[21]), .D(n29), .Q(
        n128) );
  NAND22 U192 ( .A(i_data_alures[23]), .B(n19), .Q(n133) );
  NAND22 U193 ( .A(n10), .B(i_data_rs[25]), .Q(n138) );
  NAND22 U194 ( .A(i_data_alures[28]), .B(n20), .Q(n150) );
  NAND33 U195 ( .A(n163), .B(n162), .C(n161), .Q(o_data_alusra[31]) );
endmodule


module E_fbmux5 ( i_data_rt, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fb, o_data_alusrb );
  input [31:0] i_data_rt;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fb;
  output [31:0] o_data_alusrb;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179;

  NAND33 U1 ( .A(n83), .B(n82), .C(n81), .Q(o_data_alusrb[4]) );
  NAND23 U2 ( .A(i_data_rt[4]), .B(n120), .Q(n81) );
  NAND24 U3 ( .A(i_data_rt[14]), .B(n120), .Q(n114) );
  NAND23 U4 ( .A(n179), .B(n178), .Q(n33) );
  NAND33 U5 ( .A(n113), .B(n112), .C(n111), .Q(o_data_alusrb[13]) );
  NAND23 U6 ( .A(n168), .B(n167), .Q(n43) );
  NAND33 U7 ( .A(n139), .B(n138), .C(n137), .Q(o_data_alusrb[20]) );
  CLKIN10 U8 ( .A(n27), .Q(n20) );
  INV8 U9 ( .A(n79), .Q(n15) );
  CLKIN15 U10 ( .A(n54), .Q(n173) );
  NAND26 U11 ( .A(n36), .B(n9), .Q(n90) );
  NAND24 U12 ( .A(n46), .B(i_data_rt[18]), .Q(n127) );
  NAND34 U13 ( .A(n76), .B(n77), .C(n75), .Q(o_data_alusrb[3]) );
  NAND34 U14 ( .A(n67), .B(n68), .C(n66), .Q(o_data_alusrb[0]) );
  INV12 U15 ( .A(n8), .Q(n1) );
  CLKIN15 U16 ( .A(n59), .Q(n8) );
  NAND34 U17 ( .A(n116), .B(n115), .C(n114), .Q(o_data_alusrb[14]) );
  NAND34 U18 ( .A(n73), .B(n74), .C(n72), .Q(o_data_alusrb[2]) );
  NAND24 U19 ( .A(n22), .B(n5), .Q(n58) );
  NAND24 U20 ( .A(n58), .B(i_data_rt[1]), .Q(n70) );
  INV6 U21 ( .A(n43), .Q(n44) );
  NAND34 U22 ( .A(n123), .B(n122), .C(n121), .Q(o_data_alusrb[16]) );
  NAND24 U23 ( .A(n105), .B(n107), .Q(n47) );
  NAND24 U24 ( .A(n10), .B(i_data_lwW[1]), .Q(n71) );
  CLKIN15 U25 ( .A(n63), .Q(n19) );
  AOI222 U26 ( .A(n26), .B(i_data_lwM[20]), .C(n60), .D(i_data_lwW[20]), .Q(
        n138) );
  CLKIN10 U27 ( .A(i_con_fb[2]), .Q(n130) );
  CLKIN12 U28 ( .A(n54), .Q(n23) );
  NAND24 U29 ( .A(n146), .B(n145), .Q(n38) );
  NAND33 U30 ( .A(n166), .B(n165), .C(n164), .Q(o_data_alusrb[28]) );
  NAND22 U31 ( .A(n140), .B(n35), .Q(n22) );
  CLKIN12 U32 ( .A(n65), .Q(n140) );
  NAND26 U33 ( .A(n1), .B(n140), .Q(n36) );
  INV15 U34 ( .A(n64), .Q(n26) );
  AOI222 U35 ( .A(i_data_lwM[26]), .B(n18), .C(i_data_alures[26]), .D(n175), 
        .Q(n159) );
  BUF15 U36 ( .A(n78), .Q(n54) );
  CLKIN15 U37 ( .A(n54), .Q(n24) );
  AOI222 U38 ( .A(n26), .B(i_data_lwM[30]), .C(i_data_lwW[30]), .D(n60), .Q(
        n170) );
  AOI221 U39 ( .A(n58), .B(i_data_rt[30]), .C(n173), .D(i_data_writeres[30]), 
        .Q(n172) );
  AOI222 U40 ( .A(n23), .B(i_data_writeres[14]), .C(i_data_alures[14]), .D(
        n175), .Q(n116) );
  INV15 U41 ( .A(n63), .Q(n175) );
  AOI222 U42 ( .A(n132), .B(i_data_writeres[0]), .C(i_data_alures[0]), .D(n175), .Q(n68) );
  NAND34 U43 ( .A(n86), .B(n85), .C(n84), .Q(o_data_alusrb[5]) );
  AOI222 U44 ( .A(n23), .B(i_data_writeres[16]), .C(i_data_alures[16]), .D(
        n175), .Q(n123) );
  NAND23 U45 ( .A(n17), .B(i_data_rt[9]), .Q(n98) );
  NAND23 U46 ( .A(n120), .B(i_data_rt[15]), .Q(n117) );
  CLKIN6 U47 ( .A(n49), .Q(n50) );
  NAND24 U48 ( .A(n46), .B(i_data_rt[17]), .Q(n124) );
  NAND26 U49 ( .A(n46), .B(i_data_rt[10]), .Q(n101) );
  NAND24 U50 ( .A(i_data_rt[21]), .B(n153), .Q(n141) );
  CLKIN12 U51 ( .A(n104), .Q(n153) );
  INV10 U52 ( .A(n64), .Q(n176) );
  INV10 U53 ( .A(n31), .Q(n32) );
  AOI221 U54 ( .A(i_data_lwM[7]), .B(n18), .C(i_data_lwW[7]), .D(n10), .Q(n92)
         );
  AOI220 U55 ( .A(i_data_lwM[31]), .B(n18), .C(n60), .D(i_data_lwW[31]), .Q(
        n177) );
  NAND24 U56 ( .A(n177), .B(n34), .Q(o_data_alusrb[31]) );
  CLKIN6 U57 ( .A(n40), .Q(n41) );
  NAND34 U58 ( .A(n88), .B(n89), .C(n87), .Q(o_data_alusrb[6]) );
  NAND23 U59 ( .A(i_data_rt[6]), .B(n46), .Q(n87) );
  NAND28 U60 ( .A(n50), .B(n7), .Q(o_data_alusrb[1]) );
  INV15 U61 ( .A(n94), .Q(n59) );
  CLKIN12 U62 ( .A(i_con_fb[1]), .Q(n94) );
  CLKIN6 U63 ( .A(n55), .Q(n56) );
  BUF15 U64 ( .A(n51), .Q(n61) );
  NAND24 U65 ( .A(n11), .B(n8), .Q(n12) );
  CLKIN15 U66 ( .A(n90), .Q(n174) );
  AOI221 U67 ( .A(n24), .B(i_data_writeres[27]), .C(n61), .D(i_data_lwW[27]), 
        .Q(n163) );
  NAND33 U68 ( .A(n163), .B(n162), .C(n161), .Q(o_data_alusrb[27]) );
  NAND24 U69 ( .A(n174), .B(i_data_rt[13]), .Q(n111) );
  NAND28 U70 ( .A(n39), .B(n144), .Q(o_data_alusrb[22]) );
  BUF15 U71 ( .A(n51), .Q(n62) );
  NAND28 U72 ( .A(n159), .B(n32), .Q(o_data_alusrb[26]) );
  AOI222 U73 ( .A(i_data_rt[31]), .B(n174), .C(n23), .D(i_data_writeres[31]), 
        .Q(n179) );
  NAND26 U74 ( .A(n48), .B(n106), .Q(o_data_alusrb[11]) );
  BUF15 U75 ( .A(n51), .Q(n60) );
  CLKIN3 U76 ( .A(n45), .Q(n2) );
  NAND24 U77 ( .A(n41), .B(n96), .Q(o_data_alusrb[8]) );
  AOI222 U78 ( .A(n173), .B(i_data_writeres[6]), .C(i_data_alures[6]), .D(n175), .Q(n89) );
  AOI222 U79 ( .A(i_data_lwM[5]), .B(n18), .C(n62), .D(i_data_lwW[5]), .Q(n85)
         );
  NAND24 U80 ( .A(n12), .B(n13), .Q(n57) );
  CLKIN8 U81 ( .A(i_con_fb[0]), .Q(n131) );
  NAND34 U82 ( .A(n103), .B(n102), .C(n101), .Q(o_data_alusrb[10]) );
  NAND28 U83 ( .A(n169), .B(n44), .Q(o_data_alusrb[29]) );
  NAND34 U84 ( .A(n156), .B(n155), .C(n154), .Q(o_data_alusrb[25]) );
  NAND24 U85 ( .A(n153), .B(i_data_rt[11]), .Q(n105) );
  NAND22 U86 ( .A(i_data_rt[24]), .B(n157), .Q(n150) );
  NAND24 U87 ( .A(i_data_rt[25]), .B(n157), .Q(n154) );
  NAND24 U88 ( .A(i_data_rt[0]), .B(n46), .Q(n66) );
  CLKIN15 U89 ( .A(n42), .Q(n11) );
  INV12 U90 ( .A(n64), .Q(n18) );
  AOI221 U91 ( .A(i_data_lwM[27]), .B(n26), .C(i_data_alures[27]), .D(n175), 
        .Q(n162) );
  NAND26 U92 ( .A(n160), .B(n158), .Q(n31) );
  AOI222 U93 ( .A(i_data_writeres[4]), .B(n23), .C(i_data_alures[4]), .D(n175), 
        .Q(n83) );
  NAND24 U94 ( .A(i_data_rt[23]), .B(n153), .Q(n147) );
  NAND26 U95 ( .A(n28), .B(n20), .Q(n45) );
  NAND22 U96 ( .A(i_data_lwM[1]), .B(n176), .Q(n7) );
  NAND26 U97 ( .A(n36), .B(n16), .Q(n80) );
  AOI222 U98 ( .A(i_data_writeres[13]), .B(n173), .C(i_data_alures[13]), .D(
        n175), .Q(n113) );
  NAND34 U99 ( .A(n149), .B(n148), .C(n147), .Q(o_data_alusrb[23]) );
  AOI222 U100 ( .A(n24), .B(i_data_writeres[23]), .C(i_data_lwW[23]), .D(n25), 
        .Q(n149) );
  CLKIN6 U101 ( .A(n59), .Q(n35) );
  INV4 U102 ( .A(n79), .Q(n4) );
  NAND34 U103 ( .A(n143), .B(n142), .C(n141), .Q(o_data_alusrb[21]) );
  NAND24 U104 ( .A(n30), .B(n99), .Q(o_data_alusrb[9]) );
  AOI222 U105 ( .A(n18), .B(i_data_lwM[4]), .C(n10), .D(i_data_lwW[4]), .Q(n82) );
  NAND24 U106 ( .A(n1), .B(n4), .Q(n5) );
  NAND22 U107 ( .A(n3), .B(n79), .Q(n6) );
  NAND24 U108 ( .A(n5), .B(n6), .Q(n17) );
  CLKIN2 U109 ( .A(n59), .Q(n3) );
  NAND33 U110 ( .A(n134), .B(n136), .C(n135), .Q(o_data_alusrb[19]) );
  NAND33 U111 ( .A(n152), .B(n151), .C(n150), .Q(o_data_alusrb[24]) );
  NAND34 U112 ( .A(n118), .B(n119), .C(n117), .Q(o_data_alusrb[15]) );
  NAND22 U113 ( .A(i_data_rt[22]), .B(n157), .Q(n144) );
  NAND34 U114 ( .A(n109), .B(n110), .C(n108), .Q(o_data_alusrb[12]) );
  AOI222 U115 ( .A(i_data_lwM[12]), .B(n176), .C(n62), .D(i_data_lwW[12]), .Q(
        n109) );
  NAND28 U116 ( .A(n131), .B(n130), .Q(n65) );
  NAND26 U117 ( .A(n131), .B(n130), .Q(n42) );
  CLKIN2 U118 ( .A(n59), .Q(n14) );
  NAND24 U119 ( .A(n35), .B(n15), .Q(n9) );
  CLKIN12 U120 ( .A(n104), .Q(n157) );
  BUF15 U121 ( .A(n51), .Q(n10) );
  NAND22 U122 ( .A(n65), .B(n59), .Q(n13) );
  AOI222 U123 ( .A(i_data_writeres[12]), .B(n173), .C(i_data_alures[12]), .D(
        n175), .Q(n110) );
  NAND34 U124 ( .A(n128), .B(n129), .C(n127), .Q(o_data_alusrb[18]) );
  CLKIN15 U125 ( .A(n45), .Q(n132) );
  NAND23 U126 ( .A(i_data_rt[12]), .B(n120), .Q(n108) );
  AOI222 U127 ( .A(i_data_writeres[20]), .B(n23), .C(i_data_alures[20]), .D(
        n175), .Q(n139) );
  NAND28 U128 ( .A(n11), .B(n59), .Q(n63) );
  AOI222 U129 ( .A(i_data_writeres[25]), .B(n23), .C(n62), .D(i_data_lwW[25]), 
        .Q(n156) );
  AOI221 U130 ( .A(n132), .B(i_data_writeres[2]), .C(i_data_alures[2]), .D(n19), .Q(n74) );
  AOI222 U131 ( .A(i_data_lwM[22]), .B(n26), .C(i_data_alures[22]), .D(n19), 
        .Q(n145) );
  NAND24 U132 ( .A(n14), .B(n15), .Q(n16) );
  CLKIN15 U133 ( .A(n80), .Q(n120) );
  BUF15 U134 ( .A(n51), .Q(n25) );
  AOI222 U135 ( .A(i_data_lwM[23]), .B(n26), .C(i_data_alures[23]), .D(n175), 
        .Q(n148) );
  AOI222 U136 ( .A(n26), .B(i_data_lwM[25]), .C(i_data_alures[25]), .D(n175), 
        .Q(n155) );
  NAND34 U137 ( .A(n93), .B(n92), .C(n91), .Q(o_data_alusrb[7]) );
  INV12 U138 ( .A(n140), .Q(n21) );
  INV15 U139 ( .A(n52), .Q(n51) );
  AOI221 U140 ( .A(i_data_writeres[7]), .B(n23), .C(i_data_alures[7]), .D(n175), .Q(n93) );
  NAND28 U141 ( .A(n28), .B(n27), .Q(n52) );
  CLKBU12 U142 ( .A(i_con_fb[2]), .Q(n27) );
  AOI221 U143 ( .A(i_data_rt[19]), .B(n133), .C(n2), .D(i_data_writeres[19]), 
        .Q(n136) );
  XNR21 U144 ( .A(n59), .B(n42), .Q(n133) );
  NAND24 U145 ( .A(i_data_rt[26]), .B(n157), .Q(n158) );
  AOI221 U146 ( .A(n173), .B(i_data_writeres[5]), .C(i_data_alures[5]), .D(
        n175), .Q(n86) );
  NAND22 U147 ( .A(i_data_rt[7]), .B(n174), .Q(n91) );
  CLKIN15 U148 ( .A(n65), .Q(n79) );
  NAND22 U149 ( .A(i_data_rt[28]), .B(n174), .Q(n164) );
  NAND21 U150 ( .A(n57), .B(i_data_rt[8]), .Q(n95) );
  NAND24 U151 ( .A(n174), .B(i_data_rt[20]), .Q(n137) );
  AOI222 U152 ( .A(i_data_lwM[6]), .B(n18), .C(n62), .D(i_data_lwW[6]), .Q(n88) );
  NAND22 U153 ( .A(i_data_rt[29]), .B(n174), .Q(n167) );
  INV6 U154 ( .A(n47), .Q(n48) );
  AOI222 U155 ( .A(i_data_lwM[16]), .B(n18), .C(n60), .D(i_data_lwW[16]), .Q(
        n122) );
  NAND24 U156 ( .A(i_data_rt[16]), .B(n120), .Q(n121) );
  AOI222 U157 ( .A(n18), .B(i_data_lwM[2]), .C(n61), .D(i_data_lwW[2]), .Q(n73) );
  BUF15 U158 ( .A(n57), .Q(n46) );
  AOI222 U159 ( .A(i_data_lwM[13]), .B(n18), .C(n25), .D(i_data_lwW[13]), .Q(
        n112) );
  INV6 U160 ( .A(n38), .Q(n39) );
  AOI222 U161 ( .A(n26), .B(i_data_lwM[21]), .C(i_data_alures[21]), .D(n175), 
        .Q(n142) );
  AOI221 U162 ( .A(n26), .B(i_data_lwM[28]), .C(i_data_alures[28]), .D(n175), 
        .Q(n165) );
  AOI222 U163 ( .A(i_data_lwM[3]), .B(n176), .C(n10), .D(i_data_lwW[3]), .Q(
        n76) );
  INV6 U164 ( .A(n53), .Q(n28) );
  AOI222 U165 ( .A(n176), .B(i_data_lwM[0]), .C(n10), .D(i_data_lwW[0]), .Q(
        n67) );
  NAND20 U166 ( .A(i_data_alures[30]), .B(n19), .Q(n171) );
  INV6 U167 ( .A(n29), .Q(n30) );
  NAND34 U168 ( .A(n71), .B(n69), .C(n70), .Q(n49) );
  NAND24 U169 ( .A(n97), .B(n95), .Q(n40) );
  AOI222 U170 ( .A(n132), .B(i_data_writeres[8]), .C(i_data_alures[8]), .D(n19), .Q(n97) );
  AOI222 U171 ( .A(n173), .B(i_data_writeres[15]), .C(i_data_alures[15]), .D(
        n175), .Q(n119) );
  NAND22 U172 ( .A(i_con_fb[0]), .B(n94), .Q(n53) );
  NAND21 U173 ( .A(i_data_alures[31]), .B(n175), .Q(n178) );
  AOI221 U174 ( .A(n24), .B(i_data_writeres[28]), .C(n10), .D(i_data_lwW[28]), 
        .Q(n166) );
  NAND21 U175 ( .A(n19), .B(i_data_alures[19]), .Q(n135) );
  NAND34 U176 ( .A(n125), .B(n126), .C(n124), .Q(o_data_alusrb[17]) );
  AOI222 U177 ( .A(i_data_alures[1]), .B(n19), .C(n132), .D(i_data_writeres[1]), .Q(n69) );
  NAND28 U178 ( .A(n27), .B(n56), .Q(n64) );
  AOI222 U179 ( .A(n19), .B(i_data_alures[10]), .C(n26), .D(i_data_lwM[10]), 
        .Q(n102) );
  AOI221 U180 ( .A(n62), .B(i_data_lwW[29]), .C(i_data_lwM[29]), .D(n176), .Q(
        n169) );
  AOI221 U181 ( .A(i_data_alures[29]), .B(n19), .C(i_data_writeres[29]), .D(
        n173), .Q(n168) );
  AOI222 U182 ( .A(n132), .B(i_data_writeres[9]), .C(i_data_alures[9]), .D(n19), .Q(n100) );
  AOI222 U183 ( .A(n176), .B(i_data_lwM[15]), .C(n62), .D(i_data_lwW[15]), .Q(
        n118) );
  AOI222 U184 ( .A(n18), .B(i_data_lwM[18]), .C(n60), .D(i_data_lwW[18]), .Q(
        n128) );
  AOI222 U185 ( .A(i_data_lwM[8]), .B(n176), .C(n25), .D(i_data_lwW[8]), .Q(
        n96) );
  AOI222 U186 ( .A(n26), .B(i_data_lwM[9]), .C(i_data_lwW[9]), .D(n25), .Q(n99) );
  AOI222 U187 ( .A(n26), .B(i_data_lwM[14]), .C(n25), .D(i_data_lwW[14]), .Q(
        n115) );
  AOI222 U188 ( .A(n176), .B(i_data_lwM[11]), .C(n25), .D(i_data_lwW[11]), .Q(
        n106) );
  NAND24 U189 ( .A(n100), .B(n98), .Q(n29) );
  AOI222 U190 ( .A(n24), .B(i_data_writeres[26]), .C(n60), .D(i_data_lwW[26]), 
        .Q(n160) );
  INV6 U191 ( .A(n33), .Q(n34) );
  NAND28 U192 ( .A(n35), .B(n21), .Q(n37) );
  NAND28 U193 ( .A(n36), .B(n37), .Q(n104) );
  AOI222 U194 ( .A(n24), .B(i_data_writeres[22]), .C(n61), .D(i_data_lwW[22]), 
        .Q(n146) );
  NAND31 U195 ( .A(i_con_fb[0]), .B(n130), .C(n94), .Q(n78) );
  AOI221 U196 ( .A(n24), .B(i_data_writeres[24]), .C(n62), .D(i_data_lwW[24]), 
        .Q(n152) );
  AOI222 U197 ( .A(i_data_lwM[24]), .B(n18), .C(i_data_alures[24]), .D(n175), 
        .Q(n151) );
  NAND22 U198 ( .A(n131), .B(n94), .Q(n55) );
  AOI222 U199 ( .A(i_data_writeres[11]), .B(n132), .C(i_data_alures[11]), .D(
        n19), .Q(n107) );
  AOI222 U200 ( .A(n24), .B(i_data_writeres[21]), .C(n62), .D(i_data_lwW[21]), 
        .Q(n143) );
  AOI221 U201 ( .A(n132), .B(i_data_writeres[3]), .C(i_data_alures[3]), .D(n19), .Q(n77) );
  NAND22 U202 ( .A(n17), .B(i_data_rt[2]), .Q(n72) );
  NAND22 U203 ( .A(i_data_rt[3]), .B(n17), .Q(n75) );
  NAND22 U204 ( .A(i_data_rt[5]), .B(n46), .Q(n84) );
  AOI222 U205 ( .A(n2), .B(i_data_writeres[10]), .C(n61), .D(i_data_lwW[10]), 
        .Q(n103) );
  AOI222 U206 ( .A(n2), .B(i_data_writeres[17]), .C(n61), .D(i_data_lwW[17]), 
        .Q(n126) );
  AOI222 U207 ( .A(i_data_alures[17]), .B(n175), .C(i_data_lwM[17]), .D(n176), 
        .Q(n125) );
  AOI222 U208 ( .A(i_data_writeres[18]), .B(n24), .C(i_data_alures[18]), .D(
        n175), .Q(n129) );
  AOI222 U209 ( .A(n18), .B(i_data_lwM[19]), .C(n60), .D(i_data_lwW[19]), .Q(
        n134) );
  NAND22 U210 ( .A(i_data_rt[27]), .B(n46), .Q(n161) );
  NAND33 U211 ( .A(n172), .B(n171), .C(n170), .Q(o_data_alusrb[30]) );
endmodule


module E_alubmux ( i_data_fb, i_data_imm, i_con_imm, o_data_alub );
  input [31:0] i_data_fb;
  input [31:0] i_data_imm;
  output [31:0] o_data_alub;
  input i_con_imm;
  wire   n2, n3, n5, n6, n8, n9, n11, n12, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66;

  CLKIN12 U1 ( .A(n37), .Q(o_data_alub[5]) );
  INV12 U2 ( .A(n30), .Q(o_data_alub[2]) );
  INV8 U3 ( .A(n27), .Q(o_data_alub[1]) );
  CLKIN6 U4 ( .A(n51), .Q(o_data_alub[17]) );
  CLKIN6 U5 ( .A(n52), .Q(o_data_alub[18]) );
  CLKIN6 U6 ( .A(n66), .Q(o_data_alub[31]) );
  AOI222 U7 ( .A(i_data_fb[31]), .B(n20), .C(i_data_imm[31]), .D(n16), .Q(n66)
         );
  AOI222 U8 ( .A(i_data_fb[18]), .B(n20), .C(i_data_imm[18]), .D(n15), .Q(n52)
         );
  CLKIN15 U9 ( .A(n36), .Q(o_data_alub[4]) );
  BUF12 U10 ( .A(n23), .Q(n18) );
  CLKIN6 U11 ( .A(n48), .Q(o_data_alub[16]) );
  CLKIN6 U12 ( .A(i_data_fb[9]), .Q(n12) );
  INV3 U13 ( .A(n28), .Q(n29) );
  INV12 U14 ( .A(n38), .Q(o_data_alub[6]) );
  INV6 U15 ( .A(n42), .Q(o_data_alub[10]) );
  CLKIN12 U16 ( .A(n33), .Q(o_data_alub[3]) );
  AOI222 U17 ( .A(i_data_fb[20]), .B(n20), .C(i_data_imm[20]), .D(n15), .Q(n56) );
  AOI222 U18 ( .A(i_data_fb[29]), .B(n19), .C(i_data_imm[29]), .D(n15), .Q(n64) );
  AOI222 U19 ( .A(i_data_fb[25]), .B(n19), .C(i_data_imm[25]), .D(n15), .Q(n61) );
  AOI222 U20 ( .A(i_data_fb[21]), .B(n20), .C(i_data_imm[21]), .D(n15), .Q(n57) );
  AOI222 U21 ( .A(i_data_fb[23]), .B(n20), .C(i_data_imm[23]), .D(n15), .Q(n59) );
  AOI222 U22 ( .A(n19), .B(i_data_fb[27]), .C(i_data_imm[27]), .D(n15), .Q(n62) );
  AOI222 U23 ( .A(i_data_fb[0]), .B(n19), .C(i_data_imm[0]), .D(n15), .Q(n24)
         );
  INV3 U24 ( .A(i_data_imm[13]), .Q(n9) );
  INV3 U25 ( .A(n53), .Q(n54) );
  INV3 U26 ( .A(i_data_imm[26]), .Q(n3) );
  INV3 U27 ( .A(i_data_imm[11]), .Q(n6) );
  INV6 U28 ( .A(n18), .Q(n17) );
  CLKIN6 U29 ( .A(n45), .Q(o_data_alub[15]) );
  INV12 U30 ( .A(n39), .Q(o_data_alub[7]) );
  CLKIN6 U31 ( .A(n62), .Q(o_data_alub[27]) );
  BUF2 U32 ( .A(n18), .Q(n21) );
  INV6 U33 ( .A(n18), .Q(n16) );
  BUF2 U34 ( .A(n23), .Q(n19) );
  INV3 U35 ( .A(n19), .Q(n11) );
  INV6 U36 ( .A(n55), .Q(o_data_alub[19]) );
  CLKIN6 U37 ( .A(n40), .Q(o_data_alub[8]) );
  INV6 U38 ( .A(i_data_fb[12]), .Q(n14) );
  CLKIN6 U39 ( .A(i_data_fb[13]), .Q(n8) );
  CLKIN12 U40 ( .A(n60), .Q(o_data_alub[24]) );
  CLKIN6 U41 ( .A(n63), .Q(o_data_alub[28]) );
  CLKIN6 U42 ( .A(i_con_imm), .Q(n23) );
  CLKIN6 U43 ( .A(n24), .Q(o_data_alub[0]) );
  CLKIN6 U44 ( .A(n65), .Q(o_data_alub[30]) );
  CLKIN6 U45 ( .A(n64), .Q(o_data_alub[29]) );
  INV6 U46 ( .A(i_data_fb[26]), .Q(n2) );
  NAND20 U47 ( .A(i_data_imm[1]), .B(n17), .Q(n25) );
  OAI222 U48 ( .A(n2), .B(n11), .C(n3), .D(n18), .Q(o_data_alub[26]) );
  NAND21 U49 ( .A(i_data_imm[3]), .B(n17), .Q(n31) );
  CLKIN6 U50 ( .A(n59), .Q(o_data_alub[23]) );
  CLKIN6 U51 ( .A(n61), .Q(o_data_alub[25]) );
  INV2 U52 ( .A(n31), .Q(n32) );
  INV6 U53 ( .A(i_data_fb[11]), .Q(n5) );
  CLKIN6 U54 ( .A(n44), .Q(o_data_alub[14]) );
  OAI222 U55 ( .A(n5), .B(n15), .C(n6), .D(n18), .Q(o_data_alub[11]) );
  OAI222 U56 ( .A(n8), .B(n16), .C(n9), .D(n18), .Q(o_data_alub[13]) );
  AOI222 U57 ( .A(i_data_fb[30]), .B(n19), .C(i_data_imm[30]), .D(n15), .Q(n65) );
  CLKIN6 U58 ( .A(n58), .Q(o_data_alub[22]) );
  CLKIN6 U59 ( .A(n57), .Q(o_data_alub[21]) );
  AOI222 U60 ( .A(n21), .B(i_data_fb[14]), .C(i_data_imm[14]), .D(n16), .Q(n44) );
  AOI222 U61 ( .A(i_data_fb[8]), .B(n21), .C(i_data_imm[8]), .D(n16), .Q(n40)
         );
  NAND20 U62 ( .A(i_data_imm[2]), .B(n17), .Q(n28) );
  CLKIN6 U63 ( .A(n56), .Q(o_data_alub[20]) );
  AOI222 U64 ( .A(i_data_fb[24]), .B(n19), .C(i_data_imm[24]), .D(n15), .Q(n60) );
  AOI222 U65 ( .A(n41), .B(n11), .C(n12), .D(n41), .Q(o_data_alub[9]) );
  AOI222 U66 ( .A(n14), .B(n43), .C(n43), .D(n16), .Q(o_data_alub[12]) );
  INV3 U67 ( .A(n18), .Q(n15) );
  BUF2 U68 ( .A(n23), .Q(n20) );
  BUF2 U69 ( .A(n18), .Q(n22) );
  CLKIN3 U70 ( .A(n25), .Q(n26) );
  OAI222 U71 ( .A(n26), .B(n22), .C(i_data_fb[1]), .D(n26), .Q(n27) );
  OAI222 U72 ( .A(n29), .B(n21), .C(i_data_fb[2]), .D(n29), .Q(n30) );
  OAI222 U73 ( .A(i_data_fb[3]), .B(n32), .C(n32), .D(n22), .Q(n33) );
  NAND22 U74 ( .A(i_data_imm[4]), .B(n17), .Q(n34) );
  CLKIN3 U75 ( .A(n34), .Q(n35) );
  OAI222 U76 ( .A(i_data_fb[4]), .B(n35), .C(n35), .D(n22), .Q(n36) );
  AOI222 U77 ( .A(i_data_fb[5]), .B(n22), .C(i_data_imm[5]), .D(n16), .Q(n37)
         );
  AOI222 U78 ( .A(i_data_fb[6]), .B(n22), .C(i_data_imm[6]), .D(n16), .Q(n38)
         );
  AOI222 U79 ( .A(i_data_fb[7]), .B(n21), .C(i_data_imm[7]), .D(n16), .Q(n39)
         );
  NAND22 U80 ( .A(i_data_imm[9]), .B(n16), .Q(n41) );
  AOI222 U81 ( .A(i_data_fb[10]), .B(n21), .C(i_data_imm[10]), .D(n16), .Q(n42) );
  NAND22 U82 ( .A(i_data_imm[12]), .B(n16), .Q(n43) );
  AOI222 U83 ( .A(n21), .B(i_data_fb[15]), .C(i_data_imm[15]), .D(n16), .Q(n45) );
  NAND22 U84 ( .A(i_data_imm[16]), .B(n16), .Q(n46) );
  CLKIN3 U85 ( .A(n46), .Q(n47) );
  OAI222 U86 ( .A(i_data_fb[16]), .B(n47), .C(n47), .D(n20), .Q(n48) );
  NAND22 U87 ( .A(i_data_imm[17]), .B(n17), .Q(n49) );
  CLKIN3 U88 ( .A(n49), .Q(n50) );
  OAI222 U89 ( .A(n50), .B(n20), .C(i_data_fb[17]), .D(n50), .Q(n51) );
  NAND22 U90 ( .A(i_data_imm[19]), .B(n17), .Q(n53) );
  OAI222 U91 ( .A(i_data_fb[19]), .B(n54), .C(n54), .D(n20), .Q(n55) );
  AOI222 U92 ( .A(n20), .B(i_data_fb[22]), .C(i_data_imm[22]), .D(n15), .Q(n58) );
  AOI222 U93 ( .A(i_data_fb[28]), .B(n19), .C(i_data_imm[28]), .D(n15), .Q(n63) );
endmodule


module E_rdmux ( i_data_rtE, i_data_rdE, i_con_regdst, i_con_aluPC4, 
        o_data_writeE );
  input [4:0] i_data_rtE;
  input [4:0] i_data_rdE;
  output [4:0] o_data_writeE;
  input i_con_regdst, i_con_aluPC4;
  wire   n7, n8, n9, n10, n11, n1, n2, n3, n4, n5, n6, n12;

  CLKBU12 U2 ( .A(i_con_regdst), .Q(n1) );
  INV3 U3 ( .A(i_con_aluPC4), .Q(n12) );
  NAND22 U4 ( .A(i_data_rdE[3]), .B(n1), .Q(n8) );
  NAND22 U5 ( .A(i_data_rdE[0]), .B(n1), .Q(n11) );
  NAND22 U6 ( .A(i_data_rdE[1]), .B(n1), .Q(n10) );
  NAND22 U7 ( .A(i_data_rdE[2]), .B(n1), .Q(n9) );
  OAI2110 U8 ( .A(n1), .B(n2), .C(n12), .D(n7), .Q(o_data_writeE[4]) );
  NAND20 U9 ( .A(i_data_rdE[4]), .B(n1), .Q(n7) );
  OAI2111 U10 ( .A(n1), .B(n6), .C(n12), .D(n11), .Q(o_data_writeE[0]) );
  CLKIN3 U11 ( .A(i_data_rtE[0]), .Q(n6) );
  OAI2111 U12 ( .A(n1), .B(n5), .C(n12), .D(n10), .Q(o_data_writeE[1]) );
  CLKIN3 U13 ( .A(i_data_rtE[1]), .Q(n5) );
  OAI2111 U14 ( .A(n1), .B(n4), .C(n12), .D(n9), .Q(o_data_writeE[2]) );
  CLKIN3 U15 ( .A(i_data_rtE[2]), .Q(n4) );
  INV3 U16 ( .A(i_data_rtE[4]), .Q(n2) );
  OAI2111 U17 ( .A(n1), .B(n3), .C(n12), .D(n8), .Q(o_data_writeE[3]) );
  CLKIN3 U18 ( .A(i_data_rtE[3]), .Q(n3) );
endmodule


module D_compare_DW01_cmp6_4 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162;

  NAND26 U1 ( .A(n97), .B(A[19]), .Q(n100) );
  NAND23 U2 ( .A(n47), .B(A[5]), .Q(n50) );
  NAND24 U3 ( .A(n49), .B(n50), .Q(n140) );
  NAND22 U4 ( .A(B[23]), .B(n65), .Q(n66) );
  NAND22 U5 ( .A(B[14]), .B(n36), .Q(n37) );
  NAND22 U6 ( .A(B[2]), .B(n94), .Q(n95) );
  INV3 U7 ( .A(n81), .Q(n22) );
  NAND24 U8 ( .A(B[28]), .B(n6), .Q(n7) );
  CLKIN6 U9 ( .A(A[28]), .Q(n6) );
  NAND23 U10 ( .A(n93), .B(A[2]), .Q(n96) );
  NOR23 U11 ( .A(n112), .B(n111), .Q(n107) );
  NAND26 U12 ( .A(n71), .B(n72), .Q(n153) );
  CLKIN3 U13 ( .A(B[23]), .Q(n64) );
  CLKIN12 U14 ( .A(A[5]), .Q(n48) );
  NOR23 U15 ( .A(n148), .B(n147), .Q(n143) );
  NAND22 U16 ( .A(B[27]), .B(n24), .Q(n25) );
  CLKIN10 U17 ( .A(A[29]), .Q(n52) );
  NAND26 U18 ( .A(n51), .B(A[29]), .Q(n54) );
  NAND22 U19 ( .A(n9), .B(A[17]), .Q(n12) );
  NAND24 U20 ( .A(B[13]), .B(n70), .Q(n71) );
  CLKIN12 U21 ( .A(A[13]), .Q(n70) );
  NAND23 U22 ( .A(n81), .B(A[21]), .Q(n84) );
  CLKIN4 U23 ( .A(A[21]), .Q(n82) );
  NAND24 U24 ( .A(B[11]), .B(n32), .Q(n33) );
  NAND22 U25 ( .A(A[20]), .B(n2), .Q(n3) );
  NAND22 U26 ( .A(n1), .B(B[20]), .Q(n4) );
  NAND24 U27 ( .A(n3), .B(n4), .Q(n118) );
  INV2 U28 ( .A(A[20]), .Q(n1) );
  INV3 U29 ( .A(B[20]), .Q(n2) );
  NOR24 U30 ( .A(n117), .B(n118), .Q(n113) );
  NAND28 U31 ( .A(n27), .B(A[22]), .Q(n30) );
  CLKIN12 U32 ( .A(B[22]), .Q(n27) );
  NAND24 U33 ( .A(n55), .B(A[24]), .Q(n58) );
  NAND28 U34 ( .A(n33), .B(n34), .Q(n161) );
  NAND24 U35 ( .A(n31), .B(A[11]), .Q(n34) );
  INV2 U36 ( .A(B[10]), .Q(n85) );
  NAND24 U37 ( .A(n35), .B(A[14]), .Q(n38) );
  CLKIN4 U38 ( .A(A[17]), .Q(n10) );
  CLKIN3 U39 ( .A(A[10]), .Q(n86) );
  NAND24 U40 ( .A(n11), .B(n12), .Q(n115) );
  NAND23 U41 ( .A(B[22]), .B(n28), .Q(n29) );
  CLKIN12 U42 ( .A(A[6]), .Q(n14) );
  NAND24 U43 ( .A(n13), .B(A[6]), .Q(n16) );
  NAND28 U44 ( .A(n75), .B(n76), .Q(n129) );
  NAND23 U45 ( .A(n77), .B(A[26]), .Q(n80) );
  NAND28 U46 ( .A(n15), .B(n16), .Q(n141) );
  NAND23 U47 ( .A(n39), .B(A[7]), .Q(n42) );
  NAND28 U48 ( .A(n99), .B(n100), .Q(n117) );
  NAND24 U49 ( .A(B[6]), .B(n14), .Q(n15) );
  NAND28 U50 ( .A(n29), .B(n30), .Q(n110) );
  NAND28 U51 ( .A(n53), .B(n54), .Q(n123) );
  NAND26 U52 ( .A(n43), .B(A[0]), .Q(n46) );
  NOR24 U53 ( .A(n115), .B(n116), .Q(n114) );
  CLKIN12 U54 ( .A(A[22]), .Q(n28) );
  NAND24 U55 ( .A(n121), .B(n122), .Q(n120) );
  NAND23 U56 ( .A(B[5]), .B(n48), .Q(n49) );
  CLKIN4 U57 ( .A(A[0]), .Q(n44) );
  NAND22 U58 ( .A(B[8]), .B(n90), .Q(n91) );
  CLKIN4 U59 ( .A(A[8]), .Q(n90) );
  CLKIN10 U60 ( .A(A[4]), .Q(n61) );
  NAND24 U61 ( .A(n85), .B(A[10]), .Q(n88) );
  NAND24 U62 ( .A(B[29]), .B(n52), .Q(n53) );
  NAND28 U63 ( .A(n133), .B(n134), .Q(n101) );
  NAND23 U64 ( .A(B[19]), .B(n98), .Q(n99) );
  NAND26 U65 ( .A(A[13]), .B(n69), .Q(n72) );
  CLKIN6 U66 ( .A(B[11]), .Q(n31) );
  NAND22 U67 ( .A(B[26]), .B(n78), .Q(n79) );
  NAND24 U68 ( .A(n127), .B(n128), .Q(n119) );
  NAND22 U69 ( .A(n23), .B(A[27]), .Q(n26) );
  NAND22 U70 ( .A(B[4]), .B(n61), .Q(n62) );
  INV3 U71 ( .A(B[12]), .Q(n17) );
  NAND22 U72 ( .A(n21), .B(n86), .Q(n87) );
  INV3 U73 ( .A(A[3]), .Q(n68) );
  INV3 U74 ( .A(B[18]), .Q(n59) );
  NAND23 U75 ( .A(n5), .B(A[28]), .Q(n8) );
  NAND24 U76 ( .A(n7), .B(n8), .Q(n132) );
  CLKIN3 U77 ( .A(B[28]), .Q(n5) );
  NOR24 U78 ( .A(n131), .B(n132), .Q(n127) );
  NAND21 U79 ( .A(B[17]), .B(n10), .Q(n11) );
  INV1 U80 ( .A(B[17]), .Q(n9) );
  NAND24 U81 ( .A(B[0]), .B(n44), .Q(n45) );
  INV6 U82 ( .A(B[6]), .Q(n13) );
  NOR24 U83 ( .A(n141), .B(n142), .Q(n137) );
  CLKIN6 U84 ( .A(A[14]), .Q(n36) );
  XNR22 U85 ( .A(n17), .B(A[12]), .Q(n162) );
  CLKIN6 U86 ( .A(B[0]), .Q(n43) );
  NAND21 U87 ( .A(n59), .B(A[18]), .Q(n19) );
  NAND26 U88 ( .A(B[18]), .B(n18), .Q(n20) );
  NAND24 U89 ( .A(n19), .B(n20), .Q(n116) );
  CLKIN6 U90 ( .A(A[18]), .Q(n18) );
  CLKIN12 U91 ( .A(A[7]), .Q(n40) );
  NAND28 U92 ( .A(n45), .B(n46), .Q(n145) );
  CLKIN3 U93 ( .A(n85), .Q(n21) );
  NOR23 U94 ( .A(n161), .B(n162), .Q(n157) );
  INV3 U95 ( .A(A[23]), .Q(n65) );
  NAND24 U96 ( .A(n64), .B(A[23]), .Q(n67) );
  CLKIN3 U97 ( .A(B[4]), .Q(n60) );
  NOR22 U98 ( .A(n156), .B(n155), .Q(n151) );
  CLKIN6 U99 ( .A(B[24]), .Q(n55) );
  NAND24 U100 ( .A(n103), .B(n104), .Q(n102) );
  NAND24 U101 ( .A(n57), .B(n58), .Q(n112) );
  CLKIN6 U102 ( .A(B[14]), .Q(n35) );
  NAND22 U103 ( .A(B[7]), .B(n40), .Q(n41) );
  INV2 U104 ( .A(B[29]), .Q(n51) );
  INV3 U105 ( .A(B[25]), .Q(n73) );
  CLKIN3 U106 ( .A(B[2]), .Q(n93) );
  INV2 U107 ( .A(B[21]), .Q(n81) );
  NAND24 U108 ( .A(n25), .B(n26), .Q(n131) );
  CLKIN6 U109 ( .A(B[27]), .Q(n23) );
  INV1 U110 ( .A(A[27]), .Q(n24) );
  NAND24 U111 ( .A(n73), .B(A[25]), .Q(n76) );
  CLKIN6 U112 ( .A(A[11]), .Q(n32) );
  NAND24 U113 ( .A(n60), .B(A[4]), .Q(n63) );
  NAND24 U114 ( .A(n79), .B(n80), .Q(n130) );
  NAND22 U115 ( .A(B[25]), .B(n74), .Q(n75) );
  NAND24 U116 ( .A(n37), .B(n38), .Q(n154) );
  NAND24 U117 ( .A(n41), .B(n42), .Q(n142) );
  INV1 U118 ( .A(B[7]), .Q(n39) );
  NOR24 U119 ( .A(n145), .B(n146), .Q(n144) );
  NAND22 U120 ( .A(n89), .B(A[8]), .Q(n92) );
  NAND24 U121 ( .A(n91), .B(n92), .Q(n159) );
  INV1 U122 ( .A(B[5]), .Q(n47) );
  NOR24 U123 ( .A(n139), .B(n140), .Q(n138) );
  NOR24 U124 ( .A(n123), .B(n124), .Q(n122) );
  NAND24 U125 ( .A(n157), .B(n158), .Q(n149) );
  NAND22 U126 ( .A(B[24]), .B(n56), .Q(n57) );
  CLKIN6 U127 ( .A(A[24]), .Q(n56) );
  NAND24 U128 ( .A(n62), .B(n63), .Q(n139) );
  CLKIN6 U129 ( .A(B[13]), .Q(n69) );
  CLKIN1 U130 ( .A(A[26]), .Q(n78) );
  NOR24 U131 ( .A(n109), .B(n110), .Q(n108) );
  INV3 U132 ( .A(B[19]), .Q(n97) );
  NAND24 U133 ( .A(n66), .B(n67), .Q(n111) );
  XOR22 U134 ( .A(B[16]), .B(A[16]), .Q(n156) );
  NAND22 U135 ( .A(n22), .B(n82), .Q(n83) );
  XNR22 U136 ( .A(B[3]), .B(n68), .Q(n148) );
  XOR22 U137 ( .A(B[15]), .B(A[15]), .Q(n155) );
  CLKIN6 U138 ( .A(A[25]), .Q(n74) );
  NOR24 U139 ( .A(n153), .B(n154), .Q(n152) );
  CLKIN0 U140 ( .A(B[8]), .Q(n89) );
  NAND24 U141 ( .A(n95), .B(n96), .Q(n146) );
  NAND24 U142 ( .A(n83), .B(n84), .Q(n109) );
  CLKIN6 U143 ( .A(B[26]), .Q(n77) );
  NOR24 U144 ( .A(n119), .B(n120), .Q(n103) );
  NOR24 U145 ( .A(n129), .B(n130), .Q(n128) );
  NAND24 U146 ( .A(n87), .B(n88), .Q(n160) );
  NOR24 U147 ( .A(n105), .B(n106), .Q(n104) );
  NOR24 U148 ( .A(n160), .B(n159), .Q(n158) );
  CLKIN6 U149 ( .A(A[2]), .Q(n94) );
  NAND24 U150 ( .A(n151), .B(n152), .Q(n150) );
  NOR23 U151 ( .A(n126), .B(n125), .Q(n121) );
  NAND24 U152 ( .A(n113), .B(n114), .Q(n105) );
  NAND24 U153 ( .A(n107), .B(n108), .Q(n106) );
  XOR21 U154 ( .A(B[1]), .B(A[1]), .Q(n147) );
  CLKIN6 U155 ( .A(A[19]), .Q(n98) );
  XOR22 U156 ( .A(B[9]), .B(A[9]), .Q(n124) );
  NAND24 U157 ( .A(n143), .B(n144), .Q(n135) );
  NOR24 U158 ( .A(n101), .B(n102), .Q(EQ) );
  XOR22 U159 ( .A(B[31]), .B(A[31]), .Q(n126) );
  XOR22 U160 ( .A(B[30]), .B(A[30]), .Q(n125) );
  NOR24 U161 ( .A(n135), .B(n136), .Q(n134) );
  NAND24 U162 ( .A(n137), .B(n138), .Q(n136) );
  NOR24 U163 ( .A(n150), .B(n149), .Q(n133) );
endmodule


module D_compare ( o_con_ifbranch, i_data_rs, i_data_rt, i_con_bop );
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [2:0] i_con_bop;
  output o_con_ifbranch;
  wire   equal, n3, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16;

  D_compare_DW01_cmp6_4 eq_34 ( .A(i_data_rs), .B(i_data_rt), .TC(n3), .EQ(
        equal) );
  CLKIN4 U2 ( .A(i_data_rs[31]), .Q(n5) );
  CLKIN4 U3 ( .A(equal), .Q(n9) );
  AOI2111 U4 ( .A(i_con_bop[1]), .B(n13), .C(n12), .D(n11), .Q(n14) );
  NOR21 U5 ( .A(n8), .B(n13), .Q(n16) );
  NOR21 U6 ( .A(n16), .B(n14), .Q(n1) );
  NOR24 U7 ( .A(n2), .B(n15), .Q(o_con_ifbranch) );
  INV3 U8 ( .A(n1), .Q(n2) );
  CLKIN1 U9 ( .A(n10), .Q(n12) );
  INV3 U10 ( .A(i_con_bop[2]), .Q(n13) );
  LOGIC0 U11 ( .Q(n3) );
  XNR21 U12 ( .A(i_con_bop[1]), .B(i_con_bop[2]), .Q(n4) );
  OAI212 U13 ( .A(n4), .B(n5), .C(i_con_bop[0]), .Q(n8) );
  CLKIN3 U14 ( .A(i_con_bop[1]), .Q(n7) );
  NAND22 U15 ( .A(i_con_bop[2]), .B(n5), .Q(n10) );
  CLKIN3 U16 ( .A(i_con_bop[0]), .Q(n6) );
  OAI212 U17 ( .A(n7), .B(n10), .C(n6), .Q(n11) );
  OAI222 U18 ( .A(n9), .B(n11), .C(equal), .D(n8), .Q(n15) );
endmodule


module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Efamux, i_con_Efbmux, 
        i_con_Ealuop, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread, 
        i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_bop, o_data_pc4, o_data_alures, o_data_rt, o_addr_regdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_addr_Erd, o_addr_Mrt, o_con_ifbranch );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [5:0] i_con_Ealuop;
  input [2:0] i_con_bop;
  output [31:0] o_data_pc4;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80;
  wire   [31:0] alu_o_data_AluRes;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;

  DFC3 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[0]) );
  DFC3 pipe_rt_reg_30_ ( .D(n21), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC3 pipe_rt_reg_28_ ( .D(n13), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28]) );
  DFC3 pipe_rt_reg_5_ ( .D(n43), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[5]) );
  DFC3 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  E_alu u_alu ( .o_data_AluRes(alu_o_data_AluRes), .i_data_A({
        compare_i_data_rs[31], n64, n72, compare_i_data_rs[28:26], n61, 
        compare_i_data_rs[24], n70, compare_i_data_rs[22], n15, 
        compare_i_data_rs[20:19], n67, n76, compare_i_data_rs[16], n49, n63, 
        compare_i_data_rs[13], n74, compare_i_data_rs[11:9], n16, n3, n39, n6, 
        compare_i_data_rs[4], n10, n54, n33, compare_i_data_rs[0]}), 
        .i_data_B(alu_i_data_B), .i_con_AluCtrl(alu_i_con_AluCtrl), 
        .i_data_shamt(i_data_immext[10:6]) );
  E_alu_control u_alu_control ( .o_con_AluCtrl(alu_i_con_AluCtrl), 
        .i_con_AluOp(i_con_Ealuop), .i_con_FuncCode(i_data_immext[5:0]) );
  E_famux5 u_famux5 ( .i_data_rs(i_data_rs), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fa(i_con_Efamux), .o_data_alusra(
        compare_i_data_rs) );
  E_fbmux5 u_fbmux ( .i_data_rt(i_data_rt), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fb(i_con_Efbmux), .o_data_alusrb(
        compare_i_data_rt) );
  E_alubmux u_alubmux ( .i_data_fb(compare_i_data_rt), .i_data_imm({
        i_data_immext[31:6], n1, i_data_immext[4:0]}), .i_con_imm(
        i_con_Ealusrc), .o_data_alub(alu_i_data_B) );
  E_rdmux u_rdmux ( .i_data_rtE(i_addr_rt), .i_data_rdE(i_addr_rd), 
        .i_con_regdst(i_con_Eregdst), .i_con_aluPC4(i_con_Malupc8), 
        .o_data_writeE(o_addr_Erd) );
  D_compare u_compare ( .o_con_ifbranch(o_con_ifbranch), .i_data_rs({
        compare_i_data_rs[31], n64, n72, compare_i_data_rs[28:26], n61, n30, 
        n70, compare_i_data_rs[22], n80, compare_i_data_rs[20:19], n11, 
        compare_i_data_rs[17:15], n63, compare_i_data_rs[13], n74, 
        compare_i_data_rs[11:9], n65, n59, n39, n56, compare_i_data_rs[4:3], 
        n54, compare_i_data_rs[1:0]}), .i_data_rt({compare_i_data_rt[31], n21, 
        compare_i_data_rt[29], n13, n9, n47, n8, n34, n44, n22, 
        compare_i_data_rt[21], n35, n24, n27, compare_i_data_rt[17], n78, n32, 
        n48, n50, n51, n42, compare_i_data_rt[10], n40, compare_i_data_rt[8:7], 
        n77, compare_i_data_rt[5], n19, n41, n29, compare_i_data_rt[1], n52}), 
        .i_con_bop(i_con_bop) );
  DFC1 pipe_rt_reg_11_ ( .D(n45), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11]) );
  DFC1 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC1 pipe_rt_reg_14_ ( .D(n48), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14]) );
  DFC1 pipe_rt_reg_3_ ( .D(n41), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[3]) );
  DFC1 pipe_rt_reg_8_ ( .D(n25), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[8]) );
  DFC1 pipe_rt_reg_1_ ( .D(n37), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[1]) );
  DFC1 pipe_rt_reg_27_ ( .D(n9), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27]) );
  DFC1 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC1 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC1 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC1 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC1 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC1 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC1 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC1 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC1 pipe_con_Malupc8_reg ( .D(i_con_Malupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Malupc8) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC1 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC1 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  DFC3 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC1 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC3 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC3 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC3 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC3 pipe_alures_reg_13_ ( .D(alu_o_data_AluRes[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[13]) );
  DFC1 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC1 pipe_rt_reg_22_ ( .D(n2), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC1 pipe_rt_reg_31_ ( .D(n5), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[31]) );
  DFC1 pipe_rt_reg_26_ ( .D(n4), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26]) );
  DFC1 pipe_rt_reg_9_ ( .D(n40), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[9]) );
  DFC1 pipe_rt_reg_19_ ( .D(n24), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19]) );
  DFC1 pipe_rt_reg_13_ ( .D(n50), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC1 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC1 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC1 pipe_rt_reg_2_ ( .D(n29), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[2]) );
  DFC1 pipe_rt_reg_0_ ( .D(n52), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[0]) );
  DFC1 pipe_rt_reg_12_ ( .D(n51), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12]) );
  DFC1 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC1 pipe_rt_reg_24_ ( .D(n34), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24]) );
  DFC1 pipe_alures_reg_14_ ( .D(alu_o_data_AluRes[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[14]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC1 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC1 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC1 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC1 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC1 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC1 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC1 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC1 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC1 pipe_alures_reg_15_ ( .D(alu_o_data_AluRes[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[15]) );
  DFC1 pipe_rt_reg_15_ ( .D(n32), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15]) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_rt_reg_10_ ( .D(n36), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC1 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC1 pipe_rt_reg_18_ ( .D(n27), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18]) );
  DFC1 pipe_rt_reg_25_ ( .D(n8), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25]) );
  DFC1 pipe_rt_reg_4_ ( .D(n19), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[4]) );
  DFC1 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC1 pipe_rt_reg_17_ ( .D(n17), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17]) );
  DFC1 pipe_rt_reg_6_ ( .D(n77), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[6]) );
  DFC1 pipe_rt_reg_21_ ( .D(n14), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21]) );
  DFC1 pipe_rt_reg_16_ ( .D(n78), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC1 pipe_rt_reg_23_ ( .D(n44), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23]) );
  DFC1 pipe_rt_reg_20_ ( .D(n35), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20]) );
  BUF6 U3 ( .A(compare_i_data_rt[6]), .Q(n77) );
  BUF6 U4 ( .A(compare_i_data_rt[0]), .Q(n52) );
  BUF6 U5 ( .A(compare_i_data_rt[3]), .Q(n41) );
  CLKBU4 U6 ( .A(compare_i_data_rt[14]), .Q(n48) );
  CLKIN2 U7 ( .A(compare_i_data_rt[2]), .Q(n28) );
  BUF6 U8 ( .A(compare_i_data_rt[24]), .Q(n34) );
  BUF2 U9 ( .A(i_data_immext[5]), .Q(n1) );
  INV12 U10 ( .A(compare_i_data_rs[5]), .Q(n55) );
  BUF2 U11 ( .A(n22), .Q(n2) );
  BUF4 U12 ( .A(compare_i_data_rt[11]), .Q(n42) );
  CLKIN2 U13 ( .A(compare_i_data_rt[25]), .Q(n7) );
  INV6 U14 ( .A(n28), .Q(n29) );
  CLKBU15 U15 ( .A(compare_i_data_rs[24]), .Q(n30) );
  INV6 U16 ( .A(compare_i_data_rs[23]), .Q(n69) );
  INV12 U17 ( .A(compare_i_data_rs[2]), .Q(n53) );
  CLKIN6 U18 ( .A(compare_i_data_rs[17]), .Q(n75) );
  CLKIN12 U19 ( .A(n58), .Q(n3) );
  INV12 U20 ( .A(n58), .Q(n59) );
  INV3 U21 ( .A(compare_i_data_rt[15]), .Q(n31) );
  INV12 U22 ( .A(n55), .Q(n56) );
  INV8 U23 ( .A(compare_i_data_rs[7]), .Q(n58) );
  BUF6 U24 ( .A(compare_i_data_rt[13]), .Q(n50) );
  BUF12 U25 ( .A(compare_i_data_rt[16]), .Q(n78) );
  CLKIN15 U26 ( .A(n75), .Q(n76) );
  BUF4 U27 ( .A(compare_i_data_rt[9]), .Q(n40) );
  BUF15 U28 ( .A(compare_i_data_rs[30]), .Q(n64) );
  CLKBU12 U29 ( .A(compare_i_data_rt[27]), .Q(n9) );
  BUF4 U30 ( .A(compare_i_data_rt[20]), .Q(n35) );
  CLKIN10 U31 ( .A(n79), .Q(n15) );
  INV8 U32 ( .A(n66), .Q(n67) );
  CLKIN12 U33 ( .A(n55), .Q(n6) );
  INV12 U34 ( .A(n57), .Q(n33) );
  INV12 U35 ( .A(n68), .Q(n10) );
  INV6 U36 ( .A(compare_i_data_rs[3]), .Q(n68) );
  INV3 U37 ( .A(n12), .Q(n13) );
  BUF15 U38 ( .A(compare_i_data_rs[15]), .Q(n49) );
  CLKBU12 U39 ( .A(compare_i_data_rs[8]), .Q(n16) );
  CLKIN6 U40 ( .A(n79), .Q(n80) );
  INV8 U41 ( .A(compare_i_data_rs[29]), .Q(n71) );
  INV10 U42 ( .A(compare_i_data_rs[14]), .Q(n62) );
  INV8 U43 ( .A(compare_i_data_rs[18]), .Q(n66) );
  INV6 U44 ( .A(compare_i_data_rs[25]), .Q(n60) );
  INV3 U45 ( .A(compare_i_data_rs[1]), .Q(n57) );
  BUF8 U46 ( .A(compare_i_data_rt[22]), .Q(n22) );
  BUF6 U47 ( .A(compare_i_data_rt[12]), .Q(n51) );
  CLKIN3 U48 ( .A(compare_i_data_rt[18]), .Q(n26) );
  INV3 U49 ( .A(n23), .Q(n24) );
  INV3 U50 ( .A(n7), .Q(n8) );
  BUF2 U51 ( .A(n47), .Q(n4) );
  BUF2 U52 ( .A(compare_i_data_rt[31]), .Q(n5) );
  CLKIN3 U53 ( .A(compare_i_data_rt[4]), .Q(n18) );
  CLKIN6 U54 ( .A(n20), .Q(n21) );
  CLKIN6 U55 ( .A(n66), .Q(n11) );
  INV2 U56 ( .A(compare_i_data_rt[28]), .Q(n12) );
  BUF2 U57 ( .A(compare_i_data_rt[21]), .Q(n14) );
  INV4 U58 ( .A(compare_i_data_rt[30]), .Q(n20) );
  INV15 U59 ( .A(n62), .Q(n63) );
  INV15 U60 ( .A(n69), .Q(n70) );
  INV10 U61 ( .A(compare_i_data_rs[21]), .Q(n79) );
  CLKIN2 U62 ( .A(compare_i_data_rt[19]), .Q(n23) );
  INV15 U63 ( .A(n71), .Q(n72) );
  CLKBU15 U64 ( .A(compare_i_data_rs[8]), .Q(n65) );
  BUF2 U65 ( .A(compare_i_data_rt[17]), .Q(n17) );
  CLKIN6 U66 ( .A(n18), .Q(n19) );
  CLKBU4 U67 ( .A(compare_i_data_rt[23]), .Q(n44) );
  CLKIN15 U68 ( .A(n53), .Q(n54) );
  BUF2 U69 ( .A(compare_i_data_rt[8]), .Q(n25) );
  CLKIN6 U70 ( .A(n26), .Q(n27) );
  CLKIN4 U71 ( .A(compare_i_data_rt[26]), .Q(n46) );
  CLKIN15 U72 ( .A(n73), .Q(n74) );
  INV6 U73 ( .A(n46), .Q(n47) );
  CLKIN6 U74 ( .A(n31), .Q(n32) );
  INV15 U75 ( .A(n60), .Q(n61) );
  BUF2 U76 ( .A(compare_i_data_rt[10]), .Q(n36) );
  BUF2 U77 ( .A(compare_i_data_rt[1]), .Q(n37) );
  INV6 U78 ( .A(compare_i_data_rs[6]), .Q(n38) );
  CLKIN15 U79 ( .A(n38), .Q(n39) );
  BUF2 U80 ( .A(compare_i_data_rt[5]), .Q(n43) );
  BUF2 U81 ( .A(n42), .Q(n45) );
  INV6 U82 ( .A(compare_i_data_rs[12]), .Q(n73) );
endmodule


module M_resmux ( i_data_alures, i_data_pc8, i_con_pc8, o_data_alu );
  input [31:0] i_data_alures;
  input [31:0] i_data_pc8;
  output [31:0] o_data_alu;
  input i_con_pc8;
  wire   n34, n35, n36, n37, n38, n39, n40, n43, n54, n63, n64, n65, n1, n2;

  INV3 U1 ( .A(n40), .Q(o_data_alu[3]) );
  INV3 U2 ( .A(n38), .Q(o_data_alu[5]) );
  INV3 U3 ( .A(n36), .Q(o_data_alu[7]) );
  INV3 U4 ( .A(n34), .Q(o_data_alu[9]) );
  INV3 U5 ( .A(n64), .Q(o_data_alu[10]) );
  MUX22 U6 ( .A(i_data_alures[14]), .B(i_data_pc8[14]), .S(n1), .Q(
        o_data_alu[14]) );
  MUX22 U7 ( .A(i_data_alures[18]), .B(i_data_pc8[18]), .S(n1), .Q(
        o_data_alu[18]) );
  MUX22 U8 ( .A(i_data_alures[19]), .B(i_data_pc8[19]), .S(n1), .Q(
        o_data_alu[19]) );
  MUX22 U9 ( .A(i_data_alures[22]), .B(i_data_pc8[22]), .S(i_con_pc8), .Q(
        o_data_alu[22]) );
  MUX22 U10 ( .A(i_data_alures[26]), .B(i_data_pc8[26]), .S(n1), .Q(
        o_data_alu[26]) );
  AOI220 U11 ( .A(i_data_alures[6]), .B(n2), .C(i_data_pc8[6]), .D(n1), .Q(n37) );
  MUX21 U12 ( .A(i_data_alures[23]), .B(i_data_pc8[23]), .S(i_con_pc8), .Q(
        o_data_alu[23]) );
  MUX21 U13 ( .A(i_data_alures[27]), .B(i_data_pc8[27]), .S(n1), .Q(
        o_data_alu[27]) );
  MUX21 U14 ( .A(i_data_alures[29]), .B(i_data_pc8[29]), .S(n1), .Q(
        o_data_alu[29]) );
  MUX21 U15 ( .A(i_data_alures[30]), .B(i_data_pc8[30]), .S(n1), .Q(
        o_data_alu[30]) );
  MUX21 U16 ( .A(i_data_alures[31]), .B(i_data_pc8[31]), .S(n1), .Q(
        o_data_alu[31]) );
  AOI220 U17 ( .A(i_data_alures[8]), .B(n2), .C(i_data_pc8[8]), .D(n1), .Q(n35) );
  MUX21 U18 ( .A(i_data_alures[15]), .B(i_data_pc8[15]), .S(i_con_pc8), .Q(
        o_data_alu[15]) );
  MUX21 U19 ( .A(i_data_alures[16]), .B(i_data_pc8[16]), .S(i_con_pc8), .Q(
        o_data_alu[16]) );
  MUX21 U20 ( .A(i_data_alures[20]), .B(i_data_pc8[20]), .S(i_con_pc8), .Q(
        o_data_alu[20]) );
  MUX21 U21 ( .A(i_data_alures[24]), .B(i_data_pc8[24]), .S(i_con_pc8), .Q(
        o_data_alu[24]) );
  MUX21 U22 ( .A(i_data_alures[28]), .B(i_data_pc8[28]), .S(n1), .Q(
        o_data_alu[28]) );
  AOI220 U23 ( .A(i_data_alures[11]), .B(n2), .C(i_data_pc8[11]), .D(n1), .Q(
        n63) );
  AOI220 U24 ( .A(i_data_alures[5]), .B(n2), .C(i_data_pc8[5]), .D(n1), .Q(n38) );
  AOI220 U25 ( .A(i_data_alures[10]), .B(n2), .C(i_data_pc8[10]), .D(n1), .Q(
        n64) );
  AOI220 U26 ( .A(i_data_alures[7]), .B(n2), .C(i_data_pc8[7]), .D(n1), .Q(n36) );
  AOI220 U27 ( .A(i_data_alures[9]), .B(n2), .C(i_data_pc8[9]), .D(n1), .Q(n34) );
  AOI220 U28 ( .A(i_data_alures[0]), .B(n2), .C(i_data_pc8[0]), .D(n1), .Q(n65) );
  AOI220 U29 ( .A(i_data_alures[1]), .B(n2), .C(i_data_pc8[1]), .D(n1), .Q(n54) );
  AOI220 U30 ( .A(i_data_alures[2]), .B(n2), .C(i_data_pc8[2]), .D(n1), .Q(n43) );
  AOI220 U31 ( .A(i_data_alures[4]), .B(n2), .C(i_data_pc8[4]), .D(n1), .Q(n39) );
  AOI220 U32 ( .A(i_data_alures[3]), .B(n2), .C(i_data_pc8[3]), .D(n1), .Q(n40) );
  INV3 U33 ( .A(n2), .Q(n1) );
  MUX22 U34 ( .A(i_data_alures[12]), .B(i_data_pc8[12]), .S(i_con_pc8), .Q(
        o_data_alu[12]) );
  INV3 U35 ( .A(n37), .Q(o_data_alu[6]) );
  INV3 U36 ( .A(n35), .Q(o_data_alu[8]) );
  INV3 U37 ( .A(n63), .Q(o_data_alu[11]) );
  MUX22 U38 ( .A(i_data_alures[13]), .B(i_data_pc8[13]), .S(i_con_pc8), .Q(
        o_data_alu[13]) );
  MUX22 U39 ( .A(i_data_alures[21]), .B(i_data_pc8[21]), .S(i_con_pc8), .Q(
        o_data_alu[21]) );
  MUX22 U40 ( .A(i_data_alures[25]), .B(i_data_pc8[25]), .S(n1), .Q(
        o_data_alu[25]) );
  INV3 U41 ( .A(i_con_pc8), .Q(n2) );
  INV3 U42 ( .A(n65), .Q(o_data_alu[0]) );
  INV3 U43 ( .A(n54), .Q(o_data_alu[1]) );
  INV3 U44 ( .A(n43), .Q(o_data_alu[2]) );
  INV3 U45 ( .A(n39), .Q(o_data_alu[4]) );
  MUX22 U46 ( .A(i_data_alures[17]), .B(i_data_pc8[17]), .S(i_con_pc8), .Q(
        o_data_alu[17]) );
endmodule


module mem_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  XOR21 U2 ( .A(n9), .B(n8), .Q(SUM[6]) );
  NOR21 U3 ( .A(n31), .B(n65), .Q(n66) );
  XNR21 U4 ( .A(A[12]), .B(n86), .Q(SUM[12]) );
  XNR21 U5 ( .A(n81), .B(n74), .Q(SUM[13]) );
  XNR21 U6 ( .A(n51), .B(n46), .Q(SUM[21]) );
  XNR21 U7 ( .A(n35), .B(n28), .Q(SUM[25]) );
  INV3 U8 ( .A(n31), .Q(n39) );
  INV3 U9 ( .A(n7), .Q(n9) );
  INV3 U10 ( .A(n96), .Q(n4) );
  NAND22 U11 ( .A(n97), .B(n98), .Q(n96) );
  NOR21 U12 ( .A(SUM[2]), .B(n102), .Q(n97) );
  NAND22 U13 ( .A(n64), .B(n39), .Q(n63) );
  NOR21 U14 ( .A(n65), .B(n60), .Q(n64) );
  NOR21 U15 ( .A(n10), .B(n12), .Q(n7) );
  NAND22 U16 ( .A(n7), .B(A[6]), .Q(n6) );
  NOR21 U17 ( .A(n73), .B(n74), .Q(n71) );
  NAND22 U18 ( .A(n51), .B(A[21]), .Q(n52) );
  NAND22 U19 ( .A(n35), .B(A[25]), .Q(n36) );
  NAND22 U20 ( .A(n81), .B(A[13]), .Q(n82) );
  NOR21 U21 ( .A(n63), .B(n61), .Q(n62) );
  NAND22 U22 ( .A(n67), .B(n68), .Q(n31) );
  NOR21 U23 ( .A(n69), .B(n70), .Q(n68) );
  NOR21 U24 ( .A(n75), .B(n76), .Q(n67) );
  NAND22 U25 ( .A(n71), .B(A[2]), .Q(n70) );
  INV3 U26 ( .A(n24), .Q(n23) );
  NAND31 U27 ( .A(n25), .B(n26), .C(n39), .Q(n24) );
  NOR31 U28 ( .A(n29), .B(n27), .C(n28), .Q(n26) );
  INV3 U29 ( .A(n94), .Q(n93) );
  NAND22 U30 ( .A(n95), .B(n4), .Q(n94) );
  NOR21 U31 ( .A(n2), .B(n5), .Q(n95) );
  INV3 U32 ( .A(n3), .Q(n1) );
  NAND22 U33 ( .A(A[8]), .B(n4), .Q(n3) );
  NOR21 U34 ( .A(n46), .B(n47), .Q(n50) );
  NOR21 U35 ( .A(n28), .B(n29), .Q(n34) );
  NOR21 U36 ( .A(n74), .B(n73), .Q(n80) );
  INV3 U37 ( .A(n75), .Q(n87) );
  NAND22 U38 ( .A(n42), .B(n43), .Q(n30) );
  NOR31 U39 ( .A(n47), .B(n45), .C(n46), .Q(n42) );
  NAND22 U40 ( .A(A[23]), .B(A[20]), .Q(n45) );
  NAND22 U41 ( .A(n57), .B(n58), .Q(n44) );
  NOR21 U42 ( .A(n60), .B(n61), .Q(n57) );
  INV3 U43 ( .A(n59), .Q(n58) );
  NAND22 U44 ( .A(A[19]), .B(A[16]), .Q(n59) );
  NAND31 U45 ( .A(A[12]), .B(A[15]), .C(A[3]), .Q(n76) );
  INV3 U46 ( .A(A[21]), .Q(n46) );
  INV3 U47 ( .A(A[25]), .Q(n28) );
  INV3 U48 ( .A(A[13]), .Q(n74) );
  NAND22 U49 ( .A(n99), .B(n100), .Q(n69) );
  NOR21 U50 ( .A(n77), .B(n101), .Q(n99) );
  NOR21 U51 ( .A(n10), .B(n8), .Q(n100) );
  INV3 U52 ( .A(A[7]), .Q(n101) );
  INV3 U53 ( .A(A[5]), .Q(n10) );
  INV3 U54 ( .A(A[10]), .Q(n91) );
  INV3 U55 ( .A(A[22]), .Q(n47) );
  INV3 U56 ( .A(A[26]), .Q(n29) );
  INV3 U57 ( .A(A[17]), .Q(n60) );
  INV3 U58 ( .A(A[18]), .Q(n61) );
  INV3 U59 ( .A(A[6]), .Q(n8) );
  INV3 U60 ( .A(A[9]), .Q(n2) );
  NAND22 U61 ( .A(A[27]), .B(A[24]), .Q(n27) );
  INV3 U62 ( .A(A[14]), .Q(n73) );
  NAND22 U63 ( .A(n87), .B(n4), .Q(n86) );
  INV3 U64 ( .A(n83), .Q(n81) );
  NAND22 U65 ( .A(n84), .B(n4), .Q(n83) );
  NOR21 U66 ( .A(n75), .B(n85), .Q(n84) );
  INV3 U67 ( .A(A[12]), .Q(n85) );
  INV3 U68 ( .A(n53), .Q(n51) );
  NAND22 U69 ( .A(n54), .B(n39), .Q(n53) );
  NOR21 U70 ( .A(n44), .B(n55), .Q(n54) );
  INV3 U71 ( .A(A[20]), .Q(n55) );
  INV3 U72 ( .A(n37), .Q(n35) );
  NAND22 U73 ( .A(n38), .B(n39), .Q(n37) );
  NOR21 U74 ( .A(n30), .B(n40), .Q(n38) );
  INV3 U75 ( .A(A[24]), .Q(n40) );
  INV3 U76 ( .A(n14), .Q(n13) );
  NAND22 U77 ( .A(A[3]), .B(A[2]), .Q(n14) );
  INV3 U78 ( .A(A[2]), .Q(SUM[2]) );
  XNR21 U79 ( .A(n66), .B(n60), .Q(SUM[17]) );
  INV3 U80 ( .A(n12), .Q(n11) );
  NAND22 U81 ( .A(A[4]), .B(n13), .Q(n12) );
  INV3 U82 ( .A(A[3]), .Q(n102) );
  INV3 U83 ( .A(A[4]), .Q(n77) );
  NAND22 U84 ( .A(n88), .B(n89), .Q(n75) );
  NOR21 U85 ( .A(n2), .B(n91), .Q(n88) );
  INV3 U86 ( .A(n90), .Q(n89) );
  NAND22 U87 ( .A(A[11]), .B(A[8]), .Q(n90) );
  XOR21 U88 ( .A(n36), .B(n29), .Q(SUM[26]) );
  XNR21 U89 ( .A(n1), .B(n2), .Q(SUM[9]) );
  XNR21 U90 ( .A(n11), .B(n10), .Q(SUM[5]) );
  XNR21 U91 ( .A(A[7]), .B(n6), .Q(SUM[7]) );
  XOR21 U92 ( .A(n4), .B(A[8]), .Q(SUM[8]) );
  XOR21 U93 ( .A(n92), .B(A[11]), .Q(SUM[11]) );
  NOR21 U94 ( .A(n91), .B(n94), .Q(n92) );
  XNR21 U95 ( .A(n93), .B(n91), .Q(SUM[10]) );
  XOR21 U96 ( .A(n39), .B(A[16]), .Q(SUM[16]) );
  XOR21 U97 ( .A(n78), .B(A[15]), .Q(SUM[15]) );
  NOR21 U98 ( .A(n83), .B(n79), .Q(n78) );
  INV3 U99 ( .A(n80), .Q(n79) );
  XOR21 U100 ( .A(n56), .B(A[20]), .Q(SUM[20]) );
  NOR21 U101 ( .A(n31), .B(n44), .Q(n56) );
  XOR21 U102 ( .A(n48), .B(A[23]), .Q(SUM[23]) );
  NOR21 U103 ( .A(n53), .B(n49), .Q(n48) );
  INV3 U104 ( .A(n50), .Q(n49) );
  XOR21 U105 ( .A(n41), .B(A[24]), .Q(SUM[24]) );
  NOR21 U106 ( .A(n31), .B(n30), .Q(n41) );
  XOR21 U107 ( .A(n32), .B(A[27]), .Q(SUM[27]) );
  NOR21 U108 ( .A(n37), .B(n33), .Q(n32) );
  INV3 U109 ( .A(n34), .Q(n33) );
  XOR21 U110 ( .A(n22), .B(A[29]), .Q(SUM[29]) );
  NOR21 U111 ( .A(n24), .B(n20), .Q(n22) );
  XOR21 U112 ( .A(n18), .B(A[30]), .Q(SUM[30]) );
  NOR21 U113 ( .A(n24), .B(n19), .Q(n18) );
  INV3 U114 ( .A(n17), .Q(n19) );
  XOR21 U115 ( .A(n15), .B(A[31]), .Q(SUM[31]) );
  NOR21 U116 ( .A(n24), .B(n16), .Q(n15) );
  NAND22 U117 ( .A(A[30]), .B(n17), .Q(n16) );
  XOR21 U118 ( .A(A[19]), .B(n62), .Q(SUM[19]) );
  XOR21 U119 ( .A(n23), .B(A[28]), .Q(SUM[28]) );
  XOR21 U120 ( .A(n82), .B(n73), .Q(SUM[14]) );
  XOR21 U121 ( .A(n52), .B(n47), .Q(SUM[22]) );
  XNR21 U122 ( .A(n63), .B(A[18]), .Q(SUM[18]) );
  NOR21 U123 ( .A(n20), .B(n21), .Q(n17) );
  INV3 U124 ( .A(A[29]), .Q(n21) );
  INV3 U125 ( .A(A[16]), .Q(n65) );
  INV3 U126 ( .A(A[28]), .Q(n20) );
  INV3 U127 ( .A(A[8]), .Q(n5) );
  XNR21 U128 ( .A(A[3]), .B(SUM[2]), .Q(SUM[3]) );
  XOR21 U129 ( .A(n13), .B(A[4]), .Q(SUM[4]) );
  CLKIN3 U130 ( .A(n30), .Q(n25) );
  CLKIN3 U131 ( .A(n44), .Q(n43) );
  CLKIN3 U132 ( .A(n69), .Q(n98) );
endmodule


module mem ( i_clk, i_nrst, i_data_pc4, i_data_alures, i_data_memout, 
        i_addr_regdst, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_FWmemread, i_addr_Mrt, o_data_alures, o_data_memout, 
        o_addr_regdst, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread, 
        o_addr_Wrt );
  input [31:0] i_data_pc4;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [4:0] i_addr_regdst;
  input [4:0] i_addr_Mrt;
  output [31:0] o_data_alures;
  output [31:0] o_data_memout;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Wrt;
  input i_clk, i_nrst, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite,
         i_con_FWmemread;
  output o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread;
  wire   n_Logic1_, n_Logic0_;
  wire   [31:0] pc8;
  wire   [31:0] resmux_o_data_alu;

  DFC3 pipe_rt_reg_4_ ( .D(i_addr_Mrt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(i_addr_Mrt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(i_addr_Mrt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[2]) );
  DFC3 pipe_rt_reg_0_ ( .D(i_addr_Mrt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[0]) );
  DFC3 pipe_data_alures_reg_31_ ( .D(resmux_o_data_alu[31]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[31]) );
  DFC3 pipe_data_alures_reg_30_ ( .D(resmux_o_data_alu[30]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[30]) );
  DFC3 pipe_data_alures_reg_29_ ( .D(resmux_o_data_alu[29]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[29]) );
  DFC3 pipe_data_alures_reg_28_ ( .D(resmux_o_data_alu[28]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[28]) );
  DFC3 pipe_data_alures_reg_27_ ( .D(resmux_o_data_alu[27]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[27]) );
  DFC3 pipe_data_alures_reg_26_ ( .D(resmux_o_data_alu[26]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[26]) );
  DFC3 pipe_data_alures_reg_25_ ( .D(resmux_o_data_alu[25]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[25]) );
  DFC3 pipe_data_alures_reg_24_ ( .D(resmux_o_data_alu[24]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[24]) );
  DFC3 pipe_data_alures_reg_23_ ( .D(resmux_o_data_alu[23]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[23]) );
  DFC3 pipe_data_alures_reg_22_ ( .D(resmux_o_data_alu[22]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[22]) );
  DFC3 pipe_data_alures_reg_21_ ( .D(resmux_o_data_alu[21]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[21]) );
  DFC3 pipe_data_alures_reg_20_ ( .D(resmux_o_data_alu[20]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[20]) );
  DFC3 pipe_data_alures_reg_19_ ( .D(resmux_o_data_alu[19]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[19]) );
  DFC3 pipe_data_alures_reg_18_ ( .D(resmux_o_data_alu[18]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[18]) );
  DFC3 pipe_data_alures_reg_17_ ( .D(resmux_o_data_alu[17]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[17]) );
  DFC3 pipe_data_alures_reg_16_ ( .D(resmux_o_data_alu[16]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[16]) );
  DFC3 pipe_data_alures_reg_15_ ( .D(resmux_o_data_alu[15]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[15]) );
  DFC3 pipe_data_alures_reg_14_ ( .D(resmux_o_data_alu[14]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[14]) );
  DFC3 pipe_data_alures_reg_13_ ( .D(resmux_o_data_alu[13]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[13]) );
  DFC3 pipe_data_alures_reg_12_ ( .D(resmux_o_data_alu[12]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[12]) );
  DFC3 pipe_data_alures_reg_11_ ( .D(resmux_o_data_alu[11]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[11]) );
  DFC3 pipe_data_alures_reg_10_ ( .D(resmux_o_data_alu[10]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[10]) );
  DFC3 pipe_data_alures_reg_9_ ( .D(resmux_o_data_alu[9]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[9]) );
  DFC3 pipe_data_alures_reg_8_ ( .D(resmux_o_data_alu[8]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[8]) );
  DFC3 pipe_data_alures_reg_7_ ( .D(resmux_o_data_alu[7]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[7]) );
  DFC3 pipe_data_alures_reg_6_ ( .D(resmux_o_data_alu[6]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[6]) );
  DFC3 pipe_data_alures_reg_5_ ( .D(resmux_o_data_alu[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[5]) );
  DFC3 pipe_data_alures_reg_4_ ( .D(resmux_o_data_alu[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[4]) );
  DFC3 pipe_data_alures_reg_3_ ( .D(resmux_o_data_alu[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[3]) );
  DFC3 pipe_data_alures_reg_2_ ( .D(resmux_o_data_alu[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[2]) );
  DFC3 pipe_data_alures_reg_1_ ( .D(resmux_o_data_alu[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[1]) );
  DFC3 pipe_data_alures_reg_0_ ( .D(resmux_o_data_alu[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[0]) );
  DFC3 pipe_data_memout_reg_31_ ( .D(i_data_memout[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[31]) );
  DFC3 pipe_data_memout_reg_30_ ( .D(i_data_memout[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[30]) );
  DFC3 pipe_data_memout_reg_29_ ( .D(i_data_memout[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[29]) );
  DFC3 pipe_data_memout_reg_28_ ( .D(i_data_memout[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[28]) );
  DFC3 pipe_data_memout_reg_27_ ( .D(i_data_memout[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[27]) );
  DFC3 pipe_data_memout_reg_26_ ( .D(i_data_memout[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[26]) );
  DFC3 pipe_data_memout_reg_25_ ( .D(i_data_memout[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[25]) );
  DFC3 pipe_data_memout_reg_24_ ( .D(i_data_memout[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[24]) );
  DFC3 pipe_data_memout_reg_23_ ( .D(i_data_memout[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[23]) );
  DFC3 pipe_data_memout_reg_22_ ( .D(i_data_memout[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[22]) );
  DFC3 pipe_data_memout_reg_21_ ( .D(i_data_memout[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[21]) );
  DFC3 pipe_data_memout_reg_20_ ( .D(i_data_memout[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[20]) );
  DFC3 pipe_data_memout_reg_19_ ( .D(i_data_memout[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[19]) );
  DFC3 pipe_data_memout_reg_18_ ( .D(i_data_memout[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[18]) );
  DFC3 pipe_data_memout_reg_17_ ( .D(i_data_memout[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[17]) );
  DFC3 pipe_data_memout_reg_16_ ( .D(i_data_memout[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[16]) );
  DFC3 pipe_data_memout_reg_15_ ( .D(i_data_memout[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[15]) );
  DFC3 pipe_data_memout_reg_14_ ( .D(i_data_memout[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[14]) );
  DFC3 pipe_data_memout_reg_13_ ( .D(i_data_memout[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[13]) );
  DFC3 pipe_data_memout_reg_12_ ( .D(i_data_memout[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[12]) );
  DFC3 pipe_data_memout_reg_11_ ( .D(i_data_memout[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[11]) );
  DFC3 pipe_data_memout_reg_10_ ( .D(i_data_memout[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[10]) );
  DFC3 pipe_data_memout_reg_9_ ( .D(i_data_memout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[9]) );
  DFC3 pipe_data_memout_reg_8_ ( .D(i_data_memout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[8]) );
  DFC3 pipe_data_memout_reg_7_ ( .D(i_data_memout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[7]) );
  DFC3 pipe_data_memout_reg_6_ ( .D(i_data_memout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[6]) );
  DFC3 pipe_data_memout_reg_5_ ( .D(i_data_memout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[5]) );
  DFC3 pipe_data_memout_reg_4_ ( .D(i_data_memout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[4]) );
  DFC3 pipe_data_memout_reg_3_ ( .D(i_data_memout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[3]) );
  DFC3 pipe_data_memout_reg_2_ ( .D(i_data_memout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[2]) );
  DFC3 pipe_data_memout_reg_1_ ( .D(i_data_memout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[1]) );
  DFC3 pipe_data_memout_reg_0_ ( .D(i_data_memout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[0]) );
  DFC3 pipe_addr_regdst_reg_4_ ( .D(i_addr_regdst[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[4]) );
  DFC3 pipe_addr_regdst_reg_3_ ( .D(i_addr_regdst[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[3]) );
  DFC3 pipe_addr_regdst_reg_2_ ( .D(i_addr_regdst[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[2]) );
  DFC3 pipe_addr_regdst_reg_1_ ( .D(i_addr_regdst[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[1]) );
  DFC3 pipe_addr_regdst_reg_0_ ( .D(i_addr_regdst[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[0]) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_con_FWmemread_reg ( .D(i_con_FWmemread), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_FWmemread) );
  M_resmux u_resmux ( .i_data_alures(i_data_alures), .i_data_pc8(pc8), 
        .i_con_pc8(i_con_Malupc8), .o_data_alu(resmux_o_data_alu) );
  mem_DW01_add_1 add_27 ( .A(i_data_pc4), .B({n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic1_, n_Logic0_, n_Logic0_}), .CI(n_Logic0_), .SUM(pc8) );
  DFC1 pipe_rt_reg_1_ ( .D(i_addr_Mrt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[1]) );
  LOGIC0 U3 ( .Q(n_Logic0_) );
  LOGIC1 U4 ( .Q(n_Logic1_) );
endmodule


module W_datamux ( i_data_alu, i_data_load, i_con_memtoreg, o_data_toreg );
  input [31:0] i_data_alu;
  input [31:0] i_data_load;
  output [31:0] o_data_toreg;
  input i_con_memtoreg;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n1, n2, n3, n4;

  AOI220 U1 ( .A(i_data_alu[21]), .B(n2), .C(i_data_load[21]), .D(
        i_con_memtoreg), .Q(n52) );
  AOI220 U2 ( .A(i_data_alu[22]), .B(n2), .C(i_data_load[22]), .D(
        i_con_memtoreg), .Q(n51) );
  AOI220 U3 ( .A(i_data_alu[23]), .B(n2), .C(i_data_load[23]), .D(
        i_con_memtoreg), .Q(n50) );
  AOI220 U4 ( .A(i_data_alu[0]), .B(n1), .C(i_data_load[0]), .D(i_con_memtoreg), .Q(n65) );
  AOI220 U5 ( .A(i_data_alu[2]), .B(n2), .C(i_data_load[2]), .D(i_con_memtoreg), .Q(n43) );
  AOI220 U6 ( .A(i_data_alu[3]), .B(n3), .C(i_data_load[3]), .D(i_con_memtoreg), .Q(n40) );
  AOI220 U7 ( .A(i_data_alu[4]), .B(n3), .C(i_data_load[4]), .D(i_con_memtoreg), .Q(n39) );
  AOI220 U8 ( .A(i_data_alu[5]), .B(n3), .C(i_data_load[5]), .D(i_con_memtoreg), .Q(n38) );
  AOI220 U9 ( .A(i_data_alu[6]), .B(n3), .C(i_data_load[6]), .D(i_con_memtoreg), .Q(n37) );
  AOI220 U10 ( .A(i_data_alu[7]), .B(n3), .C(i_data_load[7]), .D(
        i_con_memtoreg), .Q(n36) );
  AOI220 U11 ( .A(i_data_alu[8]), .B(n3), .C(i_data_load[8]), .D(
        i_con_memtoreg), .Q(n35) );
  AOI220 U12 ( .A(i_data_alu[9]), .B(n3), .C(i_data_load[9]), .D(
        i_con_memtoreg), .Q(n34) );
  AOI220 U13 ( .A(i_data_alu[10]), .B(n1), .C(i_data_load[10]), .D(
        i_con_memtoreg), .Q(n64) );
  AOI220 U14 ( .A(i_data_alu[11]), .B(n1), .C(i_data_load[11]), .D(
        i_con_memtoreg), .Q(n63) );
  AOI220 U15 ( .A(i_data_alu[12]), .B(n1), .C(i_data_load[12]), .D(
        i_con_memtoreg), .Q(n62) );
  AOI220 U16 ( .A(i_data_alu[13]), .B(n1), .C(i_data_load[13]), .D(
        i_con_memtoreg), .Q(n61) );
  AOI220 U17 ( .A(i_data_alu[14]), .B(n1), .C(i_data_load[14]), .D(
        i_con_memtoreg), .Q(n60) );
  AOI220 U18 ( .A(i_data_alu[15]), .B(n1), .C(i_data_load[15]), .D(
        i_con_memtoreg), .Q(n59) );
  AOI220 U19 ( .A(i_data_alu[16]), .B(n1), .C(i_data_load[16]), .D(
        i_con_memtoreg), .Q(n58) );
  AOI220 U20 ( .A(i_data_alu[24]), .B(n1), .C(i_data_load[24]), .D(
        i_con_memtoreg), .Q(n49) );
  AOI220 U21 ( .A(i_data_alu[25]), .B(n3), .C(i_data_load[25]), .D(
        i_con_memtoreg), .Q(n48) );
  AOI220 U22 ( .A(i_data_alu[26]), .B(n4), .C(i_data_load[26]), .D(
        i_con_memtoreg), .Q(n47) );
  AOI220 U23 ( .A(i_data_alu[27]), .B(n4), .C(i_data_load[27]), .D(
        i_con_memtoreg), .Q(n46) );
  AOI220 U24 ( .A(i_data_alu[28]), .B(n4), .C(i_data_load[28]), .D(
        i_con_memtoreg), .Q(n45) );
  AOI220 U25 ( .A(i_data_alu[29]), .B(n4), .C(i_data_load[29]), .D(
        i_con_memtoreg), .Q(n44) );
  AOI220 U26 ( .A(i_data_alu[30]), .B(n4), .C(i_data_load[30]), .D(
        i_con_memtoreg), .Q(n42) );
  AOI220 U27 ( .A(i_data_alu[31]), .B(n3), .C(i_data_load[31]), .D(
        i_con_memtoreg), .Q(n41) );
  AOI220 U28 ( .A(i_data_alu[17]), .B(n2), .C(i_data_load[17]), .D(
        i_con_memtoreg), .Q(n57) );
  AOI220 U29 ( .A(i_data_alu[18]), .B(n2), .C(i_data_load[18]), .D(
        i_con_memtoreg), .Q(n56) );
  AOI220 U30 ( .A(i_data_alu[19]), .B(n2), .C(i_data_load[19]), .D(
        i_con_memtoreg), .Q(n55) );
  AOI220 U31 ( .A(i_data_alu[20]), .B(n2), .C(i_data_load[20]), .D(
        i_con_memtoreg), .Q(n53) );
  BUF2 U32 ( .A(n4), .Q(n1) );
  BUF2 U33 ( .A(n4), .Q(n2) );
  BUF2 U34 ( .A(n4), .Q(n3) );
  INV3 U35 ( .A(n54), .Q(o_data_toreg[1]) );
  AOI220 U36 ( .A(i_data_alu[1]), .B(n2), .C(i_data_load[1]), .D(
        i_con_memtoreg), .Q(n54) );
  INV3 U37 ( .A(n55), .Q(o_data_toreg[19]) );
  INV3 U38 ( .A(n44), .Q(o_data_toreg[29]) );
  INV3 U39 ( .A(n42), .Q(o_data_toreg[30]) );
  INV3 U40 ( .A(n41), .Q(o_data_toreg[31]) );
  INV3 U41 ( .A(n65), .Q(o_data_toreg[0]) );
  INV3 U42 ( .A(n43), .Q(o_data_toreg[2]) );
  INV3 U43 ( .A(n40), .Q(o_data_toreg[3]) );
  INV3 U44 ( .A(n38), .Q(o_data_toreg[5]) );
  INV3 U45 ( .A(n37), .Q(o_data_toreg[6]) );
  INV3 U46 ( .A(n36), .Q(o_data_toreg[7]) );
  INV3 U47 ( .A(n35), .Q(o_data_toreg[8]) );
  INV3 U48 ( .A(n63), .Q(o_data_toreg[11]) );
  INV3 U49 ( .A(n62), .Q(o_data_toreg[12]) );
  INV3 U50 ( .A(n61), .Q(o_data_toreg[13]) );
  INV3 U51 ( .A(n60), .Q(o_data_toreg[14]) );
  INV3 U52 ( .A(n59), .Q(o_data_toreg[15]) );
  INV3 U53 ( .A(n57), .Q(o_data_toreg[17]) );
  INV3 U54 ( .A(n56), .Q(o_data_toreg[18]) );
  INV3 U55 ( .A(n51), .Q(o_data_toreg[22]) );
  INV3 U56 ( .A(n47), .Q(o_data_toreg[26]) );
  INV3 U57 ( .A(n45), .Q(o_data_toreg[28]) );
  INV3 U58 ( .A(n34), .Q(o_data_toreg[9]) );
  INV3 U59 ( .A(n58), .Q(o_data_toreg[16]) );
  INV3 U60 ( .A(n48), .Q(o_data_toreg[25]) );
  INV3 U61 ( .A(n50), .Q(o_data_toreg[23]) );
  INV3 U62 ( .A(n46), .Q(o_data_toreg[27]) );
  INV3 U63 ( .A(n39), .Q(o_data_toreg[4]) );
  INV3 U64 ( .A(n64), .Q(o_data_toreg[10]) );
  INV3 U65 ( .A(n49), .Q(o_data_toreg[24]) );
  INV3 U66 ( .A(n53), .Q(o_data_toreg[20]) );
  INV3 U67 ( .A(n52), .Q(o_data_toreg[21]) );
  INV3 U68 ( .A(i_con_memtoreg), .Q(n4) );
endmodule


module writeback ( i_data_alures, i_data_memout, i_con_Wmemtoreg, 
        o_data_regwrite );
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  output [31:0] o_data_regwrite;
  input i_con_Wmemtoreg;


  W_datamux u_datamux ( .i_data_alu(i_data_alures), .i_data_load(i_data_memout), .i_con_memtoreg(i_con_Wmemtoreg), .o_data_toreg(o_data_regwrite) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Mmemread, ex_con_Mmemwrite, ex_con_Malupc8, ex_con_Wmemtoreg,
         mem_con_Malupc8, mem_con_Wmemtoreg, wb_con_Wmemtoreg, n1,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2;
  wire   [31:0] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [31:0] id_addr_pc4;
  wire   [31:0] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] wb_data_memout;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] mem_data_alures;
  wire   [31:0] mem_data_pc4;

  fetch u_fetch ( .i_clk(clk), .i_nrst(rst_n), .i_addr_b(if_addr_b), 
        .i_addr_j({if_addr_j, n1, n1}), .i_addr_jr(id_data_jr), .i_con_b(
        if_con_b), .i_con_j(if_con_j), .i_data_instr(read_instruction), 
        .i_con_ifstall(if_con_ifstall), .o_addr_pc(instruction_address), 
        .o_addr_pc4(id_addr_pc4), .o_data_instr(id_data_instr) );
  decode u_decode ( .i_clk(clk), .i_nrst(rst_n), .i_addr_pc4(id_addr_pc4), 
        .i_data_instr(id_data_instr), .i_con_Wregwrite(id_con_Wregwrite), 
        .i_data_Wregwrite(id_data_Wregwrite), .i_addr_Wregwrite(
        id_addr_Wregwrite), .i_addr_Erd(for_o_addr_Erd), .i_addr_Mrd(
        mem_addr_regdst), .i_con_Eregwrite(ex_con_Wregwrite), 
        .i_con_Mregwrite(mem_con_Wregwrite), .i_addr_rtM(for_addr_rtM), 
        .i_addr_rtW(for_addr_rtW), .i_con_memreadM(mem_read), .i_con_memreadW(
        for_FWmemread), .i_data_Wmemout(wb_data_memout), .o_data_rs(id_data_rs), .o_data_rt(ex_data_rt), .o_addr_rd(ex_addr_rd), .o_addr_rt(ex_addr_rt), 
        .o_data_jr(id_data_jr), .o_con_jump(if_con_j), .o_addr_pc4(ex_data_pc4), .o_addr_branch(if_addr_b), .o_addr_jump({if_addr_j, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .o_con_Ealuop(ex_con_Ealuop), 
        .o_con_Ealusrc(ex_con_Ealusrc), .o_con_Eregdst(ex_con_Eregdst), 
        .o_con_Mmemread(ex_con_Mmemread), .o_con_Mmemwrite(ex_con_Mmemwrite), 
        .o_con_Malupc8(ex_con_Malupc8), .o_con_Wmemtoreg(ex_con_Wmemtoreg), 
        .o_con_Wregwrite(ex_con_Wregwrite), .o_con_ifstall(if_con_ifstall), 
        .o_con_Ebop(ex_con_bop), .o_data_signext(ex_data_immext), 
        .o_con_Efamux(for_o_con_Efamux), .o_con_Efbmux(for_o_con_Efbmux), 
        .o_data_Fmemout(for_memout) );
  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext(
        ex_data_immext), .i_addr_rt(ex_addr_rt), .i_addr_rd(ex_addr_rd), 
        .i_data_FEalures(data_address), .i_data_FMalures(mem_data_alures), 
        .i_data_FMmemout(wb_data_memout), .i_data_FWmemout(for_memout), 
        .i_con_Efamux(for_o_con_Efamux), .i_con_Efbmux(for_o_con_Efbmux), 
        .i_con_Ealuop(ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), 
        .i_con_Mmemwrite(ex_con_Mmemwrite), .i_con_Malupc8(ex_con_Malupc8), 
        .i_con_Wmemtoreg(ex_con_Wmemtoreg), .i_con_Wregwrite(ex_con_Wregwrite), 
        .i_con_bop(ex_con_bop), .o_data_pc4(mem_data_pc4), .o_data_alures(
        data_address), .o_data_rt(write_data), .o_addr_regdst(mem_addr_regdst), 
        .o_con_Mmemread(mem_read), .o_con_Mmemwrite(mem_write), 
        .o_con_Malupc8(mem_con_Malupc8), .o_con_Wmemtoreg(mem_con_Wmemtoreg), 
        .o_con_Wregwrite(mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), 
        .o_addr_Mrt(for_addr_rtM), .o_con_ifbranch(if_con_b) );
  mem u_mem ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(mem_data_pc4), 
        .i_data_alures(data_address), .i_data_memout(read_data), 
        .i_addr_regdst(mem_addr_regdst), .i_con_Malupc8(mem_con_Malupc8), 
        .i_con_Wmemtoreg(mem_con_Wmemtoreg), .i_con_Wregwrite(
        mem_con_Wregwrite), .i_con_FWmemread(ex_con_Mmemread), .i_addr_Mrt(
        for_addr_rtM), .o_data_alures(mem_data_alures), .o_data_memout(
        wb_data_memout), .o_addr_regdst(id_addr_Wregwrite), .o_con_Wmemtoreg(
        wb_con_Wmemtoreg), .o_con_Wregwrite(id_con_Wregwrite), 
        .o_con_FWmemread(for_FWmemread), .o_addr_Wrt(for_addr_rtW) );
  writeback u_writeback ( .i_data_alures(mem_data_alures), .i_data_memout(
        wb_data_memout), .i_con_Wmemtoreg(wb_con_Wmemtoreg), .o_data_regwrite(
        id_data_Wregwrite) );
  LOGIC0 U1 ( .Q(n1) );
endmodule

