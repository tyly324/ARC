`timescale 1ns / 1ps
module E_aluamux