
module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_famemout, i_data_fbmemout, i_con_Efamux, i_con_Efbmux, 
        i_con_Ealuop, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread, 
        i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_bop, o_data_alures, o_data_rt, o_addr_regdst, o_con_Mmemread, 
        o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, o_con_Wregwrite, 
        o_addr_Erd, o_addr_Mrt, o_con_ifbranch, o_data_pc4_31__BAR, 
        o_data_pc4_29_, o_data_pc4_27_, o_data_pc4_26_, o_data_pc4_25_, 
        o_data_pc4_24_, o_data_pc4_23_, o_data_pc4_22_, o_data_pc4_21_, 
        o_data_pc4_20_, o_data_pc4_19_, o_data_pc4_18_, o_data_pc4_17_, 
        o_data_pc4_16_, o_data_pc4_15_, o_data_pc4_14_, o_data_pc4_13_, 
        o_data_pc4_12_, o_data_pc4_11_, o_data_pc4_10_, o_data_pc4_9_, 
        o_data_pc4_8_, o_data_pc4_7_, o_data_pc4_6_, o_data_pc4_5_, 
        o_data_pc4_4_, o_data_pc4_3_, o_data_pc4_2_, o_data_pc4_1_, 
        o_data_pc4_0_, o_data_pc4_30__BAR, o_data_pc4_28__BAR );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_famemout;
  input [31:0] i_data_fbmemout;
  input [1:0] i_con_Efamux;
  input [1:0] i_con_Efbmux;
  input [5:0] i_con_Ealuop;
  input [2:0] i_con_bop;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch, o_data_pc4_31__BAR, o_data_pc4_29_,
         o_data_pc4_27_, o_data_pc4_26_, o_data_pc4_25_, o_data_pc4_24_,
         o_data_pc4_23_, o_data_pc4_22_, o_data_pc4_21_, o_data_pc4_20_,
         o_data_pc4_19_, o_data_pc4_18_, o_data_pc4_17_, o_data_pc4_16_,
         o_data_pc4_15_, o_data_pc4_14_, o_data_pc4_13_, o_data_pc4_12_,
         o_data_pc4_11_, o_data_pc4_10_, o_data_pc4_9_, o_data_pc4_8_,
         o_data_pc4_7_, o_data_pc4_6_, o_data_pc4_5_, o_data_pc4_4_,
         o_data_pc4_3_, o_data_pc4_2_, o_data_pc4_1_, o_data_pc4_0_,
         o_data_pc4_30__BAR, o_data_pc4_28__BAR;
  wire   compare_i_data_rt_31_, u_alu_N306, DP_OP_68_131_7244_n70,
         u_alu_DP_OP_85J3_126_1427_n379, u_alu_DP_OP_85J3_126_1427_n377,
         u_alu_DP_OP_85J3_126_1427_n374, u_alu_DP_OP_85J3_126_1427_n368,
         u_alu_ashr_4_A_17_, u_alu_ashr_4_A_16_, u_alu_ashr_4_A_9_,
         u_alu_ashr_4_A_6_, u_alu_ashr_4_A_5_, u_alu_DP_OP_83J3_124_3384_n154,
         u_alu_DP_OP_83J3_124_3384_n153, u_alu_DP_OP_83J3_124_3384_n152,
         u_alu_DP_OP_83J3_124_3384_n123, u_alu_DP_OP_83J3_124_3384_n122,
         u_alu_DP_OP_83J3_124_3384_n121, u_alu_DP_OP_83J3_124_3384_n120,
         u_alu_DP_OP_83J3_124_3384_n119, u_alu_DP_OP_83J3_124_3384_n117,
         u_alu_DP_OP_83J3_124_3384_n113, u_alu_DP_OP_83J3_124_3384_n112,
         u_alu_DP_OP_83J3_124_3384_n105, u_alu_DP_OP_83J3_124_3384_n102,
         u_alu_DP_OP_83J3_124_3384_n101, u_alu_DP_OP_83J3_124_3384_n93,
         u_alu_DP_OP_83J3_124_3384_n90, u_alu_DP_OP_83J3_124_3384_n89,
         u_alu_DP_OP_83J3_124_3384_n86, u_alu_DP_OP_83J3_124_3384_n83,
         u_alu_DP_OP_83J3_124_3384_n76, u_alu_DP_OP_83J3_124_3384_n75,
         u_alu_DP_OP_83J3_124_3384_n64, u_alu_DP_OP_83J3_124_3384_n55,
         u_alu_DP_OP_83J3_124_3384_n54, u_alu_DP_OP_83J3_124_3384_n53,
         u_alu_DP_OP_83J3_124_3384_n52, u_alu_DP_OP_83J3_124_3384_n51,
         u_alu_DP_OP_83J3_124_3384_n50, u_alu_DP_OP_83J3_124_3384_n45,
         u_alu_DP_OP_83J3_124_3384_n44, u_alu_DP_OP_83J3_124_3384_n43,
         u_alu_DP_OP_83J3_124_3384_n42, u_alu_DP_OP_83J3_124_3384_n41,
         u_alu_DP_OP_83J3_124_3384_n33, u_alu_DP_OP_83J3_124_3384_n32,
         u_alu_DP_OP_83J3_124_3384_n31, u_alu_DP_OP_83J3_124_3384_n30,
         u_alu_DP_OP_83J3_124_3384_n29, u_alu_DP_OP_83J3_124_3384_n26,
         u_alu_DP_OP_83J3_124_3384_n25, u_alu_DP_OP_83J3_124_3384_n23,
         u_alu_DP_OP_83J3_124_3384_n22, u_alu_DP_OP_83J3_124_3384_n19,
         u_alu_DP_OP_83J3_124_3384_n18, u_alu_DP_OP_83J3_124_3384_n16,
         u_alu_DP_OP_83J3_124_3384_n15, u_alu_DP_OP_83J3_124_3384_n11,
         u_alu_DP_OP_83J3_124_3384_n8, u_alu_DP_OP_83J3_124_3384_n7,
         u_alu_DP_OP_83J3_124_3384_n6, u_alu_DP_OP_83J3_124_3384_n5,
         u_alu_DP_OP_83J3_124_3384_n4, u_alu_DP_OP_83J3_124_3384_n3,
         u_alu_DP_OP_83J3_124_3384_n2, u_alu_DP_OP_83J3_124_3384_n1,
         u_alu_lt_x_11_A_31_, u_alu_lt_x_11_A_13_, u_alu_lt_x_11_A_11_,
         u_alu_lt_x_11_A_3_, u_alu_lt_x_11_A_0_, u_alu_lt_x_11_B_29_,
         u_alu_lt_x_11_B_28_, u_alu_lt_x_11_B_25_, u_alu_lt_x_11_B_24_,
         u_alu_lt_x_11_B_11_, u_alu_lt_x_11_B_1_, u_alu_lt_x_11_B_0_,
         u_alu_lt_x_11_n144, u_alu_lt_x_11_n139, u_alu_lt_x_11_n138,
         u_alu_lt_x_11_n122, u_alu_lt_x_11_n121, u_alu_lt_x_11_n119,
         u_alu_lt_x_11_n118, u_alu_lt_x_11_n117, u_alu_lt_x_11_n116,
         u_alu_lt_x_11_n115, u_alu_lt_x_11_n114, u_alu_lt_x_11_n112,
         u_alu_lt_x_11_n111, u_alu_lt_x_11_n110, u_alu_lt_x_11_n108,
         u_alu_lt_x_11_n106, u_alu_lt_x_11_n105, u_alu_lt_x_11_n104,
         u_alu_lt_x_11_n103, u_alu_lt_x_11_n102, u_alu_lt_x_11_n101,
         u_alu_lt_x_11_n100, u_alu_lt_x_11_n99, u_alu_lt_x_11_n98,
         u_alu_lt_x_11_n97, u_alu_lt_x_11_n96, u_alu_lt_x_11_n95,
         u_alu_lt_x_11_n90, u_alu_lt_x_11_n89, u_alu_lt_x_11_n88,
         u_alu_lt_x_11_n87, u_alu_lt_x_11_n86, u_alu_lt_x_11_n85,
         u_alu_lt_x_11_n84, u_alu_lt_x_11_n83, u_alu_lt_x_11_n82,
         u_alu_lt_x_11_n80, u_alu_lt_x_11_n78, u_alu_lt_x_11_n77,
         u_alu_lt_x_11_n75, u_alu_lt_x_11_n74, u_alu_lt_x_11_n71,
         u_alu_lt_x_11_n69, u_alu_lt_x_11_n68, u_alu_lt_x_11_n66,
         u_alu_lt_x_11_n64, u_alu_lt_x_11_n62, u_alu_lt_x_11_n61,
         u_alu_lt_x_11_n60, u_alu_lt_x_11_n59, u_alu_lt_x_11_n58,
         u_alu_lt_x_11_n57, u_alu_lt_x_11_n56, u_alu_lt_x_11_n55,
         u_alu_lt_x_11_n54, u_alu_lt_x_11_n53, u_alu_lt_x_11_n52,
         u_alu_lt_x_11_n51, u_alu_lt_x_11_n50, u_alu_lt_x_11_n49,
         u_alu_lt_x_11_n48, u_alu_lt_x_11_n47, u_alu_lt_x_11_n46,
         u_alu_lt_x_11_n45, u_alu_lt_x_11_n44, u_alu_lt_x_11_n43,
         u_alu_lt_x_11_n42, u_alu_lt_x_11_n41, u_alu_lt_x_11_n40,
         u_alu_lt_x_11_n39, u_alu_lt_x_11_n38, u_alu_lt_x_11_n37,
         u_alu_lt_x_11_n36, u_alu_lt_x_11_n35, u_alu_lt_x_11_n34,
         u_alu_lt_x_11_n33, u_alu_lt_x_11_n32, u_alu_lt_x_11_n31,
         u_alu_lt_x_11_n30, u_alu_lt_x_11_n29, u_alu_lt_x_11_n28,
         u_alu_lt_x_11_n27, u_alu_lt_x_11_n26, u_alu_lt_x_11_n22,
         u_alu_lt_x_11_n21, u_alu_lt_x_11_n18, u_alu_lt_x_11_n17,
         u_alu_lt_x_11_n16, u_alu_lt_x_11_n15, u_alu_lt_x_11_n14,
         u_alu_lt_x_11_n13, u_alu_lt_x_11_n12, u_alu_lt_x_11_n10,
         u_alu_lt_x_11_n9, u_alu_lt_x_11_n8, u_alu_lt_x_11_n7,
         u_alu_lt_x_11_n5, u_alu_lt_x_11_n3, u_alu_lt_x_11_n1,
         u_alu_DP_OP_84J3_125_2615_n113, u_alu_DP_OP_84J3_125_2615_n112,
         u_alu_DP_OP_84J3_125_2615_n111, u_alu_DP_OP_84J3_125_2615_n109,
         u_alu_DP_OP_84J3_125_2615_n108, u_alu_DP_OP_84J3_125_2615_n103,
         u_alu_DP_OP_84J3_125_2615_n102, u_alu_DP_OP_84J3_125_2615_n95,
         u_alu_DP_OP_84J3_125_2615_n92, u_alu_DP_OP_84J3_125_2615_n86,
         u_alu_DP_OP_84J3_125_2615_n81, u_alu_DP_OP_84J3_125_2615_n77,
         u_alu_DP_OP_84J3_125_2615_n73, u_alu_DP_OP_84J3_125_2615_n70,
         u_alu_DP_OP_84J3_125_2615_n58, u_alu_DP_OP_84J3_125_2615_n50,
         u_alu_DP_OP_84J3_125_2615_n49, u_alu_DP_OP_84J3_125_2615_n48,
         u_alu_DP_OP_84J3_125_2615_n47, u_alu_DP_OP_84J3_125_2615_n46,
         u_alu_DP_OP_84J3_125_2615_n45, u_alu_DP_OP_84J3_125_2615_n40,
         u_alu_DP_OP_84J3_125_2615_n39, u_alu_DP_OP_84J3_125_2615_n38,
         u_alu_DP_OP_84J3_125_2615_n37, u_alu_DP_OP_84J3_125_2615_n36,
         u_alu_DP_OP_84J3_125_2615_n31, u_alu_DP_OP_84J3_125_2615_n30,
         u_alu_DP_OP_84J3_125_2615_n23, u_alu_DP_OP_84J3_125_2615_n22,
         u_alu_DP_OP_84J3_125_2615_n18, u_alu_DP_OP_84J3_125_2615_n17,
         u_alu_DP_OP_84J3_125_2615_n16, u_alu_DP_OP_84J3_125_2615_n15,
         u_alu_DP_OP_84J3_125_2615_n14, u_alu_DP_OP_84J3_125_2615_n8,
         u_alu_DP_OP_84J3_125_2615_n7, u_alu_DP_OP_84J3_125_2615_n6,
         u_alu_DP_OP_84J3_125_2615_n5, u_alu_DP_OP_84J3_125_2615_n4,
         u_alu_DP_OP_84J3_125_2615_n3, u_alu_DP_OP_84J3_125_2615_n2,
         u_alu_DP_OP_84J3_125_2615_n1, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103;
  wire   [31:0] alu_o_data_AluRes;
  wire   [14:2] compare_i_data_rs;
  wire   [27:19] alu_i_data_B;
  wire   [6:1] u_alu_pre_sum_4b;
  wire   [6:0] u_alu_pre_sum_4a;
  wire   [8:1] u_alu_pre_sum_3b;
  wire   [6:0] u_alu_pre_sum_3a;

  DFC1 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC1 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC1 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC1 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC1 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC1 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_31__BAR) );
  DFC1 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_30__BAR) );
  DFC1 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_29_) );
  DFC1 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .QN(
        o_data_pc4_28__BAR) );
  DFC1 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_27_) );
  DFC1 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_26_) );
  DFC1 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_25_) );
  DFC1 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_24_) );
  DFC1 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_23_) );
  DFC1 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_22_) );
  DFC1 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_21_) );
  DFC1 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_20_) );
  DFC1 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_19_) );
  DFC1 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_18_) );
  DFC1 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_17_) );
  DFC1 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_16_) );
  DFC1 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_15_) );
  DFC1 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_14_) );
  DFC1 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_13_) );
  DFC1 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_12_) );
  DFC1 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_11_) );
  DFC1 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_10_) );
  DFC1 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_9_) );
  DFC1 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_8_) );
  DFC1 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_7_) );
  DFC1 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_6_) );
  DFC1 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_5_) );
  DFC1 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_4_) );
  DFC1 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_3_) );
  DFC1 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_2_) );
  DFC1 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_1_) );
  DFC1 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4_0_) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC1 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC1 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC1 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC1 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC1 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC1 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC1 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC1 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC1 pipe_alures_reg_15_ ( .D(alu_o_data_AluRes[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[15]) );
  DFC1 pipe_alures_reg_14_ ( .D(alu_o_data_AluRes[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[14]) );
  DFC1 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC1 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC1 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC1 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC1 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC1 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC1 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC1 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC1 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC1 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC1 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC1 pipe_rt_reg_31_ ( .D(compare_i_data_rt_31_), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC1 pipe_rt_reg_30_ ( .D(n33), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC1 pipe_rt_reg_29_ ( .D(n915), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[29])
         );
  DFC1 pipe_rt_reg_28_ ( .D(n3072), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28])
         );
  DFC1 pipe_rt_reg_27_ ( .D(n3073), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27])
         );
  DFC1 pipe_rt_reg_26_ ( .D(n3074), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26])
         );
  DFC1 pipe_rt_reg_25_ ( .D(n3075), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25])
         );
  DFC1 pipe_rt_reg_24_ ( .D(n3076), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24])
         );
  DFC1 pipe_rt_reg_23_ ( .D(n3077), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23])
         );
  DFC1 pipe_rt_reg_22_ ( .D(n3078), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22])
         );
  DFC1 pipe_rt_reg_21_ ( .D(n3079), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21])
         );
  DFC1 pipe_rt_reg_20_ ( .D(n3080), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20])
         );
  DFC1 pipe_rt_reg_19_ ( .D(n3081), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19])
         );
  DFC1 pipe_rt_reg_18_ ( .D(n913), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18])
         );
  DFC1 pipe_rt_reg_17_ ( .D(n3082), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17])
         );
  DFC1 pipe_rt_reg_16_ ( .D(n3083), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16])
         );
  DFC1 pipe_rt_reg_15_ ( .D(n3084), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15])
         );
  DFC1 pipe_rt_reg_14_ ( .D(n3085), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14])
         );
  DFC1 pipe_rt_reg_13_ ( .D(n3086), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13])
         );
  DFC1 pipe_rt_reg_12_ ( .D(n3087), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12])
         );
  DFC1 pipe_rt_reg_11_ ( .D(n3088), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11])
         );
  DFC1 pipe_rt_reg_10_ ( .D(n3089), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10])
         );
  DFC1 pipe_rt_reg_9_ ( .D(n3090), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[9]) );
  DFC1 pipe_rt_reg_8_ ( .D(n3091), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[8]) );
  DFC1 pipe_rt_reg_7_ ( .D(n3092), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[7]) );
  DFC1 pipe_rt_reg_6_ ( .D(n3093), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[6]) );
  DFC1 pipe_rt_reg_5_ ( .D(n3094), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[5]) );
  DFC1 pipe_rt_reg_4_ ( .D(n3095), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[4]) );
  DFC1 pipe_rt_reg_3_ ( .D(n3096), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[3]) );
  DFC1 pipe_rt_reg_2_ ( .D(n912), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[2]) );
  DFC1 pipe_rt_reg_1_ ( .D(n3097), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[1]) );
  DFC1 pipe_rt_reg_0_ ( .D(n3098), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[0]) );
  DFC1 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC1 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC1 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC1 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC1 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC1 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC1 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC1 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC1 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_con_Malupc8_reg ( .D(i_con_Malupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Malupc8) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U6 ( .A(u_alu_DP_OP_84J3_125_2615_n2), .B(
        u_alu_DP_OP_84J3_125_2615_n16), .Q(u_alu_pre_sum_4a[6]) );
  XNR21 u_alu_DP_OP_83J3_124_3384_U115 ( .A(u_alu_DP_OP_83J3_124_3384_n6), .B(
        u_alu_DP_OP_83J3_124_3384_n105), .Q(u_alu_pre_sum_3b[3]) );
  XNR21 u_alu_DP_OP_83J3_124_3384_U43 ( .A(u_alu_DP_OP_83J3_124_3384_n6), .B(
        u_alu_DP_OP_83J3_124_3384_n43), .Q(u_alu_pre_sum_3a[3]) );
  XNR21 u_alu_DP_OP_83J3_124_3384_U13 ( .A(u_alu_DP_OP_83J3_124_3384_n3), .B(
        n1300), .Q(u_alu_pre_sum_3a[6]) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U90 ( .A(u_alu_DP_OP_84J3_125_2615_n4), .B(
        n624), .Q(u_alu_pre_sum_4b[4]) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U102 ( .A(u_alu_DP_OP_84J3_125_2615_n5), .B(
        u_alu_DP_OP_84J3_125_2615_n95), .Q(u_alu_pre_sum_4b[3]) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U36 ( .A(u_alu_DP_OP_84J3_125_2615_n5), .B(
        u_alu_DP_OP_84J3_125_2615_n38), .Q(u_alu_pre_sum_4a[3]) );
  NOR20 u_alu_lt_x_11_U118 ( .A(u_alu_lt_x_11_n121), .B(u_alu_lt_x_11_B_1_), 
        .Q(u_alu_lt_x_11_n117) );
  NAND20 u_alu_lt_x_11_U119 ( .A(u_alu_lt_x_11_B_1_), .B(u_alu_lt_x_11_n121), 
        .Q(u_alu_lt_x_11_n118) );
  NAND20 u_alu_lt_x_11_U103 ( .A(u_alu_ashr_4_A_6_), .B(n221), .Q(
        u_alu_lt_x_11_n102) );
  NAND20 u_alu_lt_x_11_U101 ( .A(n2146), .B(n1971), .Q(u_alu_lt_x_11_n100) );
  OAI210 u_alu_lt_x_11_U76 ( .A(n2467), .B(n2482), .C(u_alu_lt_x_11_n77), .Q(
        u_alu_lt_x_11_n75) );
  OAI210 u_alu_lt_x_11_U70 ( .A(n2466), .B(n2484), .C(u_alu_lt_x_11_n71), .Q(
        u_alu_lt_x_11_n69) );
  NAND20 u_alu_lt_x_11_U61 ( .A(u_alu_ashr_4_A_17_), .B(n2516), .Q(
        u_alu_lt_x_11_n60) );
  NAND20 u_alu_lt_x_11_U43 ( .A(n1338), .B(n182), .Q(u_alu_lt_x_11_n42) );
  NAND20 u_alu_lt_x_11_U41 ( .A(u_alu_DP_OP_83J3_124_3384_n153), .B(n2780), 
        .Q(u_alu_lt_x_11_n40) );
  NAND20 u_alu_lt_x_11_U33 ( .A(u_alu_lt_x_11_B_24_), .B(u_alu_lt_x_11_n144), 
        .Q(u_alu_lt_x_11_n32) );
  OAI210 u_alu_lt_x_11_U29 ( .A(u_alu_lt_x_11_n32), .B(u_alu_lt_x_11_n29), .C(
        u_alu_lt_x_11_n30), .Q(u_alu_lt_x_11_n28) );
  NAND20 u_alu_lt_x_11_U19 ( .A(u_alu_lt_x_11_B_28_), .B(n228), .Q(
        u_alu_lt_x_11_n18) );
  OAI210 u_alu_lt_x_11_U15 ( .A(u_alu_lt_x_11_n18), .B(u_alu_lt_x_11_n15), .C(
        u_alu_lt_x_11_n16), .Q(u_alu_lt_x_11_n14) );
  OAI210 u_alu_lt_x_11_U9 ( .A(u_alu_lt_x_11_n12), .B(u_alu_lt_x_11_n9), .C(
        u_alu_lt_x_11_n10), .Q(u_alu_lt_x_11_n8) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U58 ( .A(u_alu_DP_OP_84J3_125_2615_n113), 
        .B(u_alu_DP_OP_84J3_125_2615_n48), .Q(u_alu_DP_OP_84J3_125_2615_n7) );
  XOR21 u_alu_DP_OP_84J3_125_2615_U121 ( .A(u_alu_DP_OP_84J3_125_2615_n49), 
        .B(u_alu_DP_OP_84J3_125_2615_n7), .Q(u_alu_pre_sum_4b[1]) );
  XOR21 u_alu_DP_OP_84J3_125_2615_U55 ( .A(u_alu_DP_OP_84J3_125_2615_n50), .B(
        u_alu_DP_OP_84J3_125_2615_n7), .Q(u_alu_pre_sum_4a[1]) );
  NAND22 u_alu_DP_OP_83J3_124_3384_U29 ( .A(u_alu_DP_OP_83J3_124_3384_n119), 
        .B(u_alu_DP_OP_83J3_124_3384_n30), .Q(u_alu_DP_OP_83J3_124_3384_n4) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U10 ( .A(u_alu_DP_OP_84J3_125_2615_n108), 
        .B(u_alu_DP_OP_84J3_125_2615_n15), .Q(u_alu_DP_OP_84J3_125_2615_n2) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U16 ( .A(u_alu_DP_OP_84J3_125_2615_n81), 
        .B(u_alu_DP_OP_84J3_125_2615_n109), .Q(u_alu_DP_OP_84J3_125_2615_n17)
         );
  OAI212 u_alu_DP_OP_84J3_125_2615_U57 ( .A(u_alu_DP_OP_84J3_125_2615_n50), 
        .B(u_alu_DP_OP_84J3_125_2615_n47), .C(u_alu_DP_OP_84J3_125_2615_n48), 
        .Q(u_alu_DP_OP_84J3_125_2615_n46) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U20 ( .A(u_alu_DP_OP_84J3_125_2615_n109), 
        .B(u_alu_DP_OP_84J3_125_2615_n22), .Q(u_alu_DP_OP_84J3_125_2615_n3) );
  XOR21 u_alu_DP_OP_84J3_125_2615_U14 ( .A(u_alu_DP_OP_84J3_125_2615_n3), .B(
        u_alu_DP_OP_84J3_125_2615_n23), .Q(u_alu_pre_sum_4a[5]) );
  NAND22 u_alu_DP_OP_83J3_124_3384_U47 ( .A(u_alu_DP_OP_83J3_124_3384_n121), 
        .B(u_alu_DP_OP_83J3_124_3384_n42), .Q(u_alu_DP_OP_83J3_124_3384_n6) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U32 ( .A(u_alu_DP_OP_84J3_125_2615_n81), 
        .B(u_alu_DP_OP_84J3_125_2615_n31), .Q(u_alu_DP_OP_84J3_125_2615_n4) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U51 ( .A(u_alu_DP_OP_84J3_125_2615_n112), 
        .B(u_alu_DP_OP_84J3_125_2615_n40), .Q(u_alu_DP_OP_84J3_125_2615_n6) );
  XOR21 u_alu_DP_OP_84J3_125_2615_U111 ( .A(u_alu_DP_OP_84J3_125_2615_n6), .B(
        u_alu_DP_OP_84J3_125_2615_n102), .Q(u_alu_pre_sum_4b[2]) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U41 ( .A(u_alu_DP_OP_84J3_125_2615_n111), 
        .B(u_alu_DP_OP_84J3_125_2615_n37), .Q(u_alu_DP_OP_84J3_125_2615_n5) );
  NAND22 u_alu_DP_OP_83J3_124_3384_U39 ( .A(u_alu_DP_OP_83J3_124_3384_n120), 
        .B(u_alu_DP_OP_83J3_124_3384_n33), .Q(u_alu_DP_OP_83J3_124_3384_n5) );
  NAND22 u_alu_DP_OP_83J3_124_3384_U57 ( .A(u_alu_DP_OP_83J3_124_3384_n122), 
        .B(u_alu_DP_OP_83J3_124_3384_n45), .Q(u_alu_DP_OP_83J3_124_3384_n7) );
  XOR21 u_alu_DP_OP_83J3_124_3384_U123 ( .A(u_alu_DP_OP_83J3_124_3384_n7), .B(
        u_alu_DP_OP_83J3_124_3384_n112), .Q(u_alu_pre_sum_3b[2]) );
  XOR21 u_alu_DP_OP_83J3_124_3384_U51 ( .A(u_alu_DP_OP_83J3_124_3384_n7), .B(
        u_alu_DP_OP_83J3_124_3384_n50), .Q(u_alu_pre_sum_3a[2]) );
  NOR21 u_alu_lt_x_11_U14 ( .A(u_alu_lt_x_11_n15), .B(u_alu_lt_x_11_n17), .Q(
        u_alu_lt_x_11_n13) );
  NAND22 u_alu_lt_x_11_U50 ( .A(u_alu_lt_x_11_n51), .B(u_alu_lt_x_11_n57), .Q(
        u_alu_lt_x_11_n49) );
  NOR21 u_alu_lt_x_11_U44 ( .A(u_alu_lt_x_11_n45), .B(u_alu_lt_x_11_n47), .Q(
        u_alu_lt_x_11_n43) );
  NOR21 u_alu_lt_x_11_U40 ( .A(n2780), .B(u_alu_DP_OP_83J3_124_3384_n153), .Q(
        u_alu_lt_x_11_n39) );
  NAND22 u_alu_lt_x_11_U2 ( .A(u_alu_lt_x_11_n3), .B(u_alu_lt_x_11_n33), .Q(
        u_alu_lt_x_11_n1) );
  NAND22 u_alu_lt_x_11_U96 ( .A(u_alu_lt_x_11_n97), .B(u_alu_lt_x_11_n103), 
        .Q(u_alu_lt_x_11_n95) );
  NOR21 u_alu_lt_x_11_U111 ( .A(u_alu_lt_x_11_n112), .B(u_alu_lt_x_11_n114), 
        .Q(u_alu_lt_x_11_n110) );
  AOI211 u_alu_lt_x_11_U97 ( .A(u_alu_lt_x_11_n97), .B(u_alu_lt_x_11_n104), 
        .C(u_alu_lt_x_11_n98), .Q(u_alu_lt_x_11_n96) );
  NOR21 u_alu_lt_x_11_U69 ( .A(n2486), .B(n2484), .Q(u_alu_lt_x_11_n68) );
  NOR21 u_alu_lt_x_11_U75 ( .A(u_alu_lt_x_11_n78), .B(n2482), .Q(
        u_alu_lt_x_11_n74) );
  NAND22 u_alu_lt_x_11_U67 ( .A(u_alu_lt_x_11_n68), .B(u_alu_lt_x_11_n74), .Q(
        u_alu_lt_x_11_n66) );
  NOR21 u_alu_lt_x_11_U83 ( .A(u_alu_lt_x_11_n86), .B(u_alu_lt_x_11_n84), .Q(
        u_alu_lt_x_11_n82) );
  NOR21 u_alu_lt_x_11_U89 ( .A(u_alu_lt_x_11_n90), .B(n520), .Q(
        u_alu_lt_x_11_n88) );
  NAND22 u_alu_lt_x_11_U81 ( .A(u_alu_lt_x_11_n82), .B(u_alu_lt_x_11_n88), .Q(
        u_alu_lt_x_11_n80) );
  NOR21 u_alu_lt_x_11_U65 ( .A(u_alu_lt_x_11_n66), .B(u_alu_lt_x_11_n80), .Q(
        u_alu_lt_x_11_n64) );
  AOI211 u_alu_lt_x_11_U51 ( .A(u_alu_lt_x_11_n58), .B(u_alu_lt_x_11_n51), .C(
        u_alu_lt_x_11_n52), .Q(u_alu_lt_x_11_n50) );
  AOI211 u_alu_lt_x_11_U37 ( .A(u_alu_lt_x_11_n44), .B(u_alu_lt_x_11_n37), .C(
        u_alu_lt_x_11_n38), .Q(u_alu_lt_x_11_n36) );
  NAND22 u_alu_DP_OP_84J3_125_2615_U63 ( .A(u_alu_DP_OP_84J3_125_2615_n58), 
        .B(u_alu_DP_OP_84J3_125_2615_n50), .Q(u_alu_DP_OP_84J3_125_2615_n8) );
  NAND22 u_alu_DP_OP_83J3_124_3384_U9 ( .A(u_alu_DP_OP_83J3_124_3384_n117), 
        .B(u_alu_DP_OP_83J3_124_3384_n16), .Q(u_alu_DP_OP_83J3_124_3384_n2) );
  NAND22 u_alu_DP_OP_83J3_124_3384_U15 ( .A(u_alu_DP_OP_83J3_124_3384_n89), 
        .B(n1101), .Q(u_alu_DP_OP_83J3_124_3384_n18) );
  AOI211 u_alu_DP_OP_83J3_124_3384_U16 ( .A(u_alu_DP_OP_83J3_124_3384_n90), 
        .B(n1101), .C(u_alu_DP_OP_83J3_124_3384_n83), .Q(
        u_alu_DP_OP_83J3_124_3384_n19) );
  NAND22 u_alu_DP_OP_83J3_124_3384_U64 ( .A(u_alu_DP_OP_83J3_124_3384_n123), 
        .B(u_alu_DP_OP_83J3_124_3384_n53), .Q(u_alu_DP_OP_83J3_124_3384_n8) );
  XOR21 u_alu_DP_OP_83J3_124_3384_U61 ( .A(u_alu_DP_OP_83J3_124_3384_n55), .B(
        u_alu_DP_OP_83J3_124_3384_n8), .Q(u_alu_pre_sum_3a[1]) );
  OAI212 u_alu_DP_OP_84J3_125_2615_U123 ( .A(u_alu_DP_OP_84J3_125_2615_n49), 
        .B(u_alu_DP_OP_84J3_125_2615_n47), .C(u_alu_DP_OP_84J3_125_2615_n48), 
        .Q(u_alu_DP_OP_84J3_125_2615_n103) );
  NAND20 u_alu_lt_x_11_U109 ( .A(n2025), .B(n227), .Q(u_alu_lt_x_11_n108) );
  NOR21 u_alu_lt_x_11_U42 ( .A(n182), .B(n1338), .Q(u_alu_lt_x_11_n41) );
  NOR21 u_alu_lt_x_11_U18 ( .A(n228), .B(u_alu_lt_x_11_B_28_), .Q(
        u_alu_lt_x_11_n17) );
  DFC3 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC3 pipe_alures_reg_13_ ( .D(alu_o_data_AluRes[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[13]) );
  DFC3 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC3 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  NAND23 u_alu_DP_OP_84J3_125_2615_U54 ( .A(n1336), .B(n1509), .Q(
        u_alu_DP_OP_84J3_125_2615_n40) );
  NAND21 u_alu_lt_x_11_U120 ( .A(u_alu_lt_x_11_B_0_), .B(n857), .Q(
        u_alu_lt_x_11_n119) );
  NOR21 u_alu_lt_x_11_U32 ( .A(u_alu_lt_x_11_n144), .B(n43), .Q(
        u_alu_lt_x_11_n31) );
  OAI211 u_alu_lt_x_11_U59 ( .A(u_alu_lt_x_11_n62), .B(u_alu_lt_x_11_n59), .C(
        u_alu_lt_x_11_n60), .Q(u_alu_lt_x_11_n58) );
  OAI211 u_alu_lt_x_11_U112 ( .A(u_alu_lt_x_11_n115), .B(u_alu_lt_x_11_n112), 
        .C(n2461), .Q(u_alu_lt_x_11_n111) );
  OAI211 u_alu_lt_x_11_U45 ( .A(u_alu_lt_x_11_n48), .B(u_alu_lt_x_11_n45), .C(
        u_alu_lt_x_11_n46), .Q(u_alu_lt_x_11_n44) );
  XOR21 u_alu_DP_OP_83J3_124_3384_U133 ( .A(u_alu_DP_OP_83J3_124_3384_n54), 
        .B(u_alu_DP_OP_83J3_124_3384_n8), .Q(u_alu_pre_sum_3b[1]) );
  NAND22 u_alu_lt_x_11_U13 ( .A(u_alu_DP_OP_85J3_126_1427_n368), .B(n1280), 
        .Q(u_alu_lt_x_11_n12) );
  OAI211 u_alu_lt_x_11_U53 ( .A(u_alu_lt_x_11_n56), .B(u_alu_lt_x_11_n53), .C(
        u_alu_lt_x_11_n54), .Q(u_alu_lt_x_11_n52) );
  NOR21 u_alu_lt_x_11_U102 ( .A(n221), .B(u_alu_ashr_4_A_6_), .Q(
        u_alu_lt_x_11_n101) );
  NAND22 u_alu_lt_x_11_U86 ( .A(u_alu_lt_x_11_B_11_), .B(n222), .Q(
        u_alu_lt_x_11_n85) );
  OAI210 u_alu_lt_x_11_U84 ( .A(u_alu_lt_x_11_n87), .B(u_alu_lt_x_11_n84), .C(
        u_alu_lt_x_11_n85), .Q(u_alu_lt_x_11_n83) );
  NAND22 u_alu_DP_OP_83J3_124_3384_U19 ( .A(n1101), .B(
        u_alu_DP_OP_83J3_124_3384_n23), .Q(u_alu_DP_OP_83J3_124_3384_n3) );
  XOR21 u_alu_DP_OP_84J3_125_2615_U45 ( .A(u_alu_DP_OP_84J3_125_2615_n6), .B(
        u_alu_DP_OP_84J3_125_2615_n45), .Q(u_alu_pre_sum_4a[2]) );
  NOR21 u_alu_lt_x_11_U58 ( .A(u_alu_lt_x_11_n61), .B(u_alu_lt_x_11_n59), .Q(
        u_alu_lt_x_11_n57) );
  OAI212 u_alu_lt_x_11_U117 ( .A(u_alu_lt_x_11_n117), .B(u_alu_lt_x_11_n119), 
        .C(u_alu_lt_x_11_n118), .Q(u_alu_lt_x_11_n116) );
  NAND22 u_alu_lt_x_11_U36 ( .A(u_alu_lt_x_11_n43), .B(u_alu_lt_x_11_n37), .Q(
        u_alu_lt_x_11_n35) );
  OAI211 u_alu_lt_x_11_U39 ( .A(u_alu_lt_x_11_n42), .B(u_alu_lt_x_11_n39), .C(
        u_alu_lt_x_11_n40), .Q(u_alu_lt_x_11_n38) );
  OAI211 u_alu_lt_x_11_U35 ( .A(u_alu_lt_x_11_n50), .B(u_alu_lt_x_11_n35), .C(
        u_alu_lt_x_11_n36), .Q(u_alu_lt_x_11_n34) );
  XNR21 u_alu_DP_OP_84J3_125_2615_U24 ( .A(u_alu_DP_OP_84J3_125_2615_n4), .B(
        n970), .Q(u_alu_pre_sum_4a[4]) );
  DFC1 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  NAND22 U3 ( .A(n170), .B(i_data_immext[6]), .Q(n1997) );
  NOR22 U4 ( .A(n223), .B(n1830), .Q(u_alu_lt_x_11_n112) );
  CLKBU12 U5 ( .A(i_data_immext[8]), .Q(n1362) );
  NOR31 U6 ( .A(n2188), .B(n2187), .C(n2186), .Q(n2189) );
  NOR21 U7 ( .A(n2806), .B(n2810), .Q(n2539) );
  INV3 U8 ( .A(u_alu_DP_OP_84J3_125_2615_n31), .Q(
        u_alu_DP_OP_84J3_125_2615_n86) );
  NOR21 U9 ( .A(n247), .B(n1823), .Q(n1118) );
  NOR21 U10 ( .A(n177), .B(n1332), .Q(n1695) );
  NAND22 U11 ( .A(n1545), .B(i_data_famemout[17]), .Q(n2528) );
  INV3 U12 ( .A(n815), .Q(n433) );
  NOR23 U13 ( .A(n184), .B(n92), .Q(u_alu_lt_x_11_n86) );
  INV6 U14 ( .A(n1677), .Q(n1683) );
  NOR22 U15 ( .A(n2100), .B(n2099), .Q(n2139) );
  NOR22 U16 ( .A(n2187), .B(n794), .Q(n2274) );
  NOR23 U17 ( .A(n229), .B(n2259), .Q(n2482) );
  NAND23 U18 ( .A(n2320), .B(n1364), .Q(n2020) );
  INV3 U19 ( .A(n2762), .Q(n2765) );
  INV3 U20 ( .A(n177), .Q(n45) );
  NAND33 U21 ( .A(n1598), .B(n1597), .C(n1369), .Q(n1599) );
  INV3 U22 ( .A(n1277), .Q(n1280) );
  NAND24 U23 ( .A(n1336), .B(n224), .Q(u_alu_lt_x_11_n26) );
  NOR21 U24 ( .A(u_alu_lt_x_11_n99), .B(u_alu_lt_x_11_n101), .Q(
        u_alu_lt_x_11_n97) );
  BUF6 U25 ( .A(u_alu_lt_x_11_B_24_), .Q(n43) );
  NOR21 U26 ( .A(n2931), .B(n621), .Q(u_alu_lt_x_11_n21) );
  NOR21 U27 ( .A(n2008), .B(u_alu_lt_x_11_n99), .Q(n1974) );
  NAND23 U28 ( .A(n93), .B(n184), .Q(u_alu_lt_x_11_n87) );
  NAND26 U29 ( .A(n1590), .B(n1589), .Q(u_alu_DP_OP_85J3_126_1427_n374) );
  INV3 U30 ( .A(n1588), .Q(n1589) );
  NOR22 U31 ( .A(n249), .B(n2659), .Q(n285) );
  NOR21 U32 ( .A(n2743), .B(n127), .Q(n2708) );
  NAND22 U33 ( .A(n2690), .B(n1358), .Q(n2691) );
  NAND22 U34 ( .A(n1338), .B(n1422), .Q(u_alu_DP_OP_83J3_124_3384_n23) );
  INV3 U35 ( .A(u_alu_DP_OP_83J3_124_3384_n22), .Q(n1101) );
  INV6 U36 ( .A(n2976), .Q(n3053) );
  NAND26 U37 ( .A(n2465), .B(n1294), .Q(n1296) );
  NAND24 U38 ( .A(compare_i_data_rt_31_), .B(n1369), .Q(n1275) );
  INV6 U39 ( .A(u_alu_lt_x_11_n121), .Q(n1251) );
  INV3 U40 ( .A(n54), .Q(n2946) );
  BUF2 U41 ( .A(n56), .Q(n1320) );
  NAND22 U42 ( .A(n2361), .B(n2360), .Q(n2371) );
  NAND22 U43 ( .A(u_alu_ashr_4_A_16_), .B(u_alu_DP_OP_83J3_124_3384_n154), .Q(
        u_alu_DP_OP_83J3_124_3384_n55) );
  NOR22 U44 ( .A(n2638), .B(n2575), .Q(n2576) );
  INV6 U45 ( .A(n178), .Q(n597) );
  NAND22 U46 ( .A(alu_i_data_B[20]), .B(u_alu_DP_OP_85J3_126_1427_n374), .Q(
        u_alu_DP_OP_83J3_124_3384_n33) );
  INV6 U47 ( .A(n164), .Q(n165) );
  NAND23 U48 ( .A(n638), .B(u_alu_DP_OP_84J3_125_2615_n18), .Q(
        u_alu_DP_OP_84J3_125_2615_n16) );
  XNR21 U49 ( .A(n2263), .B(n2262), .Q(n2265) );
  NOR21 U50 ( .A(n1340), .B(n1344), .Q(n2357) );
  XOR21 U51 ( .A(n1904), .B(n358), .Q(n1905) );
  AOI211 U52 ( .A(u_alu_lt_x_11_n64), .B(n137), .C(n136), .Q(n135) );
  NAND22 U53 ( .A(n2754), .B(n1717), .Q(u_alu_lt_x_11_n10) );
  NAND31 U54 ( .A(n1740), .B(n1739), .C(n1738), .Q(n1741) );
  AOI211 U55 ( .A(n1358), .B(n1697), .C(n1696), .Q(n57) );
  INV3 U56 ( .A(n1061), .Q(n2159) );
  NAND23 U57 ( .A(n954), .B(n953), .Q(n952) );
  INV3 U58 ( .A(alu_i_data_B[19]), .Q(n1332) );
  INV3 U59 ( .A(i_data_immext[3]), .Q(n981) );
  INV3 U60 ( .A(n1309), .Q(n943) );
  INV3 U61 ( .A(n309), .Q(n2829) );
  INV3 U62 ( .A(n1205), .Q(n2066) );
  NOR22 U63 ( .A(n177), .B(n3059), .Q(n1987) );
  NOR23 U64 ( .A(n120), .B(n183), .Q(n119) );
  INV3 U65 ( .A(n177), .Q(n120) );
  INV3 U66 ( .A(n122), .Q(n121) );
  NAND22 U67 ( .A(n177), .B(n1369), .Q(n122) );
  NAND22 U68 ( .A(n1362), .B(n2259), .Q(n309) );
  NAND22 U69 ( .A(n2690), .B(n1359), .Q(n287) );
  NAND22 U70 ( .A(n1334), .B(i_data_FEalures[23]), .Q(n1578) );
  INV3 U71 ( .A(n1576), .Q(n1212) );
  NAND22 U72 ( .A(n170), .B(n1367), .Q(n2408) );
  NOR23 U73 ( .A(n1392), .B(n656), .Q(n52) );
  NAND33 U74 ( .A(n1503), .B(n1504), .C(n1575), .Q(n1111) );
  NAND26 U75 ( .A(n959), .B(n1512), .Q(n1517) );
  NAND22 U76 ( .A(n1321), .B(i_data_famemout[27]), .Q(n1512) );
  NAND22 U77 ( .A(n354), .B(n352), .Q(n2873) );
  NAND22 U78 ( .A(n2675), .B(n2674), .Q(n2985) );
  INV6 U79 ( .A(n1312), .Q(n547) );
  NOR21 U80 ( .A(n2786), .B(n193), .Q(u_alu_lt_x_11_n45) );
  NOR21 U81 ( .A(u_alu_lt_x_11_n39), .B(u_alu_lt_x_11_n41), .Q(
        u_alu_lt_x_11_n37) );
  INV3 U82 ( .A(n1263), .Q(n1794) );
  NAND22 U83 ( .A(i_data_immext[3]), .B(n170), .Q(n1866) );
  INV3 U84 ( .A(n2433), .Q(n1985) );
  NAND22 U85 ( .A(n1683), .B(i_data_immext[4]), .Q(n1080) );
  INV6 U86 ( .A(i_con_Ealuop[0]), .Q(n1665) );
  INV3 U87 ( .A(n2296), .Q(n1912) );
  IMUX21 U88 ( .A(n462), .B(n2143), .S(n2139), .Q(n461) );
  NAND22 U89 ( .A(n2025), .B(n1361), .Q(n2203) );
  NAND22 U90 ( .A(n1234), .B(n2830), .Q(n1236) );
  NAND22 U91 ( .A(n93), .B(n242), .Q(n1235) );
  NAND23 U92 ( .A(u_alu_ashr_4_A_6_), .B(n2090), .Q(n929) );
  NOR22 U93 ( .A(n184), .B(n1273), .Q(n1272) );
  INV3 U94 ( .A(n2097), .Q(n213) );
  NOR22 U95 ( .A(n1367), .B(n1746), .Q(n2227) );
  NAND33 U96 ( .A(n1496), .B(n150), .C(n149), .Q(n2498) );
  NAND22 U97 ( .A(n1545), .B(i_data_famemout[16]), .Q(n150) );
  INV3 U98 ( .A(n393), .Q(n392) );
  NOR22 U99 ( .A(n1361), .B(n909), .Q(n610) );
  NAND23 U100 ( .A(n2566), .B(n2565), .Q(n2605) );
  NOR21 U101 ( .A(n1364), .B(n2639), .Q(n381) );
  NAND22 U102 ( .A(n193), .B(n2786), .Q(u_alu_lt_x_11_n46) );
  NAND22 U103 ( .A(n2835), .B(n175), .Q(n2906) );
  INV3 U104 ( .A(n172), .Q(n247) );
  INV3 U105 ( .A(n2993), .Q(n2994) );
  INV3 U106 ( .A(n703), .Q(n2631) );
  OAI2111 U107 ( .A(n704), .B(n2587), .C(n2594), .D(n183), .Q(n703) );
  NOR23 U108 ( .A(n729), .B(n2095), .Q(n2396) );
  NAND22 U109 ( .A(n2146), .B(n161), .Q(n2033) );
  NAND22 U110 ( .A(u_alu_DP_OP_83J3_124_3384_n75), .B(
        u_alu_DP_OP_83J3_124_3384_n90), .Q(n132) );
  NAND22 U111 ( .A(n1190), .B(n2857), .Q(n2927) );
  AOI311 U112 ( .A(n1356), .B(n2718), .C(n2719), .D(i_data_immext[10]), .Q(
        n2695) );
  NAND22 U113 ( .A(n1921), .B(n1948), .Q(n1928) );
  NOR21 U114 ( .A(n2631), .B(n2630), .Q(n2599) );
  NAND26 U115 ( .A(n2223), .B(n2222), .Q(n2252) );
  INV3 U116 ( .A(n2259), .Q(n664) );
  NOR21 U117 ( .A(n2482), .B(n2480), .Q(n2238) );
  NOR21 U118 ( .A(n2238), .B(n2494), .Q(n2244) );
  NOR22 U119 ( .A(n234), .B(n2026), .Q(n2029) );
  INV3 U120 ( .A(n2459), .Q(n1254) );
  INV3 U121 ( .A(n1358), .Q(n83) );
  AOI211 U122 ( .A(u_alu_lt_x_11_n28), .B(u_alu_lt_x_11_n21), .C(
        u_alu_lt_x_11_n22), .Q(n139) );
  NOR21 U123 ( .A(n177), .B(n3012), .Q(n1808) );
  NAND22 U124 ( .A(n752), .B(n751), .Q(n750) );
  NOR21 U125 ( .A(n1251), .B(n217), .Q(n1797) );
  INV12 U126 ( .A(n160), .Q(n161) );
  NAND22 U127 ( .A(n1947), .B(n1948), .Q(n1961) );
  NAND24 U128 ( .A(n1672), .B(n1724), .Q(n1730) );
  NAND22 U129 ( .A(n2021), .B(n1357), .Q(n2761) );
  NAND22 U130 ( .A(n2204), .B(n519), .Q(n2099) );
  INV3 U131 ( .A(n2227), .Q(n2056) );
  NOR23 U132 ( .A(n185), .B(n2639), .Q(n2218) );
  NOR21 U133 ( .A(n486), .B(n2946), .Q(n2234) );
  NAND33 U134 ( .A(n1302), .B(n972), .C(n1303), .Q(n1354) );
  NAND24 U135 ( .A(n631), .B(n629), .Q(n2367) );
  INV3 U136 ( .A(n328), .Q(n2516) );
  NAND23 U137 ( .A(n2549), .B(n1353), .Q(n2499) );
  NAND26 U138 ( .A(n931), .B(n930), .Q(n2550) );
  INV3 U139 ( .A(n2536), .Q(n931) );
  INV6 U140 ( .A(n193), .Q(n181) );
  NAND24 U141 ( .A(n715), .B(n717), .Q(n2762) );
  NOR23 U142 ( .A(n249), .B(n2020), .Q(n2717) );
  INV3 U143 ( .A(u_alu_DP_OP_85J3_126_1427_n377), .Q(n2780) );
  INV3 U144 ( .A(n2743), .Q(n126) );
  NOR22 U145 ( .A(u_alu_DP_OP_85J3_126_1427_n377), .B(
        u_alu_DP_OP_83J3_124_3384_n153), .Q(u_alu_DP_OP_83J3_124_3384_n15) );
  NAND22 U146 ( .A(n690), .B(n194), .Q(n2894) );
  NOR21 U147 ( .A(n2931), .B(n2855), .Q(n2861) );
  NOR22 U148 ( .A(n228), .B(n2947), .Q(n2968) );
  NAND23 U149 ( .A(n2947), .B(n228), .Q(n2993) );
  NOR21 U150 ( .A(n247), .B(n3066), .Q(n494) );
  NAND23 U151 ( .A(n2926), .B(n1307), .Q(u_alu_lt_x_11_B_28_) );
  NAND26 U152 ( .A(n2341), .B(n2340), .Q(n1299) );
  NAND23 U153 ( .A(n633), .B(n1135), .Q(n3057) );
  NAND22 U154 ( .A(n2987), .B(n1136), .Q(n1135) );
  AOI211 U155 ( .A(n1361), .B(u_alu_DP_OP_85J3_126_1427_n368), .C(n3013), .Q(
        n3016) );
  NAND22 U156 ( .A(u_alu_DP_OP_83J3_124_3384_n89), .B(
        u_alu_DP_OP_83J3_124_3384_n75), .Q(u_alu_DP_OP_83J3_124_3384_n11) );
  AOI211 U157 ( .A(n2894), .B(u_alu_lt_x_11_n26), .C(n2931), .Q(n2897) );
  INV6 U158 ( .A(n1092), .Q(n2843) );
  NOR22 U159 ( .A(n1392), .B(n656), .Q(n1305) );
  NAND22 U160 ( .A(n1861), .B(n227), .Q(n2463) );
  NOR23 U161 ( .A(n2805), .B(n2495), .Q(n1624) );
  AOI211 U162 ( .A(u_alu_lt_x_11_n89), .B(u_alu_lt_x_11_n82), .C(
        u_alu_lt_x_11_n83), .Q(n142) );
  AOI211 U163 ( .A(u_alu_lt_x_11_n116), .B(u_alu_lt_x_11_n110), .C(
        u_alu_lt_x_11_n111), .Q(n143) );
  NOR21 U164 ( .A(n140), .B(u_alu_lt_x_11_n5), .Q(u_alu_lt_x_11_n3) );
  NAND22 U165 ( .A(u_alu_lt_x_11_n21), .B(u_alu_lt_x_11_n27), .Q(n140) );
  AOI211 U166 ( .A(n1358), .B(n1697), .C(n1696), .Q(n1750) );
  NAND22 U167 ( .A(n625), .B(n1356), .Q(n1711) );
  NOR21 U168 ( .A(n1848), .B(n1854), .Q(n1828) );
  INV6 U169 ( .A(n1830), .Q(n1823) );
  NOR21 U170 ( .A(n1366), .B(n2567), .Q(n1841) );
  NOR31 U171 ( .A(n1976), .B(n1974), .C(n1975), .Q(n1973) );
  NOR21 U172 ( .A(i_data_immext[10]), .B(n1893), .Q(n1969) );
  NOR21 U173 ( .A(n1366), .B(n1360), .Q(n2955) );
  XNR21 U174 ( .A(n2185), .B(n2347), .Q(n2199) );
  INV12 U175 ( .A(n1342), .Q(n3047) );
  NAND22 U176 ( .A(n757), .B(n756), .Q(n2310) );
  NOR22 U177 ( .A(u_alu_DP_OP_83J3_124_3384_n154), .B(u_alu_ashr_4_A_16_), .Q(
        u_alu_DP_OP_83J3_124_3384_n54) );
  INV3 U178 ( .A(n2516), .Q(n993) );
  NAND22 U179 ( .A(n2660), .B(n168), .Q(n2661) );
  XNR21 U180 ( .A(n2708), .B(n2707), .Q(n2709) );
  NOR22 U181 ( .A(n541), .B(n539), .Q(n1239) );
  NAND22 U182 ( .A(n2729), .B(n1356), .Q(n2730) );
  INV3 U183 ( .A(n2751), .Q(n130) );
  NAND22 U184 ( .A(n129), .B(n2747), .Q(n124) );
  NOR23 U185 ( .A(n131), .B(n2790), .Q(n2751) );
  INV3 U186 ( .A(u_alu_lt_x_11_n40), .Q(n131) );
  AOI221 U187 ( .A(n2916), .B(n1367), .C(n824), .D(n177), .Q(n2833) );
  INV6 U188 ( .A(n1192), .Q(n2928) );
  NAND22 U189 ( .A(n1326), .B(n2881), .Q(n2882) );
  AOI211 U190 ( .A(n3033), .B(n2993), .C(n2968), .Q(n2970) );
  NOR22 U191 ( .A(n889), .B(n3007), .Q(n260) );
  INV3 U192 ( .A(n3045), .Q(n85) );
  NOR22 U193 ( .A(n3038), .B(n3032), .Q(n3044) );
  INV3 U194 ( .A(n3046), .Q(n3041) );
  NAND22 U195 ( .A(n1263), .B(n1264), .Q(n1550) );
  NOR23 U196 ( .A(i_data_FEalures[10]), .B(n1349), .Q(n438) );
  BUF2 U197 ( .A(n708), .Q(n60) );
  NAND22 U198 ( .A(n1565), .B(n1564), .Q(n1566) );
  NOR21 U199 ( .A(n2530), .B(n2532), .Q(n1565) );
  NOR21 U200 ( .A(n2533), .B(n2531), .Q(n1564) );
  BUF2 U201 ( .A(n330), .Q(n53) );
  BUF2 U202 ( .A(n1612), .Q(n65) );
  INV3 U203 ( .A(n1113), .Q(n1112) );
  NAND22 U204 ( .A(n1598), .B(n1597), .Q(n1569) );
  NAND22 U205 ( .A(n240), .B(n791), .Q(n1200) );
  NAND23 U206 ( .A(n467), .B(n1522), .Q(n1523) );
  NAND22 U207 ( .A(n1990), .B(n1356), .Q(n1991) );
  NAND22 U208 ( .A(n269), .B(n2111), .Q(n268) );
  NAND22 U209 ( .A(n1033), .B(n1344), .Q(n1032) );
  XNR21 U210 ( .A(n2272), .B(n2271), .Q(n1033) );
  XNR21 U211 ( .A(n2278), .B(n1181), .Q(n839) );
  IMUX21 U212 ( .A(n2286), .B(n2285), .S(n1320), .Q(n2293) );
  NOR21 U213 ( .A(n872), .B(n173), .Q(n2285) );
  AOI221 U214 ( .A(n1357), .B(n2603), .C(n2557), .D(n1356), .Q(n2580) );
  NOR22 U215 ( .A(n2633), .B(n597), .Q(n1105) );
  XNR21 U216 ( .A(u_alu_DP_OP_83J3_124_3384_n4), .B(
        u_alu_DP_OP_83J3_124_3384_n93), .Q(u_alu_pre_sum_3b[5]) );
  XNR21 U217 ( .A(u_alu_DP_OP_83J3_124_3384_n3), .B(
        u_alu_DP_OP_83J3_124_3384_n86), .Q(u_alu_pre_sum_3b[6]) );
  AOI211 U218 ( .A(n624), .B(u_alu_DP_OP_84J3_125_2615_n81), .C(
        u_alu_DP_OP_84J3_125_2615_n86), .Q(n846) );
  NAND31 U219 ( .A(n799), .B(n3055), .C(n796), .Q(n795) );
  XNR21 U220 ( .A(n282), .B(n1024), .Q(n281) );
  INV12 U221 ( .A(compare_i_data_rs[14]), .Q(n233) );
  NAND22 U222 ( .A(n422), .B(n168), .Q(n421) );
  NAND22 U223 ( .A(n2265), .B(n2264), .Q(n2266) );
  AOI211 U224 ( .A(n1903), .B(n179), .C(n1902), .Q(n1907) );
  NOR22 U225 ( .A(n990), .B(n1567), .Q(n3077) );
  NOR22 U226 ( .A(n1199), .B(n1523), .Q(n3072) );
  NAND22 U227 ( .A(n1201), .B(n1200), .Q(n1199) );
  NAND31 U228 ( .A(u_alu_N306), .B(n1718), .C(u_alu_lt_x_11_n10), .Q(n1745) );
  OAI2111 U229 ( .A(n3006), .B(n1767), .C(n1766), .D(n1765), .Q(
        alu_o_data_AluRes[1]) );
  AOI221 U230 ( .A(n1774), .B(n1357), .C(n1751), .D(n1356), .Q(n1767) );
  AOI221 U231 ( .A(n249), .B(n1812), .C(n1774), .D(n1356), .Q(n1806) );
  AOI211 U232 ( .A(n1357), .B(n1990), .C(n1946), .Q(n1982) );
  XNR21 U233 ( .A(n2055), .B(n2054), .Q(n2080) );
  OAI2111 U234 ( .A(n1356), .B(n2176), .C(n2157), .D(n168), .Q(n2158) );
  NAND22 U235 ( .A(n2127), .B(n179), .Q(n2160) );
  NOR31 U236 ( .A(n2214), .B(n2213), .C(n2212), .Q(n983) );
  NAND22 U237 ( .A(n2215), .B(n168), .Q(n984) );
  NOR32 U238 ( .A(n2337), .B(n2338), .C(n2336), .Q(n2381) );
  NAND22 U239 ( .A(n949), .B(n948), .Q(alu_o_data_AluRes[17]) );
  AOI211 U240 ( .A(n1345), .B(n2541), .C(n2525), .Q(n948) );
  NAND23 U241 ( .A(n536), .B(u_alu_pre_sum_4a[2]), .Q(n2890) );
  NAND23 U242 ( .A(n536), .B(u_alu_pre_sum_4a[4]), .Q(n2964) );
  NAND23 U243 ( .A(n536), .B(u_alu_pre_sum_4a[6]), .Q(n3027) );
  INV3 U244 ( .A(n2937), .Q(n1) );
  NAND22 U245 ( .A(n200), .B(n1), .Q(n3003) );
  NAND22 U246 ( .A(n158), .B(i_data_rs[8]), .Q(n2) );
  INV3 U247 ( .A(n2), .Q(n67) );
  NOR31 U248 ( .A(n2141), .B(n212), .C(n2140), .Q(n3) );
  INV3 U249 ( .A(n3), .Q(n462) );
  CLKIN0 U250 ( .A(n185), .Q(n4) );
  OAI2110 U251 ( .A(n1118), .B(n1695), .C(n200), .D(n4), .Q(n752) );
  CLKIN0 U252 ( .A(n177), .Q(n5) );
  AOI221 U253 ( .A(n2204), .B(n172), .C(n1193), .D(n5), .Q(n1747) );
  NAND22 U254 ( .A(n1117), .B(n1435), .Q(n6) );
  INV3 U255 ( .A(n6), .Q(n1594) );
  INV3 U256 ( .A(n2622), .Q(n7) );
  IMUX21 U257 ( .A(n7), .B(n2434), .S(n1361), .Q(n2556) );
  INV3 U258 ( .A(n518), .Q(n8) );
  AOI211 U259 ( .A(n2164), .B(n8), .C(u_alu_lt_x_11_n90), .Q(n2124) );
  IMUX20 U260 ( .A(n3047), .B(n174), .S(n229), .Q(n9) );
  AOI210 U261 ( .A(n180), .B(n9), .C(n2977), .Q(n2257) );
  OAI222 U262 ( .A(n1350), .B(i_data_FEalures[3]), .C(n1324), .D(
        i_data_fbmemout[3]), .Q(n10) );
  INV3 U263 ( .A(n10), .Q(n1822) );
  AOI221 U264 ( .A(n89), .B(i_data_FMalures[23]), .C(i_data_rs[23]), .D(n159), 
        .Q(n1582) );
  AOI211 U265 ( .A(n3053), .B(n1830), .C(n2607), .Q(n11) );
  NAND20 U266 ( .A(n109), .B(n2594), .Q(n12) );
  NAND22 U267 ( .A(n11), .B(n12), .Q(n108) );
  NAND20 U268 ( .A(n1681), .B(i_con_Ealuop[0]), .Q(n13) );
  OAI210 U269 ( .A(i_con_Ealuop[3]), .B(n13), .C(i_con_Ealuop[1]), .Q(n1682)
         );
  INV3 U270 ( .A(n231), .Q(n14) );
  NAND33 U271 ( .A(n2409), .B(n2408), .C(n14), .Q(n2194) );
  NAND22 U272 ( .A(n189), .B(n216), .Q(n15) );
  NAND22 U273 ( .A(n1922), .B(n15), .Q(n1949) );
  OAI222 U274 ( .A(n1324), .B(i_data_fbmemout[15]), .C(i_data_FEalures[15]), 
        .D(n1349), .Q(n16) );
  INV3 U275 ( .A(n16), .Q(n521) );
  CLKIN0 U276 ( .A(n166), .Q(n17) );
  OAI222 U277 ( .A(n185), .B(n1747), .C(n2056), .D(n17), .Q(n1882) );
  OAI212 U278 ( .A(n1359), .B(n1916), .C(n830), .Q(n18) );
  INV3 U279 ( .A(n18), .Q(n1945) );
  XNR20 U280 ( .A(n2754), .B(n290), .Q(u_alu_DP_OP_84J3_125_2615_n1) );
  CLKIN0 U281 ( .A(n2083), .Q(n19) );
  OAI210 U282 ( .A(n2124), .B(n2083), .C(n179), .Q(n20) );
  AOI211 U283 ( .A(n2082), .B(n19), .C(n20), .Q(n2086) );
  IMUX20 U284 ( .A(n3047), .B(n174), .S(n2481), .Q(n21) );
  AOI210 U285 ( .A(n180), .B(n21), .C(n2946), .Q(n2214) );
  CLKIN0 U286 ( .A(n2281), .Q(n22) );
  AOI211 U287 ( .A(n2290), .B(n22), .C(n2289), .Q(n2291) );
  NAND20 U288 ( .A(n2782), .B(n65), .Q(n23) );
  CLKIN0 U289 ( .A(n23), .Q(n3080) );
  AOI210 U290 ( .A(n2904), .B(n174), .C(n173), .Q(n2129) );
  AOI210 U291 ( .A(n2693), .B(n174), .C(n173), .Q(n1919) );
  AOI210 U292 ( .A(n217), .B(n174), .C(n173), .Q(n1754) );
  CLKIN0 U293 ( .A(n2099), .Q(n24) );
  AOI210 U294 ( .A(n316), .B(n190), .C(n24), .Q(n1152) );
  CLKIN0 U295 ( .A(n1714), .Q(n25) );
  NOR30 U296 ( .A(n1304), .B(n1715), .C(n25), .Q(n1684) );
  AOI210 U297 ( .A(n1823), .B(n174), .C(n173), .Q(n26) );
  NAND20 U298 ( .A(n1823), .B(n2643), .Q(n27) );
  IMUX20 U299 ( .A(n27), .B(n26), .S(u_alu_lt_x_11_A_3_), .Q(n1834) );
  IMUX20 U300 ( .A(n3047), .B(n174), .S(n233), .Q(n28) );
  AOI210 U301 ( .A(n180), .B(n28), .C(n2287), .Q(n2292) );
  CLKIN0 U302 ( .A(u_alu_DP_OP_83J3_124_3384_n55), .Q(n29) );
  NOR20 U303 ( .A(u_alu_DP_OP_83J3_124_3384_n54), .B(n29), .Q(
        u_alu_pre_sum_3a[0]) );
  NOR23 U304 ( .A(n145), .B(n1541), .Q(n33) );
  NOR23 U305 ( .A(n145), .B(n1541), .Q(n3071) );
  BUF6 U306 ( .A(n1372), .Q(n34) );
  NAND24 U307 ( .A(u_alu_pre_sum_3b[2]), .B(n2714), .Q(n2584) );
  NOR24 U308 ( .A(n112), .B(n111), .Q(n2641) );
  NAND26 U309 ( .A(n1208), .B(n1207), .Q(n843) );
  INV3 U310 ( .A(n1093), .Q(n35) );
  AOI212 U311 ( .A(n1958), .B(n1961), .C(n1957), .Q(n1959) );
  NOR24 U312 ( .A(n1314), .B(n1044), .Q(n1924) );
  NAND22 U313 ( .A(n3089), .B(n37), .Q(n38) );
  NAND22 U314 ( .A(n36), .B(n184), .Q(n39) );
  NAND22 U315 ( .A(n38), .B(n39), .Q(n762) );
  INV3 U316 ( .A(n3089), .Q(n36) );
  INV3 U317 ( .A(n184), .Q(n37) );
  INV15 U318 ( .A(n117), .Q(n184) );
  BUF6 U319 ( .A(n1346), .Q(n48) );
  NOR23 U320 ( .A(DP_OP_68_131_7244_n70), .B(n2481), .Q(n2483) );
  NOR22 U321 ( .A(n2481), .B(n2274), .Q(n2421) );
  NAND23 U322 ( .A(n1420), .B(n1369), .Q(n1046) );
  NAND33 U323 ( .A(n1049), .B(n1323), .C(n1045), .Q(n2778) );
  NAND23 U324 ( .A(n688), .B(n2629), .Q(u_alu_DP_OP_83J3_124_3384_n45) );
  NAND22 U325 ( .A(n2558), .B(n2629), .Q(n2596) );
  NAND23 U326 ( .A(n2610), .B(n2609), .Q(n2611) );
  NOR23 U327 ( .A(n2600), .B(n597), .Q(n2616) );
  NOR22 U328 ( .A(n1366), .B(n185), .Q(n2330) );
  IMUX20 U329 ( .A(n1920), .B(n1919), .S(n1306), .Q(n1930) );
  AOI211 U330 ( .A(n3053), .B(n2025), .C(n2647), .Q(n2648) );
  INV6 U331 ( .A(u_alu_ashr_4_A_17_), .Q(n2517) );
  NAND22 U332 ( .A(n535), .B(n1364), .Q(n2569) );
  INV6 U333 ( .A(n3039), .Q(n1298) );
  NAND33 U334 ( .A(n2785), .B(n343), .C(u_alu_DP_OP_85J3_126_1427_n374), .Q(
        n2787) );
  NAND23 U335 ( .A(n2782), .B(n295), .Q(n2785) );
  NAND22 U336 ( .A(n578), .B(n2459), .Q(n577) );
  CLKIN4 U337 ( .A(n2458), .Q(n220) );
  NAND23 U338 ( .A(u_alu_lt_x_11_B_11_), .B(n242), .Q(n340) );
  NAND24 U339 ( .A(n1007), .B(n1434), .Q(n1005) );
  NOR23 U340 ( .A(i_data_FEalures[26]), .B(n1350), .Q(n1507) );
  NOR23 U341 ( .A(n1508), .B(n1507), .Q(n1600) );
  NAND24 U342 ( .A(n2299), .B(n836), .Q(n2334) );
  NAND23 U343 ( .A(n40), .B(n41), .Q(n42) );
  NAND24 U344 ( .A(n42), .B(n424), .Q(n1176) );
  INV3 U345 ( .A(u_alu_DP_OP_83J3_124_3384_n1), .Q(n40) );
  CLKIN4 U346 ( .A(u_alu_DP_OP_83J3_124_3384_n11), .Q(n41) );
  NAND26 U347 ( .A(n2537), .B(n1353), .Q(n933) );
  XNR22 U348 ( .A(n2999), .B(n2998), .Q(n3025) );
  NOR21 U349 ( .A(i_data_FEalures[29]), .B(n1350), .Q(n508) );
  NOR21 U350 ( .A(n992), .B(n2905), .Q(n3004) );
  NOR24 U351 ( .A(n2399), .B(n2398), .Q(n2400) );
  AOI212 U352 ( .A(n2199), .B(n202), .C(n1340), .Q(n989) );
  NAND34 U353 ( .A(n2648), .B(n677), .C(n675), .Q(n674) );
  NAND22 U354 ( .A(n44), .B(n45), .Q(n46) );
  NAND23 U355 ( .A(n46), .B(n2760), .Q(n2768) );
  INV3 U356 ( .A(n2761), .Q(n44) );
  NAND26 U357 ( .A(n1707), .B(n1307), .Q(u_alu_lt_x_11_B_24_) );
  NOR21 U358 ( .A(n2595), .B(n829), .Q(n2617) );
  NAND23 U359 ( .A(n2951), .B(n1356), .Q(n636) );
  NAND26 U360 ( .A(n925), .B(n921), .Q(n2951) );
  IMUX20 U361 ( .A(n2077), .B(n2076), .S(n2406), .Q(n2078) );
  NOR23 U362 ( .A(u_alu_lt_x_11_n90), .B(n361), .Q(n2477) );
  AOI221 U363 ( .A(n2173), .B(n1359), .C(n2118), .D(n1358), .Q(n2156) );
  NAND26 U364 ( .A(n47), .B(n327), .Q(n566) );
  NAND23 U365 ( .A(n1334), .B(i_data_FEalures[17]), .Q(n2527) );
  NOR21 U366 ( .A(u_alu_DP_OP_85J3_126_1427_n377), .B(n1196), .Q(n876) );
  NOR22 U367 ( .A(n268), .B(n267), .Q(n2122) );
  NOR31 U368 ( .A(i_data_rt[9]), .B(n49), .C(n1333), .Q(n1636) );
  XNR22 U369 ( .A(n1566), .B(n328), .Q(n1479) );
  NAND26 U370 ( .A(n1665), .B(i_con_Ealuop[1]), .Q(n1677) );
  NAND26 U371 ( .A(n1079), .B(n510), .Q(n1679) );
  OAI212 U372 ( .A(n43), .B(n187), .C(n278), .Q(n2773) );
  NAND24 U373 ( .A(n2910), .B(n185), .Q(n925) );
  NAND24 U374 ( .A(i_data_famemout[15]), .B(n1321), .Q(n47) );
  INV6 U375 ( .A(n1545), .Q(n55) );
  NAND23 U376 ( .A(n158), .B(i_data_rs[15]), .Q(n1400) );
  NOR24 U377 ( .A(i_data_rt[12]), .B(n1218), .Q(n1625) );
  INV3 U378 ( .A(n1043), .Q(n49) );
  INV6 U379 ( .A(i_con_Efbmux[0]), .Q(n1043) );
  NAND24 U380 ( .A(n223), .B(n1038), .Q(n2386) );
  AOI222 U381 ( .A(n2603), .B(n1356), .C(n2625), .D(n249), .Q(n2614) );
  NAND23 U382 ( .A(n2509), .B(n249), .Q(n302) );
  AOI211 U383 ( .A(n970), .B(u_alu_DP_OP_84J3_125_2615_n81), .C(
        u_alu_DP_OP_84J3_125_2615_n86), .Q(u_alu_DP_OP_84J3_125_2615_n23) );
  NAND23 U384 ( .A(n970), .B(n206), .Q(n638) );
  NAND24 U385 ( .A(u_alu_pre_sum_3a[4]), .B(n2715), .Q(n1108) );
  NAND23 U386 ( .A(n2913), .B(n2759), .Q(n2760) );
  BUF6 U387 ( .A(n2704), .Q(n50) );
  OAI212 U388 ( .A(n187), .B(u_alu_lt_x_11_B_29_), .C(n180), .Q(n2973) );
  IMUX20 U389 ( .A(n2973), .B(n2974), .S(n1052), .Q(n2975) );
  NOR22 U390 ( .A(n1361), .B(n2059), .Q(n1881) );
  NOR23 U391 ( .A(n1618), .B(n1617), .Q(n1621) );
  BUF8 U392 ( .A(u_alu_DP_OP_83J3_124_3384_n1), .Q(n271) );
  NOR24 U393 ( .A(n227), .B(n2025), .Q(n1936) );
  NAND23 U394 ( .A(n688), .B(n1361), .Q(n771) );
  NAND24 U395 ( .A(n2694), .B(n166), .Q(n2718) );
  BUF8 U396 ( .A(n1362), .Q(n248) );
  INV3 U397 ( .A(n1867), .Q(n1037) );
  BUF6 U398 ( .A(n2136), .Q(n51) );
  NAND23 U399 ( .A(n90), .B(i_data_FMalures[19]), .Q(n816) );
  NOR23 U400 ( .A(n1361), .B(n1988), .Q(n1843) );
  NAND33 U401 ( .A(n1582), .B(n1579), .C(n1578), .Q(n1417) );
  NAND23 U402 ( .A(n2319), .B(n718), .Q(n2716) );
  NOR23 U403 ( .A(n2710), .B(n1237), .Q(n2711) );
  NOR22 U404 ( .A(i_data_fbmemout[21]), .B(n1324), .Q(n1492) );
  NOR21 U405 ( .A(i_data_fbmemout[27]), .B(n1324), .Q(n1516) );
  NAND34 U406 ( .A(n1624), .B(n1369), .C(n1623), .Q(n994) );
  NOR22 U407 ( .A(n1329), .B(n2611), .Q(n2613) );
  NOR24 U408 ( .A(n1635), .B(n450), .Q(n3090) );
  NAND33 U409 ( .A(n1901), .B(n1900), .C(n1899), .Q(n1902) );
  NAND23 U410 ( .A(n2074), .B(n1224), .Q(n1223) );
  NOR23 U411 ( .A(n1361), .B(n1941), .Q(n348) );
  NOR22 U412 ( .A(n250), .B(n1391), .Q(n1392) );
  NAND22 U413 ( .A(n1334), .B(i_data_FEalures[26]), .Q(n1575) );
  NAND22 U414 ( .A(n1334), .B(n1407), .Q(n854) );
  INV12 U415 ( .A(n453), .Q(n2406) );
  NAND24 U416 ( .A(n546), .B(n118), .Q(n157) );
  NAND23 U417 ( .A(n64), .B(n1346), .Q(n63) );
  NAND22 U418 ( .A(n1612), .B(n859), .Q(n296) );
  NAND24 U419 ( .A(n883), .B(n882), .Q(n881) );
  NAND34 U420 ( .A(n886), .B(n3000), .C(n2999), .Q(n882) );
  NAND26 U421 ( .A(n2191), .B(n2178), .Q(n54) );
  NAND24 U422 ( .A(n2191), .B(n2178), .Q(DP_OP_68_131_7244_n70) );
  NOR23 U423 ( .A(u_alu_pre_sum_3b[8]), .B(n2822), .Q(n1025) );
  NAND23 U424 ( .A(n1669), .B(n1683), .Q(n430) );
  NAND22 U425 ( .A(n226), .B(u_alu_lt_x_11_B_24_), .Q(
        u_alu_DP_OP_84J3_125_2615_n50) );
  NAND24 U426 ( .A(n2468), .B(n813), .Q(n2469) );
  NOR23 U427 ( .A(n2188), .B(n2186), .Q(n1592) );
  NAND33 U428 ( .A(n720), .B(n721), .C(n719), .Q(n723) );
  INV6 U429 ( .A(n990), .Q(n1415) );
  NAND33 U430 ( .A(n3088), .B(n1594), .C(n1593), .Q(n1153) );
  NAND28 U431 ( .A(n1582), .B(n1581), .Q(u_alu_DP_OP_85J3_126_1427_n377) );
  INV12 U432 ( .A(u_alu_ashr_4_A_9_), .Q(n162) );
  NAND26 U433 ( .A(u_alu_ashr_4_A_9_), .B(n2406), .Q(n2164) );
  INV3 U434 ( .A(n1648), .Q(n1159) );
  NAND23 U435 ( .A(n491), .B(n178), .Q(n490) );
  NAND24 U436 ( .A(n879), .B(n884), .Q(n878) );
  INV8 U437 ( .A(n580), .Q(n3076) );
  INV15 U438 ( .A(n1301), .Q(n1302) );
  INV6 U439 ( .A(n1641), .Q(n1219) );
  INV15 U440 ( .A(n250), .Q(n1545) );
  NOR23 U441 ( .A(i_data_fbmemout[14]), .B(n246), .Q(n480) );
  NOR24 U442 ( .A(n166), .B(n3060), .Q(n716) );
  NAND22 U443 ( .A(n2065), .B(n2062), .Q(n1260) );
  NAND24 U444 ( .A(n2682), .B(n969), .Q(n2683) );
  NOR33 U445 ( .A(n2681), .B(n2680), .C(n2679), .Q(n2682) );
  NAND24 U446 ( .A(n377), .B(n2759), .Q(n376) );
  NOR24 U447 ( .A(n808), .B(n1549), .Q(n3096) );
  INV15 U448 ( .A(u_alu_lt_x_11_A_3_), .Q(n223) );
  NOR22 U449 ( .A(n1492), .B(n1493), .Q(n783) );
  NAND23 U450 ( .A(n3030), .B(u_alu_lt_x_11_n12), .Q(n3038) );
  INV3 U451 ( .A(n1054), .Q(n2996) );
  OAI212 U452 ( .A(u_alu_DP_OP_84J3_125_2615_n39), .B(
        u_alu_DP_OP_84J3_125_2615_n102), .C(u_alu_DP_OP_84J3_125_2615_n40), 
        .Q(u_alu_DP_OP_84J3_125_2615_n95) );
  INV3 U453 ( .A(n233), .Q(n56) );
  NAND23 U454 ( .A(u_alu_lt_x_11_B_1_), .B(n2830), .Q(n746) );
  NAND24 U455 ( .A(n738), .B(n737), .Q(n736) );
  NOR24 U456 ( .A(n438), .B(n550), .Q(n549) );
  NAND23 U457 ( .A(n648), .B(n647), .Q(n2549) );
  NOR22 U458 ( .A(n2805), .B(n649), .Q(n648) );
  NAND23 U459 ( .A(n922), .B(n1364), .Q(n921) );
  NAND24 U460 ( .A(n1204), .B(n1203), .Q(n1202) );
  NAND24 U461 ( .A(n2634), .B(n168), .Q(n1203) );
  NAND24 U462 ( .A(n244), .B(n59), .Q(n58) );
  INV6 U463 ( .A(n58), .Q(n1635) );
  INV15 U464 ( .A(i_data_FMalures[9]), .Q(n59) );
  INV8 U465 ( .A(n115), .Q(n244) );
  INV3 U466 ( .A(n2405), .Q(n2093) );
  NAND26 U467 ( .A(n230), .B(n259), .Q(n1538) );
  INV8 U468 ( .A(n3043), .Q(n1310) );
  NAND23 U469 ( .A(n618), .B(n2893), .Q(n2860) );
  XNR21 U470 ( .A(n2814), .B(n1310), .Q(n2815) );
  NAND22 U471 ( .A(n2693), .B(n221), .Q(n1948) );
  IMUX20 U472 ( .A(n3047), .B(n174), .S(n221), .Q(n1918) );
  AOI212 U473 ( .A(n1910), .B(n1909), .C(n166), .Q(n1911) );
  NAND24 U474 ( .A(n164), .B(n100), .Q(n99) );
  INV3 U475 ( .A(u_alu_DP_OP_83J3_124_3384_n11), .Q(n100) );
  INV8 U476 ( .A(n2843), .Q(n2638) );
  NAND24 U477 ( .A(u_alu_lt_x_11_n26), .B(n2932), .Q(n788) );
  NAND24 U478 ( .A(n3031), .B(n3030), .Q(n3001) );
  NOR23 U479 ( .A(n3001), .B(n1310), .Q(n888) );
  AOI212 U480 ( .A(n2486), .B(n2485), .C(n2484), .Q(n2487) );
  NOR24 U481 ( .A(i_data_FMalures[14]), .B(n116), .Q(n482) );
  NAND23 U482 ( .A(n3039), .B(n191), .Q(n937) );
  NAND26 U483 ( .A(n413), .B(n412), .Q(n437) );
  NOR23 U484 ( .A(n249), .B(n1891), .Q(n1838) );
  NAND24 U485 ( .A(n1891), .B(n1357), .Q(n382) );
  NOR23 U486 ( .A(n507), .B(n374), .Q(n373) );
  NOR22 U487 ( .A(n1358), .B(n2938), .Q(n2872) );
  NAND28 U488 ( .A(n1416), .B(n1415), .Q(n368) );
  AOI310 U489 ( .A(n121), .B(n1604), .C(n1603), .D(n119), .Q(n1131) );
  INV6 U490 ( .A(n1476), .Q(n61) );
  INV8 U491 ( .A(n61), .Q(n62) );
  NAND24 U492 ( .A(n657), .B(n1393), .Q(n656) );
  INV15 U493 ( .A(i_data_rt[11]), .Q(n64) );
  NOR24 U494 ( .A(n275), .B(n1639), .Q(n3091) );
  NAND28 U495 ( .A(n934), .B(n1205), .Q(n1639) );
  INV8 U496 ( .A(n1630), .Q(n1348) );
  NAND23 U497 ( .A(n2911), .B(n249), .Q(n2912) );
  INV3 U498 ( .A(n53), .Q(n3081) );
  AOI222 U499 ( .A(n2075), .B(n1358), .C(n1969), .D(n1359), .Q(n1978) );
  NAND24 U500 ( .A(n807), .B(n806), .Q(n2405) );
  AOI212 U501 ( .A(n79), .B(n2404), .C(n2406), .Q(n2096) );
  NOR23 U502 ( .A(n1561), .B(n1560), .Q(n695) );
  INV8 U503 ( .A(compare_i_data_rs[7]), .Q(n160) );
  NOR23 U504 ( .A(n2810), .B(n792), .Q(n2649) );
  AOI211 U505 ( .A(n2749), .B(n208), .C(n2748), .Q(n2750) );
  NOR23 U506 ( .A(n2848), .B(n2847), .Q(n2849) );
  NAND23 U507 ( .A(n1640), .B(n1369), .Q(n1641) );
  NOR24 U508 ( .A(n481), .B(n482), .Q(n66) );
  NOR23 U509 ( .A(n481), .B(n482), .Q(n475) );
  INV6 U510 ( .A(n1442), .Q(n481) );
  XNR22 U511 ( .A(u_alu_DP_OP_83J3_124_3384_n2), .B(n601), .Q(n595) );
  NAND24 U512 ( .A(n817), .B(n816), .Q(n815) );
  INV15 U513 ( .A(n3066), .Q(n167) );
  NAND26 U514 ( .A(n167), .B(n110), .Q(n1092) );
  NAND26 U515 ( .A(n679), .B(n1822), .Q(n1867) );
  NAND24 U516 ( .A(n2110), .B(n2112), .Q(n267) );
  NAND24 U517 ( .A(n683), .B(n207), .Q(n2112) );
  NAND26 U518 ( .A(n1184), .B(n1531), .Q(n2191) );
  NOR24 U519 ( .A(n1012), .B(n304), .Q(n386) );
  NAND23 U520 ( .A(n1010), .B(n1011), .Q(n304) );
  AOI211 U521 ( .A(n1335), .B(i_data_FEalures[5]), .C(n1380), .Q(n1383) );
  NAND22 U522 ( .A(n1334), .B(i_data_FEalures[20]), .Q(n1586) );
  NAND26 U523 ( .A(n514), .B(n511), .Q(n1732) );
  NAND22 U524 ( .A(n784), .B(n783), .Q(n1494) );
  NAND23 U525 ( .A(n2910), .B(n1364), .Q(n113) );
  NOR23 U526 ( .A(n1356), .B(n2671), .Q(n1933) );
  NAND24 U527 ( .A(n504), .B(n503), .Q(n995) );
  INV3 U528 ( .A(n1042), .Q(n667) );
  NAND23 U529 ( .A(alu_i_data_B[27]), .B(n196), .Q(n2932) );
  NAND22 U530 ( .A(alu_i_data_B[27]), .B(n175), .Q(n924) );
  NOR22 U531 ( .A(n1517), .B(alu_i_data_B[27]), .Q(
        u_alu_DP_OP_84J3_125_2615_n36) );
  AOI220 U532 ( .A(n224), .B(n1337), .C(alu_i_data_B[27]), .D(n196), .Q(n720)
         );
  NOR21 U533 ( .A(n2930), .B(n2892), .Q(n2900) );
  OAI210 U534 ( .A(n971), .B(n2908), .C(n192), .Q(n2909) );
  OAI210 U535 ( .A(n173), .B(n2608), .C(alu_i_data_B[19]), .Q(n2609) );
  NOR21 U536 ( .A(u_alu_lt_x_11_n53), .B(u_alu_lt_x_11_n55), .Q(
        u_alu_lt_x_11_n51) );
  NOR23 U537 ( .A(n1359), .B(n2727), .Q(n2728) );
  NAND24 U538 ( .A(n2443), .B(n1356), .Q(n1134) );
  XOR22 U539 ( .A(n3092), .B(n160), .Q(n334) );
  NAND23 U540 ( .A(n1346), .B(i_data_rt[31]), .Q(n851) );
  NAND24 U541 ( .A(n2953), .B(n2954), .Q(n562) );
  NAND24 U542 ( .A(n2868), .B(n243), .Q(n2954) );
  NOR24 U543 ( .A(n67), .B(n1462), .Q(n1595) );
  NAND26 U544 ( .A(n581), .B(n321), .Q(n1008) );
  NAND26 U545 ( .A(n378), .B(n376), .Q(n2724) );
  NOR23 U546 ( .A(n1107), .B(n674), .Q(n961) );
  NOR24 U547 ( .A(n110), .B(n2174), .Q(n2175) );
  AOI222 U548 ( .A(n252), .B(n2729), .C(n2692), .D(n537), .Q(n540) );
  NOR23 U549 ( .A(n192), .B(n187), .Q(n1142) );
  INV12 U550 ( .A(i_data_immext[5]), .Q(n1680) );
  INV6 U551 ( .A(n2642), .Q(n205) );
  NOR24 U552 ( .A(n779), .B(n781), .Q(n68) );
  INV12 U553 ( .A(n780), .Q(n779) );
  INV15 U554 ( .A(n2813), .Q(n186) );
  NAND28 U555 ( .A(n2792), .B(n2791), .Q(n2813) );
  INV15 U556 ( .A(n1324), .Q(n240) );
  NAND34 U557 ( .A(n2796), .B(n2789), .C(n2788), .Q(n2792) );
  NOR23 U558 ( .A(n1257), .B(n1254), .Q(n1869) );
  NAND24 U559 ( .A(n2458), .B(n1258), .Q(n1257) );
  NOR24 U560 ( .A(n1030), .B(n2294), .Q(n1029) );
  NAND24 U561 ( .A(n319), .B(n70), .Q(n69) );
  INV15 U562 ( .A(n69), .Q(n912) );
  INV15 U563 ( .A(n1550), .Q(n70) );
  NOR22 U564 ( .A(n320), .B(n1297), .Q(n319) );
  NAND22 U565 ( .A(u_alu_ashr_4_A_9_), .B(n1361), .Q(n299) );
  INV6 U566 ( .A(n1076), .Q(n1075) );
  NAND23 U567 ( .A(n90), .B(i_data_FMalures[12]), .Q(n342) );
  NAND22 U568 ( .A(n89), .B(i_data_FMalures[16]), .Q(n149) );
  AOI221 U569 ( .A(n89), .B(i_data_FMalures[29]), .C(n159), .D(i_data_rs[29]), 
        .Q(n1293) );
  NAND22 U570 ( .A(n90), .B(i_data_FMalures[7]), .Q(n1386) );
  OAI222 U571 ( .A(n1749), .B(n1358), .C(n1360), .D(n626), .Q(n625) );
  NAND23 U572 ( .A(n1883), .B(n1358), .Q(n1884) );
  NAND24 U573 ( .A(n536), .B(u_alu_pre_sum_4a[1]), .Q(n2853) );
  NAND24 U574 ( .A(n536), .B(u_alu_pre_sum_4a[3]), .Q(n2924) );
  INV15 U575 ( .A(n843), .Q(n536) );
  NAND24 U576 ( .A(n728), .B(n176), .Q(n727) );
  NAND23 U577 ( .A(n74), .B(n1346), .Q(n73) );
  NAND22 U578 ( .A(n1968), .B(n253), .Q(n731) );
  INV8 U579 ( .A(n2821), .Q(n2822) );
  NAND24 U580 ( .A(n1174), .B(n1995), .Q(n681) );
  NOR23 U581 ( .A(n1356), .B(n2863), .Q(n781) );
  XNR22 U582 ( .A(u_alu_DP_OP_83J3_124_3384_n2), .B(n600), .Q(n599) );
  BUF6 U583 ( .A(n198), .Q(n71) );
  BUF4 U584 ( .A(n2795), .Q(n72) );
  NOR23 U585 ( .A(n2703), .B(n2702), .Q(n2795) );
  AOI222 U586 ( .A(n90), .B(i_data_FMalures[10]), .C(n159), .D(i_data_rs[10]), 
        .Q(n1469) );
  INV15 U587 ( .A(n73), .Q(n2530) );
  INV15 U588 ( .A(i_data_rt[17]), .Q(n74) );
  OAI212 U589 ( .A(n3006), .B(n2942), .C(n2941), .Q(n2958) );
  NAND33 U590 ( .A(n1877), .B(n1876), .C(n297), .Q(alu_o_data_AluRes[4]) );
  INV3 U591 ( .A(n1994), .Q(n75) );
  INV3 U592 ( .A(n75), .Q(n76) );
  NAND24 U593 ( .A(n1630), .B(n1451), .Q(n1994) );
  NOR23 U594 ( .A(i_data_FMalures[25]), .B(n116), .Q(n1430) );
  NOR24 U595 ( .A(n1356), .B(n3017), .Q(n3018) );
  NOR22 U596 ( .A(n1318), .B(n1339), .Q(u_alu_DP_OP_83J3_124_3384_n29) );
  INV6 U597 ( .A(n549), .Q(n548) );
  INV6 U598 ( .A(i_con_Efamux[1]), .Q(n546) );
  AOI222 U599 ( .A(n536), .B(n281), .C(n1027), .D(n1021), .Q(n1023) );
  XOR22 U600 ( .A(u_alu_DP_OP_84J3_125_2615_n1), .B(n966), .Q(n1027) );
  INV8 U601 ( .A(n250), .Q(n1319) );
  NAND22 U602 ( .A(n1335), .B(i_data_FEalures[15]), .Q(n401) );
  NAND24 U603 ( .A(n1335), .B(i_data_FEalures[3]), .Q(n737) );
  NAND22 U604 ( .A(n1334), .B(i_data_FEalures[21]), .Q(n1585) );
  NAND22 U605 ( .A(n1334), .B(i_data_FEalures[25]), .Q(n1576) );
  NAND22 U606 ( .A(n1334), .B(i_data_FEalures[16]), .Q(n2497) );
  NAND26 U607 ( .A(n515), .B(n245), .Q(n1891) );
  NOR24 U608 ( .A(n2678), .B(n3066), .Q(n2679) );
  NOR20 U609 ( .A(n62), .B(n1477), .Q(n3086) );
  NOR23 U610 ( .A(n1654), .B(n1653), .Q(n1655) );
  NAND22 U611 ( .A(n1601), .B(n1600), .Q(n1568) );
  NAND33 U612 ( .A(n1601), .B(n1600), .C(n1369), .Q(n1602) );
  NAND23 U613 ( .A(n1624), .B(n1623), .Q(n1563) );
  NAND23 U614 ( .A(n613), .B(n2009), .Q(n612) );
  NAND22 U615 ( .A(n1176), .B(n2822), .Q(n1208) );
  NOR22 U616 ( .A(n1638), .B(n1636), .Q(n807) );
  NAND23 U617 ( .A(n1062), .B(n2149), .Q(n1061) );
  INV6 U618 ( .A(n1947), .Q(n1926) );
  INV6 U619 ( .A(n2233), .Q(n77) );
  INV6 U620 ( .A(n77), .Q(n78) );
  AOI212 U621 ( .A(n1359), .B(n2298), .C(n2175), .Q(n2233) );
  NAND26 U622 ( .A(n2981), .B(n1367), .Q(n557) );
  NAND33 U623 ( .A(n1343), .B(n207), .C(n2070), .Q(n1128) );
  NAND31 U624 ( .A(n2802), .B(n2801), .C(n1369), .Q(n2803) );
  INV6 U625 ( .A(n2798), .Q(n938) );
  AOI212 U626 ( .A(n2242), .B(n2843), .C(n2241), .Q(n2247) );
  INV12 U627 ( .A(compare_i_data_rs[2]), .Q(u_alu_lt_x_11_n122) );
  NAND28 U628 ( .A(n1109), .B(n2431), .Q(n2821) );
  NAND23 U629 ( .A(u_alu_lt_x_11_B_1_), .B(n1363), .Q(n840) );
  NOR32 U630 ( .A(n170), .B(n1652), .C(n1651), .Q(n1656) );
  NAND26 U631 ( .A(n99), .B(n424), .Q(u_alu_pre_sum_3b[8]) );
  NOR22 U632 ( .A(n328), .B(u_alu_ashr_4_A_17_), .Q(
        u_alu_DP_OP_83J3_124_3384_n52) );
  INV12 U633 ( .A(n1715), .Q(n2439) );
  NOR23 U634 ( .A(i_data_fbmemout[20]), .B(n246), .Q(n1610) );
  XNR22 U635 ( .A(compare_i_data_rs[5]), .B(n3094), .Q(n337) );
  INV12 U636 ( .A(compare_i_data_rs[5]), .Q(n234) );
  NAND33 U637 ( .A(n1383), .B(n1382), .C(n1381), .Q(compare_i_data_rs[5]) );
  NOR23 U638 ( .A(n1557), .B(n1008), .Q(n1007) );
  NAND28 U639 ( .A(n849), .B(n848), .Q(compare_i_data_rt_31_) );
  AOI222 U640 ( .A(n2830), .B(n92), .C(n688), .D(n242), .Q(n2565) );
  NOR21 U641 ( .A(n2590), .B(n2589), .Q(n2591) );
  NOR22 U642 ( .A(n2880), .B(n2879), .Q(n2881) );
  CLKIN4 U643 ( .A(i_data_immext[0]), .Q(n1864) );
  NAND24 U644 ( .A(n522), .B(n451), .Q(n450) );
  NAND26 U645 ( .A(n570), .B(n569), .Q(n934) );
  NOR23 U646 ( .A(n2629), .B(n688), .Q(u_alu_DP_OP_83J3_124_3384_n44) );
  INV8 U647 ( .A(n688), .Q(n2558) );
  NAND28 U648 ( .A(n696), .B(n695), .Q(n698) );
  INV3 U649 ( .A(n2093), .Q(n79) );
  NAND24 U650 ( .A(n349), .B(n347), .Q(n1883) );
  OAI210 U651 ( .A(u_alu_DP_OP_84J3_125_2615_n39), .B(
        u_alu_DP_OP_84J3_125_2615_n45), .C(u_alu_DP_OP_84J3_125_2615_n40), .Q(
        u_alu_DP_OP_84J3_125_2615_n38) );
  INV6 U652 ( .A(n2147), .Q(n427) );
  NAND22 U653 ( .A(n2087), .B(n1356), .Q(n1226) );
  NOR23 U654 ( .A(n1972), .B(n2010), .Q(n1975) );
  NOR24 U655 ( .A(n495), .B(n493), .Q(n489) );
  NAND23 U656 ( .A(n2216), .B(n166), .Q(n2217) );
  NOR23 U657 ( .A(n646), .B(n644), .Q(n643) );
  NAND28 U658 ( .A(n2967), .B(n1353), .Q(n2295) );
  NAND23 U659 ( .A(n2295), .B(n357), .Q(n914) );
  NAND23 U660 ( .A(n2341), .B(n2340), .Q(n2369) );
  INV6 U661 ( .A(n1448), .Q(n1449) );
  NOR23 U662 ( .A(i_data_FEalures[12]), .B(n1350), .Q(n1626) );
  NAND23 U663 ( .A(n2738), .B(n168), .Q(n594) );
  AOI212 U664 ( .A(n2016), .B(n168), .C(n2015), .Q(n2051) );
  NAND23 U665 ( .A(n1346), .B(n1547), .Q(n1548) );
  NOR22 U666 ( .A(n713), .B(n712), .Q(n711) );
  AOI221 U667 ( .A(n171), .B(n205), .C(n673), .D(n177), .Q(n80) );
  NAND26 U668 ( .A(n692), .B(n1241), .Q(n699) );
  NAND34 U669 ( .A(n1169), .B(n1724), .C(n1168), .Q(n1667) );
  INV12 U670 ( .A(n1308), .Q(n1309) );
  NAND26 U671 ( .A(n105), .B(n104), .Q(n1785) );
  NOR23 U672 ( .A(n637), .B(n1471), .Q(n665) );
  INV6 U673 ( .A(n410), .Q(n1184) );
  NOR24 U674 ( .A(n170), .B(n1625), .Q(n411) );
  OAI210 U675 ( .A(n2081), .B(u_alu_lt_x_11_n90), .C(n2164), .Q(
        u_alu_lt_x_11_n89) );
  INV6 U676 ( .A(n2874), .Q(n266) );
  INV6 U677 ( .A(n2726), .Q(n211) );
  NAND24 U678 ( .A(n2725), .B(n176), .Q(n2905) );
  NAND22 U679 ( .A(n2225), .B(n1365), .Q(n2226) );
  NAND24 U680 ( .A(n1251), .B(u_alu_lt_x_11_B_1_), .Q(n2384) );
  INV6 U681 ( .A(n2538), .Q(n932) );
  NAND24 U682 ( .A(n1888), .B(n1887), .Q(n1044) );
  NOR22 U683 ( .A(n1644), .B(n1556), .Q(n3094) );
  NOR23 U684 ( .A(n170), .B(n1644), .Q(n1646) );
  NAND26 U685 ( .A(n2493), .B(n2492), .Q(n974) );
  NAND23 U686 ( .A(n1452), .B(n244), .Q(n1993) );
  NOR32 U687 ( .A(n2418), .B(n2417), .C(n2416), .Q(n2429) );
  INV12 U688 ( .A(n92), .Q(n219) );
  NAND24 U689 ( .A(n1917), .B(n1356), .Q(n423) );
  NOR23 U690 ( .A(i_data_fbmemout[13]), .B(n246), .Q(n1472) );
  NOR23 U691 ( .A(i_data_FMalures[24]), .B(n1214), .Q(n1114) );
  NOR22 U692 ( .A(n1366), .B(n2329), .Q(n81) );
  INV8 U693 ( .A(n144), .Q(n2329) );
  NAND23 U694 ( .A(n2787), .B(n2786), .Q(n2788) );
  NOR24 U695 ( .A(n1358), .B(n1773), .Q(n1696) );
  NAND22 U696 ( .A(n82), .B(n83), .Q(n84) );
  NAND24 U697 ( .A(n84), .B(n1884), .Q(n1917) );
  INV3 U698 ( .A(n1944), .Q(n82) );
  NOR22 U699 ( .A(u_alu_lt_x_11_B_24_), .B(n226), .Q(
        u_alu_DP_OP_84J3_125_2615_n49) );
  NOR22 U700 ( .A(n1361), .B(n2563), .Q(n2866) );
  INV3 U701 ( .A(n1217), .Q(n114) );
  INV6 U702 ( .A(n1189), .Q(n226) );
  XOR20 U703 ( .A(n2649), .B(n2551), .Q(n919) );
  NOR22 U704 ( .A(i_data_FEalures[27]), .B(n1350), .Q(n1515) );
  NOR23 U705 ( .A(i_data_FEalures[25]), .B(n1350), .Q(n1432) );
  AOI211 U706 ( .A(n3039), .B(n3044), .C(n3042), .Q(n3040) );
  NAND28 U707 ( .A(n938), .B(n186), .Q(n3039) );
  NOR21 U708 ( .A(n1367), .B(n68), .Q(n2242) );
  NOR24 U709 ( .A(i_data_FMalures[11]), .B(n1214), .Q(n1627) );
  NAND24 U710 ( .A(n927), .B(n926), .Q(n2910) );
  OAI210 U711 ( .A(u_alu_lt_x_11_n102), .B(u_alu_lt_x_11_n99), .C(
        u_alu_lt_x_11_n100), .Q(u_alu_lt_x_11_n98) );
  NAND24 U712 ( .A(n832), .B(n831), .Q(n835) );
  NOR23 U713 ( .A(n239), .B(n2739), .Q(n1984) );
  INV6 U714 ( .A(n1196), .Q(n2739) );
  NAND24 U715 ( .A(n748), .B(n749), .Q(n2320) );
  NAND34 U716 ( .A(n604), .B(n2629), .C(n183), .Q(n605) );
  INV12 U717 ( .A(u_alu_lt_x_11_B_1_), .Q(n217) );
  NAND26 U718 ( .A(n3071), .B(n1369), .Q(n1700) );
  NAND24 U719 ( .A(n2948), .B(n166), .Q(n2949) );
  NAND23 U720 ( .A(n978), .B(n270), .Q(n2948) );
  NAND24 U721 ( .A(n2670), .B(n1356), .Q(n2640) );
  NOR23 U722 ( .A(i_data_fbmemout[9]), .B(n246), .Q(n1638) );
  NOR22 U723 ( .A(n1358), .B(n3056), .Q(n802) );
  NAND26 U724 ( .A(n1234), .B(n1363), .Q(n573) );
  NAND28 U725 ( .A(n1091), .B(n2302), .Q(n3021) );
  NAND26 U726 ( .A(n380), .B(n379), .Q(n2670) );
  NAND22 U727 ( .A(n3043), .B(n191), .Q(n618) );
  NAND23 U728 ( .A(n3045), .B(n86), .Q(n87) );
  NAND26 U729 ( .A(n85), .B(n3041), .Q(n88) );
  NAND24 U730 ( .A(n87), .B(n88), .Q(n3069) );
  INV3 U731 ( .A(n3041), .Q(n86) );
  NOR23 U732 ( .A(n844), .B(n3069), .Q(n1020) );
  INV15 U733 ( .A(n1119), .Q(n1351) );
  NOR23 U734 ( .A(n489), .B(n488), .Q(n487) );
  NAND26 U735 ( .A(n666), .B(n665), .Q(n2223) );
  NAND24 U736 ( .A(n443), .B(n441), .Q(n1812) );
  INV12 U737 ( .A(n1790), .Q(n1352) );
  NAND22 U738 ( .A(n2704), .B(n208), .Q(n129) );
  AOI211 U739 ( .A(n2457), .B(u_alu_lt_x_11_B_1_), .C(n220), .Q(n578) );
  NAND24 U740 ( .A(n2836), .B(n1358), .Q(n1077) );
  NOR22 U741 ( .A(n1222), .B(n542), .Q(n541) );
  NAND22 U742 ( .A(n1346), .B(n1473), .Q(n1474) );
  NAND22 U743 ( .A(n1630), .B(n1419), .Q(n1420) );
  NAND22 U744 ( .A(n1630), .B(n1431), .Q(n323) );
  NOR32 U745 ( .A(n170), .B(n1637), .C(n1635), .Q(n806) );
  NAND28 U746 ( .A(n1615), .B(n1614), .Q(n330) );
  XNR22 U747 ( .A(n2826), .B(n2827), .Q(n920) );
  NAND26 U748 ( .A(n2754), .B(n357), .Q(n2937) );
  AOI212 U749 ( .A(n499), .B(n498), .C(n3006), .Q(n497) );
  NOR24 U750 ( .A(n3006), .B(n2335), .Q(n2336) );
  NOR23 U751 ( .A(n1356), .B(n2437), .Q(n608) );
  NAND22 U752 ( .A(u_alu_lt_x_11_B_25_), .B(n1361), .Q(n1126) );
  NAND24 U753 ( .A(n2868), .B(n1356), .Q(n2914) );
  NAND24 U754 ( .A(n689), .B(n1621), .Q(n607) );
  NOR24 U755 ( .A(n170), .B(n1619), .Q(n689) );
  OAI212 U756 ( .A(n1367), .B(n3019), .C(n1358), .Q(n3020) );
  INV6 U757 ( .A(n1548), .Q(n1649) );
  NAND24 U758 ( .A(n2038), .B(n506), .Q(n505) );
  NOR24 U759 ( .A(n1854), .B(n2388), .Q(n2042) );
  NOR23 U760 ( .A(i_data_FMalures[27]), .B(n198), .Q(n1513) );
  NAND24 U761 ( .A(n2209), .B(n1356), .Q(n780) );
  NOR24 U762 ( .A(n1366), .B(n2644), .Q(n2225) );
  NAND24 U763 ( .A(n560), .B(n1358), .Q(n2869) );
  NAND24 U764 ( .A(n2952), .B(n561), .Q(n560) );
  CLKIN4 U765 ( .A(n771), .Q(n770) );
  INV12 U766 ( .A(n1350), .Q(n237) );
  INV6 U767 ( .A(i_con_Efbmux[1]), .Q(n1372) );
  NOR22 U768 ( .A(n177), .B(n2567), .Q(n2571) );
  NAND24 U769 ( .A(n877), .B(n892), .Q(n880) );
  NOR22 U770 ( .A(i_data_fbmemout[1]), .B(n246), .Q(n1654) );
  NOR22 U771 ( .A(i_data_fbmemout[4]), .B(n246), .Q(n1443) );
  NOR22 U772 ( .A(i_data_fbmemout[10]), .B(n246), .Q(n1634) );
  NAND23 U773 ( .A(n2216), .B(n176), .Q(n2671) );
  NAND24 U774 ( .A(n841), .B(n840), .Q(n2216) );
  NAND33 U775 ( .A(n2711), .B(n2712), .C(n2713), .Q(alu_o_data_AluRes[22]) );
  NOR33 U776 ( .A(n170), .B(n2532), .C(n2533), .Q(n1622) );
  NAND28 U777 ( .A(n344), .B(n1353), .Q(n1339) );
  NAND26 U778 ( .A(n1191), .B(n784), .Q(n344) );
  AOI212 U779 ( .A(n1885), .B(n1356), .C(n3006), .Q(n1886) );
  NOR24 U780 ( .A(n526), .B(n524), .Q(n1885) );
  NAND28 U781 ( .A(n238), .B(n606), .Q(n604) );
  NAND23 U782 ( .A(i_con_Efbmux[0]), .B(i_con_Efbmux[1]), .Q(n1790) );
  NOR24 U783 ( .A(n1358), .B(n726), .Q(n877) );
  NAND24 U784 ( .A(u_alu_ashr_4_A_16_), .B(n1361), .Q(n669) );
  NAND23 U785 ( .A(n880), .B(n878), .Q(n261) );
  BUF6 U786 ( .A(i_data_immext[7]), .Q(n1359) );
  INV8 U787 ( .A(i_data_immext[7]), .Q(n1358) );
  INV8 U788 ( .A(i_data_immext[6]), .Q(n1356) );
  INV3 U789 ( .A(n1356), .Q(n154) );
  BUF2 U790 ( .A(i_data_immext[7]), .Q(n1360) );
  INV12 U791 ( .A(n1370), .Q(n170) );
  CLKBU15 U792 ( .A(n1370), .Q(n1369) );
  INV3 U793 ( .A(n170), .Q(n859) );
  INV12 U794 ( .A(i_con_Ealusrc), .Q(n1370) );
  BUF6 U795 ( .A(n1365), .Q(n1364) );
  INV6 U796 ( .A(n1365), .Q(n185) );
  NAND24 U797 ( .A(n1368), .B(i_data_immext[16]), .Q(n2966) );
  INV3 U798 ( .A(n2406), .Q(n218) );
  INV3 U799 ( .A(n1358), .Q(n110) );
  BUF6 U800 ( .A(i_data_immext[6]), .Q(n249) );
  NAND28 U801 ( .A(n1712), .B(n972), .Q(n3006) );
  INV12 U802 ( .A(n1362), .Q(n1361) );
  INV3 U803 ( .A(n1318), .Q(n2786) );
  NAND28 U804 ( .A(n1714), .B(n1713), .Q(n3066) );
  BUF2 U805 ( .A(u_alu_lt_x_11_A_31_), .Q(n290) );
  INV6 U806 ( .A(u_alu_lt_x_11_A_31_), .Q(n1717) );
  INV6 U807 ( .A(n1337), .Q(n3012) );
  NAND26 U808 ( .A(n1497), .B(n2497), .Q(u_alu_DP_OP_83J3_124_3384_n154) );
  INV3 U809 ( .A(n2548), .Q(n2808) );
  INV6 U810 ( .A(n1070), .Q(n2287) );
  INV3 U811 ( .A(n2439), .Q(n214) );
  INV3 U812 ( .A(n1363), .Q(n200) );
  INV6 U813 ( .A(u_alu_lt_x_11_A_0_), .Q(n857) );
  INV6 U814 ( .A(n1340), .Q(n207) );
  INV8 U815 ( .A(n2823), .Q(n1340) );
  INV3 U816 ( .A(n1353), .Q(n225) );
  INV6 U817 ( .A(n239), .Q(n183) );
  NOR24 U818 ( .A(i_data_FMalures[19]), .B(n116), .Q(n2590) );
  INV3 U819 ( .A(n2744), .Q(n127) );
  INV6 U820 ( .A(n1165), .Q(n151) );
  BUF8 U821 ( .A(n2193), .Q(n316) );
  CLKIN4 U822 ( .A(n2193), .Q(n519) );
  NOR21 U823 ( .A(n249), .B(n1366), .Q(n2759) );
  NAND22 U824 ( .A(n237), .B(n478), .Q(n477) );
  OAI212 U825 ( .A(u_alu_DP_OP_83J3_124_3384_n32), .B(n165), .C(
        u_alu_DP_OP_83J3_124_3384_n33), .Q(u_alu_DP_OP_83J3_124_3384_n93) );
  INV15 U826 ( .A(n2279), .Q(n1343) );
  NOR24 U827 ( .A(i_data_FEalures[8]), .B(n1349), .Q(n2063) );
  BUF15 U828 ( .A(n2526), .Q(n89) );
  BUF15 U829 ( .A(n2526), .Q(n90) );
  NAND24 U830 ( .A(n437), .B(n411), .Q(n410) );
  NOR33 U831 ( .A(n1068), .B(n1067), .C(n1066), .Q(n1163) );
  NAND24 U832 ( .A(n2911), .B(n767), .Q(n2953) );
  NAND24 U833 ( .A(n772), .B(n769), .Q(n2911) );
  NOR32 U834 ( .A(n170), .B(n2533), .C(n2532), .Q(n2534) );
  NAND23 U835 ( .A(n1399), .B(n1400), .Q(n565) );
  INV6 U836 ( .A(n1087), .Q(n388) );
  NAND24 U837 ( .A(n1261), .B(n2062), .Q(n2163) );
  NAND28 U838 ( .A(n1186), .B(n1185), .Q(n1261) );
  NAND24 U839 ( .A(n963), .B(n209), .Q(n757) );
  XOR22 U840 ( .A(n1937), .B(n420), .Q(n419) );
  NAND26 U841 ( .A(n1084), .B(n1456), .Q(n1863) );
  NAND23 U842 ( .A(n1086), .B(n1085), .Q(n1084) );
  CLKIN4 U843 ( .A(n1455), .Q(n1456) );
  NAND26 U844 ( .A(n1388), .B(n811), .Q(compare_i_data_rs[7]) );
  XNR22 U845 ( .A(n2896), .B(n2895), .Q(n2922) );
  NAND24 U846 ( .A(n2499), .B(n2808), .Q(n2543) );
  NAND24 U847 ( .A(n1272), .B(n2411), .Q(n660) );
  NAND26 U848 ( .A(n2137), .B(n2136), .Q(n2411) );
  NAND23 U849 ( .A(n54), .B(n1363), .Q(n670) );
  NOR31 U850 ( .A(n2488), .B(n2479), .C(n2480), .Q(n2490) );
  INV6 U851 ( .A(n203), .Q(n2834) );
  OAI212 U852 ( .A(u_alu_DP_OP_83J3_124_3384_n25), .B(n165), .C(
        u_alu_DP_OP_83J3_124_3384_n26), .Q(u_alu_DP_OP_83J3_124_3384_n86) );
  NOR23 U853 ( .A(n1364), .B(n2676), .Q(n2697) );
  NOR23 U854 ( .A(n166), .B(n2676), .Q(n306) );
  NAND24 U855 ( .A(n972), .B(n1089), .Q(n91) );
  NOR24 U856 ( .A(n320), .B(n1794), .Q(n104) );
  NOR24 U857 ( .A(i_data_FMalures[2]), .B(n198), .Q(n320) );
  NAND34 U858 ( .A(n1995), .B(n1993), .C(n655), .Q(n911) );
  NOR24 U859 ( .A(n241), .B(n274), .Q(n655) );
  NAND23 U860 ( .A(n2928), .B(n194), .Q(n721) );
  NAND26 U861 ( .A(n194), .B(n1194), .Q(n719) );
  INV15 U862 ( .A(u_alu_lt_x_11_A_13_), .Q(n229) );
  OAI210 U863 ( .A(n2365), .B(n2364), .C(n2363), .Q(n628) );
  NAND24 U864 ( .A(n2025), .B(n197), .Q(n735) );
  NOR23 U865 ( .A(n1422), .B(n1338), .Q(u_alu_DP_OP_83J3_124_3384_n22) );
  NAND26 U866 ( .A(n1143), .B(n1422), .Q(n1144) );
  NAND28 U867 ( .A(n232), .B(n1584), .Q(n1422) );
  NOR24 U868 ( .A(n224), .B(n1337), .Q(n2931) );
  INV15 U869 ( .A(n1509), .Q(n224) );
  BUF15 U870 ( .A(n93), .Q(n92) );
  NOR24 U871 ( .A(n92), .B(n231), .Q(n2394) );
  NAND24 U872 ( .A(n92), .B(n169), .Q(n672) );
  NAND20 U873 ( .A(n231), .B(n93), .Q(n383) );
  NAND28 U874 ( .A(n2409), .B(n2408), .Q(n93) );
  NOR24 U875 ( .A(n2280), .B(n94), .Q(n2563) );
  NOR24 U876 ( .A(n96), .B(n447), .Q(n94) );
  NAND24 U877 ( .A(n477), .B(n95), .Q(n447) );
  CLKIN6 U878 ( .A(n480), .Q(n95) );
  NAND24 U879 ( .A(n66), .B(n1369), .Q(n96) );
  CLKIN6 U880 ( .A(n1315), .Q(n513) );
  NAND24 U881 ( .A(n1675), .B(n1670), .Q(n1315) );
  NAND24 U882 ( .A(n98), .B(n97), .Q(n1670) );
  CLKIN3 U883 ( .A(n1016), .Q(n97) );
  NOR23 U884 ( .A(n1015), .B(n1864), .Q(n98) );
  INV6 U885 ( .A(n259), .Q(n102) );
  NAND28 U886 ( .A(n101), .B(n103), .Q(n259) );
  INV4 U887 ( .A(n1324), .Q(n101) );
  NOR24 U888 ( .A(n2001), .B(n102), .Q(n1642) );
  CLKIN4 U889 ( .A(i_data_fbmemout[7]), .Q(n103) );
  NAND28 U890 ( .A(n1785), .B(n1791), .Q(n1234) );
  CLKIN6 U891 ( .A(n777), .Q(n105) );
  NOR22 U892 ( .A(u_alu_lt_x_11_n122), .B(n1234), .Q(n2460) );
  NOR42 U893 ( .A(n1652), .B(n1654), .C(n1651), .D(n1653), .Q(n3097) );
  AOI212 U894 ( .A(n2677), .B(n203), .C(n108), .Q(n2610) );
  NAND24 U895 ( .A(n107), .B(n106), .Q(n2677) );
  AOI222 U896 ( .A(n2604), .B(n1367), .C(n2605), .D(n243), .Q(n106) );
  OAI212 U897 ( .A(n112), .B(n111), .C(n2759), .Q(n107) );
  CLKIN10 U898 ( .A(n973), .Q(n173) );
  CLKIN6 U899 ( .A(n3066), .Q(n2883) );
  OAI212 U900 ( .A(n1330), .B(n187), .C(n973), .Q(n109) );
  NOR24 U901 ( .A(n110), .B(n3066), .Q(n203) );
  OAI222 U902 ( .A(n1815), .B(n249), .C(n1356), .D(n1814), .Q(n2604) );
  AOI212 U903 ( .A(n955), .B(n956), .C(n176), .Q(n111) );
  CLKIN6 U904 ( .A(n113), .Q(n112) );
  NAND31 U905 ( .A(n1612), .B(n2782), .C(n1369), .Q(n684) );
  NOR24 U906 ( .A(n1610), .B(n1609), .Q(n2782) );
  NAND28 U907 ( .A(n114), .B(n1372), .Q(n115) );
  BUF15 U908 ( .A(n115), .Q(n116) );
  BUF15 U909 ( .A(n115), .Q(n1214) );
  NAND24 U910 ( .A(n317), .B(n1469), .Q(n117) );
  CLKIN6 U911 ( .A(n184), .Q(n231) );
  CLKIN3 U912 ( .A(i_con_Efamux[0]), .Q(n118) );
  NAND26 U913 ( .A(n1689), .B(n183), .Q(n123) );
  NAND34 U914 ( .A(n1603), .B(n1604), .C(n1369), .Q(n1689) );
  NOR24 U915 ( .A(n1432), .B(n1433), .Q(n1603) );
  NOR24 U916 ( .A(n322), .B(n1430), .Q(n1604) );
  XOR22 U917 ( .A(n130), .B(n124), .Q(n2753) );
  NOR24 U918 ( .A(n128), .B(n125), .Q(n2747) );
  OAI212 U919 ( .A(n127), .B(n2741), .C(n126), .Q(n125) );
  NOR24 U920 ( .A(n127), .B(n2742), .Q(n128) );
  OAI212 U921 ( .A(n2632), .B(n2650), .C(n2812), .Q(n2704) );
  NOR24 U922 ( .A(n2739), .B(n2740), .Q(n2790) );
  NAND33 U923 ( .A(n521), .B(n2339), .C(n1369), .Q(n2341) );
  NOR24 U924 ( .A(n1449), .B(n700), .Q(n2339) );
  CLKIN6 U925 ( .A(n132), .Q(n425) );
  OAI212 U926 ( .A(u_alu_DP_OP_83J3_124_3384_n29), .B(
        u_alu_DP_OP_83J3_124_3384_n33), .C(u_alu_DP_OP_83J3_124_3384_n30), .Q(
        u_alu_DP_OP_83J3_124_3384_n90) );
  NOR24 U927 ( .A(u_alu_DP_OP_83J3_124_3384_n15), .B(
        u_alu_DP_OP_83J3_124_3384_n22), .Q(u_alu_DP_OP_83J3_124_3384_n75) );
  OAI212 U928 ( .A(n135), .B(u_alu_lt_x_11_n1), .C(n133), .Q(u_alu_N306) );
  AOI212 U929 ( .A(u_alu_lt_x_11_n34), .B(u_alu_lt_x_11_n3), .C(n134), .Q(n133) );
  OAI212 U930 ( .A(u_alu_lt_x_11_n5), .B(n139), .C(n138), .Q(n134) );
  OAI212 U931 ( .A(u_alu_lt_x_11_n66), .B(n142), .C(n141), .Q(n136) );
  OAI212 U932 ( .A(u_alu_lt_x_11_n95), .B(n143), .C(u_alu_lt_x_11_n96), .Q(
        n137) );
  AOI211 U933 ( .A(u_alu_lt_x_11_n75), .B(u_alu_lt_x_11_n68), .C(
        u_alu_lt_x_11_n69), .Q(n141) );
  AOI211 U934 ( .A(u_alu_lt_x_11_n14), .B(u_alu_lt_x_11_n7), .C(
        u_alu_lt_x_11_n8), .Q(n138) );
  NAND24 U935 ( .A(n1700), .B(n183), .Q(n144) );
  NAND24 U936 ( .A(n147), .B(n146), .Q(n145) );
  CLKIN6 U937 ( .A(n1543), .Q(n146) );
  CLKIN6 U938 ( .A(n1542), .Q(n147) );
  NAND28 U939 ( .A(n148), .B(n2497), .Q(n2548) );
  INV6 U940 ( .A(n2498), .Q(n148) );
  NAND24 U941 ( .A(n1414), .B(n151), .Q(n990) );
  CLKIN6 U942 ( .A(n1413), .Q(n1414) );
  NAND22 U943 ( .A(n1406), .B(n1405), .Q(n1408) );
  NAND33 U944 ( .A(n1571), .B(n1279), .C(n1278), .Q(n1277) );
  NAND22 U945 ( .A(n1485), .B(n1585), .Q(n283) );
  NAND22 U946 ( .A(n90), .B(i_data_FMalures[25]), .Q(n1209) );
  INV6 U947 ( .A(u_alu_lt_x_11_n99), .Q(n613) );
  NAND34 U948 ( .A(n1614), .B(n1615), .C(n1369), .Q(n1616) );
  NAND26 U949 ( .A(n1594), .B(n1593), .Q(u_alu_lt_x_11_A_11_) );
  NOR24 U950 ( .A(n293), .B(n292), .Q(n1601) );
  OAI210 U951 ( .A(n217), .B(n2976), .C(n2518), .Q(n2519) );
  NAND24 U952 ( .A(u_alu_lt_x_11_n121), .B(n217), .Q(n529) );
  NAND24 U953 ( .A(n2409), .B(n2408), .Q(n1274) );
  INV6 U954 ( .A(n152), .Q(n1476) );
  NAND24 U955 ( .A(n2988), .B(n1357), .Q(n2302) );
  XOR22 U956 ( .A(n2935), .B(n2934), .Q(n2960) );
  INV6 U957 ( .A(n1354), .Q(n971) );
  INV6 U958 ( .A(n1491), .Q(n784) );
  NOR23 U959 ( .A(n343), .B(n2785), .Q(n2784) );
  NAND33 U960 ( .A(n2852), .B(n2854), .C(n2853), .Q(alu_o_data_AluRes[25]) );
  AOI212 U961 ( .A(n1829), .B(n1828), .C(n1340), .Q(n470) );
  OAI210 U962 ( .A(n173), .B(n1964), .C(n2146), .Q(n1965) );
  NOR24 U963 ( .A(n435), .B(n1532), .Q(n3087) );
  NAND23 U964 ( .A(n691), .B(n2897), .Q(n2899) );
  NAND33 U965 ( .A(n1200), .B(n1201), .C(n1369), .Q(n789) );
  NAND28 U966 ( .A(n280), .B(n279), .Q(n2926) );
  XOR22 U967 ( .A(n2594), .B(n330), .Q(n761) );
  OAI2112 U968 ( .A(n1340), .B(n1151), .C(n2047), .D(n2046), .Q(n2048) );
  NOR33 U969 ( .A(n170), .B(n1649), .C(n1650), .Q(n679) );
  NAND28 U970 ( .A(n2223), .B(n2222), .Q(n2259) );
  NAND23 U971 ( .A(n240), .B(n1247), .Q(n1246) );
  NOR24 U972 ( .A(n1475), .B(n637), .Q(n152) );
  NOR24 U973 ( .A(i_data_FMalures[13]), .B(n1214), .Q(n637) );
  NOR22 U974 ( .A(n199), .B(n480), .Q(n479) );
  NOR24 U975 ( .A(i_data_FEalures[23]), .B(n1350), .Q(n1165) );
  NAND23 U976 ( .A(n1786), .B(n1785), .Q(n2387) );
  INV8 U977 ( .A(n485), .Q(n2481) );
  INV6 U978 ( .A(n2810), .Q(n215) );
  NAND33 U979 ( .A(n1058), .B(n1057), .C(n1367), .Q(n1060) );
  NAND22 U980 ( .A(n1134), .B(n1356), .Q(n1057) );
  NOR21 U981 ( .A(n1535), .B(n250), .Q(n1536) );
  NOR21 U982 ( .A(n1463), .B(n250), .Q(n744) );
  NOR21 U983 ( .A(n1436), .B(n250), .Q(n1437) );
  NOR21 U984 ( .A(n1401), .B(n250), .Q(n1402) );
  NOR22 U985 ( .A(n1528), .B(n250), .Q(n2188) );
  NOR23 U986 ( .A(i_data_FMalures[0]), .B(n198), .Q(n389) );
  NOR24 U987 ( .A(i_data_FMalures[23]), .B(n198), .Q(n1000) );
  XOR22 U988 ( .A(n1833), .B(n472), .Q(n471) );
  NAND34 U989 ( .A(n1133), .B(n398), .C(n2528), .Q(n328) );
  NAND24 U990 ( .A(n1248), .B(n1246), .Q(n1556) );
  AOI212 U991 ( .A(n2026), .B(n234), .C(n735), .Q(n734) );
  CLKBU15 U992 ( .A(n1339), .Q(n193) );
  INV6 U993 ( .A(n1274), .Q(n1273) );
  NOR24 U994 ( .A(n1634), .B(n438), .Q(n2101) );
  NOR23 U995 ( .A(n2163), .B(n363), .Q(n361) );
  NOR24 U996 ( .A(n1424), .B(n1423), .Q(n1434) );
  IMUX20 U997 ( .A(n1776), .B(n1775), .S(compare_i_data_rs[2]), .Q(n1804) );
  NAND22 U998 ( .A(n1852), .B(compare_i_data_rs[2]), .Q(n1853) );
  INV15 U999 ( .A(n829), .Q(n1345) );
  NAND22 U1000 ( .A(n1351), .B(n1262), .Q(n1263) );
  NAND24 U1001 ( .A(n1612), .B(n1611), .Q(n1613) );
  NOR33 U1002 ( .A(n170), .B(n1610), .C(n1609), .Q(n1611) );
  AOI212 U1003 ( .A(n2569), .B(n2568), .C(n2766), .Q(n2570) );
  CLKIN4 U1004 ( .A(n329), .Q(n603) );
  OAI2112 U1005 ( .A(n1367), .B(n2982), .C(n1358), .D(n557), .Q(n556) );
  NAND24 U1006 ( .A(n552), .B(n2909), .Q(n551) );
  AOI212 U1007 ( .A(n168), .B(n553), .C(n2918), .Q(n552) );
  OAI222 U1008 ( .A(n249), .B(n2907), .C(n554), .D(n1356), .Q(n553) );
  NOR24 U1009 ( .A(n902), .B(n901), .Q(n2658) );
  NOR24 U1010 ( .A(i_data_FEalures[20]), .B(n1349), .Q(n1609) );
  AOI212 U1011 ( .A(n3002), .B(n888), .C(n887), .Q(n883) );
  INV6 U1012 ( .A(n607), .Q(n606) );
  OAI212 U1013 ( .A(n1356), .B(n2757), .C(n2730), .Q(n2738) );
  AOI212 U1014 ( .A(n2836), .B(n1360), .C(n2728), .Q(n2757) );
  NAND31 U1015 ( .A(n2821), .B(n207), .C(u_alu_pre_sum_3b[1]), .Q(n953) );
  NAND24 U1016 ( .A(DP_OP_68_131_7244_n70), .B(n1361), .Q(n2206) );
  INV8 U1017 ( .A(n1303), .Q(n1304) );
  NOR24 U1018 ( .A(n1302), .B(n1303), .Q(n1097) );
  OAI210 U1019 ( .A(u_alu_lt_x_11_n108), .B(u_alu_lt_x_11_n105), .C(
        u_alu_lt_x_11_n106), .Q(u_alu_lt_x_11_n104) );
  NAND24 U1020 ( .A(n893), .B(n1303), .Q(n894) );
  INV15 U1021 ( .A(n894), .Q(n1341) );
  NAND24 U1022 ( .A(n1149), .B(n1145), .Q(n1148) );
  NAND24 U1023 ( .A(n1147), .B(n1146), .Q(n1145) );
  INV6 U1024 ( .A(n1679), .Q(n514) );
  INV6 U1025 ( .A(n1639), .Q(n1185) );
  NAND24 U1026 ( .A(n2194), .B(n645), .Q(n644) );
  NAND28 U1027 ( .A(n820), .B(n819), .Q(n3023) );
  IMUX24 U1028 ( .A(n3098), .B(i_data_immext[0]), .S(n170), .Q(n2202) );
  AOI221 U1029 ( .A(n2754), .B(n200), .C(n192), .D(i_data_immext[8]), .Q(n1316) );
  NAND24 U1030 ( .A(n1579), .B(n1578), .Q(n1580) );
  NOR24 U1031 ( .A(n3022), .B(n1367), .Q(n726) );
  NAND24 U1032 ( .A(n1064), .B(n1063), .Q(n1065) );
  OAI222 U1033 ( .A(n71), .B(i_data_FMalures[2]), .C(n1348), .D(i_data_rt[2]), 
        .Q(n1792) );
  NOR24 U1034 ( .A(n153), .B(n154), .Q(n155) );
  NOR24 U1035 ( .A(n155), .B(n608), .Q(n2335) );
  INV3 U1036 ( .A(n2334), .Q(n153) );
  XNR22 U1037 ( .A(n2126), .B(n2125), .Q(n2127) );
  NAND28 U1038 ( .A(n2013), .B(n2012), .Q(n1172) );
  NAND28 U1039 ( .A(n1295), .B(n1296), .Q(n2013) );
  INV12 U1040 ( .A(n528), .Q(u_alu_lt_x_11_n121) );
  NAND23 U1041 ( .A(n810), .B(n1596), .Q(n528) );
  NAND24 U1042 ( .A(n1122), .B(n668), .Q(n2913) );
  NAND22 U1043 ( .A(n1123), .B(n176), .Q(n1122) );
  NOR24 U1044 ( .A(i_data_FEalures[19]), .B(n1349), .Q(n2589) );
  NOR24 U1045 ( .A(n564), .B(n563), .Q(n2952) );
  INV12 U1046 ( .A(n775), .Q(n564) );
  NAND23 U1047 ( .A(u_alu_ashr_4_A_5_), .B(n1363), .Q(n300) );
  NOR24 U1048 ( .A(n469), .B(n1827), .Q(n468) );
  BUF8 U1049 ( .A(n3049), .Q(n255) );
  NAND34 U1050 ( .A(n336), .B(n334), .C(n847), .Q(n332) );
  NAND24 U1051 ( .A(n906), .B(n1364), .Q(n774) );
  NAND33 U1052 ( .A(n2963), .B(n2965), .C(n2964), .Q(alu_o_data_AluRes[28]) );
  CLKBU15 U1053 ( .A(n344), .Q(n343) );
  INV6 U1054 ( .A(n1531), .Q(n1532) );
  INV3 U1055 ( .A(n2310), .Q(n2312) );
  NOR24 U1056 ( .A(n758), .B(n1626), .Q(n1531) );
  NAND33 U1057 ( .A(n1164), .B(n1163), .C(n1160), .Q(n156) );
  AOI212 U1058 ( .A(n3064), .B(n1356), .C(n3018), .Q(n3019) );
  INV8 U1059 ( .A(n731), .Q(n2039) );
  NOR22 U1060 ( .A(n732), .B(n2039), .Q(n733) );
  NOR23 U1061 ( .A(n823), .B(n822), .Q(n821) );
  NAND26 U1062 ( .A(n2087), .B(n1357), .Q(n897) );
  INV6 U1063 ( .A(n746), .Q(n2087) );
  NAND24 U1064 ( .A(n1077), .B(n1075), .Q(n2874) );
  INV3 U1065 ( .A(n1174), .Q(n241) );
  NOR24 U1066 ( .A(i_data_FMalures[17]), .B(n116), .Q(n2532) );
  NOR24 U1067 ( .A(n1608), .B(n1607), .Q(n1612) );
  NOR24 U1068 ( .A(n2406), .B(n163), .Q(u_alu_lt_x_11_n90) );
  NAND24 U1069 ( .A(n163), .B(n519), .Q(n641) );
  INV6 U1070 ( .A(n658), .Q(n2192) );
  NAND26 U1071 ( .A(n659), .B(n1104), .Q(n658) );
  NOR22 U1072 ( .A(n1717), .B(n2754), .Q(u_alu_lt_x_11_n9) );
  MUX26 U1073 ( .A(n3098), .B(i_data_immext[0]), .S(n170), .Q(
        u_alu_lt_x_11_B_0_) );
  NOR23 U1074 ( .A(n2627), .B(alu_i_data_B[20]), .Q(u_alu_lt_x_11_n47) );
  NAND28 U1075 ( .A(n1042), .B(n1858), .Q(n2025) );
  NAND34 U1076 ( .A(n1647), .B(n1648), .C(n1370), .Q(n1042) );
  NAND28 U1077 ( .A(n2273), .B(n2269), .Q(n1070) );
  NOR22 U1078 ( .A(n3034), .B(n2992), .Q(n3002) );
  NOR24 U1079 ( .A(n1971), .B(n2146), .Q(u_alu_lt_x_11_n99) );
  NOR23 U1080 ( .A(n1189), .B(n1193), .Q(n1192) );
  AOI211 U1081 ( .A(n1335), .B(i_data_FEalures[1]), .C(n1536), .Q(n1596) );
  NAND28 U1082 ( .A(n331), .B(n338), .Q(n1560) );
  NOR33 U1083 ( .A(n339), .B(n434), .C(n809), .Q(n338) );
  NOR23 U1084 ( .A(n1105), .B(n1202), .Q(n960) );
  NOR24 U1085 ( .A(n1361), .B(n2017), .Q(n2018) );
  NOR24 U1086 ( .A(n1860), .B(n667), .Q(n2017) );
  NOR33 U1087 ( .A(n1627), .B(n1628), .C(n617), .Q(n614) );
  NAND28 U1088 ( .A(n723), .B(n722), .Q(n3033) );
  CLKBU15 U1089 ( .A(n1347), .Q(n1218) );
  NOR23 U1090 ( .A(n248), .B(n909), .Q(n901) );
  AOI212 U1091 ( .A(n2844), .B(n2843), .C(n2842), .Q(n2845) );
  NAND23 U1092 ( .A(n2298), .B(n1358), .Q(n2299) );
  NOR24 U1093 ( .A(n634), .B(n1140), .Q(n3056) );
  NOR24 U1094 ( .A(n572), .B(n1932), .Q(n571) );
  INV6 U1095 ( .A(n573), .Q(n572) );
  NOR23 U1096 ( .A(i_data_FEalures[1]), .B(n1350), .Q(n1652) );
  AOI2110 U1097 ( .A(n857), .B(n2440), .C(n1788), .D(n1340), .Q(n1722) );
  NAND28 U1098 ( .A(n826), .B(n827), .Q(n1477) );
  INV6 U1099 ( .A(n1472), .Q(n826) );
  NOR23 U1100 ( .A(n2311), .B(n2310), .Q(n2316) );
  NOR24 U1101 ( .A(n2624), .B(n286), .Q(n2659) );
  INV6 U1102 ( .A(n287), .Q(n286) );
  AOI212 U1103 ( .A(n1839), .B(n249), .C(n1838), .Q(n2642) );
  NAND24 U1104 ( .A(n1308), .B(i_data_immext[5]), .Q(n1015) );
  NOR32 U1105 ( .A(i_data_immext[1]), .B(i_data_immext[0]), .C(
        i_data_immext[5]), .Q(n364) );
  NAND23 U1106 ( .A(n476), .B(n66), .Q(n2273) );
  NAND22 U1107 ( .A(n2601), .B(n1358), .Q(n2602) );
  XNR22 U1108 ( .A(n2104), .B(n2103), .Q(n2105) );
  NOR23 U1109 ( .A(n860), .B(n173), .Q(n1895) );
  NOR24 U1110 ( .A(u_alu_DP_OP_83J3_124_3384_n41), .B(
        u_alu_DP_OP_83J3_124_3384_n44), .Q(u_alu_DP_OP_83J3_124_3384_n101) );
  OAI210 U1111 ( .A(u_alu_DP_OP_83J3_124_3384_n44), .B(
        u_alu_DP_OP_83J3_124_3384_n50), .C(u_alu_DP_OP_83J3_124_3384_n45), .Q(
        u_alu_DP_OP_83J3_124_3384_n43) );
  OAI210 U1112 ( .A(u_alu_DP_OP_83J3_124_3384_n44), .B(
        u_alu_DP_OP_83J3_124_3384_n112), .C(u_alu_DP_OP_83J3_124_3384_n45), 
        .Q(u_alu_DP_OP_83J3_124_3384_n105) );
  NAND26 U1113 ( .A(n774), .B(n773), .Q(n2868) );
  NAND24 U1114 ( .A(n2504), .B(n1365), .Q(n2656) );
  INV6 U1115 ( .A(n1130), .Q(n2504) );
  AOI211 U1116 ( .A(n3039), .B(n3031), .C(n3033), .Q(n2933) );
  NAND24 U1117 ( .A(n1220), .B(n1221), .Q(n619) );
  XNR22 U1118 ( .A(n2861), .B(n2860), .Q(n2886) );
  NOR24 U1119 ( .A(n333), .B(n332), .Q(n331) );
  NAND24 U1120 ( .A(n335), .B(n337), .Q(n333) );
  NAND28 U1121 ( .A(n1867), .B(n1866), .Q(n1830) );
  INV12 U1122 ( .A(n466), .Q(n2193) );
  NAND24 U1123 ( .A(n743), .B(n1595), .Q(n466) );
  NOR22 U1124 ( .A(n185), .B(n2983), .Q(n2984) );
  NAND28 U1125 ( .A(n2136), .B(n2131), .Q(u_alu_lt_x_11_B_11_) );
  NAND28 U1126 ( .A(n2136), .B(n2131), .Q(n1104) );
  NAND28 U1127 ( .A(n615), .B(n614), .Q(n2136) );
  NOR33 U1128 ( .A(n1500), .B(n1499), .C(n1498), .Q(n1501) );
  XNR22 U1129 ( .A(n1318), .B(n1494), .Q(n1499) );
  NOR23 U1130 ( .A(n229), .B(n664), .Q(n2420) );
  NOR24 U1131 ( .A(n2208), .B(n2207), .Q(n2639) );
  NAND22 U1132 ( .A(n90), .B(i_data_FMalures[17]), .Q(n1133) );
  NAND28 U1133 ( .A(n1949), .B(n1948), .Q(n1952) );
  MUX21 U1134 ( .A(n1925), .B(n1928), .S(n1949), .Q(n415) );
  INV3 U1135 ( .A(n1008), .Q(n1006) );
  NOR23 U1136 ( .A(n2837), .B(n249), .Q(n2838) );
  AOI211 U1137 ( .A(n3053), .B(n163), .C(n2839), .Q(n2840) );
  NAND24 U1138 ( .A(n1239), .B(n1238), .Q(n1237) );
  OAI210 U1139 ( .A(n173), .B(n1764), .C(u_alu_lt_x_11_B_1_), .Q(n1765) );
  AOI212 U1140 ( .A(n1335), .B(i_data_FEalures[14]), .C(n1395), .Q(n1398) );
  AOI221 U1141 ( .A(n90), .B(i_data_FMalures[17]), .C(n159), .D(i_data_rs[17]), 
        .Q(n2529) );
  AOI221 U1142 ( .A(n89), .B(i_data_FMalures[30]), .C(n159), .D(i_data_rs[30]), 
        .Q(n1278) );
  NOR24 U1143 ( .A(n400), .B(n565), .Q(n327) );
  INV6 U1144 ( .A(n475), .Q(n448) );
  AOI212 U1145 ( .A(n2671), .B(n1356), .C(n177), .Q(n2672) );
  OAI210 U1146 ( .A(n173), .B(n2635), .C(alu_i_data_B[20]), .Q(n2636) );
  AOI220 U1147 ( .A(alu_i_data_B[20]), .B(n1367), .C(n2025), .D(n177), .Q(
        n1709) );
  NOR22 U1148 ( .A(u_alu_DP_OP_85J3_126_1427_n374), .B(alu_i_data_B[20]), .Q(
        u_alu_DP_OP_83J3_124_3384_n32) );
  NAND28 U1149 ( .A(n240), .B(n1313), .Q(n1312) );
  NAND24 U1150 ( .A(n490), .B(n487), .Q(n842) );
  AOI2111 U1151 ( .A(n1763), .B(n203), .C(n1762), .D(n1761), .Q(n1766) );
  NOR24 U1152 ( .A(n1162), .B(n1161), .Q(n1160) );
  NAND24 U1153 ( .A(n1154), .B(n1153), .Q(n1162) );
  XNR22 U1154 ( .A(n1277), .B(n33), .Q(n335) );
  NOR24 U1155 ( .A(n1359), .B(n2623), .Q(n2624) );
  AOI210 U1156 ( .A(n172), .B(n54), .C(n1880), .Q(n1710) );
  OAI222 U1157 ( .A(n1800), .B(n1340), .C(n1799), .D(n2494), .Q(n1801) );
  XNR22 U1158 ( .A(n1798), .B(n1832), .Q(n1799) );
  OAI212 U1159 ( .A(n2904), .B(n2976), .C(n2903), .Q(n2918) );
  XNR22 U1160 ( .A(n1563), .B(u_alu_DP_OP_83J3_124_3384_n154), .Q(n1498) );
  INV6 U1161 ( .A(n1000), .Q(n997) );
  INV6 U1162 ( .A(n585), .Q(n583) );
  NAND24 U1163 ( .A(n1732), .B(n1302), .Q(n1056) );
  NAND26 U1164 ( .A(n2916), .B(n172), .Q(n2147) );
  NAND26 U1165 ( .A(n1229), .B(n1228), .Q(n2916) );
  XNR22 U1166 ( .A(n2665), .B(n2654), .Q(n2662) );
  NAND24 U1167 ( .A(n727), .B(n2949), .Q(n2987) );
  INV6 U1168 ( .A(n1869), .Q(n1294) );
  INV12 U1169 ( .A(n1732), .Q(n972) );
  NAND28 U1170 ( .A(n1502), .B(n1501), .Q(n1034) );
  NAND34 U1171 ( .A(n375), .B(n373), .C(n372), .Q(n2967) );
  NAND26 U1172 ( .A(n636), .B(n2912), .Q(n2982) );
  NAND24 U1173 ( .A(n1386), .B(n1387), .Q(n812) );
  NAND33 U1174 ( .A(n1590), .B(n1587), .C(n1586), .Q(n1483) );
  AOI222 U1175 ( .A(n89), .B(i_data_FMalures[6]), .C(n1334), .D(
        i_data_FEalures[6]), .Q(n657) );
  NOR24 U1176 ( .A(n2590), .B(n2588), .Q(n1615) );
  NOR24 U1177 ( .A(i_data_FMalures[18]), .B(n116), .Q(n1619) );
  NAND24 U1178 ( .A(n939), .B(n1540), .Q(n1541) );
  AOI212 U1179 ( .A(n78), .B(n1356), .C(n2232), .Q(n2250) );
  INV3 U1180 ( .A(n1839), .Q(n1815) );
  NAND28 U1181 ( .A(n2538), .B(n1353), .Q(u_alu_ashr_4_A_17_) );
  NAND26 U1182 ( .A(n1622), .B(n2535), .Q(n2538) );
  NAND24 U1183 ( .A(n1209), .B(n1210), .Q(n1211) );
  NOR24 U1184 ( .A(n850), .B(n1371), .Q(n849) );
  NAND24 U1185 ( .A(n852), .B(n851), .Q(n850) );
  NAND23 U1186 ( .A(n2978), .B(n1356), .Q(n498) );
  AOI212 U1187 ( .A(n2424), .B(n2423), .C(n2422), .Q(n2425) );
  NOR23 U1188 ( .A(n567), .B(n2368), .Q(n2422) );
  NOR24 U1189 ( .A(n786), .B(n785), .Q(n1605) );
  NOR23 U1190 ( .A(i_data_FEalures[24]), .B(n1350), .Q(n786) );
  NAND26 U1191 ( .A(n2865), .B(n247), .Q(n775) );
  NAND24 U1192 ( .A(n898), .B(n897), .Q(n2865) );
  XNR22 U1193 ( .A(n1856), .B(n1947), .Q(n1875) );
  NAND26 U1194 ( .A(n1855), .B(n2042), .Q(n1947) );
  NOR23 U1195 ( .A(n2790), .B(n875), .Q(n2791) );
  NAND28 U1196 ( .A(n386), .B(n1014), .Q(n453) );
  NAND26 U1197 ( .A(n2102), .B(n2101), .Q(n2409) );
  NOR24 U1198 ( .A(i_data_FMalures[16]), .B(n1214), .Q(n2805) );
  NAND26 U1199 ( .A(n694), .B(n693), .Q(n692) );
  IMUX23 U1200 ( .A(n2105), .B(n2106), .S(n1343), .Q(n683) );
  CLKBU15 U1201 ( .A(n1546), .Q(n1334) );
  NOR24 U1202 ( .A(n1212), .B(n1211), .Q(n324) );
  NOR24 U1203 ( .A(i_data_FEalures[21]), .B(n1350), .Q(n1493) );
  AOI221 U1204 ( .A(u_alu_ashr_4_A_17_), .B(n2830), .C(n2829), .D(n166), .Q(
        n773) );
  NOR23 U1205 ( .A(i_data_FMalures[1]), .B(n1214), .Q(n1653) );
  NAND28 U1206 ( .A(n1602), .B(n1353), .Q(n1337) );
  NOR24 U1207 ( .A(n779), .B(n781), .Q(n2981) );
  NOR24 U1208 ( .A(n2184), .B(n2183), .Q(n2347) );
  NOR33 U1209 ( .A(n2182), .B(n213), .C(n2181), .Q(n2183) );
  NAND34 U1210 ( .A(n1642), .B(n230), .C(n1219), .Q(n1968) );
  NOR22 U1211 ( .A(u_alu_DP_OP_85J3_126_1427_n379), .B(u_alu_lt_x_11_B_25_), 
        .Q(u_alu_DP_OP_84J3_125_2615_n47) );
  INV12 U1212 ( .A(n2550), .Q(n2806) );
  NAND22 U1213 ( .A(n805), .B(n2550), .Q(n804) );
  NAND28 U1214 ( .A(n1689), .B(n1307), .Q(u_alu_lt_x_11_B_25_) );
  NOR24 U1215 ( .A(n390), .B(n389), .Q(n1087) );
  NAND34 U1216 ( .A(n762), .B(n761), .C(n759), .Q(n1478) );
  NOR24 U1217 ( .A(n1632), .B(n1633), .Q(n2102) );
  NOR33 U1218 ( .A(n1632), .B(n1634), .C(n548), .Q(n3089) );
  NOR23 U1219 ( .A(i_data_FMalures[10]), .B(n1214), .Q(n1632) );
  NOR23 U1220 ( .A(n2999), .B(n3000), .Q(n887) );
  NOR24 U1221 ( .A(i_data_FMalures[20]), .B(n1214), .Q(n1608) );
  NAND26 U1222 ( .A(n2252), .B(n229), .Q(u_alu_lt_x_11_n77) );
  INV15 U1223 ( .A(n1341), .Q(n187) );
  INV6 U1224 ( .A(n1090), .Q(n1089) );
  NOR24 U1225 ( .A(n248), .B(n2656), .Q(n2657) );
  OAI210 U1226 ( .A(n173), .B(n2521), .C(u_alu_ashr_4_A_17_), .Q(n2522) );
  OAI210 U1227 ( .A(u_alu_ashr_4_A_17_), .B(n187), .C(n278), .Q(n2520) );
  NOR23 U1228 ( .A(n1361), .B(n3012), .Q(n3013) );
  NOR24 U1229 ( .A(n1868), .B(n579), .Q(n2459) );
  NAND28 U1230 ( .A(n1070), .B(n1361), .Q(n671) );
  OAI210 U1231 ( .A(n173), .B(n2043), .C(n2204), .Q(n2047) );
  OAI210 U1232 ( .A(n187), .B(n2204), .C(n278), .Q(n2045) );
  NOR23 U1233 ( .A(n2531), .B(n2530), .Q(n2535) );
  NAND22 U1234 ( .A(n2323), .B(n1134), .Q(n1058) );
  CLKIN4 U1235 ( .A(n2323), .Q(n1093) );
  NOR33 U1236 ( .A(n1479), .B(n1480), .C(n1478), .Q(n1502) );
  NOR22 U1237 ( .A(i_data_fbmemout[30]), .B(n1324), .Q(n1542) );
  NOR22 U1238 ( .A(i_data_fbmemout[12]), .B(n1324), .Q(n758) );
  NOR22 U1239 ( .A(i_data_fbmemout[29]), .B(n1324), .Q(n507) );
  NOR22 U1240 ( .A(i_data_fbmemout[26]), .B(n1324), .Q(n1508) );
  CLKIN4 U1241 ( .A(i_con_Efamux[0]), .Q(n1018) );
  NAND34 U1242 ( .A(n1434), .B(n1006), .C(n1240), .Q(n697) );
  NAND23 U1243 ( .A(i_data_immext[1]), .B(i_data_immext[3]), .Q(n1016) );
  NAND28 U1244 ( .A(n2778), .B(n1307), .Q(u_alu_DP_OP_83J3_124_3384_n152) );
  NOR24 U1245 ( .A(n1366), .B(n2329), .Q(n2725) );
  NOR24 U1246 ( .A(n249), .B(n2988), .Q(n1140) );
  NAND26 U1247 ( .A(n305), .B(n2217), .Q(n2988) );
  CLKBU15 U1248 ( .A(n1222), .Q(n844) );
  NOR24 U1249 ( .A(n2402), .B(n502), .Q(n2279) );
  NAND34 U1250 ( .A(n2034), .B(n2033), .C(n2032), .Q(n2402) );
  NAND33 U1251 ( .A(n2397), .B(n2395), .C(n2396), .Q(n2398) );
  XNR22 U1252 ( .A(n1483), .B(n1484), .Q(n1500) );
  OAI210 U1253 ( .A(n173), .B(n1737), .C(u_alu_lt_x_11_B_0_), .Q(n1738) );
  NAND33 U1254 ( .A(u_alu_lt_x_11_B_0_), .B(n249), .C(n2830), .Q(n2074) );
  NAND23 U1255 ( .A(n1852), .B(u_alu_lt_x_11_n122), .Q(n2458) );
  OAI312 U1256 ( .A(n1794), .B(n1793), .C(n1792), .D(n1791), .Q(n1852) );
  AOI222 U1257 ( .A(n382), .B(n2672), .C(n2670), .D(n243), .Q(n378) );
  NAND24 U1258 ( .A(n384), .B(n1172), .Q(n1177) );
  NAND28 U1259 ( .A(n2013), .B(n2012), .Q(n2361) );
  NOR42 U1260 ( .A(n2318), .B(n2316), .C(n2317), .D(n2315), .Q(n2338) );
  NOR42 U1261 ( .A(n2423), .B(n2314), .C(n2313), .D(n2312), .Q(n2315) );
  XOR22 U1262 ( .A(u_alu_pre_sum_4a[0]), .B(n1176), .Q(n1147) );
  NOR33 U1263 ( .A(n895), .B(n928), .C(n896), .Q(n2863) );
  OAI212 U1264 ( .A(n2834), .B(n2870), .C(n2770), .Q(n2771) );
  NOR24 U1265 ( .A(n2768), .B(n2767), .Q(n2870) );
  OAI210 U1266 ( .A(n173), .B(n2769), .C(n43), .Q(n2770) );
  NAND24 U1267 ( .A(n1577), .B(n1426), .Q(n1167) );
  NOR24 U1268 ( .A(n1821), .B(n1037), .Q(n1038) );
  OAI212 U1269 ( .A(n1477), .B(n1476), .C(n229), .Q(n484) );
  NAND34 U1270 ( .A(n1377), .B(n1378), .C(n1376), .Q(compare_i_data_rs[2]) );
  AOI212 U1271 ( .A(n1335), .B(i_data_FEalures[2]), .C(n1375), .Q(n1378) );
  CLKIN4 U1272 ( .A(i_data_immext[1]), .Q(n980) );
  NAND28 U1273 ( .A(n994), .B(n1353), .Q(u_alu_ashr_4_A_16_) );
  NOR22 U1274 ( .A(n1865), .B(u_alu_lt_x_11_A_0_), .Q(n1256) );
  NOR24 U1275 ( .A(n1364), .B(n571), .Q(n2301) );
  CLKIN15 U1276 ( .A(n157), .Q(n158) );
  CLKIN15 U1277 ( .A(n157), .Q(n159) );
  NAND28 U1278 ( .A(n300), .B(n299), .Q(n2511) );
  AOI212 U1279 ( .A(n2884), .B(n2883), .C(n2882), .Q(n2885) );
  AOI222 U1280 ( .A(n2295), .B(n175), .C(n248), .D(u_alu_lt_x_11_B_25_), .Q(
        n2983) );
  INV3 U1281 ( .A(n2384), .Q(n1851) );
  NOR24 U1282 ( .A(n2631), .B(n701), .Q(n2812) );
  NOR24 U1283 ( .A(n605), .B(n2630), .Q(n701) );
  NAND28 U1284 ( .A(n433), .B(n432), .Q(n2594) );
  NAND28 U1285 ( .A(n1643), .B(n1997), .Q(u_alu_ashr_4_A_6_) );
  NOR24 U1286 ( .A(u_alu_lt_x_11_A_11_), .B(n2135), .Q(n2137) );
  IMUX24 U1287 ( .A(n2688), .B(n2296), .S(n245), .Q(n2555) );
  OAI210 U1288 ( .A(n173), .B(n2352), .C(n1299), .Q(n2353) );
  OAI210 U1289 ( .A(n1299), .B(n187), .C(n278), .Q(n2325) );
  NAND24 U1290 ( .A(n1299), .B(n175), .Q(n718) );
  AOI222 U1291 ( .A(u_alu_lt_x_11_B_24_), .B(n248), .C(n2947), .D(n1361), .Q(
        n2950) );
  NAND24 U1292 ( .A(n2947), .B(n172), .Q(n2655) );
  NAND28 U1293 ( .A(n2926), .B(n1353), .Q(n2947) );
  NOR23 U1294 ( .A(i_data_fbmemout[17]), .B(n246), .Q(n2533) );
  AOI212 U1295 ( .A(n632), .B(n2468), .C(n2476), .Q(n631) );
  NAND26 U1296 ( .A(n509), .B(n1606), .Q(n1707) );
  NAND28 U1297 ( .A(n1275), .B(n1353), .Q(n2754) );
  NOR23 U1298 ( .A(i_data_FMalures[7]), .B(n116), .Q(n2001) );
  CLKIN4 U1299 ( .A(n2950), .Q(n728) );
  INV15 U1300 ( .A(n162), .Q(n163) );
  NAND24 U1301 ( .A(n191), .B(n787), .Q(n3032) );
  OAI222 U1302 ( .A(n1760), .B(n2494), .C(n1340), .D(n1759), .Q(n1761) );
  AOI222 U1303 ( .A(n989), .B(n988), .C(n986), .D(n179), .Q(n985) );
  XOR22 U1304 ( .A(n2168), .B(n987), .Q(n986) );
  NOR24 U1305 ( .A(i_data_FEalures[18]), .B(n1349), .Q(n1618) );
  OAI210 U1306 ( .A(n173), .B(n2572), .C(n688), .Q(n2573) );
  AOI222 U1307 ( .A(n2252), .B(n175), .C(n248), .D(n163), .Q(n2676) );
  NAND28 U1308 ( .A(n672), .B(n671), .Q(n2694) );
  NAND28 U1309 ( .A(n1888), .B(n1887), .Q(u_alu_ashr_4_A_5_) );
  NAND24 U1310 ( .A(n1646), .B(n1645), .Q(n1888) );
  OAI212 U1311 ( .A(n187), .B(n1336), .C(n180), .Q(n2877) );
  CLKBU15 U1312 ( .A(n1354), .Q(n180) );
  XNR22 U1313 ( .A(u_alu_lt_x_11_A_31_), .B(compare_i_data_rt_31_), .Q(n847)
         );
  INV3 U1314 ( .A(n1647), .Q(n1859) );
  NAND24 U1315 ( .A(n782), .B(n1369), .Q(n2383) );
  NAND24 U1316 ( .A(n1083), .B(n1087), .Q(n782) );
  NOR23 U1317 ( .A(i_data_FMalures[26]), .B(n1214), .Q(n292) );
  AOI2112 U1318 ( .A(n417), .B(n1928), .C(n1340), .D(n1929), .Q(n416) );
  NOR33 U1319 ( .A(n1928), .B(n1927), .C(n1926), .Q(n1929) );
  NOR22 U1320 ( .A(n218), .B(n163), .Q(n2100) );
  INV6 U1321 ( .A(n2811), .Q(n1221) );
  NAND24 U1322 ( .A(n2795), .B(n2796), .Q(n2811) );
  NOR24 U1323 ( .A(n1445), .B(n1446), .Q(n1648) );
  NOR22 U1324 ( .A(i_data_FMalures[4]), .B(n116), .Q(n1446) );
  NOR24 U1325 ( .A(n803), .B(n2630), .Q(n2809) );
  NOR24 U1326 ( .A(n2594), .B(n2593), .Q(n2630) );
  XOR22 U1327 ( .A(n52), .B(n911), .Q(n1068) );
  NAND34 U1328 ( .A(n998), .B(n1001), .C(n151), .Q(n1196) );
  NOR24 U1329 ( .A(n1000), .B(n999), .Q(n998) );
  NOR24 U1330 ( .A(n2096), .B(n2396), .Q(n2181) );
  OAI212 U1331 ( .A(n166), .B(n3016), .C(n3015), .Q(n3064) );
  INV6 U1332 ( .A(u_alu_DP_OP_83J3_124_3384_n64), .Q(n164) );
  OAI212 U1333 ( .A(n165), .B(u_alu_DP_OP_83J3_124_3384_n18), .C(
        u_alu_DP_OP_83J3_124_3384_n19), .Q(n601) );
  NAND24 U1334 ( .A(n2722), .B(n2723), .Q(n2844) );
  AOI312 U1335 ( .A(n1367), .B(n249), .C(n2721), .D(n2720), .Q(n2722) );
  XOR20 U1336 ( .A(u_alu_DP_OP_83J3_124_3384_n5), .B(n165), .Q(
        u_alu_pre_sum_3b[4]) );
  NOR22 U1337 ( .A(n2470), .B(n2284), .Q(n2082) );
  INV6 U1338 ( .A(n947), .Q(n2714) );
  OAI221 U1339 ( .A(n2119), .B(n1357), .C(n2156), .D(n1356), .Q(n2120) );
  INV3 U1340 ( .A(n3002), .Q(n2999) );
  INV3 U1341 ( .A(n2359), .Q(n204) );
  NOR21 U1342 ( .A(n172), .B(n3066), .Q(n885) );
  NAND22 U1343 ( .A(n2434), .B(n1363), .Q(n2171) );
  NAND23 U1344 ( .A(n900), .B(n899), .Q(n970) );
  INV3 U1345 ( .A(n2196), .Q(n209) );
  INV3 U1346 ( .A(u_alu_DP_OP_84J3_125_2615_n30), .Q(
        u_alu_DP_OP_84J3_125_2615_n81) );
  INV3 U1347 ( .A(n1056), .Q(n1714) );
  NAND22 U1348 ( .A(u_alu_lt_x_11_B_28_), .B(n1524), .Q(
        u_alu_DP_OP_84J3_125_2615_n31) );
  INV2 U1349 ( .A(u_alu_DP_OP_83J3_124_3384_n89), .Q(
        u_alu_DP_OP_83J3_124_3384_n25) );
  INV3 U1350 ( .A(n2475), .Q(n2474) );
  INV2 U1351 ( .A(n1914), .Q(n1768) );
  NOR22 U1352 ( .A(n196), .B(n192), .Q(n621) );
  NOR22 U1353 ( .A(u_alu_DP_OP_83J3_124_3384_n29), .B(
        u_alu_DP_OP_83J3_124_3384_n32), .Q(u_alu_DP_OP_83J3_124_3384_n89) );
  INV3 U1354 ( .A(u_alu_DP_OP_84J3_125_2615_n22), .Q(
        u_alu_DP_OP_84J3_125_2615_n77) );
  NAND22 U1355 ( .A(u_alu_ashr_4_A_6_), .B(n172), .Q(n1702) );
  CLKIN6 U1356 ( .A(n2387), .Q(n1849) );
  NOR22 U1357 ( .A(n576), .B(n2005), .Q(n2464) );
  NOR21 U1358 ( .A(n221), .B(n2030), .Q(n2031) );
  NAND22 U1359 ( .A(n2259), .B(n172), .Q(n1910) );
  INV6 U1360 ( .A(n1567), .Q(n1416) );
  INV2 U1361 ( .A(n747), .Q(n3075) );
  INV3 U1362 ( .A(n1052), .Q(n1276) );
  NAND22 U1363 ( .A(n2190), .B(n1592), .Q(n485) );
  NAND24 U1364 ( .A(n574), .B(n2064), .Q(n2065) );
  INV6 U1365 ( .A(n1580), .Q(n1581) );
  NOR23 U1366 ( .A(n170), .B(n2063), .Q(n574) );
  CLKIN6 U1367 ( .A(n2000), .Q(n230) );
  NAND22 U1368 ( .A(n1321), .B(i_data_famemout[26]), .Q(n1505) );
  INV3 U1369 ( .A(n401), .Q(n400) );
  INV3 U1370 ( .A(n1297), .Q(n778) );
  CLKIN3 U1371 ( .A(n1640), .Q(n1999) );
  INV3 U1372 ( .A(n2188), .Q(n457) );
  INV3 U1373 ( .A(n2862), .Q(n2864) );
  NAND22 U1374 ( .A(i_data_immext[15]), .B(n170), .Q(n2340) );
  NAND23 U1375 ( .A(n170), .B(n1359), .Q(n2003) );
  INV2 U1376 ( .A(n1674), .Q(n946) );
  INV3 U1377 ( .A(n2330), .Q(n2432) );
  NOR23 U1378 ( .A(n1680), .B(n979), .Q(n1674) );
  INV2 U1379 ( .A(n185), .Q(n176) );
  NOR21 U1380 ( .A(n1309), .B(n1680), .Q(n1004) );
  INV12 U1381 ( .A(n1365), .Q(n166) );
  INV8 U1382 ( .A(i_data_immext[9]), .Q(n1365) );
  AOI211 U1383 ( .A(n2883), .B(n2049), .C(n2048), .Q(n2050) );
  NAND33 U1384 ( .A(n1908), .B(n1907), .C(n1906), .Q(alu_o_data_AluRes[5]) );
  AOI211 U1385 ( .A(n1813), .B(n1812), .C(n1811), .Q(n1837) );
  NAND24 U1386 ( .A(n2821), .B(n207), .Q(n947) );
  INV2 U1387 ( .A(n2939), .Q(n554) );
  AOI211 U1388 ( .A(n1819), .B(n2883), .C(n1818), .Q(n1836) );
  NOR21 U1389 ( .A(u_alu_lt_x_11_n49), .B(u_alu_lt_x_11_n35), .Q(
        u_alu_lt_x_11_n33) );
  INV12 U1390 ( .A(n3006), .Q(n168) );
  INV1 U1391 ( .A(n2288), .Q(n2282) );
  NAND21 U1392 ( .A(n2643), .B(n2644), .Q(n2646) );
  INV3 U1393 ( .A(n2462), .Q(n188) );
  INV3 U1394 ( .A(n2467), .Q(n2479) );
  INV2 U1395 ( .A(u_alu_DP_OP_83J3_124_3384_n90), .Q(
        u_alu_DP_OP_83J3_124_3384_n26) );
  INV3 U1396 ( .A(n2464), .Q(n2011) );
  INV3 U1397 ( .A(n2142), .Q(n212) );
  INV6 U1398 ( .A(u_alu_lt_x_11_n87), .Q(n2161) );
  INV3 U1399 ( .A(n2481), .Q(n486) );
  INV3 U1400 ( .A(n1280), .Q(n444) );
  NAND21 U1401 ( .A(u_alu_ashr_4_A_16_), .B(n2808), .Q(u_alu_lt_x_11_n62) );
  INV3 U1402 ( .A(n2065), .Q(n1186) );
  INV2 U1403 ( .A(n1566), .Q(n3082) );
  INV3 U1404 ( .A(n231), .Q(n620) );
  NAND26 U1405 ( .A(n1605), .B(n1369), .Q(n1188) );
  NOR22 U1406 ( .A(n455), .B(n1591), .Q(n2190) );
  INV3 U1407 ( .A(n1048), .Q(n232) );
  NOR22 U1408 ( .A(n958), .B(n957), .Q(n959) );
  INV3 U1409 ( .A(n1078), .Q(n510) );
  NAND21 U1410 ( .A(n242), .B(n172), .Q(n258) );
  INV3 U1411 ( .A(n2544), .Q(n1069) );
  INV3 U1412 ( .A(n1858), .Q(n1860) );
  NAND22 U1413 ( .A(i_data_immext[12]), .B(n170), .Q(n2178) );
  NAND22 U1414 ( .A(i_data_immext[13]), .B(n170), .Q(n2222) );
  INV3 U1415 ( .A(n1529), .Q(n1591) );
  INV3 U1416 ( .A(n177), .Q(n171) );
  INV12 U1417 ( .A(n248), .Q(n175) );
  INV12 U1418 ( .A(n1366), .Q(n177) );
  INV12 U1419 ( .A(n1367), .Q(n172) );
  INV3 U1420 ( .A(i_con_Ealuop[4]), .Q(n1662) );
  INV1 U1421 ( .A(i_data_FMalures[28]), .Q(n942) );
  INV2 U1422 ( .A(n2371), .Q(n2373) );
  NOR21 U1423 ( .A(n2494), .B(n2288), .Q(n2303) );
  NOR22 U1424 ( .A(n1716), .B(n1056), .Q(n2823) );
  NOR22 U1425 ( .A(n2479), .B(n2480), .Q(n2358) );
  NOR21 U1426 ( .A(u_alu_DP_OP_85J3_126_1427_n368), .B(n444), .Q(
        u_alu_DP_OP_84J3_125_2615_n14) );
  INV2 U1427 ( .A(n356), .Q(n351) );
  NOR21 U1428 ( .A(n2100), .B(n212), .Q(n2068) );
  INV6 U1429 ( .A(u_alu_lt_x_11_B_0_), .Q(n2440) );
  INV2 U1430 ( .A(n2420), .Q(n662) );
  NOR22 U1431 ( .A(n175), .B(n914), .Q(n356) );
  NOR22 U1432 ( .A(n223), .B(n1823), .Q(n1854) );
  INV2 U1433 ( .A(n2419), .Q(n2309) );
  INV3 U1434 ( .A(n1104), .Q(n2180) );
  NAND23 U1435 ( .A(n2204), .B(n316), .Q(n2081) );
  INV3 U1436 ( .A(n1131), .Q(n2553) );
  INV6 U1437 ( .A(alu_i_data_B[20]), .Q(n2644) );
  NOR23 U1438 ( .A(n256), .B(n2252), .Q(n2417) );
  INV2 U1439 ( .A(n1568), .Q(n3074) );
  INV6 U1440 ( .A(n1188), .Q(n509) );
  INV3 U1441 ( .A(n789), .Q(n280) );
  INV6 U1442 ( .A(n566), .Q(n567) );
  INV3 U1443 ( .A(n1215), .Q(n1650) );
  INV3 U1444 ( .A(n1465), .Q(n1266) );
  INV3 U1445 ( .A(n1620), .Q(n238) );
  NAND22 U1446 ( .A(n1587), .B(n1586), .Q(n1588) );
  INV2 U1447 ( .A(n1617), .Q(n588) );
  NAND22 U1448 ( .A(i_data_immext[14]), .B(n170), .Q(n2269) );
  INV3 U1449 ( .A(n175), .Q(n169) );
  INV3 U1450 ( .A(n1370), .Q(n1368) );
  INV6 U1451 ( .A(n1369), .Q(n199) );
  INV3 U1452 ( .A(n725), .Q(n724) );
  NAND22 U1453 ( .A(n2583), .B(n2584), .Q(n725) );
  NOR22 U1454 ( .A(n2815), .B(n597), .Q(n2816) );
  NAND22 U1455 ( .A(n918), .B(n178), .Q(n969) );
  NAND22 U1456 ( .A(n3020), .B(n167), .Q(n879) );
  NAND23 U1457 ( .A(n1093), .B(n1356), .Q(n1091) );
  INV6 U1458 ( .A(n3033), .Q(n3037) );
  NOR23 U1459 ( .A(n1358), .B(n2906), .Q(n1076) );
  INV3 U1460 ( .A(u_alu_DP_OP_84J3_125_2615_n17), .Q(n206) );
  INV3 U1461 ( .A(n3052), .Q(n798) );
  INV3 U1462 ( .A(n2313), .Q(n2311) );
  INV12 U1463 ( .A(n2494), .Q(n179) );
  NAND22 U1464 ( .A(n168), .B(n1356), .Q(n538) );
  INV3 U1465 ( .A(n2173), .Q(n2174) );
  INV2 U1466 ( .A(n2435), .Q(n837) );
  NAND26 U1467 ( .A(n464), .B(n2439), .Q(n2494) );
  INV3 U1468 ( .A(n2477), .Q(n632) );
  OAI211 U1469 ( .A(n1701), .B(n1939), .C(n185), .Q(n1706) );
  NOR23 U1470 ( .A(n1849), .B(n1848), .Q(n2038) );
  NAND22 U1471 ( .A(n3014), .B(n166), .Q(n3015) );
  OAI222 U1472 ( .A(n1699), .B(n1364), .C(n166), .D(n1698), .Q(n440) );
  INV3 U1473 ( .A(n1954), .Q(n1921) );
  NOR22 U1474 ( .A(n1056), .B(n465), .Q(n464) );
  INV3 U1475 ( .A(u_alu_DP_OP_84J3_125_2615_n14), .Q(
        u_alu_DP_OP_84J3_125_2615_n108) );
  INV3 U1476 ( .A(n2020), .Q(n2021) );
  INV6 U1477 ( .A(n2809), .Q(n2650) );
  NAND22 U1478 ( .A(u_alu_lt_x_11_n46), .B(u_alu_lt_x_11_n47), .Q(n2742) );
  BUF15 U1479 ( .A(n1341), .Q(n174) );
  INV6 U1480 ( .A(n1924), .Q(n189) );
  INV3 U1481 ( .A(n903), .Q(n902) );
  NAND24 U1482 ( .A(n1281), .B(n975), .Q(n1561) );
  NAND23 U1483 ( .A(n1070), .B(n233), .Q(n2466) );
  NAND22 U1484 ( .A(n1243), .B(n1242), .Q(n1241) );
  OAI212 U1485 ( .A(n170), .B(n368), .C(n183), .Q(n2781) );
  INV2 U1486 ( .A(n1421), .Q(n3078) );
  INV3 U1487 ( .A(n2411), .Q(n2195) );
  INV2 U1488 ( .A(n1797), .Q(n1756) );
  INV2 U1489 ( .A(n2995), .Q(n1055) );
  NAND22 U1490 ( .A(n1049), .B(n408), .Q(n1421) );
  CLKIN6 U1491 ( .A(n735), .Q(n216) );
  NAND23 U1492 ( .A(n221), .B(n2030), .Q(n2041) );
  NAND22 U1493 ( .A(n1830), .B(n223), .Q(n2461) );
  INV6 U1494 ( .A(n2929), .Q(n194) );
  NAND26 U1495 ( .A(n1707), .B(n1353), .Q(n1193) );
  INV2 U1496 ( .A(n2417), .Q(n501) );
  NAND23 U1497 ( .A(n219), .B(n620), .Q(n2097) );
  NOR22 U1498 ( .A(n977), .B(n976), .Q(n975) );
  INV2 U1499 ( .A(n567), .Q(n568) );
  INV3 U1500 ( .A(n2027), .Q(n1643) );
  NAND22 U1501 ( .A(n1639), .B(n2062), .Q(n1259) );
  NAND22 U1502 ( .A(n1323), .B(n1420), .Q(n409) );
  NAND23 U1503 ( .A(n1081), .B(n1676), .Q(n1079) );
  NAND22 U1504 ( .A(n587), .B(n588), .Q(n586) );
  INV3 U1505 ( .A(n234), .Q(n1314) );
  INV3 U1506 ( .A(n1471), .Q(n827) );
  INV2 U1507 ( .A(n1724), .Q(n1728) );
  INV3 U1508 ( .A(n2537), .Q(n930) );
  INV6 U1509 ( .A(n1524), .Q(n228) );
  NOR22 U1510 ( .A(n1266), .B(n329), .Q(n2545) );
  INV3 U1511 ( .A(n1373), .Q(n848) );
  NOR23 U1512 ( .A(n1516), .B(n1515), .Q(n1597) );
  INV2 U1513 ( .A(n2269), .Q(n2280) );
  INV3 U1514 ( .A(n342), .Q(n455) );
  INV1 U1515 ( .A(n2800), .Q(n2802) );
  NAND22 U1516 ( .A(n1080), .B(n1727), .Q(n1078) );
  INV3 U1517 ( .A(n1120), .Q(n1637) );
  INV3 U1518 ( .A(n2222), .Q(n235) );
  INV3 U1519 ( .A(n1657), .Q(n1658) );
  INV3 U1520 ( .A(n1402), .Q(n1014) );
  NOR22 U1521 ( .A(n1674), .B(n1673), .Q(n1676) );
  INV3 U1522 ( .A(n1673), .Q(n1669) );
  NAND22 U1523 ( .A(n200), .B(n185), .Q(n273) );
  NAND22 U1524 ( .A(n908), .B(n170), .Q(n1887) );
  NAND21 U1525 ( .A(n1361), .B(n201), .Q(n907) );
  INV3 U1526 ( .A(n1358), .Q(n201) );
  INV1 U1527 ( .A(i_data_FMalures[5]), .Q(n1552) );
  INV3 U1528 ( .A(i_con_Ealuop[2]), .Q(n1681) );
  BUF12 U1529 ( .A(i_data_immext[10]), .Q(n1367) );
  INV2 U1530 ( .A(i_data_rt[10]), .Q(n1629) );
  INV1 U1531 ( .A(i_data_FMalures[3]), .Q(n1216) );
  INV3 U1532 ( .A(i_con_Malupc8), .Q(n3103) );
  NAND33 U1533 ( .A(n2889), .B(n2891), .C(n2890), .Q(alu_o_data_AluRes[26]) );
  NAND33 U1534 ( .A(n2268), .B(n2267), .C(n2266), .Q(alu_o_data_AluRes[13]) );
  NAND33 U1535 ( .A(n2923), .B(n2925), .C(n2924), .Q(alu_o_data_AluRes[27]) );
  NAND32 U1536 ( .A(n2378), .B(n2377), .C(n2376), .Q(n2379) );
  NOR22 U1537 ( .A(n2816), .B(n1285), .Q(n1284) );
  NOR22 U1538 ( .A(n2582), .B(n2581), .Q(n2585) );
  NAND22 U1539 ( .A(n839), .B(n202), .Q(n838) );
  OAI212 U1540 ( .A(n1358), .B(n2870), .C(n2869), .Q(n2884) );
  NAND22 U1541 ( .A(n1172), .B(n2236), .Q(n2237) );
  NAND22 U1542 ( .A(n1106), .B(n676), .Q(n675) );
  OAI222 U1543 ( .A(n2119), .B(n1356), .C(n1357), .D(n2061), .Q(n714) );
  INV3 U1544 ( .A(n3021), .Q(n1096) );
  INV15 U1545 ( .A(n1222), .Q(n178) );
  NOR24 U1546 ( .A(n2372), .B(n2374), .Q(n1213) );
  OAI212 U1547 ( .A(n1360), .B(n2777), .C(n2883), .Q(n2700) );
  OAI212 U1548 ( .A(n1356), .B(n2641), .C(n2640), .Q(n673) );
  NAND22 U1549 ( .A(n2147), .B(n1359), .Q(n2148) );
  NAND22 U1550 ( .A(n3023), .B(n247), .Q(n892) );
  INV3 U1551 ( .A(n2574), .Q(n2575) );
  INV3 U1552 ( .A(n2333), .Q(n611) );
  OAI212 U1553 ( .A(n177), .B(n68), .C(n1360), .Q(n635) );
  AOI211 U1554 ( .A(u_alu_DP_OP_84J3_125_2615_n92), .B(n206), .C(n405), .Q(
        n404) );
  NAND22 U1555 ( .A(n403), .B(n206), .Q(n402) );
  INV3 U1556 ( .A(n525), .Q(n524) );
  INV3 U1557 ( .A(n538), .Q(n537) );
  NOR21 U1558 ( .A(n862), .B(n173), .Q(n2200) );
  INV3 U1559 ( .A(n873), .Q(n872) );
  NOR23 U1560 ( .A(n425), .B(u_alu_DP_OP_83J3_124_3384_n76), .Q(n424) );
  INV2 U1561 ( .A(u_alu_DP_OP_84J3_125_2615_n18), .Q(n405) );
  NAND22 U1562 ( .A(n837), .B(n201), .Q(n836) );
  AOI212 U1563 ( .A(n2719), .B(n2718), .C(n2766), .Q(n2720) );
  NAND22 U1564 ( .A(n1845), .B(n201), .Q(n443) );
  NAND22 U1565 ( .A(n2763), .B(n1356), .Q(n2022) );
  OAI212 U1566 ( .A(n910), .B(n187), .C(n278), .Q(n2109) );
  INV3 U1567 ( .A(n2708), .Q(n2705) );
  INV6 U1568 ( .A(n971), .Q(n973) );
  INV2 U1569 ( .A(n967), .Q(n403) );
  INV2 U1570 ( .A(n2306), .Q(n2314) );
  INV6 U1571 ( .A(n3032), .Q(n3031) );
  INV3 U1572 ( .A(n2596), .Q(n2546) );
  INV3 U1573 ( .A(n2344), .Q(n2349) );
  INV2 U1574 ( .A(n2898), .Q(n916) );
  INV3 U1575 ( .A(n2029), .Q(n1922) );
  NAND22 U1576 ( .A(n291), .B(n2041), .Q(n996) );
  NAND22 U1577 ( .A(n702), .B(n2812), .Q(n1220) );
  INV2 U1578 ( .A(u_alu_lt_x_11_n9), .Q(n3029) );
  NOR21 U1579 ( .A(n2995), .B(n2996), .Q(n2972) );
  NAND22 U1580 ( .A(n1756), .B(n1795), .Q(n1757) );
  NAND32 U1581 ( .A(n2463), .B(n2464), .C(n2462), .Q(n575) );
  NAND22 U1582 ( .A(n397), .B(n1879), .Q(n396) );
  NAND23 U1583 ( .A(n2368), .B(n567), .Q(n2424) );
  NAND23 U1584 ( .A(n660), .B(n658), .Q(n2196) );
  NAND22 U1585 ( .A(n2481), .B(n2274), .Q(n2393) );
  INV3 U1586 ( .A(n1304), .Q(n465) );
  NAND22 U1587 ( .A(n1304), .B(n1715), .Q(n1716) );
  INV3 U1588 ( .A(n2386), .Q(n1848) );
  NAND22 U1589 ( .A(u_alu_lt_x_11_B_0_), .B(n242), .Q(n1753) );
  NAND24 U1590 ( .A(n1256), .B(n2383), .Q(n1255) );
  NAND26 U1591 ( .A(u_alu_ashr_4_A_5_), .B(n234), .Q(n2462) );
  NOR22 U1592 ( .A(n1283), .B(n1282), .Q(n1281) );
  NAND23 U1593 ( .A(n1104), .B(n222), .Q(n2475) );
  NAND22 U1594 ( .A(n519), .B(n2163), .Q(n874) );
  INV2 U1595 ( .A(n2163), .Q(n2407) );
  NAND22 U1596 ( .A(n192), .B(n257), .Q(n354) );
  NAND22 U1597 ( .A(n2726), .B(n904), .Q(n903) );
  NAND23 U1598 ( .A(n1299), .B(n567), .Q(n2485) );
  INV2 U1599 ( .A(n2697), .Q(n639) );
  CLKIN6 U1600 ( .A(u_alu_DP_OP_83J3_124_3384_n152), .Q(n1143) );
  INV3 U1601 ( .A(alu_i_data_B[27]), .Q(n3058) );
  INV2 U1602 ( .A(n2033), .Q(n742) );
  INV3 U1603 ( .A(u_alu_lt_x_11_B_29_), .Q(n406) );
  INV3 U1604 ( .A(n2017), .Q(n1861) );
  INV3 U1605 ( .A(n1557), .Q(n1243) );
  INV3 U1606 ( .A(n1302), .Q(n1733) );
  INV3 U1607 ( .A(n1558), .Q(n1242) );
  INV2 U1608 ( .A(n2395), .Q(n2277) );
  NOR23 U1609 ( .A(n371), .B(n369), .Q(n915) );
  NOR24 U1610 ( .A(n3076), .B(n226), .Q(n585) );
  INV3 U1611 ( .A(u_alu_ashr_4_A_16_), .Q(n1746) );
  INV3 U1612 ( .A(n409), .Q(n408) );
  INV2 U1613 ( .A(n2025), .Q(n2040) );
  INV2 U1614 ( .A(n1569), .Q(n3073) );
  INV3 U1615 ( .A(n222), .Q(n659) );
  INV12 U1616 ( .A(n1523), .Q(n279) );
  CLKIN3 U1617 ( .A(n483), .Q(n476) );
  INV3 U1618 ( .A(n1074), .Q(n1158) );
  INV6 U1619 ( .A(n1863), .Q(n1083) );
  INV3 U1620 ( .A(n1859), .Q(n1157) );
  INV3 U1621 ( .A(n372), .Q(n371) );
  INV3 U1622 ( .A(n226), .Q(u_alu_lt_x_11_n144) );
  NAND23 U1623 ( .A(n997), .B(n1001), .Q(n1567) );
  INV6 U1624 ( .A(n1306), .Q(n221) );
  NOR21 U1625 ( .A(n1859), .B(n1159), .Q(n3095) );
  NOR23 U1626 ( .A(n586), .B(n1620), .Q(n913) );
  CLKIN6 U1627 ( .A(u_alu_DP_OP_85J3_126_1427_n374), .Q(n2627) );
  NAND22 U1628 ( .A(n1087), .B(n1370), .Q(n387) );
  CLKIN6 U1629 ( .A(n1422), .Q(n182) );
  NAND22 U1630 ( .A(n1648), .B(compare_i_data_rs[4]), .Q(n1074) );
  NAND23 U1631 ( .A(n1660), .B(n1683), .Q(n1168) );
  INV6 U1632 ( .A(n1305), .Q(n1306) );
  INV3 U1633 ( .A(n2590), .Q(n705) );
  INV3 U1634 ( .A(n1822), .Q(n1549) );
  NAND26 U1635 ( .A(n680), .B(n1544), .Q(u_alu_lt_x_11_A_3_) );
  NAND33 U1636 ( .A(n778), .B(n1369), .C(n1264), .Q(n777) );
  NAND22 U1637 ( .A(n1671), .B(n1683), .Q(n1672) );
  NOR22 U1638 ( .A(n944), .B(n965), .Q(n1081) );
  INV2 U1639 ( .A(n1866), .Q(n1821) );
  INV3 U1640 ( .A(n1997), .Q(n2028) );
  INV2 U1641 ( .A(n1791), .Q(n1784) );
  INV3 U1642 ( .A(n323), .Q(n322) );
  INV1 U1643 ( .A(n1725), .Q(n1726) );
  INV2 U1644 ( .A(n2382), .Q(n1865) );
  INV2 U1645 ( .A(n2131), .Q(n2135) );
  INV3 U1646 ( .A(n2801), .Q(n2495) );
  INV3 U1647 ( .A(n1729), .Q(n1170) );
  INV3 U1648 ( .A(n1013), .Q(n1012) );
  INV6 U1649 ( .A(n1317), .Q(n1321) );
  INV15 U1650 ( .A(n1351), .Q(n1350) );
  NAND24 U1651 ( .A(i_data_immext[11]), .B(n170), .Q(n2131) );
  INV3 U1652 ( .A(n1132), .Q(n357) );
  NAND21 U1653 ( .A(n177), .B(n1365), .Q(n1132) );
  NOR23 U1654 ( .A(n1016), .B(n1015), .Q(n944) );
  NAND23 U1655 ( .A(i_con_Efbmux[1]), .B(n1217), .Q(n1119) );
  INV2 U1656 ( .A(n34), .Q(n1333) );
  NAND22 U1657 ( .A(n1681), .B(i_con_Ealuop[5]), .Q(n531) );
  INV2 U1658 ( .A(i_data_FEalures[0]), .Q(n1085) );
  INV2 U1659 ( .A(i_data_FEalures[14]), .Q(n478) );
  INV2 U1660 ( .A(i_data_FEalures[28]), .Q(n790) );
  BUF12 U1661 ( .A(i_data_immext[10]), .Q(n1366) );
  INV3 U1662 ( .A(i_data_famemout[11]), .Q(n1436) );
  INV2 U1663 ( .A(i_data_famemout[1]), .Q(n1535) );
  INV3 U1664 ( .A(i_data_famemout[9]), .Q(n1401) );
  NAND22 U1665 ( .A(n2585), .B(n724), .Q(alu_o_data_AluRes[18]) );
  NAND33 U1666 ( .A(n2502), .B(n2503), .C(n2501), .Q(alu_o_data_AluRes[16]) );
  NOR22 U1667 ( .A(n1148), .B(n1287), .Q(n1286) );
  INV3 U1668 ( .A(n2082), .Q(n2084) );
  NOR22 U1669 ( .A(n686), .B(n685), .Q(n831) );
  NAND22 U1670 ( .A(n1021), .B(u_alu_pre_sum_4b[3]), .Q(n2925) );
  NOR22 U1671 ( .A(n1980), .B(n1979), .Q(n1981) );
  INV3 U1672 ( .A(n1177), .Q(n1030) );
  NAND22 U1673 ( .A(n2709), .B(n1345), .Q(n1238) );
  NOR22 U1674 ( .A(n555), .B(n551), .Q(n2919) );
  NOR22 U1675 ( .A(n947), .B(n2820), .Q(n1285) );
  NAND23 U1676 ( .A(n1344), .B(n207), .Q(n2317) );
  NAND22 U1677 ( .A(n298), .B(n167), .Q(n297) );
  OAI211 U1678 ( .A(n1343), .B(n1152), .C(n1150), .Q(n1151) );
  INV2 U1679 ( .A(n829), .Q(n828) );
  NAND22 U1680 ( .A(n833), .B(n168), .Q(n832) );
  NAND22 U1681 ( .A(n1172), .B(n204), .Q(n463) );
  INV3 U1682 ( .A(n1344), .Q(n202) );
  NAND22 U1683 ( .A(n1128), .B(n1127), .Q(n712) );
  INV3 U1684 ( .A(n2612), .Q(n1328) );
  INV12 U1685 ( .A(n1343), .Q(n1344) );
  INV3 U1686 ( .A(n2638), .Q(n676) );
  NOR22 U1687 ( .A(n936), .B(n2894), .Q(n935) );
  NOR22 U1688 ( .A(n251), .B(n1846), .Q(n1811) );
  INV3 U1689 ( .A(n888), .Q(n886) );
  OAI222 U1690 ( .A(n2024), .B(n1358), .C(n1359), .D(n2092), .Q(n2049) );
  INV3 U1691 ( .A(n442), .Q(n441) );
  OAI221 U1692 ( .A(n2211), .B(n1360), .C(n2092), .D(n1358), .Q(n2113) );
  NAND22 U1693 ( .A(n3021), .B(n885), .Q(n884) );
  AOI221 U1694 ( .A(n1841), .B(n1359), .C(n1840), .D(n1358), .Q(n1878) );
  NAND22 U1695 ( .A(u_alu_N306), .B(n1684), .Q(n1744) );
  MUX22 U1696 ( .A(n2601), .B(n2507), .S(n1358), .Q(n2557) );
  NAND22 U1697 ( .A(n2154), .B(n1358), .Q(n2155) );
  INV3 U1698 ( .A(n285), .Q(n284) );
  NAND21 U1699 ( .A(n2692), .B(n1357), .Q(n288) );
  INV3 U1700 ( .A(n263), .Q(n262) );
  NAND22 U1701 ( .A(n2952), .B(n2953), .Q(n822) );
  NAND22 U1702 ( .A(n2060), .B(n1359), .Q(n1943) );
  OAI211 U1703 ( .A(n229), .B(n2240), .C(n2239), .Q(n2241) );
  NOR22 U1704 ( .A(n461), .B(n458), .Q(n2144) );
  INV2 U1705 ( .A(n2367), .Q(n2167) );
  NAND22 U1706 ( .A(n404), .B(n402), .Q(u_alu_DP_OP_84J3_125_2615_n73) );
  IMUX21 U1707 ( .A(n2200), .B(n2201), .S(n2481), .Q(n2213) );
  NAND22 U1708 ( .A(n346), .B(n345), .Q(n1810) );
  NOR22 U1709 ( .A(n1773), .B(n1360), .Q(n442) );
  IMUX21 U1710 ( .A(n1754), .B(n1755), .S(u_alu_lt_x_11_n121), .Q(n1762) );
  INV3 U1711 ( .A(n2990), .Q(n496) );
  INV3 U1712 ( .A(n562), .Q(n561) );
  NAND22 U1713 ( .A(n2512), .B(n534), .Q(n2515) );
  OAI211 U1714 ( .A(n234), .B(n1895), .C(n1894), .Q(n1897) );
  INV3 U1715 ( .A(n1935), .Q(n1840) );
  NAND21 U1716 ( .A(n652), .B(n179), .Q(n1289) );
  OAI221 U1717 ( .A(n2220), .B(n249), .C(n2989), .D(n1356), .Q(n2221) );
  NAND21 U1718 ( .A(n1141), .B(n180), .Q(n2902) );
  OAI211 U1719 ( .A(n173), .B(n1898), .C(n1044), .Q(n1899) );
  INV3 U1720 ( .A(n1952), .Q(n1950) );
  NOR21 U1721 ( .A(n864), .B(n173), .Q(n1775) );
  NOR21 U1722 ( .A(n870), .B(n173), .Q(n2561) );
  NAND22 U1723 ( .A(n2358), .B(n204), .Q(n385) );
  INV3 U1724 ( .A(n610), .Q(n609) );
  AOI212 U1725 ( .A(n1947), .B(n359), .C(n216), .Q(n358) );
  AOI221 U1726 ( .A(n3052), .B(n249), .C(n3004), .D(n1356), .Q(n3005) );
  NAND22 U1727 ( .A(n1748), .B(n1361), .Q(n345) );
  NAND21 U1728 ( .A(n2913), .B(n1357), .Q(n825) );
  INV3 U1729 ( .A(n381), .Q(n380) );
  NOR22 U1730 ( .A(n1225), .B(n1223), .Q(n1229) );
  AOI211 U1731 ( .A(n1783), .B(n180), .C(n1782), .Q(n1802) );
  NOR33 U1732 ( .A(n1559), .B(n1005), .C(n1034), .Q(n694) );
  INV3 U1733 ( .A(n395), .Q(n394) );
  INV3 U1734 ( .A(n1779), .Q(n1780) );
  INV3 U1735 ( .A(n348), .Q(n347) );
  NAND22 U1736 ( .A(n2057), .B(n1363), .Q(n2058) );
  INV3 U1737 ( .A(n302), .Q(n301) );
  NOR21 U1738 ( .A(n2362), .B(n2359), .Q(n2360) );
  INV3 U1739 ( .A(n2362), .Q(n2366) );
  INV2 U1740 ( .A(n2913), .Q(n2915) );
  NAND22 U1741 ( .A(n2986), .B(n177), .Q(n633) );
  IMUX21 U1742 ( .A(n1355), .B(n91), .S(n1251), .Q(n1764) );
  INV3 U1743 ( .A(n2348), .Q(n1180) );
  NAND22 U1744 ( .A(n174), .B(n2287), .Q(n873) );
  NAND22 U1745 ( .A(n1939), .B(n245), .Q(n766) );
  NAND21 U1746 ( .A(n3053), .B(n1299), .Q(n3054) );
  NAND22 U1747 ( .A(n2505), .B(n1361), .Q(n2506) );
  NAND22 U1748 ( .A(n900), .B(n967), .Q(n624) );
  BUF12 U1749 ( .A(n180), .Q(n278) );
  NAND21 U1750 ( .A(n910), .B(n3053), .Q(n1327) );
  IMUX21 U1751 ( .A(n3047), .B(n1341), .S(n224), .Q(n2875) );
  NOR21 U1752 ( .A(n1356), .B(n3006), .Q(n252) );
  NAND22 U1753 ( .A(n982), .B(n2019), .Q(n2763) );
  INV3 U1754 ( .A(n1828), .Q(n1824) );
  IMUX21 U1755 ( .A(n3047), .B(n174), .S(n223), .Q(n1817) );
  INV2 U1756 ( .A(n869), .Q(n868) );
  NAND22 U1757 ( .A(n2162), .B(n2468), .Q(n2359) );
  NOR22 U1758 ( .A(n212), .B(n2139), .Q(n2104) );
  INV3 U1759 ( .A(n630), .Q(n629) );
  NOR21 U1760 ( .A(n2194), .B(n2141), .Q(n460) );
  IMUX21 U1761 ( .A(n1355), .B(n1342), .S(n231), .Q(n2107) );
  INV2 U1762 ( .A(n2814), .Q(n2799) );
  NAND21 U1763 ( .A(n658), .B(n2392), .Q(n2134) );
  INV3 U1764 ( .A(u_alu_DP_OP_84J3_125_2615_n8), .Q(u_alu_pre_sum_4a[0]) );
  IMUX21 U1765 ( .A(n3047), .B(n174), .S(n222), .Q(n2128) );
  NOR22 U1766 ( .A(n1687), .B(n1688), .Q(n1772) );
  NOR22 U1767 ( .A(n185), .B(n571), .Q(n2721) );
  CLKIN6 U1768 ( .A(n1035), .Q(n2388) );
  INV3 U1769 ( .A(u_alu_DP_OP_84J3_125_2615_n15), .Q(
        u_alu_DP_OP_84J3_125_2615_n70) );
  NAND22 U1770 ( .A(n2511), .B(n236), .Q(n898) );
  NAND22 U1771 ( .A(n745), .B(u_alu_DP_OP_84J3_125_2615_n103), .Q(n967) );
  INV3 U1772 ( .A(u_alu_DP_OP_84J3_125_2615_n46), .Q(
        u_alu_DP_OP_84J3_125_2615_n45) );
  NAND22 U1773 ( .A(n745), .B(u_alu_DP_OP_84J3_125_2615_n46), .Q(n899) );
  INV3 U1774 ( .A(n739), .Q(n2696) );
  INV3 U1775 ( .A(n755), .Q(n754) );
  NAND22 U1776 ( .A(n1842), .B(n272), .Q(n751) );
  INV2 U1777 ( .A(n2393), .Q(n2254) );
  INV6 U1778 ( .A(n1341), .Q(n1355) );
  OAI211 U1779 ( .A(n2649), .B(n2597), .C(n2596), .Q(n527) );
  INV3 U1780 ( .A(n353), .Q(n352) );
  NAND21 U1781 ( .A(n1341), .B(n2977), .Q(n869) );
  NOR21 U1782 ( .A(n2486), .B(n2365), .Q(n2288) );
  NAND21 U1783 ( .A(n2270), .B(n2393), .Q(n2185) );
  INV3 U1784 ( .A(n814), .Q(n813) );
  NOR21 U1785 ( .A(n1976), .B(n1972), .Q(n1937) );
  NOR23 U1786 ( .A(n2474), .B(n2161), .Q(n2468) );
  NOR22 U1787 ( .A(n2629), .B(n2558), .Q(n2597) );
  NOR21 U1788 ( .A(n2309), .B(n2308), .Q(n756) );
  INV3 U1789 ( .A(n788), .Q(n787) );
  NAND22 U1790 ( .A(n2463), .B(n2462), .Q(n2007) );
  INV3 U1791 ( .A(n874), .Q(n2403) );
  INV3 U1792 ( .A(u_alu_DP_OP_84J3_125_2615_n92), .Q(n900) );
  OAI211 U1793 ( .A(n248), .B(n2517), .C(n309), .Q(n535) );
  NAND22 U1794 ( .A(n2026), .B(n234), .Q(n291) );
  INV2 U1795 ( .A(u_alu_DP_OP_83J3_124_3384_n23), .Q(
        u_alu_DP_OP_83J3_124_3384_n83) );
  NAND28 U1796 ( .A(n1097), .B(n2439), .Q(n3049) );
  NOR22 U1797 ( .A(n857), .B(n2440), .Q(n1788) );
  INV3 U1798 ( .A(n2476), .Q(n360) );
  NAND22 U1799 ( .A(n517), .B(n516), .Q(n3014) );
  INV3 U1800 ( .A(n716), .Q(n715) );
  NAND23 U1801 ( .A(n1231), .B(n1232), .Q(n1230) );
  NOR22 U1802 ( .A(n289), .B(n2440), .Q(n1796) );
  NAND22 U1803 ( .A(n2985), .B(n176), .Q(n739) );
  NAND24 U1804 ( .A(n2466), .B(n2485), .Q(n2488) );
  NOR22 U1805 ( .A(n221), .B(n2693), .Q(n1954) );
  INV3 U1806 ( .A(u_alu_lt_x_11_n85), .Q(n2166) );
  NAND26 U1807 ( .A(n214), .B(n1097), .Q(n2976) );
  NAND20 U1808 ( .A(n1299), .B(n567), .Q(u_alu_lt_x_11_n71) );
  INV3 U1809 ( .A(n520), .Q(n518) );
  INV3 U1810 ( .A(n2466), .Q(n2365) );
  INV3 U1811 ( .A(n529), .Q(n1847) );
  NAND22 U1812 ( .A(n486), .B(n54), .Q(n2270) );
  INV3 U1813 ( .A(n1825), .Q(n1826) );
  NOR22 U1814 ( .A(n2793), .B(n2806), .Q(n792) );
  NOR21 U1815 ( .A(n2929), .B(n2856), .Q(n2828) );
  NAND24 U1816 ( .A(n1700), .B(n1353), .Q(u_alu_DP_OP_85J3_126_1427_n368) );
  NAND22 U1817 ( .A(n2164), .B(n519), .Q(n363) );
  NOR23 U1818 ( .A(n234), .B(u_alu_ashr_4_A_5_), .Q(u_alu_lt_x_11_n105) );
  NOR23 U1819 ( .A(n222), .B(u_alu_lt_x_11_B_11_), .Q(n2476) );
  NOR22 U1820 ( .A(n233), .B(n1070), .Q(n2486) );
  NOR23 U1821 ( .A(n567), .B(n1299), .Q(n2484) );
  INV3 U1822 ( .A(n2140), .Q(n2138) );
  NAND22 U1823 ( .A(n804), .B(n215), .Q(n707) );
  INV3 U1824 ( .A(n2041), .Q(n732) );
  INV3 U1825 ( .A(n1814), .Q(n1778) );
  NAND22 U1826 ( .A(n406), .B(n407), .Q(u_alu_DP_OP_84J3_125_2615_n109) );
  INV3 U1827 ( .A(n2392), .Q(n2182) );
  NOR22 U1828 ( .A(u_alu_DP_OP_84J3_125_2615_n39), .B(
        u_alu_DP_OP_84J3_125_2615_n36), .Q(n745) );
  INV3 U1829 ( .A(n306), .Q(n305) );
  INV2 U1830 ( .A(n1044), .Q(n2669) );
  INV2 U1831 ( .A(n914), .Q(n2871) );
  INV3 U1832 ( .A(n2754), .Q(n3059) );
  NOR21 U1833 ( .A(n2420), .B(n2417), .Q(n2263) );
  INV2 U1834 ( .A(u_alu_DP_OP_83J3_124_3384_n41), .Q(
        u_alu_DP_OP_83J3_124_3384_n121) );
  INV1 U1835 ( .A(n1332), .Q(n1330) );
  INV3 U1836 ( .A(n2205), .Q(n2208) );
  NOR23 U1837 ( .A(n1367), .B(n3012), .Q(n2726) );
  NAND21 U1838 ( .A(n2295), .B(n172), .Q(n2688) );
  INV3 U1839 ( .A(n2191), .Q(n794) );
  NAND22 U1840 ( .A(n664), .B(n229), .Q(n793) );
  INV2 U1841 ( .A(n2204), .Q(n190) );
  NAND22 U1842 ( .A(n1830), .B(n1363), .Q(n749) );
  INV6 U1843 ( .A(u_alu_lt_x_11_n77), .Q(n2480) );
  INV3 U1844 ( .A(n1273), .Q(n910) );
  INV6 U1845 ( .A(n2927), .Q(n191) );
  NAND22 U1846 ( .A(alu_i_data_B[27]), .B(n1517), .Q(
        u_alu_DP_OP_84J3_125_2615_n37) );
  INV3 U1847 ( .A(n764), .Q(n1777) );
  NOR22 U1848 ( .A(n225), .B(n3077), .Q(n393) );
  INV3 U1849 ( .A(n530), .Q(n1250) );
  NAND22 U1850 ( .A(u_alu_DP_OP_83J3_124_3384_n153), .B(n248), .Q(n923) );
  NAND22 U1851 ( .A(n217), .B(n1251), .Q(n1795) );
  NOR22 U1852 ( .A(n2093), .B(n730), .Q(n729) );
  INV3 U1853 ( .A(n265), .Q(n264) );
  INV3 U1854 ( .A(n1276), .Q(n407) );
  BUF6 U1855 ( .A(alu_i_data_B[27]), .Q(n192) );
  NAND21 U1856 ( .A(n2252), .B(n177), .Q(n1686) );
  NOR22 U1857 ( .A(n161), .B(n2146), .Q(n654) );
  NAND22 U1858 ( .A(n2252), .B(n256), .Q(n2275) );
  NAND32 U1859 ( .A(n2036), .B(u_alu_lt_x_11_n121), .C(n2035), .Q(n530) );
  NAND22 U1860 ( .A(n2146), .B(n1361), .Q(n748) );
  NAND32 U1861 ( .A(n2548), .B(n2549), .C(n1307), .Q(n2793) );
  NAND22 U1862 ( .A(u_alu_lt_x_11_B_25_), .B(u_alu_DP_OP_85J3_126_1427_n379), 
        .Q(u_alu_DP_OP_84J3_125_2615_n48) );
  NOR22 U1863 ( .A(n1041), .B(n1731), .Q(n893) );
  INV3 U1864 ( .A(n1494), .Q(n3079) );
  INV2 U1865 ( .A(n182), .Q(n1103) );
  NAND22 U1866 ( .A(n123), .B(n357), .Q(n2689) );
  INV3 U1867 ( .A(n2146), .Q(n1970) );
  INV2 U1868 ( .A(n2594), .Q(u_alu_lt_x_11_n139) );
  INV3 U1869 ( .A(n296), .Q(n295) );
  NAND22 U1870 ( .A(n1717), .B(n312), .Q(n1411) );
  NAND22 U1871 ( .A(n1188), .B(n1353), .Q(n1187) );
  NAND22 U1872 ( .A(u_alu_DP_OP_85J3_126_1427_n377), .B(n1353), .Q(n2740) );
  INV2 U1873 ( .A(n2629), .Q(u_alu_lt_x_11_n138) );
  NOR24 U1874 ( .A(n682), .B(n681), .Q(n2027) );
  NAND22 U1875 ( .A(n1215), .B(n1548), .Q(n808) );
  INV1 U1876 ( .A(n1606), .Q(n474) );
  INV6 U1877 ( .A(u_alu_DP_OP_85J3_126_1427_n379), .Q(n195) );
  NAND24 U1878 ( .A(n1570), .B(n1082), .Q(u_alu_lt_x_11_A_0_) );
  NOR21 U1879 ( .A(n241), .B(n855), .Q(n1996) );
  NAND22 U1880 ( .A(n437), .B(n436), .Q(n435) );
  NAND22 U1881 ( .A(n477), .B(n479), .Q(n483) );
  INV6 U1882 ( .A(n1517), .Q(n196) );
  NAND23 U1883 ( .A(n445), .B(n1322), .Q(n1323) );
  NAND22 U1884 ( .A(n513), .B(n1003), .Q(n512) );
  NAND22 U1885 ( .A(n276), .B(n2064), .Q(n275) );
  NAND22 U1886 ( .A(n445), .B(n940), .Q(n939) );
  BUF15 U1887 ( .A(n2966), .Q(n1307) );
  INV2 U1888 ( .A(n3088), .Q(n1155) );
  NAND22 U1889 ( .A(n1321), .B(i_data_famemout[30]), .Q(n1279) );
  NAND23 U1890 ( .A(n237), .B(n790), .Q(n1201) );
  INV3 U1891 ( .A(n258), .Q(n257) );
  INV3 U1892 ( .A(n945), .Q(n431) );
  INV12 U1893 ( .A(n239), .Q(n1353) );
  NOR22 U1894 ( .A(n1618), .B(n1619), .Q(n587) );
  INV3 U1895 ( .A(n452), .Q(n451) );
  NAND22 U1896 ( .A(n1993), .B(n859), .Q(n855) );
  INV3 U1897 ( .A(n1488), .Q(n623) );
  INV3 U1898 ( .A(n303), .Q(n1082) );
  INV6 U1899 ( .A(n283), .Q(n622) );
  INV3 U1900 ( .A(n399), .Q(n398) );
  NAND23 U1901 ( .A(n237), .B(n1555), .Q(n1248) );
  INV1 U1902 ( .A(n2589), .Q(n706) );
  NOR23 U1903 ( .A(i_data_FEalures[16]), .B(n1349), .Q(n2804) );
  INV3 U1904 ( .A(n273), .Q(n272) );
  NAND22 U1905 ( .A(n63), .B(n1369), .Q(n617) );
  INV3 U1906 ( .A(n507), .Q(n370) );
  NAND33 U1907 ( .A(n1398), .B(n1397), .C(n1396), .Q(compare_i_data_rs[14]) );
  NAND22 U1908 ( .A(n1427), .B(n1425), .Q(n1166) );
  OAI212 U1909 ( .A(n1658), .B(n944), .C(n1864), .Q(n1659) );
  INV3 U1910 ( .A(n294), .Q(n293) );
  CLKIN6 U1911 ( .A(n1994), .Q(n274) );
  INV3 U1912 ( .A(n1625), .Q(n436) );
  NOR23 U1913 ( .A(i_data_FEalures[7]), .B(n1350), .Q(n2000) );
  INV3 U1914 ( .A(n1116), .Q(n1115) );
  INV3 U1915 ( .A(n1461), .Q(n1462) );
  NAND22 U1916 ( .A(n2801), .B(n1369), .Q(n649) );
  INV6 U1917 ( .A(n1530), .Q(n2186) );
  INV3 U1918 ( .A(n1481), .Q(n1482) );
  NAND22 U1919 ( .A(n709), .B(n1583), .Q(n1048) );
  BUF6 U1920 ( .A(compare_i_data_rs[4]), .Q(n197) );
  NAND22 U1921 ( .A(n240), .B(i_data_fbmemout[31]), .Q(n852) );
  INV4 U1922 ( .A(n1214), .Q(n413) );
  NOR22 U1923 ( .A(i_data_fbmemout[22]), .B(n246), .Q(n1050) );
  NAND21 U1924 ( .A(n89), .B(i_data_FMalures[9]), .Q(n1010) );
  AOI211 U1925 ( .A(n1335), .B(i_data_FEalures[8]), .C(n744), .Q(n743) );
  INV2 U1926 ( .A(n2562), .Q(n2564) );
  INV3 U1927 ( .A(n2759), .Q(n2606) );
  NAND21 U1928 ( .A(n89), .B(i_data_FMalures[15]), .Q(n1399) );
  INV3 U1929 ( .A(n2766), .Q(n243) );
  NAND22 U1930 ( .A(n1319), .B(i_data_famemout[22]), .Q(n709) );
  INV3 U1931 ( .A(n313), .Q(n312) );
  INV3 U1932 ( .A(n768), .Q(n767) );
  NOR21 U1933 ( .A(i_data_fbmemout[11]), .B(n246), .Q(n616) );
  INV15 U1934 ( .A(n244), .Q(n198) );
  NAND22 U1935 ( .A(n1319), .B(i_data_famemout[18]), .Q(n1465) );
  NAND24 U1936 ( .A(n170), .B(n1362), .Q(n2062) );
  NOR22 U1937 ( .A(n246), .B(i_data_fbmemout[18]), .Q(n1620) );
  NAND21 U1938 ( .A(n89), .B(i_data_FMalures[26]), .Q(n1503) );
  NOR22 U1939 ( .A(i_data_fbmemout[24]), .B(n246), .Q(n785) );
  NOR23 U1940 ( .A(i_data_rt[2]), .B(n1218), .Q(n1297) );
  NAND22 U1941 ( .A(n90), .B(i_data_FMalures[1]), .Q(n318) );
  NOR21 U1942 ( .A(n943), .B(n1864), .Q(n367) );
  INV15 U1943 ( .A(n1352), .Q(n1324) );
  INV3 U1944 ( .A(n166), .Q(n245) );
  NAND22 U1945 ( .A(n158), .B(i_data_rs[17]), .Q(n1467) );
  NAND21 U1946 ( .A(n172), .B(n1356), .Q(n768) );
  NAND22 U1947 ( .A(n159), .B(i_data_rs[19]), .Q(n817) );
  NAND21 U1948 ( .A(n248), .B(n1364), .Q(n905) );
  NAND22 U1949 ( .A(n248), .B(n166), .Q(n2562) );
  NOR22 U1950 ( .A(i_con_Ealuop[3]), .B(n1662), .Q(n533) );
  INV6 U1951 ( .A(i_con_Efbmux[0]), .Q(n1217) );
  INV2 U1952 ( .A(i_data_FEalures[9]), .Q(n1121) );
  INV3 U1953 ( .A(i_data_FEalures[31]), .Q(n1407) );
  INV3 U1954 ( .A(i_data_rt[13]), .Q(n1473) );
  NAND32 U1955 ( .A(n985), .B(n984), .C(n983), .Q(alu_o_data_AluRes[12]) );
  NAND22 U1956 ( .A(n1286), .B(n1284), .Q(alu_o_data_AluRes[24]) );
  NOR32 U1957 ( .A(n2617), .B(n2616), .C(n2615), .Q(n2618) );
  NOR23 U1958 ( .A(n2684), .B(n2683), .Q(n2685) );
  AOI2112 U1959 ( .A(n2715), .B(u_alu_pre_sum_3a[1]), .C(n952), .D(n950), .Q(
        n949) );
  NAND33 U1960 ( .A(n1837), .B(n1835), .C(n1836), .Q(alu_o_data_AluRes[3]) );
  NAND22 U1961 ( .A(n2849), .B(n962), .Q(n2850) );
  INV3 U1962 ( .A(n678), .Q(n677) );
  NAND22 U1963 ( .A(n463), .B(n2167), .Q(n987) );
  AOI211 U1964 ( .A(n2441), .B(u_alu_ashr_4_A_16_), .C(n1094), .Q(n2451) );
  NOR22 U1965 ( .A(n2289), .B(n1177), .Q(n685) );
  NOR22 U1966 ( .A(n2494), .B(n763), .Q(n2015) );
  AOI212 U1967 ( .A(n2357), .B(n2356), .C(n2355), .Q(n2380) );
  NAND22 U1968 ( .A(n523), .B(n168), .Q(n1877) );
  NAND22 U1969 ( .A(n599), .B(n2715), .Q(n589) );
  AOI212 U1970 ( .A(n2258), .B(n2357), .C(n2257), .Q(n2267) );
  NAND22 U1971 ( .A(n2652), .B(n828), .Q(n1204) );
  NAND33 U1972 ( .A(n1967), .B(n1966), .C(n1965), .Q(n1980) );
  NAND22 U1973 ( .A(n288), .B(n284), .Q(n2660) );
  INV3 U1974 ( .A(n935), .Q(n2858) );
  NOR22 U1975 ( .A(n3066), .B(n687), .Q(n686) );
  NAND22 U1976 ( .A(n2078), .B(n426), .Q(n713) );
  INV3 U1977 ( .A(n834), .Q(n833) );
  NOR22 U1978 ( .A(n951), .B(n3006), .Q(n950) );
  NAND22 U1979 ( .A(n2113), .B(n2883), .Q(n269) );
  NAND22 U1980 ( .A(n1343), .B(n917), .Q(n1150) );
  OAI211 U1981 ( .A(n1356), .B(n2300), .C(n168), .Q(n2232) );
  INV3 U1982 ( .A(n1878), .Q(n298) );
  AOI211 U1983 ( .A(n802), .B(n1139), .C(n3066), .Q(n801) );
  XNR22 U1984 ( .A(n3041), .B(n3040), .Q(n3070) );
  NAND33 U1985 ( .A(n1873), .B(n1270), .C(n1269), .Q(n1268) );
  NOR22 U1986 ( .A(n249), .B(n1945), .Q(n1946) );
  AOI221 U1987 ( .A(n2724), .B(n1359), .C(n2844), .D(n1358), .Q(n596) );
  AOI211 U1988 ( .A(n168), .B(n2772), .C(n2771), .Q(n2819) );
  AOI212 U1989 ( .A(n2777), .B(n2843), .C(n2776), .Q(n2818) );
  NAND22 U1990 ( .A(n1810), .B(n201), .Q(n439) );
  NOR21 U1991 ( .A(n277), .B(n1897), .Q(n1900) );
  INV6 U1992 ( .A(n974), .Q(n326) );
  OAI221 U1993 ( .A(n1357), .B(n2757), .C(n2837), .D(n1356), .Q(n2772) );
  XNR21 U1994 ( .A(u_alu_DP_OP_84J3_125_2615_n2), .B(
        u_alu_DP_OP_84J3_125_2615_n73), .Q(u_alu_pre_sum_4b[6]) );
  OAI221 U1995 ( .A(n2024), .B(n1359), .C(n1935), .D(n1358), .Q(n1938) );
  NOR32 U1996 ( .A(n3056), .B(n1359), .C(n3057), .Q(n495) );
  XNR21 U1997 ( .A(n2799), .B(n1298), .Q(n2817) );
  INV3 U1998 ( .A(n497), .Q(n492) );
  INV3 U1999 ( .A(n2737), .Q(n592) );
  NAND23 U2000 ( .A(n2515), .B(n2514), .Q(n2612) );
  NAND22 U2001 ( .A(n1183), .B(n2928), .Q(n2827) );
  NOR22 U2002 ( .A(n1356), .B(n2659), .Q(n263) );
  NAND22 U2003 ( .A(n1009), .B(n2928), .Q(n2825) );
  NAND22 U2004 ( .A(n559), .B(n2917), .Q(n558) );
  IMUX21 U2005 ( .A(n2646), .B(n2645), .S(u_alu_DP_OP_85J3_126_1427_n374), .Q(
        n2647) );
  NOR31 U2006 ( .A(n1954), .B(n1953), .C(n1950), .Q(n1958) );
  INV3 U2007 ( .A(n385), .Q(n384) );
  NAND22 U2008 ( .A(n916), .B(n3043), .Q(n691) );
  NAND22 U2009 ( .A(n3043), .B(n1190), .Q(n1183) );
  NAND22 U2010 ( .A(n609), .B(n2332), .Q(n2507) );
  IMUX21 U2011 ( .A(n2130), .B(n2129), .S(u_alu_lt_x_11_A_11_), .Q(n2150) );
  XNR21 U2012 ( .A(n2351), .B(n2350), .Q(n2356) );
  NOR22 U2013 ( .A(n1358), .B(n1916), .Q(n526) );
  XOR21 U2014 ( .A(u_alu_DP_OP_84J3_125_2615_n3), .B(n846), .Q(n845) );
  INV3 U2015 ( .A(n797), .Q(n796) );
  NAND22 U2016 ( .A(n1809), .B(n1361), .Q(n349) );
  INV6 U2017 ( .A(n757), .Q(n2307) );
  OAI212 U2018 ( .A(n173), .B(n2107), .C(n910), .Q(n2111) );
  IMUX21 U2019 ( .A(n2109), .B(n2108), .S(n184), .Q(n2110) );
  XNR21 U2020 ( .A(n2256), .B(n2255), .Q(n2258) );
  NAND22 U2021 ( .A(n766), .B(n1940), .Q(n2153) );
  IMUX21 U2022 ( .A(n1963), .B(n1962), .S(n1971), .Q(n1966) );
  AOI221 U2023 ( .A(n1357), .B(n2978), .C(n2939), .D(n1356), .Q(n2942) );
  NOR21 U2024 ( .A(n866), .B(n173), .Q(n2645) );
  IMUX21 U2025 ( .A(n2045), .B(n2044), .S(n316), .Q(n2046) );
  OAI211 U2026 ( .A(n1356), .B(n2915), .C(n2914), .Q(n559) );
  NAND22 U2027 ( .A(n2954), .B(n1359), .Q(n823) );
  AOI211 U2028 ( .A(n2306), .B(n2305), .C(n2311), .Q(n2318) );
  NOR21 U2029 ( .A(n868), .B(n173), .Q(n2240) );
  IMUX21 U2030 ( .A(n1735), .B(n1734), .S(n289), .Q(n1739) );
  NOR31 U2031 ( .A(n1723), .B(n1722), .C(n1721), .Q(n1740) );
  AOI221 U2032 ( .A(n1362), .B(n1748), .C(n627), .D(n175), .Q(n626) );
  NAND21 U2033 ( .A(n3004), .B(n1357), .Q(n499) );
  INV2 U2034 ( .A(n2894), .Q(n2893) );
  IMUX21 U2035 ( .A(n1872), .B(n1871), .S(n227), .Q(n1873) );
  INV3 U2036 ( .A(n3067), .Q(n799) );
  NAND22 U2037 ( .A(n2878), .B(n1327), .Q(n2879) );
  NAND22 U2038 ( .A(n825), .B(n2914), .Q(n824) );
  OAI211 U2039 ( .A(n173), .B(n2733), .C(u_alu_DP_OP_83J3_124_3384_n153), .Q(
        n2735) );
  NOR22 U2040 ( .A(n396), .B(n394), .Q(n2059) );
  OAI211 U2041 ( .A(n173), .B(n2831), .C(u_alu_lt_x_11_B_25_), .Q(n2832) );
  NAND22 U2042 ( .A(n1706), .B(n1705), .Q(n1809) );
  NAND33 U2043 ( .A(n3011), .B(n891), .C(n890), .Q(n889) );
  NAND22 U2044 ( .A(n2156), .B(n1356), .Q(n2157) );
  OAI212 U2045 ( .A(n1825), .B(n1824), .C(n470), .Q(n469) );
  NAND22 U2046 ( .A(n1989), .B(n110), .Q(n830) );
  IMUX21 U2047 ( .A(n3047), .B(n174), .S(u_alu_lt_x_11_n122), .Q(n1783) );
  XNR21 U2048 ( .A(n527), .B(n2599), .Q(n2595) );
  NOR21 U2049 ( .A(n2025), .B(n255), .Q(n1871) );
  INV3 U2050 ( .A(n865), .Q(n864) );
  NAND22 U2051 ( .A(n278), .B(n1318), .Q(n311) );
  NAND22 U2052 ( .A(n2643), .B(n217), .Q(n1755) );
  NOR22 U2053 ( .A(n1366), .B(n428), .Q(n2075) );
  INV3 U2054 ( .A(n861), .Q(n860) );
  OAI211 U2055 ( .A(n2161), .B(n2124), .C(n2165), .Q(n1173) );
  IMUX21 U2056 ( .A(n2448), .B(n2447), .S(u_alu_DP_OP_83J3_124_3384_n154), .Q(
        n2449) );
  XNR21 U2057 ( .A(n2134), .B(n2133), .Q(n2145) );
  NAND22 U2058 ( .A(n1845), .B(n1358), .Q(n525) );
  IMUX21 U2059 ( .A(n460), .B(n2141), .S(n2140), .Q(n459) );
  NAND22 U2060 ( .A(n2643), .B(n2904), .Q(n2130) );
  INV3 U2061 ( .A(u_alu_DP_OP_84J3_125_2615_n1), .Q(n282) );
  NAND22 U2062 ( .A(n1694), .B(n753), .Q(n1844) );
  OAI212 U2063 ( .A(n271), .B(u_alu_DP_OP_83J3_124_3384_n18), .C(
        u_alu_DP_OP_83J3_124_3384_n19), .Q(n600) );
  IMUX21 U2064 ( .A(n2732), .B(n2731), .S(n2780), .Q(n2736) );
  OAI221 U2065 ( .A(n1816), .B(n1358), .C(n1896), .D(n1359), .Q(n1819) );
  IMUX21 U2066 ( .A(n3051), .B(n3050), .S(n290), .Q(n3055) );
  NAND22 U2067 ( .A(n3009), .B(n444), .Q(n890) );
  NAND22 U2068 ( .A(n1882), .B(n1362), .Q(n346) );
  NOR32 U2069 ( .A(n1826), .B(n1828), .C(n1829), .Q(n1827) );
  INV3 U2070 ( .A(n252), .Q(n251) );
  INV3 U2071 ( .A(n863), .Q(n862) );
  OAI211 U2072 ( .A(n195), .B(n2841), .C(n2840), .Q(n2842) );
  NOR21 U2073 ( .A(n2218), .B(n2219), .Q(n2989) );
  OAI212 U2074 ( .A(u_alu_DP_OP_83J3_124_3384_n25), .B(n271), .C(
        u_alu_DP_OP_83J3_124_3384_n26), .Q(n1300) );
  NOR21 U2075 ( .A(n910), .B(n255), .Q(n2108) );
  NAND21 U2076 ( .A(n2643), .B(n1924), .Q(n1894) );
  NAND22 U2077 ( .A(n3063), .B(n1138), .Q(n1137) );
  NOR21 U2078 ( .A(n2204), .B(n255), .Q(n2044) );
  XOR21 U2079 ( .A(u_alu_DP_OP_83J3_124_3384_n5), .B(n271), .Q(
        u_alu_pre_sum_3a[4]) );
  OAI211 U2080 ( .A(n1976), .B(n1975), .C(n1974), .Q(n652) );
  NAND31 U2081 ( .A(n2643), .B(n2517), .C(n2516), .Q(n2518) );
  INV3 U2082 ( .A(n867), .Q(n866) );
  OAI211 U2083 ( .A(n1720), .B(n2494), .C(n1719), .Q(n1721) );
  NOR21 U2084 ( .A(n2146), .B(n255), .Q(n1962) );
  INV3 U2085 ( .A(n871), .Q(n870) );
  INV2 U2086 ( .A(n663), .Q(n2304) );
  NAND22 U2087 ( .A(n663), .B(n2419), .Q(n2306) );
  IMUX21 U2088 ( .A(n1355), .B(n91), .S(n568), .Q(n2352) );
  IMUX21 U2089 ( .A(n91), .B(n1355), .S(n2516), .Q(n2521) );
  INV2 U2090 ( .A(n2234), .Q(n2235) );
  INV2 U2091 ( .A(n2364), .Q(n2281) );
  AOI211 U2092 ( .A(n2824), .B(n1341), .C(n971), .Q(n2841) );
  NAND22 U2093 ( .A(u_alu_lt_x_11_n13), .B(u_alu_lt_x_11_n7), .Q(
        u_alu_lt_x_11_n5) );
  INV3 U2094 ( .A(n996), .Q(n504) );
  IMUX21 U2095 ( .A(n1355), .B(n1342), .S(n289), .Q(n1737) );
  NAND22 U2096 ( .A(n1192), .B(n2857), .Q(n690) );
  NAND22 U2097 ( .A(n2669), .B(n174), .Q(n861) );
  AOI211 U2098 ( .A(n2510), .B(n2509), .C(n2606), .Q(n2442) );
  NOR21 U2099 ( .A(u_alu_ashr_4_A_16_), .B(n3049), .Q(n2448) );
  NOR22 U2100 ( .A(n2597), .B(n2546), .Q(n2551) );
  INV2 U2101 ( .A(n2671), .Q(n1892) );
  NOR22 U2102 ( .A(n177), .B(n2329), .Q(n1939) );
  INV3 U2103 ( .A(n50), .Q(n2745) );
  IMUX21 U2104 ( .A(n3047), .B(n174), .S(n227), .Q(n1857) );
  NAND22 U2105 ( .A(n174), .B(n2946), .Q(n863) );
  NAND22 U2106 ( .A(n2444), .B(n1366), .Q(n661) );
  NAND22 U2107 ( .A(n174), .B(n1782), .Q(n865) );
  NAND22 U2108 ( .A(n2604), .B(n172), .Q(n1896) );
  NOR22 U2109 ( .A(n2863), .B(n2864), .Q(n563) );
  NAND21 U2110 ( .A(n3053), .B(n2146), .Q(n2734) );
  OAI211 U2111 ( .A(u_alu_DP_OP_83J3_124_3384_n32), .B(
        u_alu_DP_OP_83J3_124_3384_n1), .C(u_alu_DP_OP_83J3_124_3384_n33), .Q(
        u_alu_DP_OP_83J3_124_3384_n31) );
  INV6 U2112 ( .A(n2053), .Q(n2012) );
  AOI211 U2113 ( .A(n2704), .B(n2663), .C(u_alu_lt_x_11_n47), .Q(n2664) );
  NAND22 U2114 ( .A(n1880), .B(n245), .Q(n395) );
  NAND21 U2115 ( .A(n174), .B(n182), .Q(n1100) );
  INV6 U2116 ( .A(n3049), .Q(n2643) );
  NOR21 U2117 ( .A(n193), .B(n3049), .Q(n2667) );
  NAND22 U2118 ( .A(n2558), .B(n174), .Q(n871) );
  INV2 U2119 ( .A(n1099), .Q(n1098) );
  IMUX21 U2120 ( .A(n1355), .B(n1342), .S(n519), .Q(n2043) );
  NOR31 U2121 ( .A(n1953), .B(n1954), .C(n1951), .Q(n741) );
  IMUX21 U2122 ( .A(n1355), .B(n1342), .S(n161), .Q(n1964) );
  NOR22 U2123 ( .A(n1849), .B(n1820), .Q(n1829) );
  OAI211 U2124 ( .A(n166), .B(n2056), .C(n2229), .Q(n2057) );
  AOI211 U2125 ( .A(n3053), .B(n1234), .C(n2559), .Q(n2560) );
  IMUX21 U2126 ( .A(n1355), .B(n1342), .S(n444), .Q(n3008) );
  NOR22 U2127 ( .A(n2011), .B(n2007), .Q(n1295) );
  IMUX21 U2128 ( .A(n3047), .B(n174), .S(n2786), .Q(n2666) );
  NAND22 U2129 ( .A(n2358), .B(n2466), .Q(n2362) );
  NAND22 U2130 ( .A(n174), .B(n2644), .Q(n867) );
  IMUX21 U2131 ( .A(n1355), .B(n91), .S(n1314), .Q(n1898) );
  IMUX21 U2132 ( .A(n3047), .B(n174), .S(n1717), .Q(n3048) );
  NAND22 U2133 ( .A(n2322), .B(n2321), .Q(n2443) );
  NOR22 U2134 ( .A(n1360), .B(n3003), .Q(n3052) );
  NOR23 U2135 ( .A(n2996), .B(n2994), .Q(n3030) );
  NOR21 U2136 ( .A(n1357), .B(n3062), .Q(n3063) );
  NAND22 U2137 ( .A(n1055), .B(n1053), .Q(n3035) );
  NOR22 U2138 ( .A(n2166), .B(n2165), .Q(n630) );
  NOR22 U2139 ( .A(n1357), .B(n1753), .Q(n2444) );
  NAND22 U2140 ( .A(n639), .B(n739), .Q(n377) );
  NOR22 U2141 ( .A(n185), .B(n2655), .Q(n2835) );
  NOR23 U2142 ( .A(n2192), .B(n2195), .Q(n2141) );
  NOR22 U2143 ( .A(n1924), .B(n1923), .Q(n1951) );
  NAND22 U2144 ( .A(n2270), .B(n2415), .Q(n2197) );
  NOR31 U2145 ( .A(n2629), .B(n688), .C(n3049), .Q(n2559) );
  OAI212 U2146 ( .A(n770), .B(n2866), .C(n185), .Q(n769) );
  INV3 U2147 ( .A(n2746), .Q(n208) );
  NAND21 U2148 ( .A(n2716), .B(n1365), .Q(n2322) );
  NOR21 U2149 ( .A(n1331), .B(n3061), .Q(n3062) );
  INV2 U2150 ( .A(n2470), .Q(n2162) );
  NOR21 U2151 ( .A(n1936), .B(n1862), .Q(n1870) );
  NOR21 U2152 ( .A(n182), .B(n91), .Q(n1099) );
  INV2 U2153 ( .A(n2421), .Q(n2276) );
  NAND22 U2154 ( .A(n2968), .B(n1054), .Q(n1053) );
  INV2 U2155 ( .A(n1891), .Q(n2673) );
  INV2 U2156 ( .A(n2422), .Q(n2342) );
  NAND22 U2157 ( .A(n2742), .B(n2741), .Q(n2706) );
  OAI211 U2158 ( .A(n2597), .B(n2632), .C(n2596), .Q(n2598) );
  OAI211 U2159 ( .A(n621), .B(u_alu_lt_x_11_n26), .C(n2932), .Q(
        u_alu_lt_x_11_n22) );
  INV2 U2160 ( .A(u_alu_DP_OP_83J3_124_3384_n44), .Q(
        u_alu_DP_OP_83J3_124_3384_n122) );
  NAND22 U2161 ( .A(n190), .B(n2406), .Q(n642) );
  NAND22 U2162 ( .A(n351), .B(n1358), .Q(n350) );
  NAND22 U2163 ( .A(n1230), .B(n1365), .Q(n982) );
  NAND22 U2164 ( .A(n2716), .B(n166), .Q(n717) );
  NAND33 U2165 ( .A(n2412), .B(n2411), .C(n2410), .Q(n2413) );
  NAND22 U2166 ( .A(n2758), .B(n166), .Q(n668) );
  NAND22 U2167 ( .A(n3014), .B(n1364), .Q(n2719) );
  NOR32 U2168 ( .A(n227), .B(n2025), .C(n188), .Q(n2454) );
  INV2 U2169 ( .A(u_alu_DP_OP_84J3_125_2615_n49), .Q(
        u_alu_DP_OP_84J3_125_2615_n58) );
  NOR22 U2170 ( .A(n1280), .B(u_alu_DP_OP_85J3_126_1427_n368), .Q(n3034) );
  NAND22 U2171 ( .A(n2871), .B(n200), .Q(n2938) );
  NAND22 U2172 ( .A(n2115), .B(n2114), .Q(n2297) );
  NOR22 U2173 ( .A(n200), .B(n2937), .Q(n353) );
  NAND22 U2174 ( .A(n964), .B(n874), .Q(n645) );
  INV2 U2175 ( .A(n2081), .Q(n1992) );
  NOR22 U2176 ( .A(n1306), .B(n2693), .Q(n1972) );
  INV1 U2177 ( .A(n2486), .Q(n2363) );
  INV3 U2178 ( .A(n2972), .Q(n210) );
  NAND22 U2179 ( .A(n670), .B(n669), .Q(n2758) );
  NAND22 U2180 ( .A(n1299), .B(n172), .Q(n755) );
  XOR21 U2181 ( .A(n2543), .B(n2539), .Q(n2542) );
  INV2 U2182 ( .A(n2463), .Q(n1862) );
  AOI211 U2183 ( .A(n2115), .B(n2114), .C(n169), .Q(n740) );
  NOR21 U2184 ( .A(n185), .B(n1685), .Q(n1688) );
  NAND21 U2185 ( .A(n2867), .B(n1364), .Q(n772) );
  NOR22 U2186 ( .A(n1251), .B(n1255), .Q(n579) );
  NOR22 U2187 ( .A(n1851), .B(n1847), .Q(n1758) );
  NOR21 U2188 ( .A(u_alu_lt_x_11_n29), .B(u_alu_lt_x_11_n31), .Q(
        u_alu_lt_x_11_n27) );
  NAND21 U2189 ( .A(u_alu_lt_x_11_n138), .B(n688), .Q(u_alu_lt_x_11_n56) );
  NAND22 U2190 ( .A(n2386), .B(n1036), .Q(n1035) );
  NOR23 U2191 ( .A(n1304), .B(n2439), .Q(n1713) );
  NOR31 U2192 ( .A(n1302), .B(n1304), .C(n2439), .Q(n1718) );
  NOR21 U2193 ( .A(n356), .B(n355), .Q(n2756) );
  NAND22 U2194 ( .A(u_alu_lt_x_11_n77), .B(n2467), .Q(n814) );
  NAND22 U2195 ( .A(n2809), .B(n707), .Q(n702) );
  NAND22 U2196 ( .A(n444), .B(u_alu_DP_OP_85J3_126_1427_n368), .Q(
        u_alu_DP_OP_84J3_125_2615_n15) );
  NOR22 U2197 ( .A(n1524), .B(u_alu_lt_x_11_B_28_), .Q(
        u_alu_DP_OP_84J3_125_2615_n30) );
  NOR22 U2198 ( .A(n876), .B(n1144), .Q(n875) );
  NAND22 U2199 ( .A(u_alu_lt_x_11_n85), .B(u_alu_lt_x_11_n86), .Q(n362) );
  INV6 U2200 ( .A(n2369), .Q(n2368) );
  NAND21 U2201 ( .A(n359), .B(n735), .Q(n1856) );
  NOR22 U2202 ( .A(n316), .B(n2204), .Q(n520) );
  NOR22 U2203 ( .A(n1715), .B(n1733), .Q(n1712) );
  NOR21 U2204 ( .A(n688), .B(u_alu_lt_x_11_n138), .Q(u_alu_lt_x_11_n55) );
  NAND22 U2205 ( .A(n2948), .B(n1364), .Q(n379) );
  AOI212 U2206 ( .A(n2461), .B(n2460), .C(u_alu_lt_x_11_n112), .Q(n2465) );
  NAND22 U2207 ( .A(n856), .B(n1251), .Q(n2457) );
  OAI221 U2208 ( .A(n1970), .B(n1367), .C(n1984), .D(n172), .Q(n1693) );
  INV1 U2209 ( .A(n2423), .Q(n2305) );
  NAND21 U2210 ( .A(u_alu_lt_x_11_B_24_), .B(n175), .Q(n1125) );
  NAND21 U2211 ( .A(n1825), .B(n2387), .Q(n1789) );
  NAND21 U2212 ( .A(u_alu_lt_x_11_B_11_), .B(n1363), .Q(n2319) );
  INV6 U2213 ( .A(u_alu_ashr_4_A_5_), .Q(n2026) );
  NAND21 U2214 ( .A(n1299), .B(n169), .Q(n927) );
  INV2 U2215 ( .A(u_alu_lt_x_11_n112), .Q(n1831) );
  INV6 U2216 ( .A(u_alu_ashr_4_A_6_), .Q(n2693) );
  INV3 U2217 ( .A(n1236), .Q(n895) );
  NAND22 U2218 ( .A(n1193), .B(n177), .Q(n1130) );
  NAND22 U2219 ( .A(n688), .B(n169), .Q(n517) );
  NAND22 U2220 ( .A(n2341), .B(n264), .Q(n2391) );
  NAND21 U2221 ( .A(n1338), .B(n1367), .Q(n1703) );
  NAND22 U2222 ( .A(n383), .B(n2097), .Q(n2098) );
  NOR22 U2223 ( .A(u_alu_DP_OP_85J3_126_1427_n374), .B(n343), .Q(n2783) );
  NAND21 U2224 ( .A(n2369), .B(n2330), .Q(n1983) );
  NAND22 U2225 ( .A(n193), .B(n172), .Q(n2296) );
  NAND22 U2226 ( .A(n2031), .B(n653), .Q(n2032) );
  INV2 U2227 ( .A(u_alu_DP_OP_83J3_124_3384_n29), .Q(
        u_alu_DP_OP_83J3_124_3384_n119) );
  NAND22 U2228 ( .A(n1044), .B(n175), .Q(n841) );
  INV2 U2229 ( .A(u_alu_DP_OP_83J3_124_3384_n15), .Q(
        u_alu_DP_OP_83J3_124_3384_n117) );
  NAND22 U2230 ( .A(n530), .B(n289), .Q(n2037) );
  AOI221 U2231 ( .A(u_alu_ashr_4_A_6_), .B(n2564), .C(n2866), .D(n245), .Q(
        n2566) );
  NAND22 U2232 ( .A(n2204), .B(n200), .Q(n1232) );
  NAND21 U2233 ( .A(n1272), .B(n2392), .Q(n2179) );
  NOR22 U2234 ( .A(n2089), .B(n1823), .Q(n1839) );
  NOR21 U2235 ( .A(n2096), .B(n2100), .Q(n2067) );
  INV2 U2236 ( .A(u_alu_DP_OP_83J3_124_3384_n32), .Q(
        u_alu_DP_OP_83J3_124_3384_n120) );
  NOR21 U2237 ( .A(n161), .B(n1970), .Q(n2008) );
  INV3 U2238 ( .A(n654), .Q(n653) );
  NAND22 U2239 ( .A(n2295), .B(n1052), .Q(n1054) );
  NOR22 U2240 ( .A(n1362), .B(n2689), .Q(n355) );
  NAND22 U2241 ( .A(n858), .B(n857), .Q(n856) );
  BUF12 U2242 ( .A(u_alu_DP_OP_83J3_124_3384_n152), .Q(n1338) );
  NAND24 U2243 ( .A(u_alu_ashr_4_A_17_), .B(n993), .Q(
        u_alu_DP_OP_83J3_124_3384_n53) );
  INV2 U2244 ( .A(u_alu_DP_OP_83J3_124_3384_n52), .Q(
        u_alu_DP_OP_83J3_124_3384_n123) );
  NOR21 U2245 ( .A(n2516), .B(u_alu_ashr_4_A_17_), .Q(u_alu_lt_x_11_n59) );
  NAND21 U2246 ( .A(n1830), .B(n2830), .Q(n341) );
  INV3 U2247 ( .A(n1235), .Q(n896) );
  NAND21 U2248 ( .A(alu_i_data_B[19]), .B(n175), .Q(n926) );
  INV3 U2249 ( .A(n1923), .Q(n359) );
  NOR21 U2250 ( .A(u_alu_lt_x_11_n139), .B(alu_i_data_B[19]), .Q(
        u_alu_lt_x_11_n53) );
  NAND22 U2251 ( .A(n1234), .B(compare_i_data_rs[2]), .Q(n1825) );
  NAND21 U2252 ( .A(alu_i_data_B[20]), .B(n1363), .Q(n1124) );
  INV2 U2253 ( .A(n163), .Q(n964) );
  NAND22 U2254 ( .A(u_alu_lt_x_11_B_1_), .B(n765), .Q(n764) );
  NAND23 U2255 ( .A(n2967), .B(n183), .Q(u_alu_lt_x_11_B_29_) );
  NAND22 U2256 ( .A(n195), .B(n123), .Q(n1195) );
  NAND22 U2257 ( .A(n2193), .B(n2062), .Q(n776) );
  NAND22 U2258 ( .A(n2406), .B(n2404), .Q(n730) );
  NAND21 U2259 ( .A(alu_i_data_B[20]), .B(n175), .Q(n978) );
  AOI212 U2260 ( .A(n1998), .B(n1997), .C(n1306), .Q(n576) );
  NAND22 U2261 ( .A(u_alu_ashr_4_A_16_), .B(n248), .Q(n270) );
  NAND22 U2262 ( .A(n567), .B(n2340), .Q(n265) );
  INV2 U2263 ( .A(n123), .Q(n2824) );
  NAND21 U2264 ( .A(n163), .B(n177), .Q(n1690) );
  OAI312 U2265 ( .A(i_con_bop[2]), .B(n1717), .C(n1410), .D(n1409), .Q(n1558)
         );
  NOR21 U2266 ( .A(n2808), .B(u_alu_ashr_4_A_16_), .Q(u_alu_lt_x_11_n61) );
  NAND22 U2267 ( .A(n3076), .B(n1166), .Q(n582) );
  OAI221 U2268 ( .A(n1863), .B(n387), .C(n859), .D(n1864), .Q(n858) );
  NAND22 U2269 ( .A(n3076), .B(n1167), .Q(n584) );
  AOI211 U2270 ( .A(n2778), .B(n183), .C(n1422), .Q(n2779) );
  NAND22 U2271 ( .A(n2146), .B(n248), .Q(n956) );
  NOR22 U2272 ( .A(n197), .B(n2025), .Q(n1923) );
  BUF12 U2273 ( .A(n1337), .Q(n1336) );
  INV6 U2274 ( .A(n161), .Q(n1971) );
  XOR22 U2275 ( .A(u_alu_DP_OP_85J3_126_1427_n379), .B(n747), .Q(n321) );
  NAND32 U2276 ( .A(n1079), .B(n1080), .C(n1730), .Q(n1041) );
  NAND22 U2277 ( .A(n474), .B(n1353), .Q(n473) );
  NAND21 U2278 ( .A(n2807), .B(n2808), .Q(n805) );
  NAND22 U2279 ( .A(n706), .B(n705), .Q(n704) );
  INV2 U2280 ( .A(n1730), .Q(n1736) );
  NOR22 U2281 ( .A(n254), .B(compare_i_data_rs[7]), .Q(n253) );
  NOR33 U2282 ( .A(n2001), .B(n1999), .C(n1538), .Q(n3092) );
  INV3 U2283 ( .A(n60), .Q(n3084) );
  INV3 U2284 ( .A(n911), .Q(n3093) );
  NAND24 U2285 ( .A(n1655), .B(n1656), .Q(n2036) );
  INV12 U2286 ( .A(u_alu_lt_x_11_A_11_), .Q(n222) );
  NAND22 U2287 ( .A(n2545), .B(n2544), .Q(n1466) );
  NOR22 U2288 ( .A(n2800), .B(n2804), .Q(n647) );
  INV2 U2289 ( .A(n934), .Q(n1311) );
  NAND22 U2290 ( .A(n1612), .B(n2782), .Q(n1484) );
  NAND24 U2291 ( .A(n1603), .B(n1604), .Q(n747) );
  AOI211 U2292 ( .A(n183), .B(n170), .C(n2432), .Q(n391) );
  NOR23 U2293 ( .A(n1051), .B(n1050), .Q(n1049) );
  INV3 U2294 ( .A(n1244), .Q(n810) );
  NOR32 U2295 ( .A(n2186), .B(n1591), .C(n456), .Q(n1533) );
  NOR21 U2296 ( .A(n1784), .B(compare_i_data_rs[2]), .Q(n1786) );
  NOR23 U2297 ( .A(n430), .B(n944), .Q(n429) );
  NOR31 U2298 ( .A(n170), .B(n1999), .C(n2000), .Q(n2002) );
  INV3 U2299 ( .A(n366), .Q(n365) );
  INV12 U2300 ( .A(n198), .Q(n445) );
  INV3 U2301 ( .A(n508), .Q(n375) );
  INV3 U2302 ( .A(n2063), .Q(n276) );
  NAND31 U2303 ( .A(n1369), .B(n1312), .C(n2586), .Q(n2587) );
  INV3 U2304 ( .A(n1214), .Q(n570) );
  INV6 U2305 ( .A(compare_i_data_rs[4]), .Q(n227) );
  NAND33 U2306 ( .A(n2529), .B(n2528), .C(n2527), .Q(n2537) );
  NAND22 U2307 ( .A(n1527), .B(n1369), .Q(n374) );
  INV3 U2308 ( .A(n616), .Q(n615) );
  INV3 U2309 ( .A(n1638), .Q(n522) );
  NAND22 U2310 ( .A(n1574), .B(n1511), .Q(n958) );
  NAND22 U2311 ( .A(n1267), .B(n1464), .Q(n329) );
  NAND22 U2312 ( .A(n457), .B(n342), .Q(n456) );
  INV3 U2313 ( .A(n1454), .Q(n390) );
  NAND22 U2314 ( .A(n1487), .B(n1486), .Q(n1488) );
  NAND22 U2315 ( .A(n1088), .B(n1457), .Q(n303) );
  INV6 U2316 ( .A(n1474), .Q(n1475) );
  INV2 U2317 ( .A(n2003), .Q(n254) );
  NOR22 U2318 ( .A(i_data_FMalures[15]), .B(n116), .Q(n700) );
  NOR22 U2319 ( .A(n1404), .B(n116), .Q(n1373) );
  INV3 U2320 ( .A(n1349), .Q(n1086) );
  NOR22 U2321 ( .A(n1349), .B(n1407), .Q(n1371) );
  NOR22 U2322 ( .A(i_data_FEalures[30]), .B(n1350), .Q(n1543) );
  NAND22 U2323 ( .A(n1674), .B(n367), .Q(n366) );
  NAND22 U2324 ( .A(n1467), .B(n2527), .Q(n399) );
  INV3 U2325 ( .A(n1418), .Q(n650) );
  NAND22 U2326 ( .A(n90), .B(i_data_FMalures[20]), .Q(n1481) );
  AOI211 U2327 ( .A(n1335), .B(i_data_FEalures[0]), .C(n1459), .Q(n1570) );
  NAND21 U2328 ( .A(n89), .B(i_data_FMalures[18]), .Q(n1267) );
  INV3 U2329 ( .A(n2088), .Q(n236) );
  NAND21 U2330 ( .A(n1864), .B(n170), .Q(n2382) );
  NAND22 U2331 ( .A(n89), .B(i_data_FMalures[8]), .Q(n1461) );
  NOR22 U2332 ( .A(i_data_fbmemout[0]), .B(n1324), .Q(n1455) );
  NAND22 U2333 ( .A(n89), .B(i_data_FMalures[2]), .Q(n1376) );
  NOR21 U2334 ( .A(n1367), .B(n1356), .Q(n1136) );
  NAND22 U2335 ( .A(n90), .B(i_data_FMalures[5]), .Q(n1381) );
  NOR22 U2336 ( .A(i_data_fbmemout[23]), .B(n1324), .Q(n1413) );
  INV12 U2337 ( .A(n2966), .Q(n239) );
  INV6 U2338 ( .A(n1545), .Q(n1317) );
  INV3 U2339 ( .A(n1047), .Q(n651) );
  NAND22 U2340 ( .A(n1335), .B(i_data_FEalures[30]), .Q(n1571) );
  NOR23 U2341 ( .A(i_data_rt[4]), .B(n1218), .Q(n1445) );
  NAND33 U2342 ( .A(n943), .B(n981), .C(n364), .Q(n1675) );
  NAND22 U2343 ( .A(n1545), .B(i_data_famemout[25]), .Q(n1429) );
  INV3 U2344 ( .A(n905), .Q(n904) );
  NOR21 U2345 ( .A(n185), .B(n248), .Q(n765) );
  NAND24 U2346 ( .A(n170), .B(n166), .Q(n2404) );
  NOR21 U2347 ( .A(n1367), .B(n1358), .Q(n2917) );
  NAND22 U2348 ( .A(n1562), .B(n314), .Q(n313) );
  INV6 U2349 ( .A(n2089), .Q(n242) );
  NAND22 U2350 ( .A(n158), .B(i_data_rs[3]), .Q(n738) );
  NAND22 U2351 ( .A(n159), .B(i_data_rs[25]), .Q(n1210) );
  INV3 U2352 ( .A(n533), .Q(n532) );
  BUF15 U2353 ( .A(n1546), .Q(n1335) );
  INV15 U2354 ( .A(n1352), .Q(n246) );
  INV2 U2355 ( .A(n1680), .Q(n908) );
  INV3 U2356 ( .A(n315), .Q(n314) );
  NOR32 U2357 ( .A(n1665), .B(i_con_Ealuop[4]), .C(n1661), .Q(n1663) );
  NOR22 U2358 ( .A(n1365), .B(n1362), .Q(n2830) );
  INV2 U2359 ( .A(i_data_rt[7]), .Q(n1537) );
  INV6 U2360 ( .A(i_data_immext[2]), .Q(n1308) );
  INV2 U2361 ( .A(i_data_famemout[7]), .Q(n1384) );
  INV2 U2362 ( .A(i_data_rt[3]), .Q(n1547) );
  INV2 U2363 ( .A(i_data_rt[26]), .Q(n1506) );
  INV2 U2364 ( .A(i_data_rt[19]), .Q(n1468) );
  INV3 U2365 ( .A(i_data_rt[22]), .Q(n1419) );
  IMUX21 U2366 ( .A(i_addr_rt[2]), .B(i_data_immext[13]), .S(i_con_Eregdst), 
        .Q(n3101) );
  INV2 U2367 ( .A(i_data_FEalures[2]), .Q(n1262) );
  INV3 U2368 ( .A(i_data_fbmemout[28]), .Q(n791) );
  INV2 U2369 ( .A(i_data_fbmemout[8]), .Q(n1206) );
  INV2 U2370 ( .A(i_data_rt[28]), .Q(n1521) );
  INV2 U2371 ( .A(i_data_FMalures[8]), .Q(n569) );
  INV2 U2372 ( .A(i_data_FMalures[12]), .Q(n412) );
  INV2 U2373 ( .A(i_data_rt[8]), .Q(n1460) );
  INV2 U2374 ( .A(i_data_FMalures[31]), .Q(n1404) );
  INV2 U2375 ( .A(i_data_rt[15]), .Q(n1447) );
  INV2 U2376 ( .A(i_data_famemout[0]), .Q(n1458) );
  INV2 U2377 ( .A(i_data_rt[24]), .Q(n1428) );
  INV2 U2378 ( .A(i_data_fbmemout[6]), .Q(n1175) );
  INV1 U2379 ( .A(i_data_FMalures[6]), .Q(n1452) );
  INV2 U2380 ( .A(i_data_FEalures[4]), .Q(n1444) );
  INV2 U2381 ( .A(i_data_immext[4]), .Q(n1678) );
  INV2 U2382 ( .A(i_data_rt[0]), .Q(n1453) );
  INV2 U2383 ( .A(i_data_rs[31]), .Q(n1403) );
  BUF15 U2384 ( .A(n1534), .Q(n250) );
  INV2 U2385 ( .A(i_data_famemout[4]), .Q(n1389) );
  INV2 U2386 ( .A(i_data_rt[29]), .Q(n1526) );
  INV1 U2387 ( .A(i_data_FMalures[29]), .Q(n941) );
  INV2 U2388 ( .A(i_data_rt[5]), .Q(n1551) );
  INV3 U2389 ( .A(i_data_FEalures[5]), .Q(n1555) );
  INV1 U2390 ( .A(i_data_FMalures[30]), .Q(n940) );
  INV2 U2391 ( .A(i_con_bop[1]), .Q(n1410) );
  INV2 U2392 ( .A(i_data_fbmemout[5]), .Q(n1247) );
  IMUX21 U2393 ( .A(i_addr_rt[0]), .B(i_data_immext[11]), .S(i_con_Eregdst), 
        .Q(n3099) );
  NAND21 U2394 ( .A(i_con_bop[1]), .B(i_con_bop[2]), .Q(n315) );
  INV2 U2395 ( .A(i_data_rt[21]), .Q(n1489) );
  INV2 U2396 ( .A(i_data_rt[14]), .Q(n1441) );
  INV2 U2397 ( .A(i_data_famemout[14]), .Q(n1394) );
  INV2 U2398 ( .A(i_data_famemout[5]), .Q(n1379) );
  INV2 U2399 ( .A(i_data_rt[23]), .Q(n1002) );
  INV2 U2400 ( .A(i_data_famemout[2]), .Q(n1374) );
  IMUX21 U2401 ( .A(i_addr_rt[4]), .B(i_data_immext[15]), .S(i_con_Eregdst), 
        .Q(n3102) );
  NAND21 U2402 ( .A(i_con_bop[0]), .B(i_con_bop[2]), .Q(n1412) );
  INV2 U2403 ( .A(i_data_rt[16]), .Q(n1495) );
  IMUX21 U2404 ( .A(i_addr_rt[3]), .B(i_data_immext[14]), .S(i_con_Eregdst), 
        .Q(n1017) );
  INV1 U2405 ( .A(i_data_FMalures[22]), .Q(n1322) );
  INV2 U2406 ( .A(i_data_rt[30]), .Q(n1539) );
  IMUX21 U2407 ( .A(i_addr_rt[1]), .B(i_data_immext[12]), .S(i_con_Eregdst), 
        .Q(n3100) );
  NOR21 U2408 ( .A(n1949), .B(n1947), .Q(n417) );
  NAND33 U2409 ( .A(n1179), .B(n1178), .C(n1182), .Q(n1181) );
  XNR22 U2410 ( .A(n1052), .B(n915), .Q(n1283) );
  BUF6 U2411 ( .A(u_alu_lt_x_11_A_13_), .Q(n256) );
  AOI212 U2412 ( .A(n2721), .B(n1357), .C(n2717), .Q(n428) );
  NAND24 U2413 ( .A(n54), .B(n2481), .Q(n2467) );
  AOI212 U2414 ( .A(n168), .B(n2453), .C(n2452), .Q(n2502) );
  CLKIN8 U2415 ( .A(n1347), .Q(n1630) );
  NAND22 U2416 ( .A(n1468), .B(n1346), .Q(n2586) );
  XNR22 U2417 ( .A(n228), .B(n3072), .Q(n1282) );
  OAI222 U2418 ( .A(n2556), .B(n1360), .C(n2623), .D(n1358), .Q(n2603) );
  AOI212 U2419 ( .A(n1360), .B(n80), .C(n2700), .Q(n2710) );
  OAI2112 U2420 ( .A(n881), .B(n844), .C(n261), .D(n260), .Q(n3024) );
  AOI222 U2421 ( .A(n2717), .B(n1366), .C(n2762), .D(n2759), .Q(n2723) );
  NOR22 U2422 ( .A(n163), .B(n2403), .Q(n2414) );
  NAND22 U2423 ( .A(n2626), .B(n262), .Q(n2634) );
  OAI222 U2424 ( .A(n1356), .B(n2907), .C(n266), .D(n154), .Q(n1325) );
  AOI212 U2425 ( .A(n2873), .B(n1358), .C(n2872), .Q(n2907) );
  AOI212 U2426 ( .A(n2261), .B(n2415), .C(n2260), .Q(n2262) );
  OAI212 U2427 ( .A(n365), .B(n1315), .C(n1683), .Q(n1664) );
  AOI221 U2428 ( .A(n1989), .B(n1358), .C(n2118), .D(n1360), .Q(n2061) );
  NOR33 U2429 ( .A(n199), .B(n1493), .C(n1492), .Q(n1191) );
  NOR24 U2430 ( .A(n2800), .B(n2804), .Q(n1623) );
  NOR31 U2431 ( .A(n1358), .B(n3066), .C(n1896), .Q(n277) );
  OAI312 U2432 ( .A(n229), .B(n1477), .C(n62), .D(n484), .Q(n759) );
  AOI212 U2433 ( .A(n2721), .B(n1356), .C(n1933), .Q(n2699) );
  INV6 U2434 ( .A(n2586), .Q(n2588) );
  NOR23 U2435 ( .A(i_data_FEalures[13]), .B(n1349), .Q(n1471) );
  BUF6 U2436 ( .A(u_alu_lt_x_11_A_0_), .Q(n289) );
  NAND24 U2437 ( .A(n431), .B(n429), .Q(n1169) );
  NAND22 U2438 ( .A(n1506), .B(n1346), .Q(n294) );
  NOR22 U2439 ( .A(n1364), .B(n1366), .Q(n2433) );
  NOR22 U2440 ( .A(u_alu_lt_x_11_B_11_), .B(n222), .Q(u_alu_lt_x_11_n84) );
  NOR22 U2441 ( .A(i_data_FEalures[22]), .B(n1349), .Q(n1051) );
  AOI222 U2442 ( .A(n3023), .B(n2917), .C(n2955), .D(n3021), .Q(n687) );
  NAND22 U2443 ( .A(n2510), .B(n301), .Q(n2512) );
  AOI221 U2444 ( .A(n177), .B(n1044), .C(n193), .D(n1366), .Q(n1685) );
  NAND22 U2445 ( .A(n308), .B(n307), .Q(alu_o_data_AluRes[29]) );
  AOI212 U2446 ( .A(u_alu_pre_sum_4a[5]), .B(n536), .C(n842), .Q(n307) );
  AOI222 U2447 ( .A(n1021), .B(n845), .C(n2991), .D(n1345), .Q(n308) );
  IMUX21 U2448 ( .A(n2876), .B(n2877), .S(n1509), .Q(n2878) );
  AOI222 U2449 ( .A(n203), .B(n2612), .C(n178), .D(n2542), .Q(n954) );
  AOI212 U2450 ( .A(u_alu_lt_x_11_A_3_), .B(n1830), .C(n2388), .Q(n2389) );
  NOR23 U2451 ( .A(i_data_FEalures[11]), .B(n1349), .Q(n1628) );
  NOR24 U2452 ( .A(i_data_FEalures[17]), .B(n1350), .Q(n2531) );
  INV3 U2453 ( .A(n310), .Q(n1880) );
  NAND22 U2454 ( .A(n2947), .B(n171), .Q(n310) );
  OAI222 U2455 ( .A(n968), .B(n311), .C(n2667), .D(n1318), .Q(n2668) );
  AOI212 U2456 ( .A(n2534), .B(n2535), .C(n239), .Q(n2536) );
  OAI312 U2457 ( .A(n2349), .B(n2348), .C(n2347), .D(n2346), .Q(n2350) );
  NAND22 U2458 ( .A(n207), .B(n2069), .Q(n1129) );
  AOI212 U2459 ( .A(n793), .B(n2421), .C(n2420), .Q(n2426) );
  NAND28 U2460 ( .A(n623), .B(n622), .Q(n1318) );
  AOI222 U2461 ( .A(i_data_FEalures[10]), .B(n1335), .C(n1319), .D(
        i_data_famemout[10]), .Q(n317) );
  NAND22 U2462 ( .A(n1245), .B(n318), .Q(n1244) );
  NAND28 U2463 ( .A(n324), .B(n1429), .Q(u_alu_DP_OP_85J3_126_1427_n379) );
  XNR22 U2464 ( .A(n2705), .B(n325), .Q(n542) );
  AOI212 U2465 ( .A(n2704), .B(n72), .C(n2706), .Q(n325) );
  AOI212 U2466 ( .A(n2550), .B(n2543), .C(n2810), .Q(n2632) );
  NAND28 U2467 ( .A(n326), .B(n179), .Q(n829) );
  XOR22 U2468 ( .A(u_alu_lt_x_11_n122), .B(n912), .Q(n336) );
  XNR22 U2469 ( .A(n3087), .B(n1533), .Q(n339) );
  OAI2112 U2470 ( .A(n185), .B(n956), .C(n341), .D(n340), .Q(n2209) );
  AOI222 U2471 ( .A(n1778), .B(n1356), .C(n1777), .D(n1357), .Q(n2567) );
  NAND33 U2472 ( .A(n2393), .B(n2392), .C(n2391), .Q(n2399) );
  INV15 U2473 ( .A(n1347), .Q(n1346) );
  NAND33 U2474 ( .A(n2191), .B(n2190), .C(n2189), .Q(n2415) );
  AOI212 U2475 ( .A(n343), .B(n183), .C(n1318), .Q(n2702) );
  AOI222 U2476 ( .A(n1883), .B(n1360), .C(n1810), .D(n1358), .Q(n1846) );
  OAI222 U2477 ( .A(n1710), .B(n245), .C(n1709), .D(n166), .Q(n1748) );
  AOI212 U2478 ( .A(n1808), .B(n176), .C(n1807), .Q(n1941) );
  OAI222 U2479 ( .A(n2873), .B(n1358), .C(n355), .D(n350), .Q(n2837) );
  NAND28 U2480 ( .A(n1599), .B(n1353), .Q(alu_i_data_B[27]) );
  OAI2112 U2481 ( .A(n2478), .B(n2477), .C(n362), .D(n360), .Q(n2491) );
  NAND28 U2482 ( .A(n2405), .B(n2404), .Q(u_alu_ashr_4_A_9_) );
  NOR24 U2483 ( .A(n1115), .B(n1437), .Q(n1593) );
  XNR22 U2484 ( .A(n368), .B(n1417), .Q(n1424) );
  NAND33 U2485 ( .A(n375), .B(n1527), .C(n370), .Q(n369) );
  NAND24 U2486 ( .A(n445), .B(n941), .Q(n372) );
  OAI212 U2487 ( .A(n213), .B(n2181), .C(n383), .Q(n2133) );
  NOR24 U2488 ( .A(n388), .B(n1863), .Q(n3098) );
  AOI222 U2489 ( .A(n1356), .B(n2508), .C(n2557), .D(n249), .Q(n951) );
  OAI222 U2490 ( .A(n2435), .B(n1360), .C(n2556), .D(n1358), .Q(n2508) );
  AOI222 U2491 ( .A(n2433), .B(n2754), .C(n392), .D(n391), .Q(n2622) );
  NAND22 U2492 ( .A(n2225), .B(n166), .Q(n397) );
  AOI212 U2493 ( .A(u_alu_DP_OP_83J3_124_3384_n51), .B(
        u_alu_DP_OP_83J3_124_3384_n101), .C(u_alu_DP_OP_83J3_124_3384_n102), 
        .Q(u_alu_DP_OP_83J3_124_3384_n1) );
  OAI212 U2494 ( .A(u_alu_DP_OP_83J3_124_3384_n41), .B(
        u_alu_DP_OP_83J3_124_3384_n45), .C(u_alu_DP_OP_83J3_124_3384_n42), .Q(
        u_alu_DP_OP_83J3_124_3384_n102) );
  OAI212 U2495 ( .A(u_alu_DP_OP_83J3_124_3384_n55), .B(
        u_alu_DP_OP_83J3_124_3384_n52), .C(u_alu_DP_OP_83J3_124_3384_n53), .Q(
        u_alu_DP_OP_83J3_124_3384_n51) );
  AOI212 U2496 ( .A(u_alu_DP_OP_84J3_125_2615_n109), .B(
        u_alu_DP_OP_84J3_125_2615_n86), .C(u_alu_DP_OP_84J3_125_2615_n77), .Q(
        u_alu_DP_OP_84J3_125_2615_n18) );
  OAI222 U2497 ( .A(n2905), .B(n1361), .C(n2089), .D(n211), .Q(n2836) );
  NAND33 U2498 ( .A(n421), .B(n418), .C(n414), .Q(alu_o_data_AluRes[6]) );
  AOI2112 U2499 ( .A(n416), .B(n415), .C(n1931), .D(n1930), .Q(n414) );
  AOI222 U2500 ( .A(n179), .B(n419), .C(n1938), .D(n2883), .Q(n418) );
  OAI212 U2501 ( .A(n2007), .B(n2006), .C(n2010), .Q(n420) );
  OAI212 U2502 ( .A(n1356), .B(n1945), .C(n423), .Q(n422) );
  AOI222 U2503 ( .A(n2843), .B(n2075), .C(n427), .D(n203), .Q(n426) );
  AOI222 U2504 ( .A(i_data_FEalures[19]), .B(n1334), .C(n1545), .D(
        i_data_famemout[19]), .Q(n432) );
  XNR22 U2505 ( .A(n223), .B(n3096), .Q(n434) );
  OAI212 U2506 ( .A(n1360), .B(n1749), .C(n439), .Q(n1774) );
  AOI222 U2507 ( .A(n1809), .B(n1362), .C(n440), .D(n200), .Q(n1749) );
  OAI212 U2508 ( .A(n1363), .B(n1772), .C(n1771), .Q(n1845) );
  OAI212 U2509 ( .A(u_alu_DP_OP_84J3_125_2615_n40), .B(
        u_alu_DP_OP_84J3_125_2615_n36), .C(u_alu_DP_OP_84J3_125_2615_n37), .Q(
        u_alu_DP_OP_84J3_125_2615_n92) );
  NAND22 U2510 ( .A(n445), .B(n942), .Q(n467) );
  NAND33 U2511 ( .A(n1072), .B(n1073), .C(n1071), .Q(compare_i_data_rs[4]) );
  AOI2112 U2512 ( .A(n1156), .B(n454), .C(n449), .D(n446), .Q(n1164) );
  XNR22 U2513 ( .A(n233), .B(n3085), .Q(n446) );
  NOR24 U2514 ( .A(n448), .B(n447), .Q(n3085) );
  XOR22 U2515 ( .A(n453), .B(n3090), .Q(n449) );
  OAI212 U2516 ( .A(i_data_rt[9]), .B(n1348), .C(n1120), .Q(n452) );
  OAI212 U2517 ( .A(n1159), .B(n1859), .C(n227), .Q(n454) );
  AOI212 U2518 ( .A(n237), .B(n1444), .C(n1443), .Q(n1647) );
  OAI212 U2519 ( .A(n2142), .B(n2143), .C(n459), .Q(n458) );
  AOI2112 U2520 ( .A(n471), .B(n179), .C(n468), .D(n1834), .Q(n1835) );
  AOI211 U2521 ( .A(n1832), .B(n2458), .C(n2460), .Q(n472) );
  NAND33 U2522 ( .A(n1187), .B(n1189), .C(n473), .Q(n1190) );
  NOR24 U2523 ( .A(n1114), .B(n1112), .Q(n1606) );
  XNR22 U2524 ( .A(n708), .B(n566), .Q(n1067) );
  IMUX21 U2525 ( .A(n2324), .B(n2325), .S(n568), .Q(n2326) );
  NAND22 U2526 ( .A(n219), .B(n231), .Q(n2165) );
  NAND33 U2527 ( .A(n496), .B(n2980), .C(n492), .Q(n488) );
  XNR22 U2528 ( .A(n210), .B(n500), .Q(n491) );
  AOI222 U2529 ( .A(n2982), .B(n494), .C(n167), .D(n635), .Q(n493) );
  OAI212 U2530 ( .A(n1310), .B(n2971), .C(n2970), .Q(n500) );
  NAND28 U2531 ( .A(n604), .B(n183), .Q(n688) );
  NAND22 U2532 ( .A(n2415), .B(n501), .Q(n2308) );
  AOI212 U2533 ( .A(n2042), .B(n505), .C(n995), .Q(n502) );
  AOI212 U2534 ( .A(n2040), .B(n227), .C(n2039), .Q(n503) );
  OAI212 U2535 ( .A(n2202), .B(n2037), .C(n2384), .Q(n506) );
  NOR24 U2536 ( .A(n1167), .B(n1166), .Q(n1189) );
  AOI212 U2537 ( .A(n512), .B(n1683), .C(n1682), .Q(n511) );
  OAI212 U2538 ( .A(n2202), .B(n175), .C(n2203), .Q(n515) );
  NAND22 U2539 ( .A(u_alu_DP_OP_83J3_124_3384_n152), .B(n175), .Q(n516) );
  NAND24 U2540 ( .A(n521), .B(n2339), .Q(n708) );
  OAI222 U2541 ( .A(n1885), .B(n1356), .C(n1846), .D(n249), .Q(n523) );
  XNR22 U2542 ( .A(n3097), .B(u_alu_lt_x_11_n121), .Q(n809) );
  AOI312 U2543 ( .A(i_con_Ealuop[1]), .B(n532), .C(n531), .D(n1665), .Q(n1725)
         );
  AOI312 U2544 ( .A(n1356), .B(n2569), .C(n2568), .D(n171), .Q(n534) );
  OAI222 U2545 ( .A(n2727), .B(n1358), .C(n2658), .D(n1360), .Q(n2692) );
  NAND22 U2546 ( .A(n543), .B(n540), .Q(n539) );
  NAND28 U2547 ( .A(n974), .B(n179), .Q(n1222) );
  AOI2111 U2548 ( .A(n1102), .B(n1103), .C(n545), .D(n544), .Q(n543) );
  OAI221 U2549 ( .A(n1101), .B(n255), .C(n2693), .D(n2976), .Q(n544) );
  AOI311 U2550 ( .A(n180), .B(n1100), .C(n1098), .D(n1143), .Q(n545) );
  NOR23 U2551 ( .A(i_con_Efamux[0]), .B(n546), .Q(n1546) );
  NOR24 U2552 ( .A(n2589), .B(n547), .Q(n1614) );
  NOR31 U2553 ( .A(n170), .B(n2588), .C(n547), .Q(n2592) );
  NOR22 U2554 ( .A(n1348), .B(i_data_rt[10]), .Q(n550) );
  AOI312 U2555 ( .A(n1227), .B(n558), .C(n556), .D(n3066), .Q(n555) );
  AOI212 U2556 ( .A(n577), .B(n2465), .C(n575), .Q(n2472) );
  NAND33 U2557 ( .A(n583), .B(n584), .C(n582), .Q(n581) );
  NAND24 U2558 ( .A(n1605), .B(n1606), .Q(n580) );
  XOR22 U2559 ( .A(n1466), .B(n913), .Q(n1480) );
  NAND33 U2560 ( .A(n598), .B(n590), .C(n589), .Q(alu_o_data_AluRes[23]) );
  AOI2112 U2561 ( .A(n2714), .B(n595), .C(n593), .D(n591), .Q(n590) );
  OAI212 U2562 ( .A(n1222), .B(n2753), .C(n592), .Q(n591) );
  OAI212 U2563 ( .A(n596), .B(n3066), .C(n594), .Q(n593) );
  NAND22 U2564 ( .A(n2752), .B(n1345), .Q(n598) );
  NOR24 U2565 ( .A(n1266), .B(n1069), .Q(n602) );
  NAND28 U2566 ( .A(n603), .B(n602), .Q(n2629) );
  AOI222 U2567 ( .A(n1358), .B(n611), .C(n2507), .D(n1360), .Q(n2437) );
  OAI312 U2568 ( .A(u_alu_lt_x_11_n99), .B(n161), .C(n1970), .D(n612), .Q(
        n2455) );
  OAI212 U2569 ( .A(n2010), .B(n2011), .C(n2455), .Q(n2053) );
  AOI212 U2570 ( .A(n1936), .B(n2462), .C(u_alu_lt_x_11_n105), .Q(n2010) );
  NAND28 U2571 ( .A(n1968), .B(n2003), .Q(n2146) );
  NAND28 U2572 ( .A(n619), .B(n186), .Q(n3043) );
  OAI221 U2573 ( .A(n1708), .B(n185), .C(n1747), .D(n176), .Q(n627) );
  AOI212 U2574 ( .A(n2367), .B(n2366), .C(n628), .Q(n2374) );
  AOI212 U2575 ( .A(n2483), .B(u_alu_lt_x_11_n77), .C(n2482), .Q(n2364) );
  OAI312 U2576 ( .A(n2218), .B(n1356), .C(n2219), .D(n247), .Q(n634) );
  AOI212 U2577 ( .A(u_alu_DP_OP_84J3_125_2615_n16), .B(
        u_alu_DP_OP_84J3_125_2615_n108), .C(u_alu_DP_OP_84J3_125_2615_n70), 
        .Q(n1024) );
  AOI222 U2578 ( .A(n1358), .B(n2724), .C(n2677), .D(n1360), .Q(n2678) );
  NAND22 U2579 ( .A(n2411), .B(n640), .Q(n646) );
  NAND22 U2580 ( .A(n2406), .B(n641), .Q(n640) );
  NAND22 U2581 ( .A(n643), .B(n642), .Q(n963) );
  NAND28 U2582 ( .A(n1261), .B(n2062), .Q(n2204) );
  NOR23 U2583 ( .A(i_data_fbmemout[16]), .B(n246), .Q(n2800) );
  NOR24 U2584 ( .A(n651), .B(n650), .Q(n1584) );
  AOI212 U2585 ( .A(n2004), .B(n2003), .C(n161), .Q(n2005) );
  NAND24 U2586 ( .A(n237), .B(n1450), .Q(n1995) );
  AOI220 U2587 ( .A(n688), .B(n1366), .C(n172), .D(n1234), .Q(n1698) );
  NAND33 U2588 ( .A(n2446), .B(n2445), .C(n661), .Q(n2574) );
  OAI211 U2589 ( .A(n2270), .B(n2417), .C(n662), .Q(n663) );
  NOR33 U2590 ( .A(n1475), .B(n199), .C(n1472), .Q(n666) );
  NAND33 U2591 ( .A(n3026), .B(n3028), .C(n3027), .Q(alu_o_data_AluRes[30]) );
  OAI212 U2592 ( .A(n2834), .B(n2701), .C(n2636), .Q(n678) );
  AOI222 U2593 ( .A(n171), .B(n205), .C(n673), .D(n177), .Q(n2701) );
  OAI212 U2594 ( .A(n1797), .B(n1796), .C(n1795), .Q(n1832) );
  AOI212 U2595 ( .A(i_data_famemout[3]), .B(n1319), .C(n736), .Q(n680) );
  NOR24 U2596 ( .A(n2028), .B(n2027), .Q(n2030) );
  NAND33 U2597 ( .A(n76), .B(n1370), .C(n1993), .Q(n682) );
  AOI212 U2598 ( .A(n684), .B(n183), .C(u_alu_DP_OP_85J3_126_1427_n374), .Q(
        n2703) );
  OAI222 U2599 ( .A(n2172), .B(n175), .C(n1363), .D(n1988), .Q(n2118) );
  AOI222 U2600 ( .A(alu_i_data_B[19]), .B(n2433), .C(n1842), .D(n245), .Q(
        n1988) );
  AOI212 U2601 ( .A(n1987), .B(n245), .C(n1986), .Q(n2172) );
  OAI212 U2602 ( .A(n1363), .B(n2117), .C(n2116), .Q(n2173) );
  AOI212 U2603 ( .A(n1912), .B(n166), .C(n1911), .Q(n2117) );
  NAND43 U2604 ( .A(n1520), .B(n1518), .C(n1573), .D(n1519), .Q(n1524) );
  NOR24 U2605 ( .A(n1561), .B(n1560), .Q(n693) );
  NOR33 U2606 ( .A(n156), .B(n697), .C(n1034), .Q(n696) );
  NAND28 U2607 ( .A(n699), .B(n698), .Q(o_con_ifbranch) );
  NAND24 U2608 ( .A(n760), .B(n1470), .Q(u_alu_lt_x_11_A_13_) );
  AOI212 U2609 ( .A(n168), .B(n714), .C(n710), .Q(n2079) );
  OAI212 U2610 ( .A(n1343), .B(n1129), .C(n711), .Q(n710) );
  AOI222 U2611 ( .A(u_alu_DP_OP_83J3_124_3384_n153), .B(n1361), .C(n169), .D(
        alu_i_data_B[19]), .Q(n3060) );
  AOI212 U2612 ( .A(n2931), .B(n2932), .C(n2930), .Q(n722) );
  AOI222 U2613 ( .A(n1356), .B(n2987), .C(n2951), .D(n1357), .Q(n3022) );
  OAI212 U2614 ( .A(n2029), .B(n734), .C(n733), .Q(n2034) );
  AOI212 U2615 ( .A(n248), .B(n2555), .C(n740), .Q(n2435) );
  IMUX21 U2616 ( .A(n1953), .B(n741), .S(n1952), .Q(n1956) );
  NOR23 U2617 ( .A(n742), .B(n2039), .Q(n1953) );
  AOI212 U2618 ( .A(n1844), .B(n1363), .C(n750), .Q(n1773) );
  OAI212 U2619 ( .A(n754), .B(n1987), .C(n185), .Q(n753) );
  NAND20 U2620 ( .A(u_alu_lt_x_11_B_11_), .B(n1361), .Q(n955) );
  AOI222 U2621 ( .A(n90), .B(i_data_FMalures[13]), .C(n158), .D(i_data_rs[13]), 
        .Q(n760) );
  XNR22 U2622 ( .A(n2014), .B(n2361), .Q(n763) );
  NAND28 U2623 ( .A(n2036), .B(n2035), .Q(u_alu_lt_x_11_B_1_) );
  AOI222 U2624 ( .A(n2331), .B(n1363), .C(n2153), .D(n1361), .Q(n2231) );
  AOI212 U2625 ( .A(n1844), .B(n200), .C(n1843), .Q(n1916) );
  NOR22 U2626 ( .A(n776), .B(n2094), .Q(n2095) );
  NAND22 U2627 ( .A(n2393), .B(n2395), .Q(n2348) );
  XNR22 U2628 ( .A(u_alu_lt_x_11_A_0_), .B(n782), .Q(n1161) );
  AOI212 U2629 ( .A(n2749), .B(n2663), .C(u_alu_lt_x_11_n47), .Q(n2654) );
  OAI212 U2630 ( .A(n2650), .B(n2649), .C(n2812), .Q(n2749) );
  AOI212 U2631 ( .A(n801), .B(n800), .C(n795), .Q(n3068) );
  OAI312 U2632 ( .A(n3006), .B(n798), .C(n154), .D(n3054), .Q(n797) );
  NAND33 U2633 ( .A(n1137), .B(n1060), .C(n1059), .Q(n800) );
  AOI212 U2634 ( .A(n604), .B(n183), .C(n2629), .Q(n803) );
  INV6 U2635 ( .A(n812), .Q(n811) );
  AOI2112 U2636 ( .A(n3022), .B(n2955), .C(n821), .D(n818), .Q(n2956) );
  OAI312 U2637 ( .A(n110), .B(n177), .C(n3023), .D(n167), .Q(n818) );
  NAND22 U2638 ( .A(n2209), .B(n1357), .Q(n819) );
  OAI212 U2639 ( .A(n2218), .B(n2219), .C(n1356), .Q(n820) );
  AOI212 U2640 ( .A(n3043), .B(n3031), .C(n3033), .Q(n2935) );
  AOI222 U2641 ( .A(n2330), .B(u_alu_DP_OP_83J3_124_3384_n152), .C(n81), .D(
        n166), .Q(n909) );
  AOI222 U2642 ( .A(n2334), .B(n1357), .C(n2300), .D(n1356), .Q(n834) );
  OAI222 U2643 ( .A(n2231), .B(n110), .C(n1358), .D(n2333), .Q(n2300) );
  AOI312 U2644 ( .A(n207), .B(n838), .C(n1032), .D(n835), .Q(n1031) );
  NOR24 U2645 ( .A(n1026), .B(n1025), .Q(n1021) );
  NOR24 U2646 ( .A(n853), .B(n1408), .Q(u_alu_lt_x_11_A_31_) );
  OAI212 U2647 ( .A(i_data_famemout[31]), .B(n55), .C(n854), .Q(n853) );
  AOI212 U2648 ( .A(u_alu_DP_OP_83J3_124_3384_n113), .B(
        u_alu_DP_OP_83J3_124_3384_n101), .C(u_alu_DP_OP_83J3_124_3384_n102), 
        .Q(u_alu_DP_OP_83J3_124_3384_n64) );
  NOR24 U2649 ( .A(n2594), .B(alu_i_data_B[19]), .Q(
        u_alu_DP_OP_83J3_124_3384_n41) );
  AOI212 U2650 ( .A(n2555), .B(n175), .C(n2554), .Q(n2623) );
  AOI221 U2651 ( .A(n3053), .B(n1070), .C(n3010), .D(n1280), .Q(n891) );
  NAND28 U2652 ( .A(n1040), .B(n1039), .Q(n1303) );
  OAI212 U2653 ( .A(n175), .B(n181), .C(n1126), .Q(n906) );
  OAI222 U2654 ( .A(n2906), .B(n1360), .C(n2905), .D(n907), .Q(n2939) );
  OAI222 U2655 ( .A(n1360), .B(n2938), .C(n3003), .D(n1358), .Q(n2978) );
  OAI221 U2656 ( .A(n3012), .B(n248), .C(n1143), .D(n175), .Q(n2867) );
  NAND22 U2657 ( .A(n2456), .B(n2455), .Q(n2473) );
  NOR22 U2658 ( .A(u_alu_lt_x_11_n9), .B(n3034), .Q(u_alu_lt_x_11_n7) );
  NAND33 U2659 ( .A(n2084), .B(n2124), .C(n2083), .Q(n2085) );
  AOI212 U2660 ( .A(n1172), .B(n1171), .C(n1173), .Q(n2125) );
  IMUX21 U2661 ( .A(n2773), .B(n2774), .S(u_alu_lt_x_11_n144), .Q(n2775) );
  INV6 U2662 ( .A(n1668), .Q(n1039) );
  INV3 U2663 ( .A(n3068), .Q(n1019) );
  AOI222 U2664 ( .A(n1545), .B(i_data_famemout[13]), .C(n1335), .D(
        i_data_FEalures[13]), .Q(n1470) );
  AOI212 U2665 ( .A(n2361), .B(n2081), .C(n520), .Q(n2054) );
  AOI212 U2666 ( .A(n1335), .B(i_data_FEalures[7]), .C(n1385), .Q(n1388) );
  NAND22 U2667 ( .A(n2002), .B(n1642), .Q(n2004) );
  NOR22 U2668 ( .A(n1362), .B(n2030), .Q(n1932) );
  AOI212 U2669 ( .A(n2812), .B(n2797), .C(n2811), .Q(n2798) );
  NAND22 U2670 ( .A(n90), .B(i_data_FMalures[3]), .Q(n1544) );
  NOR24 U2671 ( .A(n1340), .B(n2821), .Q(n2715) );
  AOI2112 U2672 ( .A(n2759), .B(n2605), .C(n2571), .D(n2570), .Q(n2637) );
  AOI212 U2673 ( .A(n2389), .B(n2390), .C(n995), .Q(n2401) );
  XNR22 U2674 ( .A(n1422), .B(n1421), .Q(n1423) );
  NOR22 U2675 ( .A(alu_i_data_B[27]), .B(n196), .Q(n2930) );
  IMUX21 U2676 ( .A(n2902), .B(n2901), .S(n196), .Q(n2903) );
  NOR21 U2677 ( .A(n1340), .B(n2821), .Q(n1146) );
  NAND28 U2678 ( .A(n1196), .B(n1307), .Q(u_alu_DP_OP_83J3_124_3384_n153) );
  AOI212 U2679 ( .A(n48), .B(n1514), .C(n1513), .Q(n1598) );
  NOR23 U2680 ( .A(n184), .B(n219), .Q(n2140) );
  NOR32 U2681 ( .A(n239), .B(n2784), .C(n2783), .Q(n2789) );
  NOR22 U2682 ( .A(n233), .B(n2563), .Q(n2423) );
  NAND24 U2683 ( .A(n2081), .B(n2164), .Q(n2470) );
  AOI212 U2684 ( .A(n2821), .B(u_alu_pre_sum_3b[8]), .C(n1340), .Q(n1207) );
  XNR22 U2685 ( .A(u_alu_pre_sum_4a[0]), .B(u_alu_pre_sum_3b[8]), .Q(n2820) );
  NOR24 U2686 ( .A(n195), .B(n123), .Q(n2929) );
  NAND24 U2687 ( .A(n123), .B(n195), .Q(n2857) );
  OAI212 U2688 ( .A(n641), .B(n2407), .C(n2406), .Q(n2412) );
  NAND33 U2689 ( .A(n2123), .B(n2122), .C(n2121), .Q(alu_o_data_AluRes[10]) );
  NAND22 U2690 ( .A(n1875), .B(n207), .Q(n1270) );
  AOI212 U2691 ( .A(n3033), .B(n3030), .C(n3035), .Q(n3000) );
  AOI212 U2692 ( .A(u_alu_DP_OP_84J3_125_2615_n73), .B(
        u_alu_DP_OP_84J3_125_2615_n108), .C(u_alu_DP_OP_84J3_125_2615_n70), 
        .Q(n966) );
  AOI211 U2693 ( .A(n1954), .B(n1953), .C(n1340), .Q(n1955) );
  NOR22 U2694 ( .A(n2295), .B(n1052), .Q(n2995) );
  NOR31 U2695 ( .A(alu_i_data_B[19]), .B(n2594), .C(n3049), .Q(n2607) );
  NOR31 U2696 ( .A(u_alu_DP_OP_85J3_126_1427_n379), .B(u_alu_lt_x_11_B_25_), 
        .C(n3049), .Q(n2839) );
  OAI212 U2697 ( .A(n2946), .B(n2976), .C(n2945), .Q(n2957) );
  IMUX21 U2698 ( .A(n2944), .B(n2943), .S(n228), .Q(n2945) );
  AOI212 U2699 ( .A(n2781), .B(n2780), .C(n2779), .Q(n2796) );
  NAND33 U2700 ( .A(n2248), .B(n2247), .C(n2246), .Q(n2249) );
  NOR21 U2701 ( .A(n2460), .B(n220), .Q(n1798) );
  NOR24 U2702 ( .A(n1198), .B(n1197), .Q(n1052) );
  NOR41 U2703 ( .A(n1804), .B(n1803), .C(n1802), .D(n1801), .Q(n1805) );
  AOI212 U2704 ( .A(n1788), .B(n1787), .C(n1851), .Q(n1820) );
  NAND33 U2705 ( .A(n51), .B(n2132), .C(n2131), .Q(n2392) );
  OAI212 U2706 ( .A(n2254), .B(n2347), .C(n2270), .Q(n2255) );
  NOR22 U2707 ( .A(n1092), .B(n1328), .Q(n1329) );
  AOI212 U2708 ( .A(n1345), .B(n2922), .C(n2921), .Q(n2923) );
  NAND28 U2709 ( .A(n1613), .B(n1353), .Q(alu_i_data_B[20]) );
  NOR21 U2710 ( .A(n3005), .B(n3006), .Q(n3007) );
  NOR32 U2711 ( .A(n2251), .B(n2249), .C(n2250), .Q(n2268) );
  OAI212 U2712 ( .A(u_alu_DP_OP_83J3_124_3384_n23), .B(
        u_alu_DP_OP_83J3_124_3384_n15), .C(u_alu_DP_OP_83J3_124_3384_n16), .Q(
        u_alu_DP_OP_83J3_124_3384_n76) );
  NOR42 U2713 ( .A(n2291), .B(n2293), .C(n2292), .D(n1029), .Q(n1028) );
  NAND28 U2714 ( .A(n972), .B(n1089), .Q(n1342) );
  IMUX21 U2715 ( .A(n187), .B(n1342), .S(u_alu_DP_OP_85J3_126_1427_n377), .Q(
        n2733) );
  AOI211 U2716 ( .A(n2875), .B(n180), .C(n3012), .Q(n2880) );
  AOI212 U2717 ( .A(n2835), .B(n248), .C(n2657), .Q(n2727) );
  XNR22 U2718 ( .A(n2193), .B(n3091), .Q(n1066) );
  XNR22 U2719 ( .A(n1517), .B(n1569), .Q(n977) );
  NAND28 U2720 ( .A(n1616), .B(n1307), .Q(alu_i_data_B[19]) );
  INV6 U2721 ( .A(n1111), .Q(n1110) );
  XNR22 U2722 ( .A(n1509), .B(n1568), .Q(n976) );
  NOR24 U2723 ( .A(n1509), .B(n1336), .Q(u_alu_DP_OP_84J3_125_2615_n39) );
  NAND28 U2724 ( .A(n1505), .B(n1110), .Q(n1509) );
  NAND22 U2725 ( .A(n2144), .B(n1344), .Q(n1064) );
  AOI212 U2726 ( .A(n1361), .B(n1882), .C(n1881), .Q(n1944) );
  AOI212 U2727 ( .A(n1271), .B(n179), .C(n1268), .Q(n1876) );
  NOR32 U2728 ( .A(n2578), .B(n2576), .C(n2577), .Q(n2579) );
  NOR21 U2729 ( .A(n1364), .B(n3060), .Q(n3061) );
  OAI311 U2730 ( .A(n2805), .B(n2804), .C(n2803), .D(n183), .Q(n2807) );
  NAND34 U2731 ( .A(n1164), .B(n1163), .C(n1160), .Q(n1559) );
  NOR33 U2732 ( .A(n1627), .B(n1628), .C(n1440), .Q(n3088) );
  OAI212 U2733 ( .A(i_data_fbmemout[11]), .B(n246), .C(n63), .Q(n1440) );
  AOI211 U2734 ( .A(n1867), .B(n1866), .C(u_alu_lt_x_11_A_3_), .Q(n1868) );
  NAND33 U2735 ( .A(n1743), .B(n1745), .C(n1744), .Q(alu_o_data_AluRes[0]) );
  AOI212 U2736 ( .A(n168), .B(n1742), .C(n1741), .Q(n1743) );
  XNR22 U2737 ( .A(n2859), .B(n2858), .Q(n2888) );
  AOI211 U2738 ( .A(n3064), .B(n1136), .C(n1359), .Q(n1059) );
  NAND43 U2739 ( .A(n1170), .B(n1724), .C(n1168), .D(n1169), .Q(n1301) );
  NOR24 U2740 ( .A(n1663), .B(n1725), .Q(n1724) );
  AOI212 U2741 ( .A(n2592), .B(n2591), .C(n239), .Q(n2593) );
  NOR32 U2742 ( .A(n857), .B(n2202), .C(n1847), .Q(n1850) );
  INV3 U2743 ( .A(n2637), .Q(n1106) );
  NAND22 U2744 ( .A(i_con_Efamux[0]), .B(i_con_Efamux[1]), .Q(n1534) );
  NAND33 U2745 ( .A(n2159), .B(n2160), .C(n2158), .Q(alu_o_data_AluRes[11]) );
  NOR22 U2746 ( .A(i_data_fbmemout[25]), .B(n246), .Q(n1433) );
  NOR23 U2747 ( .A(i_con_Efamux[1]), .B(n1018), .Q(n2526) );
  OAI212 U2748 ( .A(n2977), .B(n2976), .C(n2975), .Q(n2990) );
  NAND22 U2749 ( .A(u_alu_ashr_4_A_17_), .B(n1363), .Q(n2674) );
  AOI212 U2750 ( .A(n2985), .B(n185), .C(n2984), .Q(n3017) );
  NOR32 U2751 ( .A(n2066), .B(n1311), .C(n2065), .Q(n2094) );
  NAND22 U2752 ( .A(n1414), .B(n1369), .Q(n999) );
  NAND33 U2753 ( .A(n961), .B(n960), .C(n2653), .Q(alu_o_data_AluRes[20]) );
  AOI212 U2754 ( .A(n2505), .B(n248), .C(n2230), .Q(n2333) );
  OAI222 U2755 ( .A(n597), .B(n2552), .C(n829), .D(n919), .Q(n2582) );
  XNR22 U2756 ( .A(n2900), .B(n2899), .Q(n2920) );
  NAND22 U2757 ( .A(n2145), .B(n1343), .Q(n1063) );
  NAND33 U2758 ( .A(n2451), .B(n2450), .C(n2449), .Q(n2452) );
  AOI212 U2759 ( .A(n1364), .B(n2694), .C(n2301), .Q(n2323) );
  INV6 U2760 ( .A(n1667), .Q(n1040) );
  AOI212 U2761 ( .A(n2367), .B(n2235), .C(n2483), .Q(n2243) );
  NAND33 U2762 ( .A(n2618), .B(n2619), .C(n2620), .Q(alu_o_data_AluRes[19]) );
  AOI2112 U2763 ( .A(n207), .B(n1065), .C(n2151), .D(n2150), .Q(n1062) );
  OAI212 U2764 ( .A(n2834), .B(n2637), .C(n2573), .Q(n2577) );
  INV6 U2765 ( .A(n2498), .Q(n1497) );
  NOR24 U2766 ( .A(n1679), .B(n1730), .Q(n1715) );
  NOR24 U2767 ( .A(n933), .B(n932), .Q(n2810) );
  AOI212 U2768 ( .A(n1345), .B(n2888), .C(n2887), .Q(n2889) );
  OAI212 U2769 ( .A(n2662), .B(n829), .C(n2661), .Q(n2684) );
  NAND33 U2770 ( .A(n2381), .B(n2380), .C(n2379), .Q(alu_o_data_AluRes[15]) );
  AOI212 U2771 ( .A(n3044), .B(n3043), .C(n3042), .Q(n3045) );
  AOI212 U2772 ( .A(n159), .B(i_data_rs[20]), .C(n1482), .Q(n1590) );
  AOI212 U2773 ( .A(n1345), .B(n2962), .C(n2961), .Q(n2963) );
  AOI212 U2774 ( .A(n1345), .B(n3025), .C(n3024), .Q(n3026) );
  NAND42 U2775 ( .A(n179), .B(n2243), .C(n2238), .D(n2237), .Q(n2248) );
  AOI212 U2776 ( .A(n1345), .B(n2851), .C(n2850), .Q(n2852) );
  OAI212 U2777 ( .A(n2846), .B(n3006), .C(n2845), .Q(n2847) );
  AOI2112 U2778 ( .A(n3070), .B(n1345), .C(n1020), .D(n1019), .Q(n1022) );
  NAND33 U2779 ( .A(n2687), .B(n2685), .C(n2686), .Q(alu_o_data_AluRes[21]) );
  OAI212 U2780 ( .A(n1222), .B(n2960), .C(n2959), .Q(n2961) );
  NOR32 U2781 ( .A(n2957), .B(n2958), .C(n2956), .Q(n2959) );
  INV15 U2782 ( .A(n1351), .Q(n1349) );
  OAI212 U2783 ( .A(n2833), .B(n2834), .C(n2832), .Q(n2848) );
  INV3 U2784 ( .A(n1563), .Q(n3083) );
  NOR21 U2785 ( .A(n2423), .B(n2309), .Q(n2272) );
  NOR21 U2786 ( .A(u_alu_lt_x_11_n105), .B(n188), .Q(n1890) );
  NAND22 U2787 ( .A(n2275), .B(n2395), .Q(n2256) );
  NAND30 U2788 ( .A(n2643), .B(n229), .C(n2977), .Q(n2239) );
  IMUX21 U2789 ( .A(n1345), .B(n178), .S(n2500), .Q(n2501) );
  NAND22 U2790 ( .A(n2540), .B(n2543), .Q(n2500) );
  NAND22 U2791 ( .A(n2496), .B(u_alu_DP_OP_83J3_124_3384_n154), .Q(n2540) );
  NAND22 U2792 ( .A(n2052), .B(n2164), .Q(n2055) );
  INV3 U2793 ( .A(u_alu_lt_x_11_n90), .Q(n2052) );
  NOR21 U2794 ( .A(n2161), .B(n2470), .Q(n1171) );
  INV3 U2795 ( .A(n247), .Q(n1138) );
  NOR21 U2796 ( .A(n1299), .B(n255), .Q(n2324) );
  AOI221 U2797 ( .A(n2154), .B(n1359), .C(n2060), .D(n1358), .Q(n2119) );
  NOR21 U2798 ( .A(u_alu_lt_x_11_B_0_), .B(n3049), .Q(n1735) );
  OAI220 U2799 ( .A(n1366), .B(n217), .C(n2517), .D(n177), .Q(n1691) );
  NAND22 U2800 ( .A(n2643), .B(n2693), .Q(n1920) );
  NOR20 U2801 ( .A(n177), .B(n249), .Q(n2862) );
  INV3 U2802 ( .A(n2857), .Q(n2856) );
  NAND22 U2803 ( .A(i_con_Ealuop[5]), .B(i_con_Ealuop[0]), .Q(n1727) );
  NOR21 U2804 ( .A(i_con_bop[2]), .B(n1562), .Q(n1240) );
  INV3 U2805 ( .A(i_data_fbmemout[19]), .Q(n1313) );
  INV3 U2806 ( .A(i_data_rt[27]), .Q(n1514) );
  NAND22 U2807 ( .A(n1346), .B(n1521), .Q(n1522) );
  INV3 U2808 ( .A(i_data_rt[25]), .Q(n1431) );
  INV3 U2809 ( .A(i_con_bop[0]), .Q(n1562) );
  INV3 U2810 ( .A(i_data_famemout[12]), .Q(n1528) );
  NOR21 U2811 ( .A(i_data_rt[1]), .B(n1347), .Q(n1651) );
  INV3 U2812 ( .A(i_data_rt[6]), .Q(n1451) );
  OAI222 U2813 ( .A(n1096), .B(n1095), .C(n2976), .D(n2440), .Q(n1094) );
  OAI212 U2814 ( .A(n190), .B(n2976), .C(n2775), .Q(n2776) );
  INV3 U2815 ( .A(u_alu_DP_OP_84J3_125_2615_n47), .Q(
        u_alu_DP_OP_84J3_125_2615_n113) );
  NAND22 U2816 ( .A(n1675), .B(n1683), .Q(n965) );
  INV3 U2817 ( .A(i_data_fbmemout[2]), .Q(n1265) );
  NOR21 U2818 ( .A(n195), .B(u_alu_lt_x_11_B_25_), .Q(u_alu_lt_x_11_n29) );
  NAND22 U2819 ( .A(n2916), .B(n1233), .Q(n1227) );
  INV3 U2820 ( .A(n2252), .Q(n2977) );
  NOR21 U2821 ( .A(n235), .B(n256), .Q(n2253) );
  NAND22 U2822 ( .A(n1346), .B(n1526), .Q(n1527) );
  NOR21 U2823 ( .A(n163), .B(n255), .Q(n2076) );
  NAND22 U2824 ( .A(n1630), .B(n1453), .Q(n1454) );
  NAND22 U2825 ( .A(n159), .B(i_data_rs[9]), .Q(n1011) );
  NOR31 U2826 ( .A(n2282), .B(n2281), .C(n2494), .Q(n2283) );
  NAND31 U2827 ( .A(n167), .B(n110), .C(n177), .Q(n1095) );
  NAND22 U2828 ( .A(n2227), .B(n242), .Q(n2228) );
  AOI211 U2829 ( .A(n172), .B(n910), .C(n1808), .Q(n1699) );
  NAND31 U2830 ( .A(n688), .B(n1364), .C(n172), .Q(n2152) );
  OAI212 U2831 ( .A(n1358), .B(n2756), .C(n2691), .Q(n2729) );
  NAND22 U2832 ( .A(n2758), .B(n1365), .Q(n2509) );
  NOR21 U2833 ( .A(n1357), .B(n3017), .Q(n2986) );
  AOI211 U2834 ( .A(n249), .B(n2874), .C(n2838), .Q(n2846) );
  OAI2111 U2835 ( .A(n1729), .B(n1728), .C(n1727), .D(n1726), .Q(n1731) );
  AOI212 U2836 ( .A(n2490), .B(n2491), .C(n2489), .Q(n2492) );
  NAND22 U2837 ( .A(n1346), .B(n1629), .Q(n1631) );
  NAND22 U2838 ( .A(n159), .B(i_data_rs[16]), .Q(n1496) );
  NAND22 U2839 ( .A(n90), .B(i_data_FMalures[21]), .Q(n1486) );
  NAND22 U2840 ( .A(n90), .B(i_data_FMalures[27]), .Q(n1510) );
  NAND22 U2841 ( .A(n1334), .B(i_data_FEalures[27]), .Q(n1574) );
  NAND22 U2842 ( .A(n90), .B(i_data_FMalures[28]), .Q(n1518) );
  NAND22 U2843 ( .A(n90), .B(i_data_FMalures[22]), .Q(n1418) );
  NAND22 U2844 ( .A(n89), .B(i_data_FMalures[24]), .Q(n1425) );
  NOR21 U2845 ( .A(n1374), .B(n250), .Q(n1375) );
  NOR21 U2846 ( .A(n1384), .B(n250), .Q(n1385) );
  NOR21 U2847 ( .A(n1379), .B(n250), .Q(n1380) );
  NAND22 U2848 ( .A(n89), .B(i_data_FMalures[0]), .Q(n1457) );
  NAND22 U2849 ( .A(n90), .B(i_data_FMalures[11]), .Q(n1435) );
  NAND22 U2850 ( .A(n90), .B(i_data_FMalures[14]), .Q(n1396) );
  AOI221 U2851 ( .A(n89), .B(i_data_FMalures[4]), .C(n158), .D(i_data_rs[4]), 
        .Q(n1072) );
  NAND22 U2852 ( .A(n2438), .B(n180), .Q(n2441) );
  OAI212 U2853 ( .A(n248), .B(n2229), .C(n2228), .Q(n2230) );
  AOI221 U2854 ( .A(n1070), .B(n2330), .C(n2433), .D(n1338), .Q(n1940) );
  NAND22 U2855 ( .A(n163), .B(n218), .Q(n2142) );
  NOR31 U2856 ( .A(n1359), .B(n3066), .C(n1779), .Q(n1723) );
  NAND22 U2857 ( .A(n54), .B(n2330), .Q(n1879) );
  NAND22 U2858 ( .A(n2457), .B(u_alu_lt_x_11_B_1_), .Q(n1258) );
  NAND22 U2859 ( .A(n2625), .B(n1356), .Q(n2626) );
  NAND22 U2860 ( .A(n2511), .B(n166), .Q(n2568) );
  NAND22 U2861 ( .A(n1230), .B(n166), .Q(n2510) );
  OAI212 U2862 ( .A(n2658), .B(n1358), .C(n2602), .Q(n2625) );
  NOR21 U2863 ( .A(n185), .B(n1361), .Q(n2090) );
  NOR21 U2864 ( .A(n1361), .B(n2689), .Q(n2554) );
  NAND22 U2865 ( .A(alu_i_data_B[27]), .B(n172), .Q(n991) );
  NAND22 U2866 ( .A(n3039), .B(n1190), .Q(n1009) );
  NAND22 U2867 ( .A(n946), .B(n1675), .Q(n945) );
  AOI2112 U2868 ( .A(n1309), .B(n1680), .C(i_data_immext[3]), .D(n980), .Q(
        n1673) );
  AOI212 U2869 ( .A(n2430), .B(n2429), .C(n2428), .Q(n2431) );
  NAND22 U2870 ( .A(n1631), .B(n1369), .Q(n1633) );
  OAI212 U2871 ( .A(i_data_FMalures[21]), .B(n198), .C(n1490), .Q(n1491) );
  NAND22 U2872 ( .A(n1334), .B(i_data_FEalures[28]), .Q(n1573) );
  NAND22 U2873 ( .A(n1335), .B(i_data_FEalures[29]), .Q(n1572) );
  NAND22 U2874 ( .A(n1335), .B(i_data_FEalures[24]), .Q(n1577) );
  NAND22 U2875 ( .A(n1335), .B(i_data_FEalures[11]), .Q(n1116) );
  NAND22 U2876 ( .A(n1352), .B(n1175), .Q(n1174) );
  NAND22 U2877 ( .A(n1335), .B(i_data_FEalures[4]), .Q(n1071) );
  NAND31 U2878 ( .A(n3023), .B(n2955), .C(n2883), .Q(n2210) );
  AOI221 U2879 ( .A(n1841), .B(n1358), .C(n1780), .D(n1359), .Q(n1781) );
  IMUX21 U2880 ( .A(n2714), .B(n2715), .S(u_alu_pre_sum_3a[0]), .Q(n2503) );
  NAND22 U2881 ( .A(n2817), .B(n1345), .Q(n1149) );
  AOI211 U2882 ( .A(n3035), .B(u_alu_lt_x_11_n12), .C(n3034), .Q(n3036) );
  NOR21 U2883 ( .A(n2494), .B(n1213), .Q(n2376) );
  OAI212 U2884 ( .A(n222), .B(n2180), .C(n2179), .Q(n2184) );
  OAI212 U2885 ( .A(n2172), .B(n1363), .C(n2171), .Q(n2298) );
  NAND31 U2886 ( .A(n2883), .B(n1358), .C(n177), .Q(n2328) );
  AOI211 U2887 ( .A(n1857), .B(n180), .C(n2040), .Q(n1874) );
  AOI221 U2888 ( .A(n2673), .B(n1357), .C(n1892), .D(n1356), .Q(n1893) );
  NAND22 U2889 ( .A(u_alu_ashr_4_A_17_), .B(n2330), .Q(n2114) );
  NAND22 U2890 ( .A(n2553), .B(n166), .Q(n2115) );
  OAI222 U2891 ( .A(n1942), .B(n1361), .C(n1362), .D(n1941), .Q(n2060) );
  OAI212 U2892 ( .A(n1363), .B(n2059), .C(n2058), .Q(n2154) );
  NAND22 U2893 ( .A(n2504), .B(n166), .Q(n2229) );
  NOR21 U2894 ( .A(n1357), .B(n2863), .Q(n2091) );
  NAND22 U2895 ( .A(n2444), .B(n172), .Q(n1779) );
  OAI212 U2896 ( .A(n3006), .B(n2580), .C(n2579), .Q(n2581) );
  NOR21 U2897 ( .A(n1367), .B(n2287), .Q(n1701) );
  OAI222 U2898 ( .A(n219), .B(n2432), .C(n2558), .D(n1985), .Q(n1807) );
  OAI222 U2899 ( .A(n3058), .B(n172), .C(n2180), .D(n1367), .Q(n1842) );
  OAI212 U2900 ( .A(n177), .B(n2824), .C(n1690), .Q(n1913) );
  NAND22 U2901 ( .A(n2295), .B(n1367), .Q(n1909) );
  NAND22 U2902 ( .A(u_alu_lt_x_11_B_0_), .B(n2830), .Q(n2019) );
  OAI311 U2903 ( .A(n2696), .B(n2697), .C(n1356), .D(n2695), .Q(n2698) );
  OAI212 U2904 ( .A(n2614), .B(n3006), .C(n2613), .Q(n2615) );
  OAI212 U2905 ( .A(n2656), .B(n1361), .C(n2506), .Q(n2601) );
  OAI212 U2906 ( .A(n2655), .B(n245), .C(n2226), .Q(n2505) );
  NAND31 U2907 ( .A(alu_i_data_B[19]), .B(n1364), .C(n177), .Q(n2169) );
  NAND22 U2908 ( .A(n2755), .B(n166), .Q(n2170) );
  OAI222 U2909 ( .A(n1364), .B(n2203), .C(n2202), .D(n2562), .Q(n2219) );
  NAND31 U2910 ( .A(n1260), .B(n1259), .C(n1363), .Q(n2205) );
  NAND22 U2911 ( .A(n1302), .B(n1736), .Q(n1090) );
  NAND22 U2912 ( .A(n245), .B(n249), .Q(n2088) );
  BUF6 U2913 ( .A(n1362), .Q(n1363) );
  OAI212 U2914 ( .A(n2806), .B(n2793), .C(n215), .Q(n2794) );
  OAI212 U2915 ( .A(u_alu_lt_x_11_n105), .B(n2454), .C(n2464), .Q(n2456) );
  NAND31 U2916 ( .A(n1996), .B(n1995), .C(n76), .Q(n1998) );
  OAI212 U2917 ( .A(n2821), .B(n1176), .C(n207), .Q(n1026) );
  INV3 U2918 ( .A(n1556), .Q(n1645) );
  OAI2111 U2919 ( .A(i_con_bop[1]), .B(i_con_bop[2]), .C(n1717), .D(n1562), 
        .Q(n1409) );
  NAND22 U2920 ( .A(n1334), .B(i_data_FEalures[18]), .Q(n2544) );
  NAND22 U2921 ( .A(n1334), .B(i_data_FEalures[22]), .Q(n1583) );
  OAI312 U2922 ( .A(i_con_bop[1]), .B(n1717), .C(n1412), .D(n1411), .Q(n1557)
         );
  NAND22 U2923 ( .A(n1335), .B(i_data_FEalures[12]), .Q(n1530) );
  NOR21 U2924 ( .A(n1458), .B(n250), .Q(n1459) );
  INV3 U2925 ( .A(i_data_FEalures[6]), .Q(n1450) );
  NAND22 U2926 ( .A(n1351), .B(n1121), .Q(n1120) );
  NAND22 U2927 ( .A(n1335), .B(i_data_FEalures[9]), .Q(n1013) );
  INV3 U2928 ( .A(n1816), .Q(n1763) );
  INV3 U2929 ( .A(n57), .Q(n1751) );
  OAI212 U2930 ( .A(n2638), .B(n2211), .C(n2210), .Q(n2212) );
  NAND22 U2931 ( .A(n2643), .B(n2946), .Q(n2201) );
  OAI212 U2932 ( .A(n1356), .B(n78), .C(n2177), .Q(n2215) );
  NAND22 U2933 ( .A(n2176), .B(n1356), .Q(n2177) );
  NOR21 U2934 ( .A(n2483), .B(n2234), .Q(n2168) );
  NAND22 U2935 ( .A(n2198), .B(n1344), .Q(n988) );
  NAND22 U2936 ( .A(n1831), .B(n2461), .Q(n1833) );
  AOI211 U2937 ( .A(n1817), .B(n180), .C(n1823), .Q(n1818) );
  NAND22 U2938 ( .A(n2513), .B(n172), .Q(n1816) );
  NOR21 U2939 ( .A(n1357), .B(n3006), .Q(n1813) );
  NAND22 U2940 ( .A(n1031), .B(n1028), .Q(alu_o_data_AluRes[14]) );
  NAND22 U2941 ( .A(n2290), .B(n2283), .Q(n2294) );
  NAND22 U2942 ( .A(n2643), .B(n2287), .Q(n2286) );
  NAND22 U2943 ( .A(n2367), .B(n2358), .Q(n2290) );
  INV3 U2944 ( .A(n2303), .Q(n2289) );
  OAI212 U2945 ( .A(n2308), .B(n2307), .C(n2304), .Q(n2271) );
  INV3 U2946 ( .A(n2345), .Q(n1182) );
  NAND22 U2947 ( .A(n1180), .B(n2184), .Q(n1178) );
  NAND22 U2948 ( .A(n2183), .B(n1180), .Q(n1179) );
  NOR21 U2949 ( .A(n2343), .B(n2349), .Q(n2278) );
  OAI212 U2950 ( .A(n3006), .B(n1806), .C(n1805), .Q(alu_o_data_AluRes[2]) );
  INV3 U2951 ( .A(n1847), .Q(n1787) );
  NOR21 U2952 ( .A(n3066), .B(n1781), .Q(n1803) );
  NAND22 U2953 ( .A(n2643), .B(n1782), .Q(n1776) );
  INV3 U2954 ( .A(n1234), .Q(n1782) );
  NAND22 U2955 ( .A(n2051), .B(n2050), .Q(alu_o_data_AluRes[8]) );
  NOR21 U2956 ( .A(n1992), .B(n520), .Q(n2014) );
  OAI212 U2957 ( .A(n2061), .B(n1356), .C(n1991), .Q(n2016) );
  NAND22 U2958 ( .A(n3103), .B(n3101), .Q(o_addr_Erd[2]) );
  NAND22 U2959 ( .A(n3103), .B(n3102), .Q(o_addr_Erd[4]) );
  NAND22 U2960 ( .A(n1905), .B(n207), .Q(n1906) );
  NAND22 U2961 ( .A(n189), .B(n1922), .Q(n1904) );
  NAND22 U2962 ( .A(n1969), .B(n203), .Q(n1901) );
  AOI211 U2963 ( .A(n1296), .B(n2463), .C(n1936), .Q(n1889) );
  OAI212 U2964 ( .A(n1356), .B(n1917), .C(n1886), .Q(n1908) );
  INV3 U2965 ( .A(n2317), .Q(n2264) );
  INV3 U2966 ( .A(n2270), .Q(n2260) );
  INV3 U2967 ( .A(n2307), .Q(n2261) );
  NAND22 U2968 ( .A(n2245), .B(n2244), .Q(n2246) );
  INV3 U2969 ( .A(n2243), .Q(n2245) );
  OAI212 U2970 ( .A(n2354), .B(n2834), .C(n2224), .Q(n2251) );
  NAND31 U2971 ( .A(n2361), .B(n2236), .C(n2244), .Q(n2224) );
  NOR21 U2972 ( .A(n2234), .B(n2359), .Q(n2236) );
  NAND31 U2973 ( .A(n2574), .B(n2883), .C(n1358), .Q(n2450) );
  OAI212 U2974 ( .A(n1357), .B(n2437), .C(n2436), .Q(n2453) );
  NAND22 U2975 ( .A(n2508), .B(n1357), .Q(n2436) );
  NAND31 U2976 ( .A(n2524), .B(n2523), .C(n2522), .Q(n2525) );
  NAND31 U2977 ( .A(n3065), .B(n2843), .C(n177), .Q(n2523) );
  AOI211 U2978 ( .A(n2520), .B(n993), .C(n2519), .Q(n2524) );
  INV3 U2979 ( .A(n2499), .Q(n2496) );
  OAI212 U2980 ( .A(n2494), .B(n2080), .C(n2079), .Q(alu_o_data_AluRes[9]) );
  INV3 U2981 ( .A(n2072), .Q(n1127) );
  AOI211 U2982 ( .A(n2071), .B(n180), .C(n964), .Q(n2072) );
  NAND31 U2983 ( .A(n2736), .B(n2735), .C(n2734), .Q(n2737) );
  INV3 U2984 ( .A(n2747), .Q(n2748) );
  NAND22 U2985 ( .A(n2795), .B(n2744), .Q(n2746) );
  OAI212 U2986 ( .A(n2231), .B(n1358), .C(n2155), .Q(n2176) );
  AOI211 U2987 ( .A(n2128), .B(n180), .C(n2904), .Q(n2151) );
  NAND22 U2988 ( .A(n2141), .B(n2194), .Q(n2143) );
  OAI2111 U2989 ( .A(n1360), .B(n2242), .C(n2148), .D(n2883), .Q(n2149) );
  NOR21 U2990 ( .A(n2476), .B(n2166), .Q(n2126) );
  NAND22 U2991 ( .A(n2819), .B(n2818), .Q(n1287) );
  NAND22 U2992 ( .A(n1190), .B(n2928), .Q(n2814) );
  NAND22 U2993 ( .A(n1023), .B(n1022), .Q(alu_o_data_AluRes[31]) );
  NOR21 U2994 ( .A(n185), .B(n1316), .Q(n1331) );
  INV3 U2995 ( .A(n3057), .Q(n1139) );
  AOI211 U2996 ( .A(n3048), .B(n180), .C(n3059), .Q(n3067) );
  OAI212 U2997 ( .A(n3038), .B(n3037), .C(n3036), .Q(n3042) );
  NAND22 U2998 ( .A(n3029), .B(u_alu_lt_x_11_n10), .Q(n3046) );
  NAND22 U2999 ( .A(n2373), .B(n2375), .Q(n2377) );
  INV3 U3000 ( .A(n2372), .Q(n2375) );
  NAND31 U3001 ( .A(n2371), .B(n2374), .C(n2372), .Q(n2378) );
  NAND22 U3002 ( .A(n2370), .B(n2485), .Q(n2372) );
  INV3 U3003 ( .A(n2484), .Q(n2370) );
  OAI212 U3004 ( .A(n2638), .B(n2354), .C(n2353), .Q(n2355) );
  NAND22 U3005 ( .A(n2221), .B(n172), .Q(n2354) );
  INV3 U3006 ( .A(n2988), .Q(n2220) );
  AOI211 U3007 ( .A(n2345), .B(n2344), .C(n2343), .Q(n2346) );
  NOR21 U3008 ( .A(n233), .B(n2287), .Q(n2343) );
  OAI212 U3009 ( .A(n2277), .B(n2276), .C(n2275), .Q(n2345) );
  NAND22 U3010 ( .A(n2287), .B(n233), .Q(n2344) );
  NAND22 U3011 ( .A(n2342), .B(n2391), .Q(n2351) );
  OAI212 U3012 ( .A(n2328), .B(n2327), .C(n2326), .Q(n2337) );
  INV3 U3013 ( .A(n3065), .Q(n2327) );
  OAI212 U3014 ( .A(n35), .B(n1356), .C(n1134), .Q(n3065) );
  NOR21 U3015 ( .A(n2422), .B(n2418), .Q(n2313) );
  INV3 U3016 ( .A(n1874), .Q(n1269) );
  NAND22 U3017 ( .A(n1770), .B(n1363), .Q(n1771) );
  NAND22 U3018 ( .A(n1769), .B(n1768), .Q(n1770) );
  NAND22 U3019 ( .A(n1913), .B(n1364), .Q(n1769) );
  OAI212 U3020 ( .A(n1982), .B(n3006), .C(n1981), .Q(alu_o_data_AluRes[7]) );
  OAI212 U3021 ( .A(n1978), .B(n3066), .C(n1977), .Q(n1979) );
  OAI212 U3022 ( .A(n1291), .B(n1290), .C(n1288), .Q(n1977) );
  AOI211 U3023 ( .A(n1291), .B(n1973), .C(n1289), .Q(n1288) );
  INV3 U3024 ( .A(n1974), .Q(n1290) );
  NAND22 U3025 ( .A(n1296), .B(n1292), .Q(n1291) );
  NOR21 U3026 ( .A(n2007), .B(n1972), .Q(n1292) );
  OAI212 U3027 ( .A(n1961), .B(n1960), .C(n1959), .Q(n1967) );
  NAND22 U3028 ( .A(n1956), .B(n1955), .Q(n1957) );
  NAND22 U3029 ( .A(n1951), .B(n1953), .Q(n1960) );
  OAI212 U3030 ( .A(n110), .B(n1944), .C(n1943), .Q(n1990) );
  NAND22 U3031 ( .A(n2120), .B(n168), .Q(n2121) );
  NAND22 U3032 ( .A(n2297), .B(n248), .Q(n2116) );
  OAI212 U3033 ( .A(n1985), .B(n1984), .C(n1983), .Q(n1986) );
  INV3 U3034 ( .A(n2153), .Q(n1942) );
  NAND22 U3035 ( .A(n2138), .B(n2194), .Q(n2103) );
  NAND22 U3036 ( .A(n2023), .B(n172), .Q(n2092) );
  NAND22 U3037 ( .A(n2022), .B(n2761), .Q(n2023) );
  OAI212 U3038 ( .A(n2865), .B(n2091), .C(n172), .Q(n2211) );
  NAND22 U3039 ( .A(n2086), .B(n2085), .Q(n2123) );
  NAND22 U3040 ( .A(u_alu_lt_x_11_n87), .B(n2165), .Q(n2083) );
  INV3 U3041 ( .A(n2361), .Q(n2284) );
  OAI212 U3042 ( .A(n1750), .B(n1356), .C(n1711), .Q(n1742) );
  OAI222 U3043 ( .A(n1772), .B(n175), .C(n1692), .D(n248), .Q(n1697) );
  AOI221 U3044 ( .A(n1691), .B(n1364), .C(n1913), .D(n166), .Q(n1692) );
  AOI211 U3045 ( .A(n1909), .B(n1686), .C(n176), .Q(n1687) );
  NOR21 U3046 ( .A(u_alu_lt_x_11_n105), .B(n1936), .Q(u_alu_lt_x_11_n103) );
  NOR21 U3047 ( .A(n1052), .B(u_alu_lt_x_11_B_29_), .Q(u_alu_lt_x_11_n15) );
  NAND22 U3048 ( .A(u_alu_pre_sum_3a[2]), .B(n2715), .Q(n2583) );
  NAND22 U3049 ( .A(n2443), .B(n243), .Q(n2445) );
  NAND22 U3050 ( .A(n2320), .B(n166), .Q(n2321) );
  INV3 U3051 ( .A(n2442), .Q(n2446) );
  OAI212 U3052 ( .A(u_alu_lt_x_11_n138), .B(n2561), .C(n2560), .Q(n2578) );
  NAND22 U3053 ( .A(n2331), .B(n200), .Q(n2332) );
  OAI212 U3054 ( .A(n245), .B(n211), .C(n2152), .Q(n2331) );
  INV3 U3055 ( .A(n2551), .Q(n2547) );
  NAND22 U3056 ( .A(n1704), .B(n245), .Q(n1705) );
  NAND22 U3057 ( .A(n1703), .B(n1702), .Q(n1704) );
  NAND22 U3058 ( .A(n1693), .B(n176), .Q(n1694) );
  OAI212 U3059 ( .A(n1361), .B(n2117), .C(n1915), .Q(n1989) );
  AOI221 U3060 ( .A(n1914), .B(n175), .C(n1913), .D(n242), .Q(n1915) );
  NOR21 U3061 ( .A(n1985), .B(n2517), .Q(n1914) );
  INV3 U3062 ( .A(n1296), .Q(n2006) );
  INV3 U3063 ( .A(n2009), .Q(n1976) );
  NAND22 U3064 ( .A(n205), .B(n177), .Q(n1935) );
  NAND22 U3065 ( .A(n1934), .B(n172), .Q(n2024) );
  INV3 U3066 ( .A(n2699), .Q(n1934) );
  NAND22 U3067 ( .A(n1928), .B(n1927), .Q(n1925) );
  INV3 U3068 ( .A(n1951), .Q(n1927) );
  OAI212 U3069 ( .A(n1851), .B(n1850), .C(n2038), .Q(n1855) );
  AOI211 U3070 ( .A(n1918), .B(n180), .C(n2693), .Q(n1931) );
  NAND22 U3071 ( .A(n2628), .B(n2663), .Q(n2651) );
  INV3 U3072 ( .A(u_alu_lt_x_11_n47), .Q(n2628) );
  INV3 U3073 ( .A(n1108), .Q(n1107) );
  NAND22 U3074 ( .A(u_alu_pre_sum_3b[4]), .B(n2714), .Q(n2653) );
  OAI212 U3075 ( .A(n2920), .B(n844), .C(n2919), .Q(n2921) );
  INV3 U3076 ( .A(n1142), .Q(n1141) );
  INV3 U3077 ( .A(u_alu_lt_x_11_B_11_), .Q(n2904) );
  OAI212 U3078 ( .A(n1298), .B(n2898), .C(n2897), .Q(n2895) );
  NAND22 U3079 ( .A(n191), .B(u_alu_lt_x_11_n26), .Q(n2898) );
  INV3 U3080 ( .A(n2900), .Q(n2896) );
  INV3 U3081 ( .A(n2932), .Q(n2892) );
  INV3 U3082 ( .A(u_alu_DP_OP_84J3_125_2615_n36), .Q(
        u_alu_DP_OP_84J3_125_2615_n111) );
  OAI212 U3083 ( .A(n2886), .B(n844), .C(n2885), .Q(n2887) );
  NAND22 U3084 ( .A(n168), .B(n1325), .Q(n1326) );
  OAI212 U3085 ( .A(n2766), .B(n2765), .C(n2764), .Q(n2767) );
  NAND22 U3086 ( .A(n2763), .B(n2862), .Q(n2764) );
  INV3 U3087 ( .A(n937), .Q(n936) );
  INV3 U3088 ( .A(n2861), .Q(n2859) );
  INV3 U3089 ( .A(u_alu_lt_x_11_n26), .Q(n2855) );
  NAND22 U3090 ( .A(n1021), .B(u_alu_pre_sum_4b[2]), .Q(n2891) );
  INV3 U3091 ( .A(u_alu_DP_OP_84J3_125_2615_n103), .Q(
        u_alu_DP_OP_84J3_125_2615_n102) );
  INV3 U3092 ( .A(u_alu_DP_OP_84J3_125_2615_n39), .Q(
        u_alu_DP_OP_84J3_125_2615_n112) );
  INV3 U3093 ( .A(n2936), .Q(n2934) );
  NAND22 U3094 ( .A(n2997), .B(n2993), .Q(n2936) );
  INV3 U3095 ( .A(n2968), .Q(n2997) );
  NAND22 U3096 ( .A(n1021), .B(u_alu_pre_sum_4b[4]), .Q(n2965) );
  NAND22 U3097 ( .A(u_alu_pre_sum_3a[6]), .B(n2715), .Q(n2712) );
  NAND22 U3098 ( .A(u_alu_pre_sum_3b[6]), .B(n2714), .Q(n2713) );
  OAI212 U3099 ( .A(n177), .B(n2699), .C(n2698), .Q(n2777) );
  AOI211 U3100 ( .A(n2749), .B(n72), .C(n2706), .Q(n2707) );
  NAND22 U3101 ( .A(u_alu_DP_OP_83J3_124_3384_n152), .B(n182), .Q(n2744) );
  INV3 U3102 ( .A(n1144), .Q(n2743) );
  NAND22 U3103 ( .A(n2513), .B(n1366), .Q(n2514) );
  OAI222 U3104 ( .A(n1753), .B(n1356), .C(n1752), .D(n249), .Q(n2513) );
  INV3 U3105 ( .A(n1777), .Q(n1752) );
  NAND22 U3106 ( .A(n2170), .B(n2169), .Q(n2434) );
  NAND22 U3107 ( .A(u_alu_pre_sum_3a[3]), .B(n2715), .Q(n2619) );
  INV3 U3108 ( .A(u_alu_DP_OP_83J3_124_3384_n51), .Q(
        u_alu_DP_OP_83J3_124_3384_n50) );
  NAND22 U3109 ( .A(u_alu_pre_sum_3b[3]), .B(n2714), .Q(n2620) );
  INV3 U3110 ( .A(u_alu_DP_OP_83J3_124_3384_n113), .Q(
        u_alu_DP_OP_83J3_124_3384_n112) );
  INV3 U3111 ( .A(n929), .Q(n928) );
  OAI212 U3112 ( .A(n1298), .B(n2971), .C(n2970), .Q(n2969) );
  NAND22 U3113 ( .A(n3031), .B(n2993), .Q(n2971) );
  NAND22 U3114 ( .A(n924), .B(n923), .Q(n922) );
  OAI212 U3115 ( .A(n1298), .B(n3001), .C(n3000), .Q(n2998) );
  INV3 U3116 ( .A(n1195), .Q(n1194) );
  INV3 U3117 ( .A(u_alu_lt_x_11_n12), .Q(n2992) );
  NAND22 U3118 ( .A(n1021), .B(u_alu_pre_sum_4b[6]), .Q(n3028) );
  NAND22 U3119 ( .A(u_alu_lt_x_11_B_29_), .B(n1276), .Q(
        u_alu_DP_OP_84J3_125_2615_n22) );
  XOR21 U3120 ( .A(n2665), .B(n2664), .Q(n918) );
  INV3 U3121 ( .A(n2206), .Q(n2207) );
  NAND22 U3122 ( .A(n1234), .B(n242), .Q(n1814) );
  NAND22 U3123 ( .A(n1361), .B(n1365), .Q(n2089) );
  OAI212 U3124 ( .A(n2669), .B(n2976), .C(n2668), .Q(n2680) );
  NOR21 U3125 ( .A(n193), .B(n187), .Q(n968) );
  AOI211 U3126 ( .A(n2666), .B(n180), .C(n181), .Q(n2681) );
  OAI212 U3127 ( .A(n248), .B(n2622), .C(n2621), .Q(n2690) );
  NAND31 U3128 ( .A(n2755), .B(n248), .C(n176), .Q(n2621) );
  INV3 U3129 ( .A(n991), .Q(n2755) );
  NAND22 U3130 ( .A(n2627), .B(alu_i_data_B[20]), .Q(n2663) );
  NAND22 U3131 ( .A(n2741), .B(u_alu_lt_x_11_n46), .Q(n2665) );
  NAND22 U3132 ( .A(n181), .B(n1318), .Q(n2741) );
  NAND22 U3133 ( .A(u_alu_pre_sum_3a[5]), .B(n2715), .Q(n2686) );
  NAND22 U3134 ( .A(u_alu_pre_sum_3b[5]), .B(n2714), .Q(n2687) );
  NAND22 U3135 ( .A(n920), .B(n178), .Q(n962) );
  NAND22 U3136 ( .A(n177), .B(n249), .Q(n2766) );
  BUF6 U3137 ( .A(i_data_immext[6]), .Q(n1357) );
  NAND22 U3138 ( .A(n1125), .B(n1124), .Q(n1123) );
  NAND22 U3139 ( .A(n1230), .B(n236), .Q(n1228) );
  INV3 U3140 ( .A(n2018), .Q(n1231) );
  NAND22 U3141 ( .A(n2511), .B(n2073), .Q(n1224) );
  INV3 U3142 ( .A(n1226), .Q(n1225) );
  NAND22 U3143 ( .A(n2809), .B(n2794), .Q(n2797) );
  INV3 U3144 ( .A(n2828), .Q(n2826) );
  OAI212 U3145 ( .A(n2488), .B(n2364), .C(n2487), .Q(n2489) );
  NAND22 U3146 ( .A(n2475), .B(u_alu_lt_x_11_n87), .Q(n2478) );
  OAI212 U3147 ( .A(n2472), .B(n2473), .C(n2471), .Q(n2493) );
  NOR31 U3148 ( .A(n2469), .B(n2488), .C(n2470), .Q(n2471) );
  NAND22 U3149 ( .A(n2030), .B(n1306), .Q(n2009) );
  NAND22 U3150 ( .A(n1021), .B(u_alu_pre_sum_4b[1]), .Q(n2854) );
  OAI212 U3151 ( .A(u_alu_DP_OP_83J3_124_3384_n52), .B(
        u_alu_DP_OP_83J3_124_3384_n54), .C(u_alu_DP_OP_83J3_124_3384_n53), .Q(
        u_alu_DP_OP_83J3_124_3384_n113) );
  OAI222 U3152 ( .A(n1677), .B(n1657), .C(n1665), .D(n1662), .Q(n1729) );
  INV3 U3153 ( .A(n1004), .Q(n1003) );
  NAND22 U3154 ( .A(n1670), .B(n1669), .Q(n1671) );
  OAI212 U3155 ( .A(n1666), .B(n1665), .C(n1664), .Q(n1668) );
  AOI211 U3156 ( .A(n1681), .B(i_con_Ealuop[3]), .C(i_con_Ealuop[5]), .Q(n1666) );
  NAND22 U3157 ( .A(n1659), .B(n1678), .Q(n1660) );
  NAND22 U3158 ( .A(i_data_immext[1]), .B(n1309), .Q(n1657) );
  NAND22 U3159 ( .A(i_con_Ealuop[2]), .B(i_con_Ealuop[3]), .Q(n1661) );
  NAND22 U3160 ( .A(n981), .B(n980), .Q(n979) );
  NAND22 U3161 ( .A(u_alu_DP_OP_83J3_124_3384_n153), .B(
        u_alu_DP_OP_85J3_126_1427_n377), .Q(u_alu_DP_OP_83J3_124_3384_n16) );
  NAND22 U3162 ( .A(n1339), .B(n1318), .Q(u_alu_DP_OP_83J3_124_3384_n30) );
  NAND22 U3163 ( .A(alu_i_data_B[19]), .B(n2594), .Q(
        u_alu_DP_OP_83J3_124_3384_n42) );
  INV3 U3164 ( .A(n1046), .Q(n1045) );
  OAI212 U3165 ( .A(n2427), .B(n2426), .C(n2425), .Q(n2428) );
  NAND22 U3166 ( .A(n2424), .B(n2419), .Q(n2427) );
  NAND22 U3167 ( .A(n2419), .B(n2415), .Q(n2416) );
  NAND22 U3168 ( .A(n2563), .B(n233), .Q(n2419) );
  INV3 U3169 ( .A(n2424), .Q(n2418) );
  OAI212 U3170 ( .A(n2414), .B(n2413), .C(n209), .Q(n2430) );
  NAND31 U3171 ( .A(n184), .B(n2409), .C(n2408), .Q(n2410) );
  OAI212 U3172 ( .A(n2402), .B(n2401), .C(n2400), .Q(n1109) );
  NAND22 U3173 ( .A(n2253), .B(n2223), .Q(n2395) );
  AOI211 U3174 ( .A(n2287), .B(n233), .C(n2394), .Q(n2397) );
  NOR21 U3175 ( .A(n1438), .B(n1439), .Q(n2132) );
  INV3 U3176 ( .A(n2178), .Q(n2187) );
  NAND22 U3177 ( .A(n1249), .B(n1252), .Q(n2390) );
  INV3 U3178 ( .A(n1253), .Q(n1252) );
  NAND22 U3179 ( .A(n2386), .B(n2387), .Q(n1253) );
  OAI212 U3180 ( .A(n1250), .B(n2385), .C(n2384), .Q(n1249) );
  NAND31 U3181 ( .A(n2383), .B(n2382), .C(u_alu_lt_x_11_A_0_), .Q(n2385) );
  NAND22 U3182 ( .A(i_data_immext[1]), .B(n170), .Q(n2035) );
  INV3 U3183 ( .A(n1853), .Q(n1036) );
  NAND22 U3184 ( .A(n1309), .B(n170), .Q(n1791) );
  NAND22 U3185 ( .A(i_data_immext[4]), .B(n170), .Q(n1858) );
  NAND22 U3186 ( .A(n1346), .B(n1495), .Q(n2801) );
  NAND22 U3187 ( .A(n1346), .B(n1489), .Q(n1490) );
  NAND22 U3188 ( .A(n1319), .B(i_data_famemout[21]), .Q(n1487) );
  NAND22 U3189 ( .A(n158), .B(i_data_rs[21]), .Q(n1485) );
  NAND22 U3190 ( .A(n1545), .B(i_data_famemout[20]), .Q(n1587) );
  NOR21 U3191 ( .A(i_data_rt[20]), .B(n1347), .Q(n1607) );
  NAND22 U3192 ( .A(n158), .B(i_data_rs[18]), .Q(n1464) );
  NAND22 U3193 ( .A(n158), .B(i_data_rs[26]), .Q(n1504) );
  INV3 U3194 ( .A(n1510), .Q(n957) );
  NAND22 U3195 ( .A(n158), .B(i_data_rs[27]), .Q(n1511) );
  NAND22 U3196 ( .A(n159), .B(i_data_rs[28]), .Q(n1519) );
  NAND22 U3197 ( .A(n1319), .B(i_data_famemout[28]), .Q(n1520) );
  INV3 U3198 ( .A(n1293), .Q(n1197) );
  NAND22 U3199 ( .A(n1525), .B(n1572), .Q(n1198) );
  NAND22 U3200 ( .A(n1319), .B(i_data_famemout[29]), .Q(n1525) );
  NAND22 U3201 ( .A(n158), .B(i_data_rs[22]), .Q(n1047) );
  NAND22 U3202 ( .A(n1319), .B(i_data_famemout[23]), .Q(n1579) );
  NAND22 U3203 ( .A(n1346), .B(n1002), .Q(n1001) );
  NAND22 U3204 ( .A(n1346), .B(n1428), .Q(n1113) );
  NAND22 U3205 ( .A(n1319), .B(i_data_famemout[24]), .Q(n1427) );
  NAND22 U3206 ( .A(n158), .B(i_data_rs[24]), .Q(n1426) );
  NAND22 U3207 ( .A(n89), .B(n1404), .Q(n1405) );
  NAND22 U3208 ( .A(n159), .B(n1403), .Q(n1406) );
  NAND22 U3209 ( .A(n158), .B(i_data_rs[2]), .Q(n1377) );
  NAND22 U3210 ( .A(n1352), .B(n1265), .Q(n1264) );
  NAND22 U3211 ( .A(n159), .B(i_data_rs[12]), .Q(n1529) );
  NAND22 U3212 ( .A(n48), .B(n1539), .Q(n1540) );
  NAND22 U3213 ( .A(n1346), .B(n1537), .Q(n1640) );
  NAND22 U3214 ( .A(n158), .B(i_data_rs[7]), .Q(n1387) );
  NAND22 U3215 ( .A(n1554), .B(n1553), .Q(n1644) );
  NAND22 U3216 ( .A(n244), .B(n1552), .Q(n1553) );
  NAND22 U3217 ( .A(n1346), .B(n1551), .Q(n1554) );
  NAND22 U3218 ( .A(n158), .B(i_data_rs[5]), .Q(n1382) );
  NAND22 U3219 ( .A(n244), .B(n1216), .Q(n1215) );
  NAND22 U3220 ( .A(n159), .B(i_data_rs[1]), .Q(n1245) );
  NAND22 U3221 ( .A(n158), .B(i_data_rs[0]), .Q(n1088) );
  OAI212 U3222 ( .A(n1439), .B(n1438), .C(n1155), .Q(n1154) );
  INV3 U3223 ( .A(n1593), .Q(n1438) );
  INV3 U3224 ( .A(n1594), .Q(n1439) );
  NAND22 U3225 ( .A(n159), .B(i_data_rs[11]), .Q(n1117) );
  NAND22 U3226 ( .A(n1346), .B(n1460), .Q(n2064) );
  NAND22 U3227 ( .A(n1352), .B(n1206), .Q(n1205) );
  INV3 U3228 ( .A(i_data_famemout[8]), .Q(n1463) );
  NAND22 U3229 ( .A(n1346), .B(n1447), .Q(n1448) );
  NAND22 U3230 ( .A(n159), .B(i_data_rs[6]), .Q(n1393) );
  INV3 U3231 ( .A(i_data_famemout[6]), .Q(n1391) );
  NAND22 U3232 ( .A(n1346), .B(n1441), .Q(n1442) );
  NAND22 U3233 ( .A(n158), .B(i_data_rs[14]), .Q(n1397) );
  NOR21 U3234 ( .A(n1394), .B(n250), .Q(n1395) );
  NAND22 U3235 ( .A(n1158), .B(n1157), .Q(n1156) );
  INV3 U3236 ( .A(n1390), .Q(n1073) );
  NOR21 U3237 ( .A(n1389), .B(n250), .Q(n1390) );
  NOR21 U3238 ( .A(i_data_rt[18]), .B(n1347), .Q(n1617) );
  XNR21 U3239 ( .A(n1758), .B(n1788), .Q(n1759) );
  XNR21 U3240 ( .A(n1796), .B(n1757), .Q(n1760) );
  XNR21 U3241 ( .A(n2197), .B(n2307), .Q(n2198) );
  XNR21 U3242 ( .A(n1789), .B(n1820), .Q(n1800) );
  NAND22 U3243 ( .A(n1017), .B(n3103), .Q(o_addr_Erd[3]) );
  XNR21 U3244 ( .A(n1890), .B(n1889), .Q(n1903) );
  IMUX20 U3245 ( .A(n174), .B(n3047), .S(u_alu_DP_OP_83J3_124_3384_n154), .Q(
        n2438) );
  XNR21 U3246 ( .A(n2540), .B(n2539), .Q(n2541) );
  IMUX20 U3247 ( .A(n3047), .B(n174), .S(n2406), .Q(n2071) );
  XNR21 U3248 ( .A(n2095), .B(n2067), .Q(n2070) );
  XNR21 U3249 ( .A(n2099), .B(n2068), .Q(n2069) );
  NOR20 U3250 ( .A(u_alu_DP_OP_83J3_124_3384_n153), .B(n3049), .Q(n2731) );
  OAI210 U3251 ( .A(n187), .B(u_alu_DP_OP_83J3_124_3384_n153), .C(n180), .Q(
        n2732) );
  XNR21 U3252 ( .A(n2751), .B(n2750), .Q(n2752) );
  IMUX20 U3253 ( .A(n1355), .B(n91), .S(n226), .Q(n2769) );
  OAI210 U3254 ( .A(n187), .B(n2754), .C(n180), .Q(n3050) );
  NOR20 U3255 ( .A(n2754), .B(n3049), .Q(n3051) );
  OAI210 U3256 ( .A(n2025), .B(n187), .C(n180), .Q(n1872) );
  XNR21 U3257 ( .A(n1870), .B(n2006), .Q(n1271) );
  OAI210 U3258 ( .A(n2146), .B(n187), .C(n180), .Q(n1963) );
  NAND20 U3259 ( .A(n1718), .B(u_alu_lt_x_11_n9), .Q(n1719) );
  XNR21 U3260 ( .A(n289), .B(u_alu_lt_x_11_B_0_), .Q(n1720) );
  NAND20 U3261 ( .A(u_alu_lt_x_11_B_29_), .B(n1052), .Q(u_alu_lt_x_11_n16) );
  NAND20 U3262 ( .A(alu_i_data_B[20]), .B(n2627), .Q(u_alu_lt_x_11_n48) );
  NAND20 U3263 ( .A(alu_i_data_B[19]), .B(u_alu_lt_x_11_n139), .Q(
        u_alu_lt_x_11_n54) );
  NOR20 U3264 ( .A(n2481), .B(n54), .Q(u_alu_lt_x_11_n78) );
  NAND20 U3265 ( .A(u_alu_lt_x_11_n122), .B(n1234), .Q(u_alu_lt_x_11_n115) );
  NOR20 U3266 ( .A(n1234), .B(u_alu_lt_x_11_n122), .Q(u_alu_lt_x_11_n114) );
  IMUX20 U3267 ( .A(n187), .B(n1342), .S(n2629), .Q(n2572) );
  XNR21 U3268 ( .A(n2651), .B(n2749), .Q(n2652) );
  XNR21 U3269 ( .A(n2651), .B(n2745), .Q(n2633) );
  IMUX20 U3270 ( .A(n187), .B(n91), .S(u_alu_DP_OP_85J3_126_1427_n374), .Q(
        n2635) );
  NOR20 U3271 ( .A(n177), .B(n1358), .Q(n1233) );
  IMUX20 U3272 ( .A(n1355), .B(n1342), .S(n1517), .Q(n2908) );
  NOR20 U3273 ( .A(alu_i_data_B[27]), .B(n3049), .Q(n2901) );
  NOR20 U3274 ( .A(n1336), .B(n3049), .Q(n2876) );
  NOR20 U3275 ( .A(u_alu_lt_x_11_B_28_), .B(n3049), .Q(n2943) );
  OAI210 U3276 ( .A(n187), .B(u_alu_lt_x_11_B_28_), .C(n180), .Q(n2944) );
  OAI210 U3277 ( .A(n173), .B(n2940), .C(u_alu_lt_x_11_B_28_), .Q(n2941) );
  IMUX20 U3278 ( .A(n1355), .B(n91), .S(n1524), .Q(n2940) );
  OAI210 U3279 ( .A(n1338), .B(n187), .C(n180), .Q(n1102) );
  IMUX20 U3280 ( .A(n187), .B(n1342), .S(n2594), .Q(n2608) );
  XNR21 U3281 ( .A(n2599), .B(n2598), .Q(n2600) );
  OAI210 U3282 ( .A(n971), .B(n2979), .C(u_alu_lt_x_11_B_29_), .Q(n2980) );
  IMUX20 U3283 ( .A(n1342), .B(n1355), .S(n1052), .Q(n2979) );
  NOR20 U3284 ( .A(u_alu_lt_x_11_B_29_), .B(n3049), .Q(n2974) );
  XNR21 U3285 ( .A(n210), .B(n2969), .Q(n2991) );
  OAI210 U3286 ( .A(n187), .B(u_alu_DP_OP_85J3_126_1427_n368), .C(n180), .Q(
        n3009) );
  NOR20 U3287 ( .A(u_alu_DP_OP_85J3_126_1427_n368), .B(n3049), .Q(n3010) );
  OAI210 U3288 ( .A(n971), .B(n3008), .C(u_alu_DP_OP_85J3_126_1427_n368), .Q(
        n3011) );
  NAND20 U3289 ( .A(n1361), .B(n1358), .Q(n992) );
  NAND20 U3290 ( .A(n1339), .B(n1361), .Q(n2675) );
  IMUX20 U3291 ( .A(n187), .B(n1342), .S(u_alu_DP_OP_85J3_126_1427_n379), .Q(
        n2831) );
  NOR20 U3292 ( .A(n249), .B(n185), .Q(n2073) );
  XNR21 U3293 ( .A(n2826), .B(n2825), .Q(n2851) );
  OAI210 U3294 ( .A(i_data_fbmemout[2]), .B(n246), .C(n1369), .Q(n1793) );
  XNR21 U3295 ( .A(n316), .B(n2204), .Q(n917) );
  NAND28 U3296 ( .A(n1372), .B(n1043), .Q(n1347) );
  OAI210 U3297 ( .A(u_alu_ashr_4_A_16_), .B(n187), .C(n180), .Q(n2447) );
  AOI220 U3298 ( .A(n247), .B(u_alu_ashr_4_A_16_), .C(u_alu_lt_x_11_B_0_), .D(
        n177), .Q(n1708) );
  XNR21 U3299 ( .A(n2632), .B(n2547), .Q(n2552) );
  NAND20 U3300 ( .A(u_alu_lt_x_11_B_25_), .B(n195), .Q(u_alu_lt_x_11_n30) );
  XNR21 U3301 ( .A(n2181), .B(n2098), .Q(n2106) );
  XNR21 U3302 ( .A(u_alu_DP_OP_83J3_124_3384_n4), .B(
        u_alu_DP_OP_83J3_124_3384_n31), .Q(u_alu_pre_sum_3a[5]) );
  NAND20 U3303 ( .A(n1044), .B(n234), .Q(u_alu_lt_x_11_n106) );
  NOR20 U3304 ( .A(n43), .B(n255), .Q(n2774) );
  XNR21 U3305 ( .A(n2934), .B(n2933), .Q(n2962) );
  NAND22 U3306 ( .A(n3103), .B(n3100), .Q(o_addr_Erd[1]) );
  OAI210 U3307 ( .A(u_alu_lt_x_11_B_0_), .B(n187), .C(n180), .Q(n1734) );
  NAND22 U3308 ( .A(n3103), .B(n3099), .Q(o_addr_Erd[0]) );
  OAI210 U3309 ( .A(n163), .B(n187), .C(n180), .Q(n2077) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_addr_Rt, i_con_RegWr, 
        i_addr_Rd, i_data_Rd, o_data_Rs, o_data_Rt );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rt;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr;
  wire   n5, n6, n9, n11, n13, n15, n16, n17, n18, n20, n21, n22, n23, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n1, n2, n3, n4, n7, n8, n10, n12, n14, n19, n24,
         n33, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608;
  wire   [1023:0] regs;

  DFEC1 regs_reg_31__31_ ( .D(n147), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1023]) );
  DFEC1 regs_reg_31__30_ ( .D(n145), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(n143), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(n141), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(n139), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(n137), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(n135), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(n133), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(n132), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(n129), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(n127), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(n125), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(n124), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(n121), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(n119), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(n117), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(n115), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(n113), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(n111), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(n109), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(n107), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(n105), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(n103), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(n101), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(n99), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(n97), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(n95), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(n93), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(n91), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(n89), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(n87), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(n85), .E(n31), .C(i_clk), .RN(i_rst_n), .Q(
        regs[992]) );
  DFEC1 regs_reg_30__31_ ( .D(n147), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(n145), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(n143), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(n141), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(n139), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(n137), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(n135), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(n133), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(n131), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(n129), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(n127), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(n125), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(n123), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(n121), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(n119), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(n117), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(n115), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(n113), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(n111), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(n109), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(n107), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(n105), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(n103), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(n101), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(n99), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(n97), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(n95), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(n93), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(n91), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(n89), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(n87), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(n85), .E(n30), .C(i_clk), .RN(i_rst_n), .Q(
        regs[960]) );
  DFEC1 regs_reg_29__31_ ( .D(n147), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(n145), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(n143), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(n141), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[956]) );
  DFEC1 regs_reg_29__27_ ( .D(n139), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(n137), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(n135), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(n133), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(n131), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(n129), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(n127), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(n125), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(n123), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(n121), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(n119), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(n117), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(n115), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(n113), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(n111), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(n109), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(n107), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(n105), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(n103), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(n101), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(n99), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(n97), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(n95), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(n93), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(n91), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(n89), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(n87), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(n85), .E(n29), .C(i_clk), .RN(i_rst_n), .Q(
        regs[928]) );
  DFEC1 regs_reg_28__31_ ( .D(n147), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(n145), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(n143), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(n141), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(n139), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(n137), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(n135), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(n133), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(n132), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(n129), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(n127), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(n125), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(n124), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(n121), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(n119), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(n117), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(n115), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(n113), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(n111), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(n109), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(n107), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(n105), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(n103), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(n101), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(n99), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(n97), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(n95), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(n93), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(n91), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(n89), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(n87), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(n85), .E(n28), .C(i_clk), .RN(i_rst_n), .Q(
        regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(n147), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(n145), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(n143), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(n141), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(n139), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(n137), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(n135), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(n133), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(n131), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(n129), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(n127), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(n125), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(n123), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(n121), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(n119), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(n117), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(n115), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(n113), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(n111), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(n109), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(n107), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(n105), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(n103), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(n101), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(n99), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(n97), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(n95), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(n93), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(n91), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(n89), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(n87), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(n85), .E(n27), .C(i_clk), .RN(i_rst_n), .Q(
        regs[864]) );
  DFEC1 regs_reg_26__31_ ( .D(n147), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(n145), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(n143), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(n141), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(n139), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(n137), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(n135), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(n133), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(n132), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(n129), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(n127), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(n125), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(n124), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(n121), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(n119), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(n117), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(n115), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(n113), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(n111), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(n109), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(n107), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(n105), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(n103), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(n101), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(n99), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(n97), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(n95), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(n93), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(n91), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(n89), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(n87), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(n85), .E(n26), .C(i_clk), .RN(i_rst_n), .Q(
        regs[832]) );
  DFEC1 regs_reg_25__31_ ( .D(n147), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(n145), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(n143), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(n141), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(n139), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(n137), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(n135), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(n133), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(n132), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(n129), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(n127), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(n125), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(n124), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(n121), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(n119), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(n117), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(n115), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(n113), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(n111), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(n109), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(n107), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(n105), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(n103), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(n101), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(n99), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(n97), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(n95), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(n93), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(n91), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(n89), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(n87), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(n85), .E(n25), .C(i_clk), .RN(i_rst_n), .Q(
        regs[800]) );
  DFEC1 regs_reg_24__31_ ( .D(n147), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(n145), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(n143), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(n141), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(n139), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(n137), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(n135), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(n133), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(n131), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(n129), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(n127), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(n125), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(n123), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(n121), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(n119), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(n117), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(n115), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(n113), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(n111), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(n109), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(n107), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(n105), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(n103), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(n101), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(n99), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(n97), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(n95), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(n93), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(n91), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(n89), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(n87), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(n85), .E(n23), .C(i_clk), .RN(i_rst_n), .Q(
        regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(n148), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(n146), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(n144), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(n142), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(n140), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(n138), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(n136), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(n134), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(n131), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(n130), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(n128), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(n126), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(n123), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(n122), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(n120), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(n118), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(n116), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(n114), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(n112), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(n110), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(n108), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(n106), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(n104), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(n102), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(n100), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(n98), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(n96), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(n94), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(n92), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(n90), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(n88), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(n86), .E(n22), .C(i_clk), .RN(i_rst_n), .Q(
        regs[736]) );
  DFEC1 regs_reg_22__31_ ( .D(n147), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(n145), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(n143), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(n141), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(n139), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(n137), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(n135), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(n133), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(n131), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(n129), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(n127), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(n125), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(n123), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(n121), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(n119), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(n117), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(n115), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(n113), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(n111), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(n109), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(n107), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(n105), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(n103), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(n101), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(n99), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(n97), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(n95), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(n93), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(n91), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(n89), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(n87), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(n85), .E(n21), .C(i_clk), .RN(i_rst_n), .Q(
        regs[704]) );
  DFEC1 regs_reg_21__31_ ( .D(n148), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(n146), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(n144), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(n142), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(n140), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(n138), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(n136), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(n134), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(n131), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(n130), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(n128), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(n125), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(n123), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(n121), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(n119), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(n117), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(n116), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(n114), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(n112), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(n110), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(n108), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(n106), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(n104), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(n101), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(n99), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(n97), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(n95), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(n93), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(n91), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(n89), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(n87), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(n85), .E(n20), .C(i_clk), .RN(i_rst_n), .Q(
        regs[672]) );
  DFEC1 regs_reg_20__31_ ( .D(n148), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(n146), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(n144), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(n142), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(n140), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(n138), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(n136), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(n134), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(n131), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(n130), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(n128), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(n126), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(n123), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(n122), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(n120), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(n118), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(n116), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(n114), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(n112), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(n110), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(n108), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(n106), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(n104), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(n102), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(n100), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(n98), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(n96), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(n94), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(n92), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(n90), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(n88), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(n86), .E(n18), .C(i_clk), .RN(i_rst_n), .Q(
        regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(n147), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(n145), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(n143), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(n141), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(n139), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(n137), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(n135), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(n133), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(n131), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(n129), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(n127), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(n125), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(n123), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(n121), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(n119), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(n117), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(n115), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(n113), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(n111), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(n109), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(n107), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(n105), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(n103), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(n101), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(n99), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(n97), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(n95), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(n93), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(n91), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(n89), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(n87), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(n85), .E(n17), .C(i_clk), .RN(i_rst_n), .Q(
        regs[608]) );
  DFEC1 regs_reg_18__31_ ( .D(n147), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(n145), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(n143), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(n141), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(n139), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(n137), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(n135), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(n133), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(n131), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(n129), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(n127), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(n126), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(n123), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(n122), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(n120), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(n118), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(n115), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(n113), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(n111), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(n109), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(n107), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(n105), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(n103), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(n102), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(n100), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(n98), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(n96), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(n94), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(n92), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(n90), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(n88), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(n86), .E(n16), .C(i_clk), .RN(i_rst_n), .Q(
        regs[576]) );
  DFEC1 regs_reg_17__31_ ( .D(n148), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(n146), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(n144), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(n142), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(n140), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(n138), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(n136), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(n134), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(n131), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(n130), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(n128), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(n126), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(n123), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(n122), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(n120), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(n118), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(n116), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(n114), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(n112), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(n110), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(n108), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(n106), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(n104), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(n102), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(n100), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(n98), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(n96), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(n94), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(n92), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(n90), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(n88), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(n86), .E(n15), .C(i_clk), .RN(i_rst_n), .Q(
        regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(n147), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(n145), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(n143), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(n141), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(n139), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(n137), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(n135), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(n133), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(n131), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(n129), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(n127), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(n125), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(n123), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(n121), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(n119), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(n117), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(n115), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(n113), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(n111), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(n109), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(n107), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(n105), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(n103), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(n101), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(n99), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(n97), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(n95), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(n93), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(n91), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(n89), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(n87), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(n85), .E(n13), .C(i_clk), .RN(i_rst_n), .Q(
        regs[512]) );
  DFEC1 regs_reg_15__31_ ( .D(n147), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(i_data_Rd[30]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(i_data_Rd[29]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(i_data_Rd[28]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(i_data_Rd[27]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(i_data_Rd[26]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(i_data_Rd[25]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(i_data_Rd[24]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(n131), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(i_data_Rd[22]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(n127), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(n125), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(n124), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(n121), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(n119), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(n117), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(n115), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(n111), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(n109), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(n107), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(n105), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(n103), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(n101), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(n99), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(n97), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(n95), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(n93), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(n91), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(n89), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(n87), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(n85), .E(n11), .C(i_clk), .RN(i_rst_n), .Q(
        regs[480]) );
  DFEC1 regs_reg_14__31_ ( .D(n148), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(i_data_Rd[30]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(i_data_Rd[29]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(i_data_Rd[28]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(i_data_Rd[27]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(i_data_Rd[26]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(i_data_Rd[25]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(i_data_Rd[24]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(n132), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(i_data_Rd[22]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(n128), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(n126), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(n123), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(n122), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(n120), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(n118), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(n116), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(n112), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(n110), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(n108), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(n106), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(n104), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(n102), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(n100), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(n98), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(n96), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(n94), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(n92), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(n90), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(n88), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(n86), .E(n9), .C(i_clk), .RN(i_rst_n), .Q(
        regs[448]) );
  DFEC1 regs_reg_13__31_ ( .D(n147), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(i_data_Rd[30]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(i_data_Rd[29]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(i_data_Rd[28]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[444]) );
  DFEC1 regs_reg_13__27_ ( .D(i_data_Rd[27]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(i_data_Rd[26]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(i_data_Rd[25]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(i_data_Rd[24]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(n131), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(i_data_Rd[22]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(n127), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(n125), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(n124), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(n121), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(n119), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(n117), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(n115), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(n111), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(n109), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(n107), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(n105), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(n103), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(n101), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(n99), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(n97), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(n95), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(n93), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(n91), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(n89), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(n87), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(n85), .E(n6), .C(i_clk), .RN(i_rst_n), .Q(
        regs[416]) );
  DFEC1 regs_reg_12__31_ ( .D(n148), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(i_data_Rd[30]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(i_data_Rd[29]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(i_data_Rd[28]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(i_data_Rd[27]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(i_data_Rd[26]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(i_data_Rd[25]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(i_data_Rd[24]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(n132), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(i_data_Rd[22]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(n128), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(n126), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(n123), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(n122), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(n120), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(n118), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(n116), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(n112), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(n110), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(n108), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(n106), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(n104), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(n102), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(n100), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(n98), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(n96), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(n94), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(n92), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(n90), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(n88), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(n86), .E(n5), .C(i_clk), .RN(i_rst_n), .Q(
        regs[384]) );
  DFEC1 regs_reg_11__31_ ( .D(n147), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(i_data_Rd[30]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(i_data_Rd[29]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(i_data_Rd[28]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(i_data_Rd[27]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(i_data_Rd[26]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(i_data_Rd[25]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(i_data_Rd[24]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(n131), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(i_data_Rd[22]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(n127), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(n125), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(n124), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(n121), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(n119), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(n117), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(n115), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(n111), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(n109), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(n107), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(n105), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(n103), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(n101), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(n99), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(n97), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(n95), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(n93), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(n91), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(n89), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(n87), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(n85), .E(n44), .C(i_clk), .RN(i_rst_n), .Q(
        regs[352]) );
  DFEC1 regs_reg_10__31_ ( .D(n148), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(i_data_Rd[30]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(i_data_Rd[29]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(i_data_Rd[28]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(i_data_Rd[27]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(i_data_Rd[26]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(i_data_Rd[25]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(i_data_Rd[24]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(n132), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(i_data_Rd[22]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(n128), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(n126), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(n123), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(n122), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(n120), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(n118), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(n116), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(n112), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(n110), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(n108), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(n106), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(n104), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(n102), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(n100), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(n98), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(n96), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(n94), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(n92), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(n90), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(n88), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(n86), .E(n43), .C(i_clk), .RN(i_rst_n), .Q(
        regs[320]) );
  DFEC1 regs_reg_9__31_ ( .D(n147), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(n146), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(n144), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(n142), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(n140), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(n138), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(n136), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(n134), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(n131), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(n130), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(n127), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(n125), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(n124), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(n121), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(n119), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(n117), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(n115), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(n114), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(n111), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(n109), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(n107), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(n105), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(n103), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(n101), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(n99), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(n97), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(n95), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(n93), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(n91), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(n89), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(n87), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(n85), .E(n42), .C(i_clk), .RN(i_rst_n), .Q(
        regs[288]) );
  DFEC1 regs_reg_8__31_ ( .D(n148), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(n145), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(n143), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(n141), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(n139), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(n137), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(n135), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(n133), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(n132), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(n129), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(n128), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(n126), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(n123), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(n122), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(n120), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(n118), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(n116), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(n113), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(n112), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(n110), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(n108), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(n106), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(n104), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(n102), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(n100), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(n98), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(n96), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(n94), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(n92), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(n90), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(n88), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(n86), .E(n41), .C(i_clk), .RN(i_rst_n), .Q(
        regs[256]) );
  DFEC1 regs_reg_7__31_ ( .D(n148), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(n146), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(n144), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(n142), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(n140), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(n138), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(n136), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(n134), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(n132), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(n130), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(n128), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(n126), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(n124), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(n122), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(n120), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(n118), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(n116), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(n114), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(n112), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(n110), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(n108), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(n106), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(n104), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(n102), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(n100), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(n98), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(n96), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(n94), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(n92), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(n90), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(n88), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(n86), .E(n40), .C(i_clk), .RN(i_rst_n), .Q(
        regs[224]) );
  DFEC1 regs_reg_6__31_ ( .D(n148), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(n146), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(n144), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(n142), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(n140), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(n138), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(n136), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(n134), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(n132), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(n130), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(n128), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(n126), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(n124), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(n122), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(n120), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(n118), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(n116), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(n114), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(n112), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(n110), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(n108), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(n106), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(n104), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(n102), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(n100), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(n98), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(n96), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(n94), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(n92), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(n90), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(n88), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(n86), .E(n39), .C(i_clk), .RN(i_rst_n), .Q(
        regs[192]) );
  DFEC1 regs_reg_5__31_ ( .D(n148), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(n146), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(n144), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(n142), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[188]) );
  DFEC1 regs_reg_5__27_ ( .D(n140), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(n138), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(n136), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(n134), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(n132), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(n130), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(n128), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(n126), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(n124), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(n122), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(n120), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(n118), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(n116), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(n114), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(n112), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(n110), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(n108), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(n106), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(n104), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(n102), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(n100), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(n98), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(n96), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(n94), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(n92), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(n90), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(n88), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(n86), .E(n38), .C(i_clk), .RN(i_rst_n), .Q(
        regs[160]) );
  DFEC1 regs_reg_4__31_ ( .D(n148), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(n146), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(n144), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(n142), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(n140), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(n138), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(n136), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(n134), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(n132), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(n130), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(n128), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(n126), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(n124), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(n122), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(n120), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(n118), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(n116), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(n114), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(n112), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(n110), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(n108), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(n106), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(n104), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(n102), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(n100), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(n98), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(n96), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(n94), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(n92), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(n90), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(n88), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(n86), .E(n37), .C(i_clk), .RN(i_rst_n), .Q(
        regs[128]) );
  DFEC1 regs_reg_3__31_ ( .D(n148), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(n146), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(n144), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(n142), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(n140), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(n138), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(n136), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(n134), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(n132), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(n130), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(n128), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(n126), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(n124), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(n122), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(n120), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(n118), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(n116), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(n114), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(n112), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(n110), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(n108), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(n106), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(n104), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(n102), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(n100), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(n98), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(n96), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(n94), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(n92), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(n90), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(n88), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(n86), .E(n36), .C(i_clk), .RN(i_rst_n), .Q(
        regs[96]) );
  DFEC1 regs_reg_2__31_ ( .D(n148), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(n146), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(n144), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(n142), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(n140), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(n138), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(n136), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(n134), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(n132), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(n130), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(n128), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(n126), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(n124), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(n122), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(n120), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(n118), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(n116), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(n114), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(n112), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(n110), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(n108), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(n106), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(n104), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(n102), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(n100), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(n98), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(n96), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(n94), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(n92), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(n90), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(n88), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(n86), .E(n35), .C(i_clk), .RN(i_rst_n), .Q(
        regs[64]) );
  DFEC1 regs_reg_1__31_ ( .D(n148), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(n146), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(n144), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(n142), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(n140), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(n138), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(n136), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(n134), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(n132), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(n130), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(n128), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(n126), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(n124), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(n122), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(n120), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(n118), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(n116), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(n114), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(n112), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(n110), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(n108), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(n106), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(n104), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(n102), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(n100), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(n98), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(n96), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(n94), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(n92), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(n90), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(n88), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(n86), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[32]) );
  DFEC1 regs_reg_0__31_ ( .D(n148), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(n146), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(n144), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(n142), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(n140), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(n138), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(n136), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(n134), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(n132), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(n130), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(n128), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(n126), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(n124), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(n122), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(n120), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(n118), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(n116), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(n114), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(n112), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(n110), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(n108), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(n106), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(n104), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(n102), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(n100), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(n98), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(n96), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(n94), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(n92), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(n90), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(n88), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(n86), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(regs[0]) );
  NOR31 U2 ( .A(i_addr_Rt[1]), .B(i_addr_Rt[2]), .C(n876), .Q(n1582) );
  NAND22 U3 ( .A(i_addr_Rt[0]), .B(i_addr_Rt[1]), .Q(n875) );
  INV3 U4 ( .A(i_addr_Rt[2]), .Q(n874) );
  NOR21 U5 ( .A(i_addr_Rd[4]), .B(n1596), .Q(n1597) );
  BUF8 U6 ( .A(n861), .Q(n56) );
  BUF8 U7 ( .A(n858), .Q(n12) );
  BUF6 U8 ( .A(n69), .Q(n58) );
  NOR32 U9 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[2]), .C(n151), .Q(n861) );
  BUF8 U10 ( .A(n859), .Q(n66) );
  CLKBU12 U11 ( .A(n862), .Q(n65) );
  BUF8 U12 ( .A(n856), .Q(n76) );
  BUF6 U13 ( .A(n1582), .Q(n33) );
  BUF6 U14 ( .A(n1585), .Q(n55) );
  CLKBU12 U15 ( .A(n1580), .Q(n2) );
  INV3 U16 ( .A(n67), .Q(n1598) );
  NOR21 U17 ( .A(n68), .B(i_addr_Rd[3]), .Q(n67) );
  INV3 U18 ( .A(n1597), .Q(n68) );
  NAND22 U19 ( .A(n1597), .B(i_addr_Rd[3]), .Q(n1608) );
  BUF8 U20 ( .A(i_addr_Rd[0]), .Q(n73) );
  INV3 U21 ( .A(n74), .Q(n1602) );
  INV3 U22 ( .A(n73), .Q(n1603) );
  BUF6 U23 ( .A(i_addr_Rd[2]), .Q(n75) );
  NAND31 U24 ( .A(n75), .B(n1603), .C(n1602), .Q(n1601) );
  NAND31 U25 ( .A(n73), .B(n75), .C(n1602), .Q(n1607) );
  NAND31 U26 ( .A(n74), .B(n75), .C(n1603), .Q(n1606) );
  NAND31 U27 ( .A(n73), .B(n74), .C(n75), .Q(n1605) );
  NAND41 U28 ( .A(n867), .B(n866), .C(n865), .D(n864), .Q(n868) );
  NAND41 U29 ( .A(n197), .B(n196), .C(n195), .D(n194), .Q(n198) );
  NAND41 U30 ( .A(n158), .B(n157), .C(n156), .D(n155), .Q(n166) );
  INV3 U31 ( .A(n160), .Q(n849) );
  NOR22 U32 ( .A(i_addr_Rt[3]), .B(i_addr_Rt[4]), .Q(n1591) );
  NOR22 U33 ( .A(i_addr_Rt[4]), .B(n882), .Q(n1571) );
  NOR31 U34 ( .A(i_addr_Rt[0]), .B(i_addr_Rt[2]), .C(n877), .Q(n1585) );
  AOI220 U35 ( .A(n7), .B(regs[351]), .C(n1584), .D(regs[287]), .Q(n1566) );
  AOI220 U36 ( .A(n7), .B(regs[322]), .C(n1584), .D(regs[258]), .Q(n928) );
  AOI220 U37 ( .A(n7), .B(regs[320]), .C(n1584), .D(regs[256]), .Q(n883) );
  NOR31 U38 ( .A(i_addr_Rt[0]), .B(n877), .C(n874), .Q(n1581) );
  BUF2 U39 ( .A(i_data_Rd[2]), .Q(n90) );
  BUF2 U40 ( .A(i_data_Rd[2]), .Q(n89) );
  BUF2 U41 ( .A(i_data_Rd[17]), .Q(n120) );
  BUF2 U42 ( .A(i_data_Rd[17]), .Q(n119) );
  BUF2 U43 ( .A(i_data_Rd[16]), .Q(n118) );
  BUF2 U44 ( .A(i_data_Rd[16]), .Q(n117) );
  BUF2 U45 ( .A(i_data_Rd[7]), .Q(n100) );
  BUF2 U46 ( .A(i_data_Rd[7]), .Q(n99) );
  BUF2 U47 ( .A(i_data_Rd[20]), .Q(n126) );
  BUF2 U48 ( .A(i_data_Rd[20]), .Q(n125) );
  BUF2 U49 ( .A(i_data_Rd[23]), .Q(n132) );
  BUF2 U50 ( .A(i_data_Rd[23]), .Q(n131) );
  BUF2 U51 ( .A(i_data_Rd[0]), .Q(n86) );
  BUF2 U52 ( .A(i_data_Rd[0]), .Q(n85) );
  BUF2 U53 ( .A(i_data_Rd[1]), .Q(n88) );
  BUF2 U54 ( .A(i_data_Rd[1]), .Q(n87) );
  BUF2 U55 ( .A(i_data_Rd[3]), .Q(n92) );
  BUF2 U56 ( .A(i_data_Rd[3]), .Q(n91) );
  BUF2 U57 ( .A(i_data_Rd[4]), .Q(n94) );
  BUF2 U58 ( .A(i_data_Rd[4]), .Q(n93) );
  BUF2 U59 ( .A(i_data_Rd[5]), .Q(n96) );
  BUF2 U60 ( .A(i_data_Rd[5]), .Q(n95) );
  BUF2 U61 ( .A(i_data_Rd[6]), .Q(n98) );
  BUF2 U62 ( .A(i_data_Rd[6]), .Q(n97) );
  BUF2 U63 ( .A(i_data_Rd[8]), .Q(n102) );
  BUF2 U64 ( .A(i_data_Rd[8]), .Q(n101) );
  BUF2 U65 ( .A(i_data_Rd[9]), .Q(n104) );
  BUF2 U66 ( .A(i_data_Rd[9]), .Q(n103) );
  BUF2 U67 ( .A(i_data_Rd[10]), .Q(n106) );
  BUF2 U68 ( .A(i_data_Rd[10]), .Q(n105) );
  BUF2 U69 ( .A(i_data_Rd[11]), .Q(n108) );
  BUF2 U70 ( .A(i_data_Rd[11]), .Q(n107) );
  BUF2 U71 ( .A(i_data_Rd[12]), .Q(n110) );
  BUF2 U72 ( .A(i_data_Rd[12]), .Q(n109) );
  BUF2 U73 ( .A(i_data_Rd[13]), .Q(n112) );
  BUF2 U74 ( .A(i_data_Rd[13]), .Q(n111) );
  BUF2 U75 ( .A(i_data_Rd[15]), .Q(n116) );
  BUF2 U76 ( .A(i_data_Rd[15]), .Q(n115) );
  BUF2 U77 ( .A(i_data_Rd[18]), .Q(n122) );
  BUF2 U78 ( .A(i_data_Rd[18]), .Q(n121) );
  BUF2 U79 ( .A(i_data_Rd[21]), .Q(n128) );
  BUF2 U80 ( .A(i_data_Rd[21]), .Q(n127) );
  BUF2 U81 ( .A(i_data_Rd[31]), .Q(n148) );
  BUF2 U82 ( .A(i_data_Rd[31]), .Q(n147) );
  BUF2 U83 ( .A(i_data_Rd[19]), .Q(n123) );
  BUF2 U84 ( .A(i_data_Rd[19]), .Q(n124) );
  NOR24 U85 ( .A(i_addr_Rt[2]), .B(n875), .Q(n1583) );
  CLKBU15 U86 ( .A(n1583), .Q(n10) );
  NOR33 U87 ( .A(i_addr_Rt[1]), .B(n876), .C(n874), .Q(n1578) );
  NOR32 U88 ( .A(i_addr_Rt[0]), .B(i_addr_Rt[1]), .C(i_addr_Rt[2]), .Q(n1584)
         );
  BUF6 U89 ( .A(n1584), .Q(n4) );
  NOR22 U90 ( .A(n154), .B(n153), .Q(n862) );
  NOR23 U91 ( .A(n875), .B(n874), .Q(n1579) );
  BUF6 U92 ( .A(n1579), .Q(n1) );
  BUF8 U93 ( .A(n858), .Q(n62) );
  BUF8 U94 ( .A(n858), .Q(n52) );
  INV12 U95 ( .A(n70), .Q(n71) );
  NOR22 U96 ( .A(n882), .B(n889), .Q(n1573) );
  NOR42 U97 ( .A(n73), .B(n74), .C(n75), .D(n1604), .Q(n13) );
  NOR42 U98 ( .A(n75), .B(n74), .C(n1603), .D(n1604), .Q(n15) );
  NOR42 U99 ( .A(n73), .B(n75), .C(n1602), .D(n1604), .Q(n16) );
  NOR42 U100 ( .A(n75), .B(n1602), .C(n1603), .D(n1604), .Q(n17) );
  NOR42 U101 ( .A(n73), .B(n75), .C(n1608), .D(n1602), .Q(n43) );
  NOR42 U102 ( .A(n75), .B(n1603), .C(n1608), .D(n1602), .Q(n44) );
  NOR42 U103 ( .A(n73), .B(n74), .C(n75), .D(n1598), .Q(n32) );
  NOR42 U104 ( .A(n74), .B(n73), .C(n75), .D(n1608), .Q(n41) );
  NOR42 U105 ( .A(n73), .B(n75), .C(n1602), .D(n1598), .Q(n35) );
  NOR42 U106 ( .A(n74), .B(n75), .C(n1603), .D(n1608), .Q(n42) );
  NOR42 U107 ( .A(n75), .B(n74), .C(n1603), .D(n1598), .Q(n34) );
  NOR42 U108 ( .A(n75), .B(n1602), .C(n1603), .D(n1598), .Q(n36) );
  NOR42 U109 ( .A(n73), .B(n74), .C(n75), .D(n1599), .Q(n23) );
  NOR42 U110 ( .A(n75), .B(n74), .C(n1603), .D(n1599), .Q(n25) );
  NOR42 U111 ( .A(n73), .B(n75), .C(n1602), .D(n1599), .Q(n26) );
  NOR42 U112 ( .A(n75), .B(n1602), .C(n1603), .D(n1599), .Q(n27) );
  NOR22 U113 ( .A(n1598), .B(n1607), .Q(n38) );
  NOR22 U114 ( .A(n1598), .B(n1606), .Q(n39) );
  NOR22 U115 ( .A(n1601), .B(n1598), .Q(n37) );
  NOR22 U116 ( .A(n1605), .B(n1598), .Q(n40) );
  NOR22 U117 ( .A(n1605), .B(n1604), .Q(n22) );
  AOI220 U118 ( .A(n66), .B(regs[893]), .C(n12), .D(regs[829]), .Q(n802) );
  AOI220 U119 ( .A(n66), .B(regs[617]), .C(n62), .D(regs[553]), .Q(n372) );
  AOI220 U120 ( .A(n66), .B(regs[360]), .C(n62), .D(regs[296]), .Q(n336) );
  AOI220 U121 ( .A(n66), .B(regs[872]), .C(n62), .D(regs[808]), .Q(n340) );
  AOI220 U122 ( .A(n66), .B(regs[616]), .C(n62), .D(regs[552]), .Q(n350) );
  AOI220 U123 ( .A(n66), .B(regs[871]), .C(n62), .D(regs[807]), .Q(n318) );
  AOI220 U124 ( .A(n66), .B(regs[615]), .C(n62), .D(regs[551]), .Q(n328) );
  AOI220 U125 ( .A(n66), .B(regs[614]), .C(n62), .D(regs[550]), .Q(n306) );
  AOI220 U126 ( .A(n66), .B(regs[877]), .C(n62), .D(regs[813]), .Q(n450) );
  AOI220 U127 ( .A(n66), .B(regs[364]), .C(n62), .D(regs[300]), .Q(n424) );
  AOI220 U128 ( .A(n66), .B(regs[620]), .C(n52), .D(regs[556]), .Q(n438) );
  AOI220 U129 ( .A(n66), .B(regs[363]), .C(n62), .D(regs[299]), .Q(n402) );
  AOI220 U130 ( .A(n66), .B(regs[619]), .C(n62), .D(regs[555]), .Q(n416) );
  AOI220 U131 ( .A(n66), .B(regs[362]), .C(n62), .D(regs[298]), .Q(n380) );
  AOI220 U132 ( .A(n66), .B(regs[874]), .C(n62), .D(regs[810]), .Q(n384) );
  AOI220 U133 ( .A(n66), .B(regs[618]), .C(n62), .D(regs[554]), .Q(n394) );
  AOI220 U134 ( .A(n66), .B(regs[356]), .C(n52), .D(regs[292]), .Q(n248) );
  AOI220 U135 ( .A(n66), .B(regs[868]), .C(n52), .D(regs[804]), .Q(n252) );
  AOI220 U136 ( .A(n66), .B(regs[867]), .C(n52), .D(regs[803]), .Q(n230) );
  AOI220 U137 ( .A(n66), .B(regs[611]), .C(n52), .D(regs[547]), .Q(n240) );
  INV15 U138 ( .A(n70), .Q(n72) );
  AOI220 U139 ( .A(n66), .B(regs[365]), .C(n52), .D(regs[301]), .Q(n446) );
  BUF12 U140 ( .A(n1585), .Q(n7) );
  BUF12 U141 ( .A(n1582), .Q(n8) );
  BUF6 U142 ( .A(n1580), .Q(n24) );
  NOR21 U143 ( .A(i_addr_Rs[2]), .B(n153), .Q(n860) );
  BUF15 U144 ( .A(n861), .Q(n3) );
  NAND41 U145 ( .A(n821), .B(n820), .C(n819), .D(n818), .Q(n827) );
  NAND41 U146 ( .A(n835), .B(n834), .C(n833), .D(n832), .Q(n836) );
  NAND41 U147 ( .A(n825), .B(n824), .C(n823), .D(n822), .Q(n826) );
  NAND41 U148 ( .A(n1261), .B(n1260), .C(n1259), .D(n1258), .Q(n1262) );
  NAND41 U149 ( .A(n1213), .B(n1212), .C(n1211), .D(n1210), .Q(n1219) );
  NAND41 U150 ( .A(n1235), .B(n1234), .C(n1233), .D(n1232), .Q(n1241) );
  NAND41 U151 ( .A(n1245), .B(n1244), .C(n1243), .D(n1242), .Q(n1251) );
  NAND41 U152 ( .A(n1257), .B(n1256), .C(n1255), .D(n1254), .Q(n1263) );
  NAND41 U153 ( .A(n1201), .B(n1200), .C(n1199), .D(n1198), .Q(n1207) );
  NAND41 U154 ( .A(n1205), .B(n1204), .C(n1203), .D(n1202), .Q(n1206) );
  NAND41 U155 ( .A(n1217), .B(n1216), .C(n1215), .D(n1214), .Q(n1218) );
  NAND41 U156 ( .A(n1589), .B(n1588), .C(n1587), .D(n1586), .Q(n1590) );
  NAND41 U157 ( .A(n1223), .B(n1222), .C(n1221), .D(n1220), .Q(n1229) );
  NAND41 U158 ( .A(n1227), .B(n1226), .C(n1225), .D(n1224), .Q(n1228) );
  AOI221 U159 ( .A(n82), .B(regs[448]), .C(n1580), .D(regs[384]), .Q(n885) );
  AOI221 U160 ( .A(n82), .B(regs[450]), .C(n1580), .D(regs[386]), .Q(n930) );
  AOI221 U161 ( .A(n82), .B(regs[449]), .C(n1580), .D(regs[385]), .Q(n908) );
  BUF12 U162 ( .A(n860), .Q(n79) );
  BUF12 U163 ( .A(n1578), .Q(n81) );
  BUF6 U164 ( .A(n1580), .Q(n59) );
  BUF6 U165 ( .A(n1584), .Q(n45) );
  NAND41 U166 ( .A(n843), .B(n842), .C(n841), .D(n840), .Q(n851) );
  NAND41 U167 ( .A(n1191), .B(n1190), .C(n1189), .D(n1188), .Q(n1197) );
  NAND41 U168 ( .A(n1195), .B(n1194), .C(n1193), .D(n1192), .Q(n1196) );
  NAND41 U169 ( .A(n1267), .B(n1266), .C(n1265), .D(n1264), .Q(n1273) );
  NAND41 U170 ( .A(n1279), .B(n1278), .C(n1277), .D(n1276), .Q(n1285) );
  NAND41 U171 ( .A(n1249), .B(n1248), .C(n1247), .D(n1246), .Q(n1250) );
  NAND41 U172 ( .A(n1161), .B(n1160), .C(n1159), .D(n1158), .Q(n1162) );
  NAND41 U173 ( .A(n1157), .B(n1156), .C(n1155), .D(n1154), .Q(n1163) );
  NAND41 U174 ( .A(n1183), .B(n1182), .C(n1181), .D(n1180), .Q(n1184) );
  NAND41 U175 ( .A(n1179), .B(n1178), .C(n1177), .D(n1176), .Q(n1185) );
  NAND41 U176 ( .A(n1173), .B(n1172), .C(n1171), .D(n1170), .Q(n1174) );
  NAND41 U177 ( .A(n1169), .B(n1168), .C(n1167), .D(n1166), .Q(n1175) );
  AOI220 U178 ( .A(n48), .B(regs[985]), .C(n1580), .D(regs[921]), .Q(n1432) );
  AOI220 U179 ( .A(n84), .B(regs[476]), .C(n1580), .D(regs[412]), .Q(n1502) );
  AOI220 U180 ( .A(n83), .B(regs[477]), .C(n1580), .D(regs[413]), .Q(n1524) );
  BUF6 U181 ( .A(n1584), .Q(n47) );
  BUF8 U182 ( .A(n1578), .Q(n49) );
  NOR22 U183 ( .A(n1606), .B(n1599), .Q(n30) );
  BUF12 U184 ( .A(n79), .Q(n14) );
  BUF12 U185 ( .A(n861), .Q(n46) );
  NOR22 U186 ( .A(n1601), .B(n1599), .Q(n28) );
  BUF12 U187 ( .A(n69), .Q(n50) );
  NOR22 U188 ( .A(n1601), .B(n1604), .Q(n18) );
  NOR22 U189 ( .A(n1606), .B(n1604), .Q(n21) );
  NOR22 U190 ( .A(n1607), .B(n1604), .Q(n20) );
  BUF6 U191 ( .A(n1579), .Q(n53) );
  NOR22 U192 ( .A(n1607), .B(n1599), .Q(n29) );
  BUF6 U193 ( .A(n1579), .Q(n19) );
  NOR24 U194 ( .A(i_addr_Rs[2]), .B(n152), .Q(n858) );
  BUF12 U195 ( .A(n857), .Q(n69) );
  NAND33 U196 ( .A(i_con_RegWr), .B(i_addr_Rd[4]), .C(n1600), .Q(n1604) );
  INV3 U197 ( .A(i_addr_Rt[0]), .Q(n876) );
  NAND41 U198 ( .A(n993), .B(n992), .C(n991), .D(n990), .Q(n999) );
  NAND41 U199 ( .A(n997), .B(n996), .C(n995), .D(n994), .Q(n998) );
  NAND41 U200 ( .A(n1015), .B(n1014), .C(n1013), .D(n1012), .Q(n1021) );
  NAND41 U201 ( .A(n1019), .B(n1018), .C(n1017), .D(n1016), .Q(n1020) );
  NAND41 U202 ( .A(n981), .B(n980), .C(n979), .D(n978), .Q(n987) );
  NAND41 U203 ( .A(n1003), .B(n1002), .C(n1001), .D(n1000), .Q(n1009) );
  NAND41 U204 ( .A(n985), .B(n984), .C(n983), .D(n982), .Q(n986) );
  NAND41 U205 ( .A(n1007), .B(n1006), .C(n1005), .D(n1004), .Q(n1008) );
  BUF12 U206 ( .A(n79), .Q(n51) );
  BUF12 U207 ( .A(n76), .Q(n57) );
  BUF6 U208 ( .A(n1581), .Q(n83) );
  INV6 U209 ( .A(n863), .Q(n70) );
  BUF6 U210 ( .A(n1581), .Q(n82) );
  BUF6 U211 ( .A(n1581), .Q(n84) );
  BUF12 U212 ( .A(n66), .Q(n54) );
  NOR22 U213 ( .A(n154), .B(n152), .Q(n863) );
  BUF6 U214 ( .A(n1581), .Q(n48) );
  NOR21 U215 ( .A(n150), .B(n149), .Q(n857) );
  NOR22 U216 ( .A(i_addr_Rt[3]), .B(n889), .Q(n1593) );
  INV3 U217 ( .A(i_addr_Rt[4]), .Q(n889) );
  INV3 U218 ( .A(i_addr_Rt[3]), .Q(n882) );
  NAND22 U219 ( .A(n795), .B(n794), .Q(o_data_Rs[28]) );
  NAND22 U220 ( .A(n817), .B(n816), .Q(o_data_Rs[29]) );
  BUF12 U221 ( .A(n79), .Q(n63) );
  BUF12 U222 ( .A(n76), .Q(n60) );
  BUF12 U223 ( .A(n76), .Q(n64) );
  BUF12 U224 ( .A(n69), .Q(n77) );
  NOR22 U225 ( .A(n1605), .B(n1599), .Q(n31) );
  NAND22 U226 ( .A(n151), .B(n150), .Q(n153) );
  INV3 U227 ( .A(i_addr_Rt[1]), .Q(n877) );
  BUF15 U228 ( .A(i_addr_Rd[1]), .Q(n74) );
  NAND22 U229 ( .A(n873), .B(n872), .Q(o_data_Rs[31]) );
  NAND22 U230 ( .A(n685), .B(n684), .Q(o_data_Rs[23]) );
  NAND22 U231 ( .A(n223), .B(n222), .Q(o_data_Rs[2]) );
  NAND41 U232 ( .A(n1433), .B(n1432), .C(n1431), .D(n1430), .Q(n1439) );
  NAND41 U233 ( .A(n1455), .B(n1454), .C(n1453), .D(n1452), .Q(n1461) );
  NAND41 U234 ( .A(n1491), .B(n1490), .C(n1489), .D(n1488), .Q(n1492) );
  NAND41 U235 ( .A(n1469), .B(n1468), .C(n1467), .D(n1466), .Q(n1470) );
  AOI221 U236 ( .A(n71), .B(regs[946]), .C(n65), .D(regs[914]), .Q(n558) );
  AOI221 U237 ( .A(n72), .B(regs[420]), .C(n65), .D(regs[388]), .Q(n246) );
  AOI221 U238 ( .A(n861), .B(regs[325]), .C(n63), .D(regs[261]), .Q(n269) );
  AOI221 U239 ( .A(n72), .B(regs[932]), .C(n65), .D(regs[900]), .Q(n250) );
  AOI221 U240 ( .A(n71), .B(regs[434]), .C(n65), .D(regs[402]), .Q(n554) );
  AOI221 U241 ( .A(n71), .B(regs[690]), .C(n65), .D(regs[658]), .Q(n568) );
  AOI221 U242 ( .A(n72), .B(regs[419]), .C(n65), .D(regs[387]), .Q(n224) );
  AOI221 U243 ( .A(n72), .B(regs[180]), .C(n65), .D(regs[148]), .Q(n608) );
  AOI221 U244 ( .A(n66), .B(regs[355]), .C(n52), .D(regs[291]), .Q(n226) );
  AOI221 U245 ( .A(n72), .B(regs[692]), .C(n65), .D(regs[660]), .Q(n612) );
  AOI221 U246 ( .A(n72), .B(regs[675]), .C(n65), .D(regs[643]), .Q(n238) );
  AOI221 U247 ( .A(n72), .B(regs[163]), .C(n65), .D(regs[131]), .Q(n234) );
  AOI221 U248 ( .A(n66), .B(regs[99]), .C(n52), .D(regs[35]), .Q(n236) );
  AOI221 U249 ( .A(n71), .B(regs[436]), .C(n65), .D(regs[404]), .Q(n598) );
  AOI221 U250 ( .A(n72), .B(regs[931]), .C(n65), .D(regs[899]), .Q(n228) );
  AOI221 U251 ( .A(n71), .B(regs[435]), .C(n65), .D(regs[403]), .Q(n576) );
  AOI221 U252 ( .A(n71), .B(regs[179]), .C(n65), .D(regs[147]), .Q(n586) );
  BUF12 U253 ( .A(n66), .Q(n78) );
  BUF12 U254 ( .A(n66), .Q(n61) );
  BUF12 U255 ( .A(i_data_Rd[29]), .Q(n144) );
  BUF12 U256 ( .A(i_data_Rd[28]), .Q(n142) );
  BUF12 U257 ( .A(i_data_Rd[14]), .Q(n114) );
  BUF12 U258 ( .A(i_data_Rd[30]), .Q(n145) );
  BUF12 U259 ( .A(i_data_Rd[29]), .Q(n143) );
  BUF12 U260 ( .A(i_data_Rd[24]), .Q(n134) );
  BUF12 U261 ( .A(i_data_Rd[27]), .Q(n140) );
  BUF12 U262 ( .A(i_data_Rd[27]), .Q(n139) );
  BUF12 U263 ( .A(i_data_Rd[26]), .Q(n137) );
  BUF12 U264 ( .A(i_data_Rd[25]), .Q(n135) );
  BUF12 U265 ( .A(i_data_Rd[24]), .Q(n133) );
  BUF12 U266 ( .A(i_data_Rd[22]), .Q(n129) );
  BUF12 U267 ( .A(i_data_Rd[26]), .Q(n138) );
  BUF12 U268 ( .A(i_data_Rd[14]), .Q(n113) );
  BUF12 U269 ( .A(i_data_Rd[22]), .Q(n130) );
  BUF12 U270 ( .A(i_data_Rd[25]), .Q(n136) );
  BUF12 U271 ( .A(i_data_Rd[28]), .Q(n141) );
  BUF12 U272 ( .A(i_data_Rd[30]), .Q(n146) );
  INV3 U273 ( .A(i_addr_Rd[3]), .Q(n1600) );
  AOI221 U274 ( .A(n84), .B(regs[220]), .C(n1580), .D(regs[156]), .Q(n1512) );
  AOI221 U275 ( .A(n83), .B(regs[720]), .C(n2), .D(regs[656]), .Q(n1244) );
  AOI221 U276 ( .A(n82), .B(regs[732]), .C(n1580), .D(regs[668]), .Q(n1508) );
  AOI221 U277 ( .A(n82), .B(regs[710]), .C(n1580), .D(regs[646]), .Q(n1024) );
  AOI221 U278 ( .A(n48), .B(regs[733]), .C(n1580), .D(regs[669]), .Q(n1530) );
  AOI221 U279 ( .A(n48), .B(regs[986]), .C(n2), .D(regs[922]), .Q(n1454) );
  AOI221 U280 ( .A(n83), .B(regs[721]), .C(n2), .D(regs[657]), .Q(n1266) );
  AOI221 U281 ( .A(n83), .B(regs[221]), .C(n1580), .D(regs[157]), .Q(n1534) );
  AOI221 U282 ( .A(n1579), .B(regs[994]), .C(n81), .D(regs[930]), .Q(n927) );
  AOI221 U283 ( .A(n1579), .B(regs[480]), .C(n81), .D(regs[416]), .Q(n886) );
  AOI221 U284 ( .A(n1579), .B(regs[224]), .C(n81), .D(regs[160]), .Q(n897) );
  AOI221 U285 ( .A(n1), .B(regs[737]), .C(n81), .D(regs[673]), .Q(n915) );
  AOI221 U286 ( .A(n1579), .B(regs[481]), .C(n81), .D(regs[417]), .Q(n909) );
  AOI221 U287 ( .A(n1579), .B(regs[993]), .C(n81), .D(regs[929]), .Q(n905) );
  AOI221 U288 ( .A(n1579), .B(regs[482]), .C(n81), .D(regs[418]), .Q(n931) );
  AOI221 U289 ( .A(n1579), .B(regs[225]), .C(n81), .D(regs[161]), .Q(n919) );
  AOI221 U290 ( .A(n71), .B(regs[178]), .C(n80), .D(regs[146]), .Q(n564) );
  AOI221 U291 ( .A(n71), .B(regs[947]), .C(n80), .D(regs[915]), .Q(n580) );
  AOI221 U292 ( .A(n71), .B(regs[691]), .C(n80), .D(regs[659]), .Q(n590) );
  AOI221 U293 ( .A(n56), .B(regs[862]), .C(n79), .D(regs[798]), .Q(n823) );
  AOI221 U294 ( .A(n3), .B(regs[578]), .C(n79), .D(regs[514]), .Q(n217) );
  AOI221 U295 ( .A(n69), .B(regs[995]), .C(n57), .D(regs[963]), .Q(n231) );
  AOI221 U296 ( .A(n69), .B(regs[1011]), .C(n57), .D(regs[979]), .Q(n583) );
  AOI221 U297 ( .A(n69), .B(regs[483]), .C(n57), .D(regs[451]), .Q(n227) );
  AOI221 U298 ( .A(n56), .B(regs[95]), .C(n79), .D(regs[31]), .Q(n853) );
  AOI221 U299 ( .A(n46), .B(regs[66]), .C(n79), .D(regs[2]), .Q(n213) );
  AOI221 U300 ( .A(n69), .B(regs[756]), .C(n57), .D(regs[724]), .Q(n615) );
  AOI221 U301 ( .A(n56), .B(regs[863]), .C(n79), .D(regs[799]), .Q(n845) );
  AOI221 U302 ( .A(n56), .B(regs[351]), .C(n79), .D(regs[287]), .Q(n841) );
  AOI221 U303 ( .A(n69), .B(regs[996]), .C(n57), .D(regs[964]), .Q(n253) );
  AOI221 U304 ( .A(n56), .B(regs[94]), .C(n79), .D(regs[30]), .Q(n829) );
  AOI221 U305 ( .A(n56), .B(regs[350]), .C(n79), .D(regs[286]), .Q(n819) );
  AOI221 U306 ( .A(n69), .B(regs[1010]), .C(n57), .D(regs[978]), .Q(n561) );
  AOI221 U307 ( .A(n46), .B(regs[322]), .C(n79), .D(regs[258]), .Q(n203) );
  AOI221 U308 ( .A(n56), .B(regs[606]), .C(n79), .D(regs[542]), .Q(n833) );
  AOI221 U309 ( .A(n56), .B(regs[607]), .C(n79), .D(regs[543]), .Q(n865) );
  AOI221 U310 ( .A(n54), .B(regs[97]), .C(n858), .D(regs[33]), .Q(n192) );
  AOI221 U311 ( .A(n46), .B(regs[65]), .C(n79), .D(regs[1]), .Q(n191) );
  AOI221 U312 ( .A(n69), .B(regs[1006]), .C(n60), .D(regs[974]), .Q(n473) );
  AOI221 U313 ( .A(n54), .B(regs[609]), .C(n858), .D(regs[545]), .Q(n196) );
  AOI221 U314 ( .A(n46), .B(regs[577]), .C(n79), .D(regs[513]), .Q(n195) );
  AOI221 U315 ( .A(n69), .B(regs[494]), .C(n60), .D(regs[462]), .Q(n469) );
  AOI221 U316 ( .A(n46), .B(regs[576]), .C(n79), .D(regs[512]), .Q(n173) );
  AOI221 U317 ( .A(n54), .B(regs[352]), .C(n858), .D(regs[288]), .Q(n157) );
  AOI221 U318 ( .A(n69), .B(regs[739]), .C(n57), .D(regs[707]), .Q(n241) );
  AOI221 U319 ( .A(n54), .B(regs[608]), .C(n858), .D(regs[544]), .Q(n174) );
  AOI221 U320 ( .A(n69), .B(regs[495]), .C(n60), .D(regs[463]), .Q(n491) );
  AOI221 U321 ( .A(n46), .B(regs[832]), .C(n79), .D(regs[768]), .Q(n162) );
  AOI221 U322 ( .A(n69), .B(regs[1007]), .C(n60), .D(regs[975]), .Q(n495) );
  AOI221 U323 ( .A(n46), .B(regs[64]), .C(n79), .D(regs[0]), .Q(n168) );
  AOI221 U324 ( .A(n69), .B(regs[239]), .C(n60), .D(regs[207]), .Q(n501) );
  AOI221 U325 ( .A(n54), .B(regs[96]), .C(n858), .D(regs[32]), .Q(n169) );
  AOI221 U326 ( .A(n69), .B(regs[244]), .C(n57), .D(regs[212]), .Q(n611) );
  AOI221 U327 ( .A(n46), .B(regs[321]), .C(n79), .D(regs[257]), .Q(n181) );
  AOI221 U328 ( .A(n54), .B(regs[353]), .C(n858), .D(regs[289]), .Q(n182) );
  AOI221 U329 ( .A(n69), .B(regs[237]), .C(n60), .D(regs[205]), .Q(n457) );
  AOI221 U330 ( .A(n69), .B(regs[749]), .C(n60), .D(regs[717]), .Q(n461) );
  AOI221 U331 ( .A(n54), .B(regs[865]), .C(n858), .D(regs[801]), .Q(n186) );
  AOI221 U332 ( .A(n69), .B(regs[227]), .C(n57), .D(regs[195]), .Q(n237) );
  AOI221 U333 ( .A(n46), .B(regs[320]), .C(n79), .D(regs[256]), .Q(n156) );
  AOI221 U334 ( .A(n69), .B(regs[750]), .C(n60), .D(regs[718]), .Q(n483) );
  AOI221 U335 ( .A(n46), .B(regs[833]), .C(n79), .D(regs[769]), .Q(n185) );
  AOI221 U336 ( .A(n69), .B(regs[484]), .C(n57), .D(regs[452]), .Q(n249) );
  NOR22 U337 ( .A(n1608), .B(n1606), .Q(n9) );
  NOR22 U338 ( .A(n1608), .B(n1605), .Q(n11) );
  NOR22 U339 ( .A(n1608), .B(n1607), .Q(n6) );
  BUF12 U340 ( .A(n862), .Q(n80) );
  NOR22 U341 ( .A(n1608), .B(n1601), .Q(n5) );
  NAND33 U342 ( .A(i_addr_Rd[4]), .B(i_con_RegWr), .C(i_addr_Rd[3]), .Q(n1599)
         );
  CLKIN6 U343 ( .A(i_addr_Rs[0]), .Q(n150) );
  INV2 U344 ( .A(i_con_RegWr), .Q(n1596) );
  AOI221 U345 ( .A(n10), .B(regs[97]), .C(n8), .D(regs[33]), .Q(n917) );
  AOI221 U346 ( .A(n82), .B(regs[193]), .C(n1580), .D(regs[129]), .Q(n918) );
  AOI221 U347 ( .A(n10), .B(regs[609]), .C(n8), .D(regs[545]), .Q(n913) );
  AOI221 U348 ( .A(n82), .B(regs[705]), .C(n1580), .D(regs[641]), .Q(n914) );
  AOI221 U349 ( .A(n10), .B(regs[353]), .C(n8), .D(regs[289]), .Q(n907) );
  AOI221 U350 ( .A(n82), .B(regs[197]), .C(n24), .D(regs[133]), .Q(n1006) );
  AOI221 U351 ( .A(n82), .B(regs[709]), .C(n24), .D(regs[645]), .Q(n1002) );
  AOI221 U352 ( .A(n82), .B(regs[453]), .C(n24), .D(regs[389]), .Q(n996) );
  AOI221 U353 ( .A(n82), .B(regs[196]), .C(n24), .D(regs[132]), .Q(n984) );
  AOI221 U354 ( .A(n82), .B(regs[708]), .C(n24), .D(regs[644]), .Q(n980) );
  AOI221 U355 ( .A(n10), .B(regs[356]), .C(n8), .D(regs[292]), .Q(n973) );
  AOI221 U356 ( .A(n82), .B(regs[452]), .C(n2), .D(regs[388]), .Q(n974) );
  AOI221 U357 ( .A(n10), .B(regs[868]), .C(n8), .D(regs[804]), .Q(n969) );
  AOI221 U358 ( .A(n82), .B(regs[964]), .C(n2), .D(regs[900]), .Q(n970) );
  AOI221 U359 ( .A(n7), .B(regs[67]), .C(n47), .D(regs[3]), .Q(n960) );
  AOI221 U360 ( .A(n10), .B(regs[99]), .C(n8), .D(regs[35]), .Q(n961) );
  AOI221 U361 ( .A(n82), .B(regs[195]), .C(n2), .D(regs[131]), .Q(n962) );
  AOI221 U362 ( .A(n10), .B(regs[611]), .C(n8), .D(regs[547]), .Q(n957) );
  AOI221 U363 ( .A(n82), .B(regs[707]), .C(n24), .D(regs[643]), .Q(n958) );
  AOI221 U364 ( .A(n10), .B(regs[355]), .C(n8), .D(regs[291]), .Q(n951) );
  AOI221 U365 ( .A(n10), .B(regs[867]), .C(n8), .D(regs[803]), .Q(n947) );
  AOI221 U366 ( .A(n82), .B(regs[963]), .C(n59), .D(regs[899]), .Q(n948) );
  AOI221 U367 ( .A(n19), .B(regs[230]), .C(n49), .D(regs[166]), .Q(n1029) );
  AOI221 U368 ( .A(n53), .B(regs[742]), .C(n49), .D(regs[678]), .Q(n1025) );
  AOI221 U369 ( .A(n82), .B(regs[454]), .C(n24), .D(regs[390]), .Q(n1018) );
  AOI221 U370 ( .A(n1), .B(regs[486]), .C(n1578), .D(regs[422]), .Q(n1019) );
  AOI221 U371 ( .A(n1), .B(regs[998]), .C(n1578), .D(regs[934]), .Q(n1015) );
  AOI221 U372 ( .A(n55), .B(regs[332]), .C(n4), .D(regs[268]), .Q(n1148) );
  AOI221 U373 ( .A(n84), .B(regs[460]), .C(n59), .D(regs[396]), .Q(n1150) );
  AOI221 U374 ( .A(n19), .B(regs[492]), .C(n49), .D(regs[428]), .Q(n1151) );
  AOI221 U375 ( .A(n55), .B(regs[844]), .C(n4), .D(regs[780]), .Q(n1144) );
  AOI221 U376 ( .A(n48), .B(regs[972]), .C(n2), .D(regs[908]), .Q(n1146) );
  AOI221 U377 ( .A(n19), .B(regs[1004]), .C(n49), .D(regs[940]), .Q(n1147) );
  AOI221 U378 ( .A(n10), .B(regs[96]), .C(n8), .D(regs[32]), .Q(n895) );
  AOI221 U379 ( .A(n82), .B(regs[192]), .C(n1580), .D(regs[128]), .Q(n896) );
  AOI221 U380 ( .A(regs[576]), .B(n7), .C(regs[512]), .D(n47), .Q(n890) );
  AOI221 U381 ( .A(n10), .B(regs[352]), .C(n8), .D(regs[288]), .Q(n884) );
  AOI221 U382 ( .A(n7), .B(regs[832]), .C(n45), .D(regs[768]), .Q(n878) );
  AOI221 U383 ( .A(n7), .B(regs[333]), .C(n45), .D(regs[269]), .Q(n1170) );
  AOI221 U384 ( .A(n83), .B(regs[209]), .C(n2), .D(regs[145]), .Q(n1270) );
  AOI221 U385 ( .A(n7), .B(regs[66]), .C(n47), .D(regs[2]), .Q(n938) );
  AOI221 U386 ( .A(n10), .B(regs[98]), .C(n8), .D(regs[34]), .Q(n939) );
  AOI221 U387 ( .A(n82), .B(regs[194]), .C(n24), .D(regs[130]), .Q(n940) );
  AOI221 U388 ( .A(n10), .B(regs[610]), .C(n8), .D(regs[546]), .Q(n935) );
  AOI221 U389 ( .A(n82), .B(regs[706]), .C(n2), .D(regs[642]), .Q(n936) );
  AOI221 U390 ( .A(n1), .B(regs[738]), .C(n81), .D(regs[674]), .Q(n937) );
  AOI221 U391 ( .A(n10), .B(regs[354]), .C(n8), .D(regs[290]), .Q(n929) );
  AOI221 U392 ( .A(n10), .B(regs[866]), .C(n8), .D(regs[802]), .Q(n925) );
  AOI221 U393 ( .A(n7), .B(regs[82]), .C(n4), .D(regs[18]), .Q(n1290) );
  AOI221 U394 ( .A(n10), .B(regs[114]), .C(n8), .D(regs[50]), .Q(n1291) );
  AOI221 U395 ( .A(n84), .B(regs[210]), .C(n24), .D(regs[146]), .Q(n1292) );
  AOI221 U396 ( .A(n1579), .B(regs[242]), .C(n1578), .D(regs[178]), .Q(n1293)
         );
  AOI221 U397 ( .A(n10), .B(regs[626]), .C(n8), .D(regs[562]), .Q(n1287) );
  AOI221 U398 ( .A(n84), .B(regs[722]), .C(n24), .D(regs[658]), .Q(n1288) );
  AOI221 U399 ( .A(n19), .B(regs[754]), .C(n81), .D(regs[690]), .Q(n1289) );
  AOI221 U400 ( .A(n10), .B(regs[370]), .C(n8), .D(regs[306]), .Q(n1281) );
  AOI221 U401 ( .A(n1579), .B(regs[498]), .C(n1578), .D(regs[434]), .Q(n1283)
         );
  AOI221 U402 ( .A(n7), .B(regs[87]), .C(n47), .D(regs[23]), .Q(n1400) );
  AOI221 U403 ( .A(n84), .B(regs[215]), .C(n24), .D(regs[151]), .Q(n1402) );
  AOI221 U404 ( .A(n1), .B(regs[247]), .C(n49), .D(regs[183]), .Q(n1403) );
  AOI221 U405 ( .A(n7), .B(regs[599]), .C(n47), .D(regs[535]), .Q(n1396) );
  AOI221 U406 ( .A(n84), .B(regs[727]), .C(n24), .D(regs[663]), .Q(n1398) );
  AOI221 U407 ( .A(n1), .B(regs[759]), .C(n81), .D(regs[695]), .Q(n1399) );
  AOI221 U408 ( .A(n7), .B(regs[343]), .C(n47), .D(regs[279]), .Q(n1390) );
  AOI221 U409 ( .A(n1), .B(regs[503]), .C(n1578), .D(regs[439]), .Q(n1393) );
  AOI221 U410 ( .A(n1), .B(regs[1015]), .C(n1578), .D(regs[951]), .Q(n1389) );
  AOI221 U411 ( .A(n7), .B(regs[83]), .C(n4), .D(regs[19]), .Q(n1312) );
  AOI221 U412 ( .A(n10), .B(regs[115]), .C(n8), .D(regs[51]), .Q(n1313) );
  AOI221 U413 ( .A(n84), .B(regs[211]), .C(n59), .D(regs[147]), .Q(n1314) );
  AOI221 U414 ( .A(n1579), .B(regs[243]), .C(n1578), .D(regs[179]), .Q(n1315)
         );
  AOI221 U415 ( .A(n10), .B(regs[627]), .C(n8), .D(regs[563]), .Q(n1309) );
  AOI221 U416 ( .A(n84), .B(regs[723]), .C(n59), .D(regs[659]), .Q(n1310) );
  AOI221 U417 ( .A(n1), .B(regs[755]), .C(n81), .D(regs[691]), .Q(n1311) );
  AOI221 U418 ( .A(n7), .B(regs[339]), .C(n4), .D(regs[275]), .Q(n1302) );
  AOI221 U419 ( .A(n10), .B(regs[371]), .C(n8), .D(regs[307]), .Q(n1303) );
  AOI221 U420 ( .A(n84), .B(regs[467]), .C(n59), .D(regs[403]), .Q(n1304) );
  AOI221 U421 ( .A(n1579), .B(regs[499]), .C(n1578), .D(regs[435]), .Q(n1305)
         );
  AOI221 U422 ( .A(n10), .B(regs[883]), .C(n8), .D(regs[819]), .Q(n1299) );
  AOI221 U423 ( .A(n84), .B(regs[979]), .C(n24), .D(regs[915]), .Q(n1300) );
  AOI221 U424 ( .A(n1579), .B(regs[1011]), .C(n1578), .D(regs[947]), .Q(n1301)
         );
  AOI221 U425 ( .A(n7), .B(regs[86]), .C(n4), .D(regs[22]), .Q(n1378) );
  AOI221 U426 ( .A(n84), .B(regs[214]), .C(n24), .D(regs[150]), .Q(n1380) );
  AOI221 U427 ( .A(n1), .B(regs[246]), .C(n81), .D(regs[182]), .Q(n1381) );
  AOI221 U428 ( .A(n7), .B(regs[598]), .C(n4), .D(regs[534]), .Q(n1374) );
  AOI221 U429 ( .A(n84), .B(regs[726]), .C(n24), .D(regs[662]), .Q(n1376) );
  AOI221 U430 ( .A(n1), .B(regs[758]), .C(n81), .D(regs[694]), .Q(n1377) );
  AOI221 U431 ( .A(n7), .B(regs[342]), .C(n47), .D(regs[278]), .Q(n1368) );
  AOI221 U432 ( .A(n1), .B(regs[502]), .C(n1578), .D(regs[438]), .Q(n1371) );
  AOI221 U433 ( .A(n10), .B(regs[116]), .C(n8), .D(regs[52]), .Q(n1335) );
  AOI221 U434 ( .A(n84), .B(regs[212]), .C(n59), .D(regs[148]), .Q(n1336) );
  AOI221 U435 ( .A(n53), .B(regs[244]), .C(n49), .D(regs[180]), .Q(n1337) );
  AOI221 U436 ( .A(n10), .B(regs[628]), .C(n8), .D(regs[564]), .Q(n1331) );
  AOI221 U437 ( .A(n84), .B(regs[724]), .C(n59), .D(regs[660]), .Q(n1332) );
  AOI221 U438 ( .A(n53), .B(regs[756]), .C(n81), .D(regs[692]), .Q(n1333) );
  AOI221 U439 ( .A(n10), .B(regs[372]), .C(n8), .D(regs[308]), .Q(n1325) );
  AOI221 U440 ( .A(n84), .B(regs[468]), .C(n59), .D(regs[404]), .Q(n1326) );
  AOI221 U441 ( .A(n53), .B(regs[500]), .C(n1578), .D(regs[436]), .Q(n1327) );
  AOI221 U442 ( .A(n10), .B(regs[884]), .C(n8), .D(regs[820]), .Q(n1321) );
  AOI221 U443 ( .A(n84), .B(regs[980]), .C(n59), .D(regs[916]), .Q(n1322) );
  AOI221 U444 ( .A(n1579), .B(regs[1012]), .C(n1578), .D(regs[948]), .Q(n1323)
         );
  AOI221 U445 ( .A(n10), .B(regs[117]), .C(n8), .D(regs[53]), .Q(n1357) );
  AOI221 U446 ( .A(n84), .B(regs[213]), .C(n59), .D(regs[149]), .Q(n1358) );
  AOI221 U447 ( .A(n19), .B(regs[245]), .C(n81), .D(regs[181]), .Q(n1359) );
  AOI221 U448 ( .A(n10), .B(regs[629]), .C(n8), .D(regs[565]), .Q(n1353) );
  AOI221 U449 ( .A(n84), .B(regs[725]), .C(n59), .D(regs[661]), .Q(n1354) );
  AOI221 U450 ( .A(n19), .B(regs[757]), .C(n81), .D(regs[693]), .Q(n1355) );
  AOI221 U451 ( .A(n10), .B(regs[373]), .C(n8), .D(regs[309]), .Q(n1347) );
  AOI221 U452 ( .A(n84), .B(regs[469]), .C(n59), .D(regs[405]), .Q(n1348) );
  AOI221 U453 ( .A(n19), .B(regs[501]), .C(n1578), .D(regs[437]), .Q(n1349) );
  AOI221 U454 ( .A(n10), .B(regs[885]), .C(n8), .D(regs[821]), .Q(n1343) );
  AOI221 U455 ( .A(n84), .B(regs[981]), .C(n59), .D(regs[917]), .Q(n1344) );
  AOI221 U456 ( .A(n19), .B(regs[1013]), .C(n1578), .D(regs[949]), .Q(n1345)
         );
  AOI221 U457 ( .A(n7), .B(regs[94]), .C(n45), .D(regs[30]), .Q(n1554) );
  AOI221 U458 ( .A(n7), .B(regs[606]), .C(n45), .D(regs[542]), .Q(n1550) );
  AOI221 U459 ( .A(n7), .B(regs[350]), .C(n45), .D(regs[286]), .Q(n1544) );
  AOI221 U460 ( .A(n1579), .B(regs[510]), .C(n49), .D(regs[446]), .Q(n1547) );
  AOI221 U461 ( .A(n1581), .B(regs[990]), .C(n2), .D(regs[926]), .Q(n1542) );
  AOI221 U462 ( .A(n1), .B(regs[1022]), .C(n81), .D(regs[958]), .Q(n1543) );
  AOI221 U463 ( .A(n7), .B(regs[607]), .C(n47), .D(regs[543]), .Q(n1574) );
  AOI220 U464 ( .A(n1579), .B(regs[767]), .C(n49), .D(regs[703]), .Q(n1577) );
  AOI221 U465 ( .A(n1579), .B(regs[511]), .C(n49), .D(regs[447]), .Q(n1569) );
  AOI221 U466 ( .A(n7), .B(regs[863]), .C(n47), .D(regs[799]), .Q(n1562) );
  AOI221 U467 ( .A(n1579), .B(regs[1023]), .C(n49), .D(regs[959]), .Q(n1565)
         );
  AOI221 U468 ( .A(n19), .B(regs[231]), .C(n49), .D(regs[167]), .Q(n1051) );
  AOI221 U469 ( .A(n53), .B(regs[743]), .C(n49), .D(regs[679]), .Q(n1047) );
  AOI221 U470 ( .A(n55), .B(regs[327]), .C(n47), .D(regs[263]), .Q(n1038) );
  AOI221 U471 ( .A(n83), .B(regs[455]), .C(n2), .D(regs[391]), .Q(n1040) );
  AOI221 U472 ( .A(n19), .B(regs[487]), .C(n49), .D(regs[423]), .Q(n1041) );
  AOI221 U473 ( .A(n55), .B(regs[839]), .C(n47), .D(regs[775]), .Q(n1034) );
  AOI221 U474 ( .A(n53), .B(regs[999]), .C(n49), .D(regs[935]), .Q(n1037) );
  AOI221 U475 ( .A(n53), .B(regs[232]), .C(n49), .D(regs[168]), .Q(n1073) );
  AOI221 U476 ( .A(n53), .B(regs[744]), .C(n49), .D(regs[680]), .Q(n1069) );
  AOI221 U477 ( .A(n55), .B(regs[328]), .C(n47), .D(regs[264]), .Q(n1060) );
  AOI221 U478 ( .A(n84), .B(regs[456]), .C(n2), .D(regs[392]), .Q(n1062) );
  AOI221 U479 ( .A(n53), .B(regs[488]), .C(n49), .D(regs[424]), .Q(n1063) );
  AOI221 U480 ( .A(n53), .B(regs[1000]), .C(n49), .D(regs[936]), .Q(n1059) );
  AOI221 U481 ( .A(n53), .B(regs[233]), .C(n49), .D(regs[169]), .Q(n1095) );
  AOI221 U482 ( .A(n53), .B(regs[745]), .C(n49), .D(regs[681]), .Q(n1091) );
  AOI221 U483 ( .A(n55), .B(regs[329]), .C(n4), .D(regs[265]), .Q(n1082) );
  AOI221 U484 ( .A(n53), .B(regs[489]), .C(n49), .D(regs[425]), .Q(n1085) );
  AOI221 U485 ( .A(n53), .B(regs[1001]), .C(n49), .D(regs[937]), .Q(n1081) );
  AOI221 U486 ( .A(n48), .B(regs[202]), .C(n2), .D(regs[138]), .Q(n1116) );
  AOI221 U487 ( .A(n53), .B(regs[234]), .C(n49), .D(regs[170]), .Q(n1117) );
  AOI221 U488 ( .A(n83), .B(regs[714]), .C(n2), .D(regs[650]), .Q(n1112) );
  AOI221 U489 ( .A(n19), .B(regs[746]), .C(n49), .D(regs[682]), .Q(n1113) );
  AOI221 U490 ( .A(n55), .B(regs[330]), .C(n45), .D(regs[266]), .Q(n1104) );
  AOI221 U491 ( .A(n53), .B(regs[490]), .C(n49), .D(regs[426]), .Q(n1107) );
  AOI221 U492 ( .A(n53), .B(regs[1002]), .C(n49), .D(regs[938]), .Q(n1103) );
  AOI221 U493 ( .A(n55), .B(regs[75]), .C(n4), .D(regs[11]), .Q(n1136) );
  AOI221 U494 ( .A(n48), .B(regs[203]), .C(n2), .D(regs[139]), .Q(n1138) );
  AOI221 U495 ( .A(n53), .B(regs[235]), .C(n49), .D(regs[171]), .Q(n1139) );
  AOI221 U496 ( .A(n48), .B(regs[715]), .C(n2), .D(regs[651]), .Q(n1134) );
  AOI221 U497 ( .A(n53), .B(regs[747]), .C(n49), .D(regs[683]), .Q(n1135) );
  AOI221 U498 ( .A(n55), .B(regs[331]), .C(n4), .D(regs[267]), .Q(n1126) );
  AOI221 U499 ( .A(n83), .B(regs[459]), .C(n2), .D(regs[395]), .Q(n1128) );
  AOI221 U500 ( .A(n19), .B(regs[491]), .C(n49), .D(regs[427]), .Q(n1129) );
  AOI221 U501 ( .A(n55), .B(regs[843]), .C(n4), .D(regs[779]), .Q(n1122) );
  AOI221 U502 ( .A(n84), .B(regs[971]), .C(n2), .D(regs[907]), .Q(n1124) );
  AOI221 U503 ( .A(n53), .B(regs[1003]), .C(n49), .D(regs[939]), .Q(n1125) );
  AOI221 U504 ( .A(n55), .B(regs[88]), .C(n45), .D(regs[24]), .Q(n1422) );
  AOI221 U505 ( .A(n48), .B(regs[216]), .C(n2), .D(regs[152]), .Q(n1424) );
  AOI221 U506 ( .A(n1579), .B(regs[248]), .C(n81), .D(regs[184]), .Q(n1425) );
  AOI221 U507 ( .A(n55), .B(regs[600]), .C(n45), .D(regs[536]), .Q(n1418) );
  AOI221 U508 ( .A(n48), .B(regs[728]), .C(n2), .D(regs[664]), .Q(n1420) );
  AOI221 U509 ( .A(n19), .B(regs[760]), .C(n81), .D(regs[696]), .Q(n1421) );
  AOI221 U510 ( .A(n55), .B(regs[344]), .C(n45), .D(regs[280]), .Q(n1412) );
  AOI221 U511 ( .A(n48), .B(regs[472]), .C(n2), .D(regs[408]), .Q(n1414) );
  AOI221 U512 ( .A(n1579), .B(regs[504]), .C(n81), .D(regs[440]), .Q(n1415) );
  AOI221 U513 ( .A(n1), .B(regs[252]), .C(n81), .D(regs[188]), .Q(n1513) );
  AOI221 U514 ( .A(n1), .B(regs[764]), .C(n81), .D(regs[700]), .Q(n1509) );
  AOI221 U515 ( .A(n55), .B(regs[348]), .C(n45), .D(regs[284]), .Q(n1500) );
  AOI221 U516 ( .A(n19), .B(regs[1020]), .C(n1578), .D(regs[956]), .Q(n1499)
         );
  AOI221 U517 ( .A(n1), .B(regs[253]), .C(n81), .D(regs[189]), .Q(n1535) );
  AOI221 U518 ( .A(n1), .B(regs[765]), .C(n81), .D(regs[701]), .Q(n1531) );
  AOI221 U519 ( .A(n55), .B(regs[349]), .C(n45), .D(regs[285]), .Q(n1522) );
  AOI221 U520 ( .A(n1), .B(regs[509]), .C(n81), .D(regs[445]), .Q(n1525) );
  AOI221 U521 ( .A(n48), .B(regs[989]), .C(n2), .D(regs[925]), .Q(n1520) );
  AOI221 U522 ( .A(n1), .B(regs[1021]), .C(n81), .D(regs[957]), .Q(n1521) );
  AOI221 U523 ( .A(n48), .B(regs[217]), .C(n2), .D(regs[153]), .Q(n1446) );
  AOI221 U524 ( .A(n1), .B(regs[249]), .C(n81), .D(regs[185]), .Q(n1447) );
  AOI221 U525 ( .A(n55), .B(regs[601]), .C(n47), .D(regs[537]), .Q(n1440) );
  AOI221 U526 ( .A(n48), .B(regs[729]), .C(n2), .D(regs[665]), .Q(n1442) );
  AOI221 U527 ( .A(n53), .B(regs[761]), .C(n81), .D(regs[697]), .Q(n1443) );
  AOI221 U528 ( .A(n55), .B(regs[345]), .C(n45), .D(regs[281]), .Q(n1434) );
  AOI221 U529 ( .A(n48), .B(regs[473]), .C(n2), .D(regs[409]), .Q(n1436) );
  AOI221 U530 ( .A(n53), .B(regs[251]), .C(n81), .D(regs[187]), .Q(n1491) );
  AOI221 U531 ( .A(n55), .B(regs[603]), .C(n45), .D(regs[539]), .Q(n1484) );
  AOI221 U532 ( .A(n53), .B(regs[763]), .C(n81), .D(regs[699]), .Q(n1487) );
  AOI221 U533 ( .A(n55), .B(regs[347]), .C(n45), .D(regs[283]), .Q(n1478) );
  AOI221 U534 ( .A(n53), .B(regs[507]), .C(n1578), .D(regs[443]), .Q(n1481) );
  AOI221 U535 ( .A(n55), .B(regs[859]), .C(n45), .D(regs[795]), .Q(n1474) );
  AOI221 U536 ( .A(n53), .B(regs[1019]), .C(n1578), .D(regs[955]), .Q(n1477)
         );
  AOI221 U537 ( .A(n19), .B(regs[250]), .C(n81), .D(regs[186]), .Q(n1469) );
  AOI221 U538 ( .A(n55), .B(regs[602]), .C(n4), .D(regs[538]), .Q(n1462) );
  AOI221 U539 ( .A(n19), .B(regs[762]), .C(n81), .D(regs[698]), .Q(n1465) );
  AOI221 U540 ( .A(n55), .B(regs[346]), .C(n45), .D(regs[282]), .Q(n1456) );
  AOI221 U541 ( .A(n19), .B(regs[506]), .C(n1578), .D(regs[442]), .Q(n1459) );
  AOI221 U542 ( .A(n55), .B(regs[858]), .C(n1584), .D(regs[794]), .Q(n1452) );
  NOR32 U543 ( .A(i_addr_Rt[0]), .B(i_addr_Rt[1]), .C(n874), .Q(n1580) );
  AOI221 U544 ( .A(n77), .B(regs[736]), .C(n76), .D(regs[704]), .Q(n175) );
  AOI221 U545 ( .A(n71), .B(regs[160]), .C(n80), .D(regs[128]), .Q(n167) );
  AOI221 U546 ( .A(n77), .B(regs[224]), .C(n76), .D(regs[192]), .Q(n170) );
  AOI221 U547 ( .A(n71), .B(regs[928]), .C(n65), .D(regs[896]), .Q(n161) );
  AOI221 U548 ( .A(n54), .B(regs[864]), .C(n858), .D(regs[800]), .Q(n163) );
  AOI221 U549 ( .A(n77), .B(regs[480]), .C(n76), .D(regs[448]), .Q(n158) );
  AOI221 U550 ( .A(n77), .B(regs[758]), .C(n76), .D(regs[726]), .Q(n659) );
  AOI221 U551 ( .A(n78), .B(regs[118]), .C(n12), .D(regs[54]), .Q(n654) );
  AOI221 U552 ( .A(n77), .B(regs[246]), .C(n76), .D(regs[214]), .Q(n655) );
  AOI221 U553 ( .A(n72), .B(regs[950]), .C(n80), .D(regs[918]), .Q(n646) );
  AOI221 U554 ( .A(n78), .B(regs[886]), .C(n12), .D(regs[822]), .Q(n648) );
  AOI221 U555 ( .A(n72), .B(regs[438]), .C(n65), .D(regs[406]), .Q(n642) );
  AOI221 U556 ( .A(n78), .B(regs[374]), .C(n12), .D(regs[310]), .Q(n644) );
  AOI221 U557 ( .A(n72), .B(regs[674]), .C(n80), .D(regs[642]), .Q(n216) );
  AOI221 U558 ( .A(n72), .B(regs[930]), .C(n65), .D(regs[898]), .Q(n206) );
  AOI221 U559 ( .A(n3), .B(regs[834]), .C(n79), .D(regs[770]), .Q(n207) );
  AOI221 U560 ( .A(n71), .B(regs[418]), .C(n80), .D(regs[386]), .Q(n202) );
  AOI221 U561 ( .A(n54), .B(regs[354]), .C(n858), .D(regs[290]), .Q(n204) );
  AOI221 U562 ( .A(n77), .B(regs[482]), .C(n76), .D(regs[450]), .Q(n205) );
  AOI221 U563 ( .A(n77), .B(regs[737]), .C(n76), .D(regs[705]), .Q(n197) );
  AOI221 U564 ( .A(n71), .B(regs[161]), .C(n80), .D(regs[129]), .Q(n190) );
  AOI221 U565 ( .A(n77), .B(regs[225]), .C(n76), .D(regs[193]), .Q(n193) );
  AOI221 U566 ( .A(n71), .B(regs[929]), .C(n80), .D(regs[897]), .Q(n184) );
  AOI221 U567 ( .A(n77), .B(regs[993]), .C(n76), .D(regs[961]), .Q(n187) );
  AOI221 U568 ( .A(n77), .B(regs[481]), .C(n76), .D(regs[449]), .Q(n183) );
  AOI221 U569 ( .A(n72), .B(regs[693]), .C(n65), .D(regs[661]), .Q(n634) );
  AOI221 U570 ( .A(n72), .B(regs[181]), .C(n65), .D(regs[149]), .Q(n630) );
  AOI221 U571 ( .A(n72), .B(regs[949]), .C(n65), .D(regs[917]), .Q(n624) );
  AOI221 U572 ( .A(n72), .B(regs[437]), .C(n65), .D(regs[405]), .Q(n620) );
  AOI221 U573 ( .A(n77), .B(regs[252]), .C(n76), .D(regs[220]), .Q(n787) );
  AOI221 U574 ( .A(n71), .B(regs[956]), .C(n65), .D(regs[924]), .Q(n778) );
  AOI221 U575 ( .A(n77), .B(regs[508]), .C(n76), .D(regs[476]), .Q(n777) );
  AOI221 U576 ( .A(n58), .B(regs[1018]), .C(n76), .D(regs[986]), .Q(n737) );
  AOI221 U577 ( .A(n58), .B(regs[506]), .C(n76), .D(regs[474]), .Q(n733) );
  AOI221 U578 ( .A(n71), .B(regs[191]), .C(n80), .D(regs[159]), .Q(n852) );
  AOI221 U579 ( .A(n77), .B(regs[255]), .C(n76), .D(regs[223]), .Q(n855) );
  AOI221 U580 ( .A(n71), .B(regs[699]), .C(n65), .D(regs[667]), .Q(n766) );
  AOI221 U581 ( .A(n77), .B(regs[763]), .C(n76), .D(regs[731]), .Q(n769) );
  AOI221 U582 ( .A(n77), .B(regs[251]), .C(n76), .D(regs[219]), .Q(n765) );
  AOI221 U583 ( .A(n77), .B(regs[507]), .C(n76), .D(regs[475]), .Q(n755) );
  AOI221 U584 ( .A(n72), .B(regs[953]), .C(n80), .D(regs[921]), .Q(n712) );
  AOI221 U585 ( .A(n72), .B(regs[441]), .C(n80), .D(regs[409]), .Q(n708) );
  AOI221 U586 ( .A(n77), .B(regs[248]), .C(n76), .D(regs[216]), .Q(n699) );
  AOI221 U587 ( .A(n71), .B(regs[952]), .C(n65), .D(regs[920]), .Q(n690) );
  AOI221 U588 ( .A(n77), .B(regs[1016]), .C(n76), .D(regs[984]), .Q(n693) );
  AOI221 U589 ( .A(n77), .B(regs[504]), .C(n76), .D(regs[472]), .Q(n689) );
  AOI221 U590 ( .A(n77), .B(regs[759]), .C(n76), .D(regs[727]), .Q(n681) );
  AOI221 U591 ( .A(n77), .B(regs[247]), .C(n76), .D(regs[215]), .Q(n677) );
  AOI221 U592 ( .A(n71), .B(regs[951]), .C(n65), .D(regs[919]), .Q(n668) );
  AOI221 U593 ( .A(n77), .B(regs[1015]), .C(n76), .D(regs[983]), .Q(n671) );
  AOI221 U594 ( .A(n78), .B(regs[375]), .C(n12), .D(regs[311]), .Q(n666) );
  AOI221 U595 ( .A(n77), .B(regs[503]), .C(n76), .D(regs[471]), .Q(n667) );
  AOI221 U596 ( .A(n50), .B(regs[1021]), .C(n76), .D(regs[989]), .Q(n803) );
  AOI221 U597 ( .A(n77), .B(regs[509]), .C(n76), .D(regs[477]), .Q(n799) );
  AOI221 U598 ( .A(n3), .B(regs[579]), .C(n63), .D(regs[515]), .Q(n239) );
  AOI221 U599 ( .A(n46), .B(regs[67]), .C(n63), .D(regs[3]), .Q(n235) );
  AOI221 U600 ( .A(n3), .B(regs[835]), .C(n63), .D(regs[771]), .Q(n229) );
  AOI221 U601 ( .A(n3), .B(regs[323]), .C(n63), .D(regs[259]), .Q(n225) );
  AOI221 U602 ( .A(n3), .B(regs[596]), .C(n51), .D(regs[532]), .Q(n613) );
  AOI221 U603 ( .A(n78), .B(regs[628]), .C(n52), .D(regs[564]), .Q(n614) );
  AOI221 U604 ( .A(n3), .B(regs[84]), .C(n51), .D(regs[20]), .Q(n609) );
  AOI221 U605 ( .A(n78), .B(regs[116]), .C(n52), .D(regs[52]), .Q(n610) );
  AOI221 U606 ( .A(n861), .B(regs[852]), .C(n51), .D(regs[788]), .Q(n603) );
  AOI221 U607 ( .A(n78), .B(regs[884]), .C(n52), .D(regs[820]), .Q(n604) );
  AOI221 U608 ( .A(n69), .B(regs[1012]), .C(n57), .D(regs[980]), .Q(n605) );
  AOI221 U609 ( .A(n3), .B(regs[340]), .C(n51), .D(regs[276]), .Q(n599) );
  AOI221 U610 ( .A(n54), .B(regs[372]), .C(n52), .D(regs[308]), .Q(n600) );
  AOI221 U611 ( .A(n77), .B(regs[500]), .C(n57), .D(regs[468]), .Q(n601) );
  AOI221 U612 ( .A(n3), .B(regs[589]), .C(n51), .D(regs[525]), .Q(n459) );
  AOI221 U613 ( .A(n54), .B(regs[621]), .C(n52), .D(regs[557]), .Q(n460) );
  AOI221 U614 ( .A(n3), .B(regs[77]), .C(n51), .D(regs[13]), .Q(n455) );
  AOI221 U615 ( .A(n61), .B(regs[109]), .C(n62), .D(regs[45]), .Q(n456) );
  AOI221 U616 ( .A(n72), .B(regs[941]), .C(n65), .D(regs[909]), .Q(n448) );
  AOI221 U617 ( .A(n3), .B(regs[845]), .C(n51), .D(regs[781]), .Q(n449) );
  AOI221 U618 ( .A(n58), .B(regs[1005]), .C(n60), .D(regs[973]), .Q(n451) );
  AOI221 U619 ( .A(n72), .B(regs[429]), .C(n80), .D(regs[397]), .Q(n444) );
  AOI221 U620 ( .A(n3), .B(regs[333]), .C(n51), .D(regs[269]), .Q(n445) );
  AOI221 U621 ( .A(n58), .B(regs[493]), .C(n60), .D(regs[461]), .Q(n447) );
  AOI221 U622 ( .A(n46), .B(regs[591]), .C(n63), .D(regs[527]), .Q(n503) );
  AOI221 U623 ( .A(n61), .B(regs[623]), .C(n62), .D(regs[559]), .Q(n504) );
  AOI221 U624 ( .A(n58), .B(regs[751]), .C(n60), .D(regs[719]), .Q(n505) );
  AOI221 U625 ( .A(n3), .B(regs[79]), .C(n63), .D(regs[15]), .Q(n499) );
  AOI221 U626 ( .A(n61), .B(regs[111]), .C(n62), .D(regs[47]), .Q(n500) );
  AOI221 U627 ( .A(n71), .B(regs[943]), .C(n65), .D(regs[911]), .Q(n492) );
  AOI221 U628 ( .A(n861), .B(regs[847]), .C(n63), .D(regs[783]), .Q(n493) );
  AOI221 U629 ( .A(n61), .B(regs[879]), .C(n62), .D(regs[815]), .Q(n494) );
  AOI221 U630 ( .A(n56), .B(regs[335]), .C(n63), .D(regs[271]), .Q(n489) );
  AOI221 U631 ( .A(n61), .B(regs[367]), .C(n62), .D(regs[303]), .Q(n490) );
  AOI221 U632 ( .A(n3), .B(regs[585]), .C(n14), .D(regs[521]), .Q(n371) );
  AOI221 U633 ( .A(n50), .B(regs[745]), .C(n64), .D(regs[713]), .Q(n373) );
  AOI221 U634 ( .A(n56), .B(regs[73]), .C(n14), .D(regs[9]), .Q(n367) );
  AOI221 U635 ( .A(n66), .B(regs[105]), .C(n52), .D(regs[41]), .Q(n368) );
  AOI221 U636 ( .A(n50), .B(regs[233]), .C(n64), .D(regs[201]), .Q(n369) );
  AOI221 U637 ( .A(n71), .B(regs[937]), .C(n65), .D(regs[905]), .Q(n360) );
  AOI221 U638 ( .A(n861), .B(regs[841]), .C(n14), .D(regs[777]), .Q(n361) );
  AOI221 U639 ( .A(n54), .B(regs[873]), .C(n52), .D(regs[809]), .Q(n362) );
  AOI221 U640 ( .A(n50), .B(regs[1001]), .C(n64), .D(regs[969]), .Q(n363) );
  AOI221 U641 ( .A(n71), .B(regs[425]), .C(n65), .D(regs[393]), .Q(n356) );
  AOI221 U642 ( .A(n3), .B(regs[329]), .C(n14), .D(regs[265]), .Q(n357) );
  AOI221 U643 ( .A(n61), .B(regs[361]), .C(n52), .D(regs[297]), .Q(n358) );
  AOI221 U644 ( .A(n50), .B(regs[489]), .C(n64), .D(regs[457]), .Q(n359) );
  AOI221 U645 ( .A(n71), .B(regs[677]), .C(n65), .D(regs[645]), .Q(n282) );
  AOI221 U646 ( .A(n46), .B(regs[581]), .C(n63), .D(regs[517]), .Q(n283) );
  AOI221 U647 ( .A(n78), .B(regs[613]), .C(n52), .D(regs[549]), .Q(n284) );
  AOI221 U648 ( .A(n50), .B(regs[741]), .C(n57), .D(regs[709]), .Q(n285) );
  AOI221 U649 ( .A(n71), .B(regs[165]), .C(n65), .D(regs[133]), .Q(n278) );
  AOI221 U650 ( .A(n46), .B(regs[69]), .C(n63), .D(regs[5]), .Q(n279) );
  AOI221 U651 ( .A(n78), .B(regs[101]), .C(n52), .D(regs[37]), .Q(n280) );
  AOI221 U652 ( .A(n50), .B(regs[229]), .C(n57), .D(regs[197]), .Q(n281) );
  AOI221 U653 ( .A(n71), .B(regs[933]), .C(n65), .D(regs[901]), .Q(n272) );
  AOI221 U654 ( .A(n3), .B(regs[837]), .C(n63), .D(regs[773]), .Q(n273) );
  AOI221 U655 ( .A(n78), .B(regs[869]), .C(n52), .D(regs[805]), .Q(n274) );
  AOI221 U656 ( .A(n50), .B(regs[997]), .C(n57), .D(regs[965]), .Q(n275) );
  AOI221 U657 ( .A(n71), .B(regs[421]), .C(n65), .D(regs[389]), .Q(n268) );
  AOI221 U658 ( .A(n78), .B(regs[357]), .C(n52), .D(regs[293]), .Q(n270) );
  AOI221 U659 ( .A(n50), .B(regs[485]), .C(n57), .D(regs[453]), .Q(n271) );
  AOI221 U660 ( .A(n3), .B(regs[582]), .C(n79), .D(regs[518]), .Q(n305) );
  AOI221 U661 ( .A(n50), .B(regs[742]), .C(n64), .D(regs[710]), .Q(n307) );
  AOI221 U662 ( .A(n46), .B(regs[70]), .C(n79), .D(regs[6]), .Q(n301) );
  AOI221 U663 ( .A(n78), .B(regs[102]), .C(n62), .D(regs[38]), .Q(n302) );
  AOI221 U664 ( .A(n50), .B(regs[230]), .C(n64), .D(regs[198]), .Q(n303) );
  AOI221 U665 ( .A(n71), .B(regs[934]), .C(n80), .D(regs[902]), .Q(n294) );
  AOI221 U666 ( .A(n78), .B(regs[870]), .C(n62), .D(regs[806]), .Q(n296) );
  AOI221 U667 ( .A(n50), .B(regs[998]), .C(n64), .D(regs[966]), .Q(n297) );
  AOI221 U668 ( .A(n71), .B(regs[422]), .C(n80), .D(regs[390]), .Q(n290) );
  AOI221 U669 ( .A(n78), .B(regs[358]), .C(n62), .D(regs[294]), .Q(n292) );
  AOI221 U670 ( .A(n50), .B(regs[486]), .C(n64), .D(regs[454]), .Q(n293) );
  AOI221 U671 ( .A(n3), .B(regs[586]), .C(n14), .D(regs[522]), .Q(n393) );
  AOI221 U672 ( .A(n50), .B(regs[746]), .C(n64), .D(regs[714]), .Q(n395) );
  AOI221 U673 ( .A(n56), .B(regs[74]), .C(n14), .D(regs[10]), .Q(n389) );
  AOI221 U674 ( .A(n66), .B(regs[106]), .C(n62), .D(regs[42]), .Q(n390) );
  AOI221 U675 ( .A(n50), .B(regs[234]), .C(n64), .D(regs[202]), .Q(n391) );
  AOI221 U676 ( .A(n71), .B(regs[938]), .C(n65), .D(regs[906]), .Q(n382) );
  AOI221 U677 ( .A(n3), .B(regs[842]), .C(n14), .D(regs[778]), .Q(n383) );
  AOI221 U678 ( .A(n50), .B(regs[1002]), .C(n64), .D(regs[970]), .Q(n385) );
  AOI221 U679 ( .A(n71), .B(regs[426]), .C(n65), .D(regs[394]), .Q(n378) );
  AOI221 U680 ( .A(n56), .B(regs[330]), .C(n14), .D(regs[266]), .Q(n379) );
  AOI221 U681 ( .A(n50), .B(regs[490]), .C(n64), .D(regs[458]), .Q(n381) );
  AOI221 U682 ( .A(n71), .B(regs[676]), .C(n65), .D(regs[644]), .Q(n260) );
  AOI221 U683 ( .A(n46), .B(regs[580]), .C(n63), .D(regs[516]), .Q(n261) );
  AOI221 U684 ( .A(n78), .B(regs[612]), .C(n52), .D(regs[548]), .Q(n262) );
  AOI221 U685 ( .A(n50), .B(regs[740]), .C(n57), .D(regs[708]), .Q(n263) );
  AOI221 U686 ( .A(n71), .B(regs[164]), .C(n65), .D(regs[132]), .Q(n256) );
  AOI221 U687 ( .A(n46), .B(regs[68]), .C(n63), .D(regs[4]), .Q(n257) );
  AOI221 U688 ( .A(n78), .B(regs[100]), .C(n52), .D(regs[36]), .Q(n258) );
  AOI221 U689 ( .A(n50), .B(regs[228]), .C(n57), .D(regs[196]), .Q(n259) );
  AOI221 U690 ( .A(n3), .B(regs[836]), .C(n63), .D(regs[772]), .Q(n251) );
  AOI221 U691 ( .A(n3), .B(regs[324]), .C(n63), .D(regs[260]), .Q(n247) );
  AOI221 U692 ( .A(n3), .B(regs[595]), .C(n51), .D(regs[531]), .Q(n591) );
  AOI221 U693 ( .A(n54), .B(regs[627]), .C(n52), .D(regs[563]), .Q(n592) );
  AOI221 U694 ( .A(n77), .B(regs[755]), .C(n57), .D(regs[723]), .Q(n593) );
  AOI221 U695 ( .A(n56), .B(regs[83]), .C(n51), .D(regs[19]), .Q(n587) );
  AOI221 U696 ( .A(n54), .B(regs[115]), .C(n52), .D(regs[51]), .Q(n588) );
  AOI221 U697 ( .A(n77), .B(regs[243]), .C(n57), .D(regs[211]), .Q(n589) );
  AOI221 U698 ( .A(n56), .B(regs[851]), .C(n51), .D(regs[787]), .Q(n581) );
  AOI221 U699 ( .A(n54), .B(regs[883]), .C(n52), .D(regs[819]), .Q(n582) );
  AOI221 U700 ( .A(n56), .B(regs[339]), .C(n51), .D(regs[275]), .Q(n577) );
  AOI221 U701 ( .A(n54), .B(regs[371]), .C(n52), .D(regs[307]), .Q(n578) );
  AOI221 U702 ( .A(n77), .B(regs[499]), .C(n57), .D(regs[467]), .Q(n579) );
  AOI221 U703 ( .A(n56), .B(regs[590]), .C(n51), .D(regs[526]), .Q(n481) );
  AOI221 U704 ( .A(n54), .B(regs[622]), .C(n52), .D(regs[558]), .Q(n482) );
  AOI221 U705 ( .A(n56), .B(regs[78]), .C(n51), .D(regs[14]), .Q(n477) );
  AOI221 U706 ( .A(n54), .B(regs[110]), .C(n52), .D(regs[46]), .Q(n478) );
  AOI221 U707 ( .A(n77), .B(regs[238]), .C(n60), .D(regs[206]), .Q(n479) );
  AOI221 U708 ( .A(n71), .B(regs[942]), .C(n80), .D(regs[910]), .Q(n470) );
  AOI221 U709 ( .A(n861), .B(regs[846]), .C(n51), .D(regs[782]), .Q(n471) );
  AOI221 U710 ( .A(n78), .B(regs[878]), .C(n62), .D(regs[814]), .Q(n472) );
  AOI221 U711 ( .A(n71), .B(regs[430]), .C(n80), .D(regs[398]), .Q(n466) );
  AOI221 U712 ( .A(n3), .B(regs[334]), .C(n51), .D(regs[270]), .Q(n467) );
  AOI221 U713 ( .A(n61), .B(regs[366]), .C(n62), .D(regs[302]), .Q(n468) );
  AOI221 U714 ( .A(n56), .B(regs[594]), .C(n51), .D(regs[530]), .Q(n569) );
  AOI221 U715 ( .A(n54), .B(regs[626]), .C(n52), .D(regs[562]), .Q(n570) );
  AOI221 U716 ( .A(n77), .B(regs[754]), .C(n57), .D(regs[722]), .Q(n571) );
  AOI221 U717 ( .A(n56), .B(regs[82]), .C(n51), .D(regs[18]), .Q(n565) );
  AOI221 U718 ( .A(n61), .B(regs[114]), .C(n52), .D(regs[50]), .Q(n566) );
  AOI221 U719 ( .A(n77), .B(regs[242]), .C(n57), .D(regs[210]), .Q(n567) );
  AOI221 U720 ( .A(n3), .B(regs[850]), .C(n51), .D(regs[786]), .Q(n559) );
  AOI221 U721 ( .A(n61), .B(regs[882]), .C(n52), .D(regs[818]), .Q(n560) );
  AOI221 U722 ( .A(n56), .B(regs[338]), .C(n51), .D(regs[274]), .Q(n555) );
  AOI221 U723 ( .A(n61), .B(regs[370]), .C(n52), .D(regs[306]), .Q(n556) );
  AOI221 U724 ( .A(n77), .B(regs[498]), .C(n57), .D(regs[466]), .Q(n557) );
  AOI221 U725 ( .A(n46), .B(regs[593]), .C(n63), .D(regs[529]), .Q(n547) );
  AOI221 U726 ( .A(n61), .B(regs[625]), .C(n62), .D(regs[561]), .Q(n548) );
  AOI221 U727 ( .A(n58), .B(regs[753]), .C(n60), .D(regs[721]), .Q(n549) );
  AOI221 U728 ( .A(n46), .B(regs[81]), .C(n63), .D(regs[17]), .Q(n543) );
  AOI221 U729 ( .A(n61), .B(regs[113]), .C(n62), .D(regs[49]), .Q(n544) );
  AOI221 U730 ( .A(n58), .B(regs[241]), .C(n60), .D(regs[209]), .Q(n545) );
  AOI221 U731 ( .A(n72), .B(regs[945]), .C(n80), .D(regs[913]), .Q(n536) );
  AOI221 U732 ( .A(n46), .B(regs[849]), .C(n63), .D(regs[785]), .Q(n537) );
  AOI221 U733 ( .A(n61), .B(regs[881]), .C(n62), .D(regs[817]), .Q(n538) );
  AOI221 U734 ( .A(n58), .B(regs[1009]), .C(n60), .D(regs[977]), .Q(n539) );
  AOI221 U735 ( .A(n72), .B(regs[433]), .C(n80), .D(regs[401]), .Q(n532) );
  AOI221 U736 ( .A(n46), .B(regs[337]), .C(n63), .D(regs[273]), .Q(n533) );
  AOI221 U737 ( .A(n61), .B(regs[369]), .C(n62), .D(regs[305]), .Q(n534) );
  AOI221 U738 ( .A(n58), .B(regs[497]), .C(n60), .D(regs[465]), .Q(n535) );
  AOI221 U739 ( .A(n72), .B(regs[679]), .C(n80), .D(regs[647]), .Q(n326) );
  AOI221 U740 ( .A(n3), .B(regs[583]), .C(n79), .D(regs[519]), .Q(n327) );
  AOI221 U741 ( .A(n50), .B(regs[743]), .C(n64), .D(regs[711]), .Q(n329) );
  AOI221 U742 ( .A(n72), .B(regs[167]), .C(n80), .D(regs[135]), .Q(n322) );
  AOI221 U743 ( .A(n3), .B(regs[71]), .C(n79), .D(regs[7]), .Q(n323) );
  AOI221 U744 ( .A(n66), .B(regs[103]), .C(n62), .D(regs[39]), .Q(n324) );
  AOI221 U745 ( .A(n50), .B(regs[231]), .C(n64), .D(regs[199]), .Q(n325) );
  AOI221 U746 ( .A(n72), .B(regs[935]), .C(n80), .D(regs[903]), .Q(n316) );
  AOI221 U747 ( .A(n3), .B(regs[839]), .C(n79), .D(regs[775]), .Q(n317) );
  AOI221 U748 ( .A(n50), .B(regs[999]), .C(n64), .D(regs[967]), .Q(n319) );
  AOI221 U749 ( .A(n72), .B(regs[423]), .C(n80), .D(regs[391]), .Q(n312) );
  AOI221 U750 ( .A(n3), .B(regs[327]), .C(n79), .D(regs[263]), .Q(n313) );
  AOI221 U751 ( .A(n66), .B(regs[359]), .C(n62), .D(regs[295]), .Q(n314) );
  AOI221 U752 ( .A(n50), .B(regs[487]), .C(n64), .D(regs[455]), .Q(n315) );
  AOI221 U753 ( .A(n3), .B(regs[587]), .C(n14), .D(regs[523]), .Q(n415) );
  AOI221 U754 ( .A(n58), .B(regs[747]), .C(n64), .D(regs[715]), .Q(n417) );
  AOI221 U755 ( .A(n3), .B(regs[75]), .C(n14), .D(regs[11]), .Q(n411) );
  AOI221 U756 ( .A(n66), .B(regs[107]), .C(n52), .D(regs[43]), .Q(n412) );
  AOI221 U757 ( .A(n58), .B(regs[235]), .C(n64), .D(regs[203]), .Q(n413) );
  AOI221 U758 ( .A(n72), .B(regs[939]), .C(n65), .D(regs[907]), .Q(n404) );
  AOI221 U759 ( .A(n3), .B(regs[843]), .C(n14), .D(regs[779]), .Q(n405) );
  AOI221 U760 ( .A(n61), .B(regs[875]), .C(n62), .D(regs[811]), .Q(n406) );
  AOI221 U761 ( .A(n58), .B(regs[1003]), .C(n64), .D(regs[971]), .Q(n407) );
  AOI221 U762 ( .A(n71), .B(regs[427]), .C(n65), .D(regs[395]), .Q(n400) );
  AOI221 U763 ( .A(n3), .B(regs[331]), .C(n14), .D(regs[267]), .Q(n401) );
  AOI221 U764 ( .A(n50), .B(regs[491]), .C(n64), .D(regs[459]), .Q(n403) );
  AOI221 U765 ( .A(n72), .B(regs[684]), .C(n80), .D(regs[652]), .Q(n436) );
  AOI221 U766 ( .A(n3), .B(regs[588]), .C(n51), .D(regs[524]), .Q(n437) );
  AOI221 U767 ( .A(n58), .B(regs[748]), .C(n60), .D(regs[716]), .Q(n439) );
  AOI221 U768 ( .A(n72), .B(regs[172]), .C(n80), .D(regs[140]), .Q(n432) );
  AOI221 U769 ( .A(n3), .B(regs[76]), .C(n51), .D(regs[12]), .Q(n433) );
  AOI221 U770 ( .A(n66), .B(regs[108]), .C(n52), .D(regs[44]), .Q(n434) );
  AOI221 U771 ( .A(n58), .B(regs[236]), .C(n60), .D(regs[204]), .Q(n435) );
  AOI221 U772 ( .A(n72), .B(regs[940]), .C(n80), .D(regs[908]), .Q(n426) );
  AOI221 U773 ( .A(n3), .B(regs[844]), .C(n51), .D(regs[780]), .Q(n427) );
  AOI221 U774 ( .A(n54), .B(regs[876]), .C(n52), .D(regs[812]), .Q(n428) );
  AOI221 U775 ( .A(n58), .B(regs[1004]), .C(n60), .D(regs[972]), .Q(n429) );
  AOI221 U776 ( .A(n72), .B(regs[428]), .C(n80), .D(regs[396]), .Q(n422) );
  AOI221 U777 ( .A(n3), .B(regs[332]), .C(n51), .D(regs[268]), .Q(n423) );
  AOI221 U778 ( .A(n58), .B(regs[492]), .C(n60), .D(regs[460]), .Q(n425) );
  AOI221 U779 ( .A(n72), .B(regs[680]), .C(n80), .D(regs[648]), .Q(n348) );
  AOI221 U780 ( .A(n3), .B(regs[584]), .C(n79), .D(regs[520]), .Q(n349) );
  AOI221 U781 ( .A(n50), .B(regs[744]), .C(n64), .D(regs[712]), .Q(n351) );
  AOI221 U782 ( .A(n72), .B(regs[168]), .C(n80), .D(regs[136]), .Q(n344) );
  AOI221 U783 ( .A(n3), .B(regs[72]), .C(n79), .D(regs[8]), .Q(n345) );
  AOI221 U784 ( .A(n66), .B(regs[104]), .C(n62), .D(regs[40]), .Q(n346) );
  AOI221 U785 ( .A(n50), .B(regs[232]), .C(n64), .D(regs[200]), .Q(n347) );
  AOI221 U786 ( .A(n72), .B(regs[936]), .C(n80), .D(regs[904]), .Q(n338) );
  AOI221 U787 ( .A(n3), .B(regs[840]), .C(n79), .D(regs[776]), .Q(n339) );
  AOI221 U788 ( .A(n50), .B(regs[1000]), .C(n64), .D(regs[968]), .Q(n341) );
  AOI221 U789 ( .A(n72), .B(regs[424]), .C(n80), .D(regs[392]), .Q(n334) );
  AOI221 U790 ( .A(n3), .B(regs[328]), .C(n79), .D(regs[264]), .Q(n335) );
  AOI221 U791 ( .A(n50), .B(regs[488]), .C(n64), .D(regs[456]), .Q(n337) );
  AOI221 U792 ( .A(n46), .B(regs[592]), .C(n63), .D(regs[528]), .Q(n525) );
  AOI221 U793 ( .A(n61), .B(regs[624]), .C(n62), .D(regs[560]), .Q(n526) );
  AOI221 U794 ( .A(n58), .B(regs[752]), .C(n60), .D(regs[720]), .Q(n527) );
  NOR24 U795 ( .A(n171), .B(i_addr_Rs[3]), .Q(n869) );
  INV3 U796 ( .A(i_addr_Rs[4]), .Q(n171) );
  NOR24 U797 ( .A(i_addr_Rs[3]), .B(i_addr_Rs[4]), .Q(n870) );
  AOI221 U798 ( .A(n46), .B(regs[80]), .C(n63), .D(regs[16]), .Q(n521) );
  AOI221 U799 ( .A(n61), .B(regs[112]), .C(n62), .D(regs[48]), .Q(n522) );
  AOI221 U800 ( .A(n58), .B(regs[240]), .C(n60), .D(regs[208]), .Q(n523) );
  AOI221 U801 ( .A(n72), .B(regs[944]), .C(n80), .D(regs[912]), .Q(n514) );
  AOI221 U802 ( .A(n46), .B(regs[848]), .C(n63), .D(regs[784]), .Q(n515) );
  AOI221 U803 ( .A(n61), .B(regs[880]), .C(n62), .D(regs[816]), .Q(n516) );
  AOI221 U804 ( .A(n58), .B(regs[1008]), .C(n60), .D(regs[976]), .Q(n517) );
  NAND22 U805 ( .A(i_addr_Rs[4]), .B(i_addr_Rs[3]), .Q(n160) );
  NOR24 U806 ( .A(n159), .B(i_addr_Rs[4]), .Q(n850) );
  INV3 U807 ( .A(i_addr_Rs[3]), .Q(n159) );
  AOI221 U808 ( .A(n46), .B(regs[336]), .C(n63), .D(regs[272]), .Q(n511) );
  AOI221 U809 ( .A(n61), .B(regs[368]), .C(n62), .D(regs[304]), .Q(n512) );
  AOI221 U810 ( .A(n58), .B(regs[496]), .C(n60), .D(regs[464]), .Q(n513) );
  AOI221 U811 ( .A(n7), .B(regs[324]), .C(n47), .D(regs[260]), .Q(n972) );
  AOI221 U812 ( .A(n7), .B(regs[323]), .C(n47), .D(regs[259]), .Q(n950) );
  AOI221 U813 ( .A(n82), .B(regs[451]), .C(n24), .D(regs[387]), .Q(n952) );
  AOI221 U814 ( .A(n7), .B(regs[835]), .C(n47), .D(regs[771]), .Q(n946) );
  AOI221 U815 ( .A(n1579), .B(regs[992]), .C(n49), .D(regs[928]), .Q(n881) );
  AOI221 U816 ( .A(n7), .B(regs[335]), .C(n4), .D(regs[271]), .Q(n1214) );
  AOI221 U817 ( .A(n7), .B(regs[337]), .C(n4), .D(regs[273]), .Q(n1258) );
  AOI221 U818 ( .A(n7), .B(regs[334]), .C(n45), .D(regs[270]), .Q(n1192) );
  AOI221 U819 ( .A(n84), .B(regs[983]), .C(n24), .D(regs[919]), .Q(n1388) );
  AOI221 U820 ( .A(n10), .B(regs[886]), .C(n8), .D(regs[822]), .Q(n1365) );
  AOI221 U821 ( .A(n53), .B(regs[1014]), .C(n1578), .D(regs[950]), .Q(n1367)
         );
  AOI221 U822 ( .A(n83), .B(regs[199]), .C(n2), .D(regs[135]), .Q(n1050) );
  AOI221 U823 ( .A(n48), .B(regs[711]), .C(n2), .D(regs[647]), .Q(n1046) );
  AOI221 U824 ( .A(n82), .B(regs[200]), .C(n2), .D(regs[136]), .Q(n1072) );
  AOI221 U825 ( .A(n48), .B(regs[712]), .C(n2), .D(regs[648]), .Q(n1068) );
  AOI221 U826 ( .A(n48), .B(regs[201]), .C(n2), .D(regs[137]), .Q(n1094) );
  AOI221 U827 ( .A(n84), .B(regs[713]), .C(n2), .D(regs[649]), .Q(n1090) );
  AOI221 U828 ( .A(n1581), .B(regs[457]), .C(n2), .D(regs[393]), .Q(n1084) );
  AOI221 U829 ( .A(n48), .B(regs[458]), .C(n2), .D(regs[394]), .Q(n1106) );
  AOI221 U830 ( .A(n1), .B(regs[1016]), .C(n1578), .D(regs[952]), .Q(n1411) );
  AOI221 U831 ( .A(n1), .B(regs[508]), .C(n81), .D(regs[444]), .Q(n1503) );
  AOI221 U832 ( .A(n55), .B(regs[860]), .C(n47), .D(regs[796]), .Q(n1496) );
  AOI221 U833 ( .A(n55), .B(regs[861]), .C(n45), .D(regs[797]), .Q(n1518) );
  AOI221 U834 ( .A(n1579), .B(regs[505]), .C(n81), .D(regs[441]), .Q(n1437) );
  AOI221 U835 ( .A(n72), .B(regs[190]), .C(n80), .D(regs[158]), .Q(n828) );
  AOI221 U836 ( .A(n58), .B(regs[1022]), .C(n76), .D(regs[990]), .Q(n825) );
  AOI221 U837 ( .A(n58), .B(regs[510]), .C(n76), .D(regs[478]), .Q(n821) );
  AOI221 U838 ( .A(n58), .B(regs[250]), .C(n76), .D(regs[218]), .Q(n743) );
  AOI221 U839 ( .A(n54), .B(regs[639]), .C(n858), .D(regs[575]), .Q(n866) );
  AOI221 U840 ( .A(n72), .B(regs[701]), .C(n65), .D(regs[669]), .Q(n810) );
  AOI221 U841 ( .A(n7), .B(regs[836]), .C(n47), .D(regs[772]), .Q(n968) );
  AOI221 U842 ( .A(n48), .B(regs[198]), .C(n24), .D(regs[134]), .Q(n1028) );
  AOI221 U843 ( .A(n83), .B(regs[208]), .C(n2), .D(regs[144]), .Q(n1248) );
  AOI221 U844 ( .A(n84), .B(regs[984]), .C(n24), .D(regs[920]), .Q(n1410) );
  AOI221 U845 ( .A(n1579), .B(regs[1017]), .C(n81), .D(regs[953]), .Q(n1433)
         );
  AOI221 U846 ( .A(n1579), .B(regs[1018]), .C(n81), .D(regs[954]), .Q(n1455)
         );
  AOI221 U847 ( .A(n50), .B(regs[762]), .C(n76), .D(regs[730]), .Q(n747) );
  AOI221 U848 ( .A(n58), .B(regs[760]), .C(n76), .D(regs[728]), .Q(n703) );
  AOI221 U849 ( .A(regs[736]), .B(n19), .C(regs[672]), .D(n49), .Q(n893) );
  AOI221 U850 ( .A(n58), .B(regs[766]), .C(n76), .D(regs[734]), .Q(n835) );
  AOI221 U851 ( .A(n50), .B(regs[764]), .C(n76), .D(regs[732]), .Q(n791) );
  AOI221 U852 ( .A(n50), .B(regs[511]), .C(n76), .D(regs[479]), .Q(n843) );
  AOI221 U853 ( .A(n50), .B(regs[249]), .C(n76), .D(regs[217]), .Q(n721) );
  AOI221 U854 ( .A(n58), .B(regs[253]), .C(n76), .D(regs[221]), .Q(n809) );
  AOI221 U855 ( .A(n83), .B(regs[222]), .C(n59), .D(regs[158]), .Q(n1556) );
  AOI221 U856 ( .A(n82), .B(regs[734]), .C(n59), .D(regs[670]), .Q(n1552) );
  AOI221 U857 ( .A(n55), .B(regs[862]), .C(n45), .D(regs[798]), .Q(n1540) );
  AOI221 U858 ( .A(n55), .B(regs[93]), .C(n45), .D(regs[29]), .Q(n1532) );
  AOI221 U859 ( .A(n48), .B(regs[731]), .C(n2), .D(regs[667]), .Q(n1486) );
  AOI221 U860 ( .A(n48), .B(regs[730]), .C(n2), .D(regs[666]), .Q(n1464) );
  AOI220 U861 ( .A(n861), .B(regs[838]), .C(n79), .D(regs[774]), .Q(n295) );
  AOI220 U862 ( .A(n861), .B(regs[326]), .C(n79), .D(regs[262]), .Q(n291) );
  NOR21 U863 ( .A(i_addr_Rs[0]), .B(n149), .Q(n856) );
  AOI221 U864 ( .A(n1573), .B(n999), .C(n1571), .D(n998), .Q(n1011) );
  AOI221 U865 ( .A(n1573), .B(n1021), .C(n1571), .D(n1020), .Q(n1033) );
  AOI221 U866 ( .A(n1593), .B(n1163), .C(n1591), .D(n1162), .Q(n1164) );
  AOI221 U867 ( .A(n1573), .B(n1153), .C(n1571), .D(n1152), .Q(n1165) );
  AOI221 U868 ( .A(n1573), .B(n1241), .C(n1571), .D(n1240), .Q(n1253) );
  AOI221 U869 ( .A(n1573), .B(n1175), .C(n1571), .D(n1174), .Q(n1187) );
  AOI221 U870 ( .A(n1573), .B(n1219), .C(n1571), .D(n1218), .Q(n1231) );
  AOI221 U871 ( .A(n1573), .B(n1263), .C(n1571), .D(n1262), .Q(n1275) );
  AOI221 U872 ( .A(n1593), .B(n1207), .C(n1591), .D(n1206), .Q(n1208) );
  AOI221 U873 ( .A(n1573), .B(n1285), .C(n1571), .D(n1284), .Q(n1297) );
  AOI221 U874 ( .A(n1573), .B(n1549), .C(n1571), .D(n1548), .Q(n1561) );
  AOI221 U875 ( .A(n1573), .B(n1572), .C(n1571), .D(n1570), .Q(n1595) );
  AOI221 U876 ( .A(n1573), .B(n1043), .C(n1571), .D(n1042), .Q(n1055) );
  AOI221 U877 ( .A(n1573), .B(n1065), .C(n1571), .D(n1064), .Q(n1077) );
  AOI221 U878 ( .A(n1573), .B(n1087), .C(n1571), .D(n1086), .Q(n1099) );
  AOI221 U879 ( .A(n1593), .B(n1119), .C(n1591), .D(n1118), .Q(n1120) );
  AOI221 U880 ( .A(n1573), .B(n1109), .C(n1571), .D(n1108), .Q(n1121) );
  AOI221 U881 ( .A(n1593), .B(n1141), .C(n1591), .D(n1140), .Q(n1142) );
  AOI221 U882 ( .A(n1573), .B(n1131), .C(n1571), .D(n1130), .Q(n1143) );
  AOI221 U883 ( .A(n177), .B(n870), .C(n869), .D(n176), .Q(n178) );
  AOI221 U884 ( .A(n166), .B(n850), .C(n849), .D(n165), .Q(n179) );
  AOI220 U885 ( .A(n69), .B(regs[992]), .C(n76), .D(regs[960]), .Q(n164) );
  AOI221 U886 ( .A(n661), .B(n870), .C(n869), .D(n660), .Q(n662) );
  AOI221 U887 ( .A(n651), .B(n850), .C(n849), .D(n650), .Q(n663) );
  AOI220 U888 ( .A(n69), .B(regs[738]), .C(n76), .D(regs[706]), .Q(n219) );
  AOI220 U889 ( .A(n69), .B(regs[226]), .C(n76), .D(regs[194]), .Q(n215) );
  AOI220 U890 ( .A(n69), .B(regs[994]), .C(n76), .D(regs[962]), .Q(n209) );
  AOI221 U891 ( .A(n199), .B(n870), .C(n869), .D(n198), .Q(n200) );
  AOI221 U892 ( .A(n189), .B(n850), .C(n849), .D(n188), .Q(n201) );
  AOI221 U893 ( .A(n639), .B(n870), .C(n869), .D(n638), .Q(n640) );
  AOI220 U894 ( .A(n69), .B(regs[757]), .C(n76), .D(regs[725]), .Q(n637) );
  AOI220 U895 ( .A(n69), .B(regs[245]), .C(n76), .D(regs[213]), .Q(n633) );
  AOI221 U896 ( .A(n629), .B(n850), .C(n849), .D(n628), .Q(n641) );
  AOI220 U897 ( .A(n69), .B(regs[1013]), .C(n76), .D(regs[981]), .Q(n627) );
  AOI220 U898 ( .A(n69), .B(regs[501]), .C(n76), .D(regs[469]), .Q(n623) );
  AOI221 U899 ( .A(n837), .B(n870), .C(n869), .D(n836), .Q(n838) );
  AOI220 U900 ( .A(n69), .B(regs[254]), .C(n76), .D(regs[222]), .Q(n831) );
  AOI221 U901 ( .A(n827), .B(n850), .C(n849), .D(n826), .Q(n839) );
  AOI221 U902 ( .A(n793), .B(n870), .C(n869), .D(n792), .Q(n794) );
  AOI221 U903 ( .A(n783), .B(n850), .C(n849), .D(n782), .Q(n795) );
  AOI220 U904 ( .A(n69), .B(regs[1020]), .C(n76), .D(regs[988]), .Q(n781) );
  AOI221 U905 ( .A(n749), .B(n870), .C(n869), .D(n748), .Q(n750) );
  AOI221 U906 ( .A(n739), .B(n850), .C(n849), .D(n738), .Q(n751) );
  AOI221 U907 ( .A(n871), .B(n870), .C(n869), .D(n868), .Q(n872) );
  AOI221 U908 ( .A(n851), .B(n850), .C(n849), .D(n848), .Q(n873) );
  AOI220 U909 ( .A(n69), .B(regs[1023]), .C(n76), .D(regs[991]), .Q(n847) );
  AOI221 U910 ( .A(n771), .B(n870), .C(n869), .D(n770), .Q(n772) );
  AOI221 U911 ( .A(n761), .B(n850), .C(n849), .D(n760), .Q(n773) );
  AOI220 U912 ( .A(n69), .B(regs[1019]), .C(n76), .D(regs[987]), .Q(n759) );
  AOI221 U913 ( .A(n727), .B(n870), .C(n869), .D(n726), .Q(n728) );
  AOI220 U914 ( .A(n69), .B(regs[761]), .C(n76), .D(regs[729]), .Q(n725) );
  AOI221 U915 ( .A(n717), .B(n850), .C(n849), .D(n716), .Q(n729) );
  AOI220 U916 ( .A(n69), .B(regs[1017]), .C(n76), .D(regs[985]), .Q(n715) );
  AOI220 U917 ( .A(n69), .B(regs[505]), .C(n76), .D(regs[473]), .Q(n711) );
  AOI221 U918 ( .A(n705), .B(n870), .C(n869), .D(n704), .Q(n706) );
  AOI221 U919 ( .A(n695), .B(n850), .C(n849), .D(n694), .Q(n707) );
  AOI221 U920 ( .A(n683), .B(n870), .C(n869), .D(n682), .Q(n684) );
  AOI221 U921 ( .A(n673), .B(n850), .C(n849), .D(n672), .Q(n685) );
  AOI221 U922 ( .A(n815), .B(n870), .C(n869), .D(n814), .Q(n816) );
  AOI220 U923 ( .A(n69), .B(regs[765]), .C(n76), .D(regs[733]), .Q(n813) );
  AOI221 U924 ( .A(n805), .B(n850), .C(n849), .D(n804), .Q(n817) );
  AOI221 U925 ( .A(n243), .B(n870), .C(n869), .D(n242), .Q(n244) );
  AOI221 U926 ( .A(n233), .B(n850), .C(n849), .D(n232), .Q(n245) );
  AOI221 U927 ( .A(n617), .B(n870), .C(n869), .D(n616), .Q(n618) );
  AOI221 U928 ( .A(n607), .B(n850), .C(n849), .D(n606), .Q(n619) );
  AOI221 U929 ( .A(n463), .B(n870), .C(n869), .D(n462), .Q(n464) );
  AOI221 U930 ( .A(n453), .B(n850), .C(n849), .D(n452), .Q(n465) );
  AOI221 U931 ( .A(n507), .B(n870), .C(n869), .D(n506), .Q(n508) );
  AOI221 U932 ( .A(n497), .B(n850), .C(n849), .D(n496), .Q(n509) );
  AOI221 U933 ( .A(n375), .B(n870), .C(n869), .D(n374), .Q(n376) );
  AOI221 U934 ( .A(n365), .B(n850), .C(n849), .D(n364), .Q(n377) );
  AOI221 U935 ( .A(n287), .B(n870), .C(n869), .D(n286), .Q(n288) );
  AOI221 U936 ( .A(n277), .B(n850), .C(n849), .D(n276), .Q(n289) );
  AOI221 U937 ( .A(n309), .B(n870), .C(n869), .D(n308), .Q(n310) );
  AOI221 U938 ( .A(n299), .B(n850), .C(n849), .D(n298), .Q(n311) );
  AOI221 U939 ( .A(n397), .B(n870), .C(n869), .D(n396), .Q(n398) );
  AOI221 U940 ( .A(n387), .B(n850), .C(n849), .D(n386), .Q(n399) );
  AOI221 U941 ( .A(n265), .B(n870), .C(n869), .D(n264), .Q(n266) );
  AOI221 U942 ( .A(n255), .B(n850), .C(n849), .D(n254), .Q(n267) );
  AOI221 U943 ( .A(n595), .B(n870), .C(n869), .D(n594), .Q(n596) );
  AOI221 U944 ( .A(n585), .B(n850), .C(n849), .D(n584), .Q(n597) );
  AOI221 U945 ( .A(n485), .B(n870), .C(n869), .D(n484), .Q(n486) );
  AOI221 U946 ( .A(n475), .B(n850), .C(n849), .D(n474), .Q(n487) );
  AOI221 U947 ( .A(n573), .B(n870), .C(n869), .D(n572), .Q(n574) );
  AOI221 U948 ( .A(n563), .B(n850), .C(n849), .D(n562), .Q(n575) );
  AOI221 U949 ( .A(n551), .B(n870), .C(n869), .D(n550), .Q(n552) );
  AOI221 U950 ( .A(n541), .B(n850), .C(n849), .D(n540), .Q(n553) );
  AOI221 U951 ( .A(n331), .B(n870), .C(n869), .D(n330), .Q(n332) );
  AOI221 U952 ( .A(n321), .B(n850), .C(n849), .D(n320), .Q(n333) );
  AOI221 U953 ( .A(n419), .B(n870), .C(n869), .D(n418), .Q(n420) );
  AOI221 U954 ( .A(n409), .B(n850), .C(n849), .D(n408), .Q(n421) );
  AOI221 U955 ( .A(n441), .B(n870), .C(n869), .D(n440), .Q(n442) );
  AOI221 U956 ( .A(n431), .B(n850), .C(n849), .D(n430), .Q(n443) );
  AOI221 U957 ( .A(n353), .B(n870), .C(n869), .D(n352), .Q(n354) );
  AOI221 U958 ( .A(n343), .B(n850), .C(n849), .D(n342), .Q(n355) );
  AOI221 U959 ( .A(n529), .B(n870), .C(n869), .D(n528), .Q(n530) );
  AOI221 U960 ( .A(n519), .B(n850), .C(n849), .D(n518), .Q(n531) );
  NAND22 U961 ( .A(n923), .B(n922), .Q(o_data_Rt[1]) );
  AOI221 U962 ( .A(n1593), .B(n921), .C(n1591), .D(n920), .Q(n922) );
  NAND41 U963 ( .A(n919), .B(n918), .C(n917), .D(n916), .Q(n920) );
  AOI221 U964 ( .A(n7), .B(regs[65]), .C(n45), .D(regs[1]), .Q(n916) );
  NAND41 U965 ( .A(n915), .B(n914), .C(n913), .D(n912), .Q(n921) );
  AOI221 U966 ( .A(n7), .B(regs[577]), .C(n47), .D(regs[513]), .Q(n912) );
  AOI221 U967 ( .A(n1573), .B(n911), .C(n1571), .D(n910), .Q(n923) );
  NAND41 U968 ( .A(n909), .B(n908), .C(n907), .D(n906), .Q(n910) );
  AOI221 U969 ( .A(n7), .B(regs[321]), .C(n1584), .D(regs[257]), .Q(n906) );
  NAND41 U970 ( .A(n905), .B(n904), .C(n903), .D(n902), .Q(n911) );
  AOI221 U971 ( .A(n7), .B(regs[833]), .C(n4), .D(regs[769]), .Q(n902) );
  AOI221 U972 ( .A(n10), .B(regs[865]), .C(n8), .D(regs[801]), .Q(n903) );
  AOI221 U973 ( .A(n82), .B(regs[961]), .C(n1580), .D(regs[897]), .Q(n904) );
  NAND22 U974 ( .A(n1011), .B(n1010), .Q(o_data_Rt[5]) );
  AOI221 U975 ( .A(n1593), .B(n1009), .C(n1591), .D(n1008), .Q(n1010) );
  AOI221 U976 ( .A(n7), .B(regs[69]), .C(n47), .D(regs[5]), .Q(n1004) );
  AOI221 U977 ( .A(n10), .B(regs[101]), .C(n8), .D(regs[37]), .Q(n1005) );
  AOI221 U978 ( .A(n1), .B(regs[229]), .C(n49), .D(regs[165]), .Q(n1007) );
  AOI221 U979 ( .A(n7), .B(regs[581]), .C(n47), .D(regs[517]), .Q(n1000) );
  AOI221 U980 ( .A(n10), .B(regs[613]), .C(n8), .D(regs[549]), .Q(n1001) );
  AOI221 U981 ( .A(n1), .B(regs[741]), .C(n81), .D(regs[677]), .Q(n1003) );
  AOI221 U982 ( .A(n7), .B(regs[325]), .C(n47), .D(regs[261]), .Q(n994) );
  AOI221 U983 ( .A(n10), .B(regs[357]), .C(n8), .D(regs[293]), .Q(n995) );
  AOI221 U984 ( .A(n1), .B(regs[485]), .C(n1578), .D(regs[421]), .Q(n997) );
  AOI221 U985 ( .A(n7), .B(regs[837]), .C(n47), .D(regs[773]), .Q(n990) );
  AOI221 U986 ( .A(n10), .B(regs[869]), .C(n8), .D(regs[805]), .Q(n991) );
  AOI221 U987 ( .A(n82), .B(regs[965]), .C(n24), .D(regs[901]), .Q(n992) );
  AOI221 U988 ( .A(n1), .B(regs[997]), .C(n1578), .D(regs[933]), .Q(n993) );
  NAND22 U989 ( .A(n989), .B(n988), .Q(o_data_Rt[4]) );
  AOI221 U990 ( .A(n1593), .B(n987), .C(n1591), .D(n986), .Q(n988) );
  AOI221 U991 ( .A(n7), .B(regs[68]), .C(n47), .D(regs[4]), .Q(n982) );
  AOI221 U992 ( .A(n10), .B(regs[100]), .C(n8), .D(regs[36]), .Q(n983) );
  AOI221 U993 ( .A(n1), .B(regs[228]), .C(n81), .D(regs[164]), .Q(n985) );
  AOI221 U994 ( .A(n7), .B(regs[580]), .C(n47), .D(regs[516]), .Q(n978) );
  AOI221 U995 ( .A(n10), .B(regs[612]), .C(n8), .D(regs[548]), .Q(n979) );
  AOI221 U996 ( .A(n1), .B(regs[740]), .C(n81), .D(regs[676]), .Q(n981) );
  AOI221 U997 ( .A(n1573), .B(n977), .C(n1571), .D(n976), .Q(n989) );
  NAND41 U998 ( .A(n975), .B(n974), .C(n973), .D(n972), .Q(n976) );
  AOI221 U999 ( .A(n1), .B(regs[484]), .C(n1578), .D(regs[420]), .Q(n975) );
  NAND41 U1000 ( .A(n971), .B(n970), .C(n969), .D(n968), .Q(n977) );
  AOI221 U1001 ( .A(n1), .B(regs[996]), .C(n1578), .D(regs[932]), .Q(n971) );
  NAND22 U1002 ( .A(n967), .B(n966), .Q(o_data_Rt[3]) );
  AOI221 U1003 ( .A(n1593), .B(n965), .C(n1591), .D(n964), .Q(n966) );
  NAND41 U1004 ( .A(n963), .B(n962), .C(n961), .D(n960), .Q(n964) );
  AOI221 U1005 ( .A(n1), .B(regs[227]), .C(n81), .D(regs[163]), .Q(n963) );
  NAND41 U1006 ( .A(n959), .B(n958), .C(n957), .D(n956), .Q(n965) );
  AOI221 U1007 ( .A(n7), .B(regs[579]), .C(n47), .D(regs[515]), .Q(n956) );
  AOI221 U1008 ( .A(n1), .B(regs[739]), .C(n81), .D(regs[675]), .Q(n959) );
  AOI221 U1009 ( .A(n1573), .B(n955), .C(n1571), .D(n954), .Q(n967) );
  NAND41 U1010 ( .A(n953), .B(n952), .C(n951), .D(n950), .Q(n954) );
  AOI221 U1011 ( .A(n1), .B(regs[483]), .C(n1578), .D(regs[419]), .Q(n953) );
  NAND41 U1012 ( .A(n949), .B(n948), .C(n947), .D(n946), .Q(n955) );
  AOI221 U1013 ( .A(n1), .B(regs[995]), .C(n1578), .D(regs[931]), .Q(n949) );
  NAND22 U1014 ( .A(n1033), .B(n1032), .Q(o_data_Rt[6]) );
  AOI221 U1015 ( .A(n1593), .B(n1031), .C(n1591), .D(n1030), .Q(n1032) );
  NAND41 U1016 ( .A(n1029), .B(n1028), .C(n1027), .D(n1026), .Q(n1030) );
  AOI221 U1017 ( .A(n55), .B(regs[70]), .C(n47), .D(regs[6]), .Q(n1026) );
  AOI221 U1018 ( .A(n10), .B(regs[102]), .C(n33), .D(regs[38]), .Q(n1027) );
  NAND41 U1019 ( .A(n1025), .B(n1024), .C(n1023), .D(n1022), .Q(n1031) );
  AOI221 U1020 ( .A(n55), .B(regs[582]), .C(n45), .D(regs[518]), .Q(n1022) );
  AOI221 U1021 ( .A(n10), .B(regs[614]), .C(n33), .D(regs[550]), .Q(n1023) );
  AOI221 U1022 ( .A(n7), .B(regs[326]), .C(n47), .D(regs[262]), .Q(n1016) );
  AOI221 U1023 ( .A(n10), .B(regs[358]), .C(n8), .D(regs[294]), .Q(n1017) );
  AOI221 U1024 ( .A(n7), .B(regs[838]), .C(n47), .D(regs[774]), .Q(n1012) );
  AOI221 U1025 ( .A(n10), .B(regs[870]), .C(n8), .D(regs[806]), .Q(n1013) );
  AOI221 U1026 ( .A(n82), .B(regs[966]), .C(n24), .D(regs[902]), .Q(n1014) );
  NAND22 U1027 ( .A(n1165), .B(n1164), .Q(o_data_Rt[12]) );
  AOI221 U1028 ( .A(n7), .B(regs[76]), .C(n45), .D(regs[12]), .Q(n1158) );
  AOI221 U1029 ( .A(n1583), .B(regs[108]), .C(n33), .D(regs[44]), .Q(n1159) );
  AOI221 U1030 ( .A(n83), .B(regs[204]), .C(n2), .D(regs[140]), .Q(n1160) );
  AOI221 U1031 ( .A(n19), .B(regs[236]), .C(n81), .D(regs[172]), .Q(n1161) );
  AOI221 U1032 ( .A(n7), .B(regs[588]), .C(n45), .D(regs[524]), .Q(n1154) );
  AOI221 U1033 ( .A(n10), .B(regs[620]), .C(n33), .D(regs[556]), .Q(n1155) );
  AOI221 U1034 ( .A(n83), .B(regs[716]), .C(n2), .D(regs[652]), .Q(n1156) );
  AOI221 U1035 ( .A(n19), .B(regs[748]), .C(n81), .D(regs[684]), .Q(n1157) );
  NAND41 U1036 ( .A(n1151), .B(n1150), .C(n1149), .D(n1148), .Q(n1152) );
  AOI221 U1037 ( .A(n10), .B(regs[364]), .C(n33), .D(regs[300]), .Q(n1149) );
  NAND41 U1038 ( .A(n1147), .B(n1146), .C(n1145), .D(n1144), .Q(n1153) );
  AOI221 U1039 ( .A(n10), .B(regs[876]), .C(n33), .D(regs[812]), .Q(n1145) );
  NAND22 U1040 ( .A(n901), .B(n900), .Q(o_data_Rt[0]) );
  AOI221 U1041 ( .A(n1593), .B(n899), .C(n1591), .D(n898), .Q(n900) );
  NAND41 U1042 ( .A(n897), .B(n896), .C(n895), .D(n894), .Q(n898) );
  AOI221 U1043 ( .A(n7), .B(regs[64]), .C(n47), .D(regs[0]), .Q(n894) );
  NAND41 U1044 ( .A(n893), .B(n892), .C(n891), .D(n890), .Q(n899) );
  AOI221 U1045 ( .A(regs[608]), .B(n10), .C(regs[544]), .D(n8), .Q(n891) );
  AOI221 U1046 ( .A(regs[704]), .B(n84), .C(regs[640]), .D(n59), .Q(n892) );
  AOI221 U1047 ( .A(n1573), .B(n888), .C(n1571), .D(n887), .Q(n901) );
  NAND41 U1048 ( .A(n886), .B(n885), .C(n884), .D(n883), .Q(n887) );
  NAND41 U1049 ( .A(n881), .B(n880), .C(n879), .D(n878), .Q(n888) );
  AOI221 U1050 ( .A(n10), .B(regs[864]), .C(n8), .D(regs[800]), .Q(n879) );
  AOI221 U1051 ( .A(n84), .B(regs[960]), .C(n59), .D(regs[896]), .Q(n880) );
  NAND22 U1052 ( .A(n1253), .B(n1252), .Q(o_data_Rt[16]) );
  AOI221 U1053 ( .A(n1593), .B(n1251), .C(n1591), .D(n1250), .Q(n1252) );
  AOI221 U1054 ( .A(n7), .B(regs[80]), .C(n45), .D(regs[16]), .Q(n1246) );
  AOI221 U1055 ( .A(n1583), .B(regs[112]), .C(n33), .D(regs[48]), .Q(n1247) );
  AOI221 U1056 ( .A(n53), .B(regs[240]), .C(n81), .D(regs[176]), .Q(n1249) );
  AOI221 U1057 ( .A(n7), .B(regs[592]), .C(n4), .D(regs[528]), .Q(n1242) );
  AOI221 U1058 ( .A(n10), .B(regs[624]), .C(n33), .D(regs[560]), .Q(n1243) );
  AOI221 U1059 ( .A(n53), .B(regs[752]), .C(n81), .D(regs[688]), .Q(n1245) );
  NAND41 U1060 ( .A(n1239), .B(n1238), .C(n1237), .D(n1236), .Q(n1240) );
  AOI221 U1061 ( .A(n7), .B(regs[336]), .C(n47), .D(regs[272]), .Q(n1236) );
  AOI221 U1062 ( .A(n1583), .B(regs[368]), .C(n33), .D(regs[304]), .Q(n1237)
         );
  AOI221 U1063 ( .A(n83), .B(regs[464]), .C(n2), .D(regs[400]), .Q(n1238) );
  AOI221 U1064 ( .A(n53), .B(regs[496]), .C(n81), .D(regs[432]), .Q(n1239) );
  AOI221 U1065 ( .A(n7), .B(regs[848]), .C(n4), .D(regs[784]), .Q(n1232) );
  AOI221 U1066 ( .A(n1583), .B(regs[880]), .C(n33), .D(regs[816]), .Q(n1233)
         );
  AOI221 U1067 ( .A(n83), .B(regs[976]), .C(n2), .D(regs[912]), .Q(n1234) );
  AOI221 U1068 ( .A(n19), .B(regs[1008]), .C(n81), .D(regs[944]), .Q(n1235) );
  NAND22 U1069 ( .A(n1187), .B(n1186), .Q(o_data_Rt[13]) );
  AOI221 U1070 ( .A(n1593), .B(n1185), .C(n1591), .D(n1184), .Q(n1186) );
  AOI221 U1071 ( .A(n7), .B(regs[77]), .C(n45), .D(regs[13]), .Q(n1180) );
  AOI221 U1072 ( .A(n1583), .B(regs[109]), .C(n33), .D(regs[45]), .Q(n1181) );
  AOI221 U1073 ( .A(n83), .B(regs[205]), .C(n2), .D(regs[141]), .Q(n1182) );
  AOI221 U1074 ( .A(n19), .B(regs[237]), .C(n81), .D(regs[173]), .Q(n1183) );
  AOI221 U1075 ( .A(n7), .B(regs[589]), .C(n45), .D(regs[525]), .Q(n1176) );
  AOI221 U1076 ( .A(n10), .B(regs[621]), .C(n33), .D(regs[557]), .Q(n1177) );
  AOI221 U1077 ( .A(n83), .B(regs[717]), .C(n2), .D(regs[653]), .Q(n1178) );
  AOI221 U1078 ( .A(n19), .B(regs[749]), .C(n81), .D(regs[685]), .Q(n1179) );
  AOI221 U1079 ( .A(n1583), .B(regs[365]), .C(n33), .D(regs[301]), .Q(n1171)
         );
  AOI221 U1080 ( .A(n83), .B(regs[461]), .C(n2), .D(regs[397]), .Q(n1172) );
  AOI221 U1081 ( .A(n19), .B(regs[493]), .C(n81), .D(regs[429]), .Q(n1173) );
  AOI221 U1082 ( .A(n7), .B(regs[845]), .C(n45), .D(regs[781]), .Q(n1166) );
  AOI221 U1083 ( .A(n1583), .B(regs[877]), .C(n33), .D(regs[813]), .Q(n1167)
         );
  AOI221 U1084 ( .A(n83), .B(regs[973]), .C(n2), .D(regs[909]), .Q(n1168) );
  AOI221 U1085 ( .A(n19), .B(regs[1005]), .C(n81), .D(regs[941]), .Q(n1169) );
  NAND22 U1086 ( .A(n1231), .B(n1230), .Q(o_data_Rt[15]) );
  AOI221 U1087 ( .A(n1593), .B(n1229), .C(n1591), .D(n1228), .Q(n1230) );
  AOI221 U1088 ( .A(n7), .B(regs[79]), .C(n4), .D(regs[15]), .Q(n1224) );
  AOI221 U1089 ( .A(n1583), .B(regs[111]), .C(n33), .D(regs[47]), .Q(n1225) );
  AOI221 U1090 ( .A(n83), .B(regs[207]), .C(n2), .D(regs[143]), .Q(n1226) );
  AOI221 U1091 ( .A(n19), .B(regs[239]), .C(n81), .D(regs[175]), .Q(n1227) );
  AOI221 U1092 ( .A(n7), .B(regs[591]), .C(n4), .D(regs[527]), .Q(n1220) );
  AOI221 U1093 ( .A(n10), .B(regs[623]), .C(n33), .D(regs[559]), .Q(n1221) );
  AOI221 U1094 ( .A(n83), .B(regs[719]), .C(n2), .D(regs[655]), .Q(n1222) );
  AOI221 U1095 ( .A(n19), .B(regs[751]), .C(n81), .D(regs[687]), .Q(n1223) );
  AOI221 U1096 ( .A(n1583), .B(regs[367]), .C(n33), .D(regs[303]), .Q(n1215)
         );
  AOI221 U1097 ( .A(n83), .B(regs[463]), .C(n59), .D(regs[399]), .Q(n1216) );
  AOI221 U1098 ( .A(n19), .B(regs[495]), .C(n81), .D(regs[431]), .Q(n1217) );
  AOI221 U1099 ( .A(n7), .B(regs[847]), .C(n4), .D(regs[783]), .Q(n1210) );
  AOI221 U1100 ( .A(n1583), .B(regs[879]), .C(n33), .D(regs[815]), .Q(n1211)
         );
  AOI221 U1101 ( .A(n83), .B(regs[975]), .C(n2), .D(regs[911]), .Q(n1212) );
  AOI221 U1102 ( .A(n19), .B(regs[1007]), .C(n81), .D(regs[943]), .Q(n1213) );
  NAND22 U1103 ( .A(n1275), .B(n1274), .Q(o_data_Rt[17]) );
  AOI221 U1104 ( .A(n1593), .B(n1273), .C(n1591), .D(n1272), .Q(n1274) );
  NAND41 U1105 ( .A(n1271), .B(n1270), .C(n1269), .D(n1268), .Q(n1272) );
  AOI221 U1106 ( .A(n7), .B(regs[81]), .C(n47), .D(regs[17]), .Q(n1268) );
  AOI221 U1107 ( .A(n1583), .B(regs[113]), .C(n33), .D(regs[49]), .Q(n1269) );
  AOI221 U1108 ( .A(n53), .B(regs[241]), .C(n81), .D(regs[177]), .Q(n1271) );
  AOI221 U1109 ( .A(n7), .B(regs[593]), .C(n45), .D(regs[529]), .Q(n1264) );
  AOI221 U1110 ( .A(n10), .B(regs[625]), .C(n33), .D(regs[561]), .Q(n1265) );
  AOI221 U1111 ( .A(n53), .B(regs[753]), .C(n81), .D(regs[689]), .Q(n1267) );
  AOI221 U1112 ( .A(n1583), .B(regs[369]), .C(n33), .D(regs[305]), .Q(n1259)
         );
  AOI221 U1113 ( .A(n83), .B(regs[465]), .C(n2), .D(regs[401]), .Q(n1260) );
  AOI221 U1114 ( .A(n53), .B(regs[497]), .C(n81), .D(regs[433]), .Q(n1261) );
  AOI221 U1115 ( .A(n7), .B(regs[849]), .C(n4), .D(regs[785]), .Q(n1254) );
  AOI221 U1116 ( .A(n1583), .B(regs[881]), .C(n33), .D(regs[817]), .Q(n1255)
         );
  AOI221 U1117 ( .A(n83), .B(regs[977]), .C(n2), .D(regs[913]), .Q(n1256) );
  AOI221 U1118 ( .A(n53), .B(regs[1009]), .C(n81), .D(regs[945]), .Q(n1257) );
  NAND22 U1119 ( .A(n1209), .B(n1208), .Q(o_data_Rt[14]) );
  AOI221 U1120 ( .A(n7), .B(regs[78]), .C(n4), .D(regs[14]), .Q(n1202) );
  AOI221 U1121 ( .A(n1583), .B(regs[110]), .C(n33), .D(regs[46]), .Q(n1203) );
  AOI221 U1122 ( .A(n83), .B(regs[206]), .C(n2), .D(regs[142]), .Q(n1204) );
  AOI221 U1123 ( .A(n19), .B(regs[238]), .C(n81), .D(regs[174]), .Q(n1205) );
  AOI221 U1124 ( .A(n7), .B(regs[590]), .C(n4), .D(regs[526]), .Q(n1198) );
  AOI221 U1125 ( .A(n10), .B(regs[622]), .C(n33), .D(regs[558]), .Q(n1199) );
  AOI221 U1126 ( .A(n83), .B(regs[718]), .C(n2), .D(regs[654]), .Q(n1200) );
  AOI221 U1127 ( .A(n19), .B(regs[750]), .C(n81), .D(regs[686]), .Q(n1201) );
  AOI221 U1128 ( .A(n1573), .B(n1197), .C(n1571), .D(n1196), .Q(n1209) );
  AOI221 U1129 ( .A(n1583), .B(regs[366]), .C(n33), .D(regs[302]), .Q(n1193)
         );
  AOI221 U1130 ( .A(n83), .B(regs[462]), .C(n2), .D(regs[398]), .Q(n1194) );
  AOI221 U1131 ( .A(n19), .B(regs[494]), .C(n81), .D(regs[430]), .Q(n1195) );
  AOI221 U1132 ( .A(n7), .B(regs[846]), .C(n45), .D(regs[782]), .Q(n1188) );
  AOI221 U1133 ( .A(n1583), .B(regs[878]), .C(n33), .D(regs[814]), .Q(n1189)
         );
  AOI221 U1134 ( .A(n83), .B(regs[974]), .C(n2), .D(regs[910]), .Q(n1190) );
  AOI221 U1135 ( .A(n19), .B(regs[1006]), .C(n81), .D(regs[942]), .Q(n1191) );
  NAND22 U1136 ( .A(n945), .B(n944), .Q(o_data_Rt[2]) );
  AOI221 U1137 ( .A(n1593), .B(n943), .C(n1591), .D(n942), .Q(n944) );
  NAND41 U1138 ( .A(n941), .B(n940), .C(n939), .D(n938), .Q(n942) );
  AOI221 U1139 ( .A(n1), .B(regs[226]), .C(n1578), .D(regs[162]), .Q(n941) );
  NAND41 U1140 ( .A(n937), .B(n936), .C(n935), .D(n934), .Q(n943) );
  AOI221 U1141 ( .A(n7), .B(regs[578]), .C(n47), .D(regs[514]), .Q(n934) );
  AOI221 U1142 ( .A(n1573), .B(n933), .C(n1571), .D(n932), .Q(n945) );
  NAND41 U1143 ( .A(n931), .B(n930), .C(n929), .D(n928), .Q(n932) );
  NAND41 U1144 ( .A(n927), .B(n926), .C(n925), .D(n924), .Q(n933) );
  AOI221 U1145 ( .A(n7), .B(regs[834]), .C(n45), .D(regs[770]), .Q(n924) );
  AOI221 U1146 ( .A(n82), .B(regs[962]), .C(n1580), .D(regs[898]), .Q(n926) );
  NAND22 U1147 ( .A(n1297), .B(n1296), .Q(o_data_Rt[18]) );
  AOI221 U1148 ( .A(n1593), .B(n1295), .C(n1591), .D(n1294), .Q(n1296) );
  NAND41 U1149 ( .A(n1293), .B(n1292), .C(n1291), .D(n1290), .Q(n1294) );
  NAND41 U1150 ( .A(n1289), .B(n1288), .C(n1287), .D(n1286), .Q(n1295) );
  AOI221 U1151 ( .A(n7), .B(regs[594]), .C(n4), .D(regs[530]), .Q(n1286) );
  NAND41 U1152 ( .A(n1283), .B(n1282), .C(n1281), .D(n1280), .Q(n1284) );
  AOI221 U1153 ( .A(n7), .B(regs[338]), .C(n4), .D(regs[274]), .Q(n1280) );
  AOI221 U1154 ( .A(n84), .B(regs[466]), .C(n24), .D(regs[402]), .Q(n1282) );
  AOI221 U1155 ( .A(n7), .B(regs[850]), .C(n45), .D(regs[786]), .Q(n1276) );
  AOI221 U1156 ( .A(n1583), .B(regs[882]), .C(n33), .D(regs[818]), .Q(n1277)
         );
  AOI221 U1157 ( .A(n83), .B(regs[978]), .C(n2), .D(regs[914]), .Q(n1278) );
  AOI221 U1158 ( .A(n53), .B(regs[1010]), .C(n81), .D(regs[946]), .Q(n1279) );
  NAND22 U1159 ( .A(n1407), .B(n1406), .Q(o_data_Rt[23]) );
  AOI221 U1160 ( .A(n1593), .B(n1405), .C(n1591), .D(n1404), .Q(n1406) );
  NAND41 U1161 ( .A(n1403), .B(n1402), .C(n1401), .D(n1400), .Q(n1404) );
  AOI221 U1162 ( .A(n10), .B(regs[119]), .C(n8), .D(regs[55]), .Q(n1401) );
  NAND41 U1163 ( .A(n1399), .B(n1398), .C(n1397), .D(n1396), .Q(n1405) );
  AOI221 U1164 ( .A(n10), .B(regs[631]), .C(n8), .D(regs[567]), .Q(n1397) );
  AOI221 U1165 ( .A(n1573), .B(n1395), .C(n1571), .D(n1394), .Q(n1407) );
  NAND41 U1166 ( .A(n1393), .B(n1392), .C(n1391), .D(n1390), .Q(n1394) );
  AOI221 U1167 ( .A(n10), .B(regs[375]), .C(n8), .D(regs[311]), .Q(n1391) );
  AOI221 U1168 ( .A(n84), .B(regs[471]), .C(n24), .D(regs[407]), .Q(n1392) );
  NAND41 U1169 ( .A(n1389), .B(n1388), .C(n1387), .D(n1386), .Q(n1395) );
  AOI221 U1170 ( .A(n7), .B(regs[855]), .C(n1584), .D(regs[791]), .Q(n1386) );
  AOI221 U1171 ( .A(n10), .B(regs[887]), .C(n8), .D(regs[823]), .Q(n1387) );
  NAND22 U1172 ( .A(n1319), .B(n1318), .Q(o_data_Rt[19]) );
  AOI221 U1173 ( .A(n1593), .B(n1317), .C(n1591), .D(n1316), .Q(n1318) );
  NAND41 U1174 ( .A(n1315), .B(n1314), .C(n1313), .D(n1312), .Q(n1316) );
  NAND41 U1175 ( .A(n1311), .B(n1310), .C(n1309), .D(n1308), .Q(n1317) );
  AOI221 U1176 ( .A(n7), .B(regs[595]), .C(n4), .D(regs[531]), .Q(n1308) );
  AOI221 U1177 ( .A(n1573), .B(n1307), .C(n1571), .D(n1306), .Q(n1319) );
  NAND41 U1178 ( .A(n1305), .B(n1304), .C(n1303), .D(n1302), .Q(n1306) );
  NAND41 U1179 ( .A(n1301), .B(n1300), .C(n1299), .D(n1298), .Q(n1307) );
  AOI221 U1180 ( .A(n7), .B(regs[851]), .C(n4), .D(regs[787]), .Q(n1298) );
  NAND22 U1181 ( .A(n1385), .B(n1384), .Q(o_data_Rt[22]) );
  AOI221 U1182 ( .A(n1593), .B(n1383), .C(n1591), .D(n1382), .Q(n1384) );
  NAND41 U1183 ( .A(n1381), .B(n1380), .C(n1379), .D(n1378), .Q(n1382) );
  AOI221 U1184 ( .A(n10), .B(regs[118]), .C(n8), .D(regs[54]), .Q(n1379) );
  NAND41 U1185 ( .A(n1377), .B(n1376), .C(n1375), .D(n1374), .Q(n1383) );
  AOI221 U1186 ( .A(n10), .B(regs[630]), .C(n8), .D(regs[566]), .Q(n1375) );
  AOI221 U1187 ( .A(n1573), .B(n1373), .C(n1571), .D(n1372), .Q(n1385) );
  NAND41 U1188 ( .A(n1371), .B(n1370), .C(n1369), .D(n1368), .Q(n1372) );
  AOI221 U1189 ( .A(n10), .B(regs[374]), .C(n8), .D(regs[310]), .Q(n1369) );
  AOI221 U1190 ( .A(n84), .B(regs[470]), .C(n24), .D(regs[406]), .Q(n1370) );
  NAND41 U1191 ( .A(n1367), .B(n1366), .C(n1365), .D(n1364), .Q(n1373) );
  AOI221 U1192 ( .A(n7), .B(regs[854]), .C(n47), .D(regs[790]), .Q(n1364) );
  AOI221 U1193 ( .A(n84), .B(regs[982]), .C(n59), .D(regs[918]), .Q(n1366) );
  NAND22 U1194 ( .A(n1341), .B(n1340), .Q(o_data_Rt[20]) );
  AOI221 U1195 ( .A(n1593), .B(n1339), .C(n1591), .D(n1338), .Q(n1340) );
  NAND41 U1196 ( .A(n1337), .B(n1336), .C(n1335), .D(n1334), .Q(n1338) );
  AOI221 U1197 ( .A(n7), .B(regs[84]), .C(n4), .D(regs[20]), .Q(n1334) );
  NAND41 U1198 ( .A(n1333), .B(n1332), .C(n1331), .D(n1330), .Q(n1339) );
  AOI221 U1199 ( .A(n7), .B(regs[596]), .C(n47), .D(regs[532]), .Q(n1330) );
  AOI221 U1200 ( .A(n1573), .B(n1329), .C(n1571), .D(n1328), .Q(n1341) );
  NAND41 U1201 ( .A(n1327), .B(n1326), .C(n1325), .D(n1324), .Q(n1328) );
  AOI221 U1202 ( .A(n7), .B(regs[340]), .C(n47), .D(regs[276]), .Q(n1324) );
  NAND41 U1203 ( .A(n1323), .B(n1322), .C(n1321), .D(n1320), .Q(n1329) );
  AOI221 U1204 ( .A(n7), .B(regs[852]), .C(n4), .D(regs[788]), .Q(n1320) );
  NAND22 U1205 ( .A(n1363), .B(n1362), .Q(o_data_Rt[21]) );
  AOI221 U1206 ( .A(n1593), .B(n1361), .C(n1591), .D(n1360), .Q(n1362) );
  NAND41 U1207 ( .A(n1359), .B(n1358), .C(n1357), .D(n1356), .Q(n1360) );
  AOI221 U1208 ( .A(n7), .B(regs[85]), .C(n4), .D(regs[21]), .Q(n1356) );
  NAND41 U1209 ( .A(n1355), .B(n1354), .C(n1353), .D(n1352), .Q(n1361) );
  AOI221 U1210 ( .A(n7), .B(regs[597]), .C(n45), .D(regs[533]), .Q(n1352) );
  AOI221 U1211 ( .A(n1573), .B(n1351), .C(n1571), .D(n1350), .Q(n1363) );
  NAND41 U1212 ( .A(n1349), .B(n1348), .C(n1347), .D(n1346), .Q(n1350) );
  AOI221 U1213 ( .A(n7), .B(regs[341]), .C(n4), .D(regs[277]), .Q(n1346) );
  NAND41 U1214 ( .A(n1345), .B(n1344), .C(n1343), .D(n1342), .Q(n1351) );
  AOI221 U1215 ( .A(n7), .B(regs[853]), .C(n4), .D(regs[789]), .Q(n1342) );
  NAND22 U1216 ( .A(n1561), .B(n1560), .Q(o_data_Rt[30]) );
  AOI221 U1217 ( .A(n1593), .B(n1559), .C(n1591), .D(n1558), .Q(n1560) );
  NAND41 U1218 ( .A(n1557), .B(n1556), .C(n1555), .D(n1554), .Q(n1558) );
  AOI221 U1219 ( .A(n10), .B(regs[126]), .C(n8), .D(regs[62]), .Q(n1555) );
  AOI221 U1220 ( .A(n1579), .B(regs[254]), .C(n49), .D(regs[190]), .Q(n1557)
         );
  NAND41 U1221 ( .A(n1553), .B(n1552), .C(n1551), .D(n1550), .Q(n1559) );
  AOI221 U1222 ( .A(n10), .B(regs[638]), .C(n8), .D(regs[574]), .Q(n1551) );
  AOI221 U1223 ( .A(n1), .B(regs[766]), .C(n49), .D(regs[702]), .Q(n1553) );
  NAND41 U1224 ( .A(n1547), .B(n1546), .C(n1545), .D(n1544), .Q(n1548) );
  AOI221 U1225 ( .A(n10), .B(regs[382]), .C(n8), .D(regs[318]), .Q(n1545) );
  AOI221 U1226 ( .A(n1581), .B(regs[478]), .C(n59), .D(regs[414]), .Q(n1546)
         );
  NAND41 U1227 ( .A(n1543), .B(n1542), .C(n1541), .D(n1540), .Q(n1549) );
  AOI221 U1228 ( .A(n1583), .B(regs[894]), .C(n8), .D(regs[830]), .Q(n1541) );
  NAND22 U1229 ( .A(n1595), .B(n1594), .Q(o_data_Rt[31]) );
  AOI221 U1230 ( .A(n1593), .B(n1592), .C(n1591), .D(n1590), .Q(n1594) );
  AOI221 U1231 ( .A(n7), .B(regs[95]), .C(n4), .D(regs[31]), .Q(n1586) );
  AOI221 U1232 ( .A(n1583), .B(regs[127]), .C(n33), .D(regs[63]), .Q(n1587) );
  AOI221 U1233 ( .A(n83), .B(regs[223]), .C(n2), .D(regs[159]), .Q(n1588) );
  AOI221 U1234 ( .A(n19), .B(regs[255]), .C(n81), .D(regs[191]), .Q(n1589) );
  NAND41 U1235 ( .A(n1577), .B(n1576), .C(n1575), .D(n1574), .Q(n1592) );
  AOI221 U1236 ( .A(n10), .B(regs[639]), .C(n8), .D(regs[575]), .Q(n1575) );
  AOI221 U1237 ( .A(n48), .B(regs[735]), .C(n59), .D(regs[671]), .Q(n1576) );
  NAND41 U1238 ( .A(n1569), .B(n1568), .C(n1567), .D(n1566), .Q(n1570) );
  AOI221 U1239 ( .A(n10), .B(regs[383]), .C(n8), .D(regs[319]), .Q(n1567) );
  AOI221 U1240 ( .A(n1581), .B(regs[479]), .C(n59), .D(regs[415]), .Q(n1568)
         );
  NAND41 U1241 ( .A(n1565), .B(n1564), .C(n1563), .D(n1562), .Q(n1572) );
  AOI221 U1242 ( .A(n10), .B(regs[895]), .C(n8), .D(regs[831]), .Q(n1563) );
  AOI221 U1243 ( .A(n82), .B(regs[991]), .C(n59), .D(regs[927]), .Q(n1564) );
  NAND22 U1244 ( .A(n1055), .B(n1054), .Q(o_data_Rt[7]) );
  AOI221 U1245 ( .A(n1593), .B(n1053), .C(n1591), .D(n1052), .Q(n1054) );
  NAND41 U1246 ( .A(n1051), .B(n1050), .C(n1049), .D(n1048), .Q(n1052) );
  AOI221 U1247 ( .A(n55), .B(regs[71]), .C(n47), .D(regs[7]), .Q(n1048) );
  AOI221 U1248 ( .A(n10), .B(regs[103]), .C(n33), .D(regs[39]), .Q(n1049) );
  NAND41 U1249 ( .A(n1047), .B(n1046), .C(n1045), .D(n1044), .Q(n1053) );
  AOI221 U1250 ( .A(n55), .B(regs[583]), .C(n45), .D(regs[519]), .Q(n1044) );
  AOI221 U1251 ( .A(n10), .B(regs[615]), .C(n33), .D(regs[551]), .Q(n1045) );
  NAND41 U1252 ( .A(n1041), .B(n1040), .C(n1039), .D(n1038), .Q(n1042) );
  AOI221 U1253 ( .A(n10), .B(regs[359]), .C(n33), .D(regs[295]), .Q(n1039) );
  NAND41 U1254 ( .A(n1037), .B(n1036), .C(n1035), .D(n1034), .Q(n1043) );
  AOI221 U1255 ( .A(n10), .B(regs[871]), .C(n33), .D(regs[807]), .Q(n1035) );
  AOI221 U1256 ( .A(n48), .B(regs[967]), .C(n2), .D(regs[903]), .Q(n1036) );
  NAND22 U1257 ( .A(n1077), .B(n1076), .Q(o_data_Rt[8]) );
  AOI221 U1258 ( .A(n1593), .B(n1075), .C(n1591), .D(n1074), .Q(n1076) );
  NAND41 U1259 ( .A(n1073), .B(n1072), .C(n1071), .D(n1070), .Q(n1074) );
  AOI221 U1260 ( .A(n55), .B(regs[72]), .C(n1584), .D(regs[8]), .Q(n1070) );
  AOI221 U1261 ( .A(n10), .B(regs[104]), .C(n33), .D(regs[40]), .Q(n1071) );
  NAND41 U1262 ( .A(n1069), .B(n1068), .C(n1067), .D(n1066), .Q(n1075) );
  AOI221 U1263 ( .A(n55), .B(regs[584]), .C(n47), .D(regs[520]), .Q(n1066) );
  AOI221 U1264 ( .A(n10), .B(regs[616]), .C(n33), .D(regs[552]), .Q(n1067) );
  NAND41 U1265 ( .A(n1063), .B(n1062), .C(n1061), .D(n1060), .Q(n1064) );
  AOI221 U1266 ( .A(n10), .B(regs[360]), .C(n33), .D(regs[296]), .Q(n1061) );
  NAND41 U1267 ( .A(n1059), .B(n1058), .C(n1057), .D(n1056), .Q(n1065) );
  AOI221 U1268 ( .A(n55), .B(regs[840]), .C(n1584), .D(regs[776]), .Q(n1056)
         );
  AOI221 U1269 ( .A(n10), .B(regs[872]), .C(n33), .D(regs[808]), .Q(n1057) );
  AOI221 U1270 ( .A(n83), .B(regs[968]), .C(n2), .D(regs[904]), .Q(n1058) );
  NAND22 U1271 ( .A(n1099), .B(n1098), .Q(o_data_Rt[9]) );
  AOI221 U1272 ( .A(n1593), .B(n1097), .C(n1591), .D(n1096), .Q(n1098) );
  NAND41 U1273 ( .A(n1095), .B(n1094), .C(n1093), .D(n1092), .Q(n1096) );
  AOI221 U1274 ( .A(n55), .B(regs[73]), .C(n1584), .D(regs[9]), .Q(n1092) );
  AOI221 U1275 ( .A(n10), .B(regs[105]), .C(n33), .D(regs[41]), .Q(n1093) );
  NAND41 U1276 ( .A(n1091), .B(n1090), .C(n1089), .D(n1088), .Q(n1097) );
  AOI221 U1277 ( .A(n55), .B(regs[585]), .C(n4), .D(regs[521]), .Q(n1088) );
  AOI221 U1278 ( .A(n10), .B(regs[617]), .C(n33), .D(regs[553]), .Q(n1089) );
  NAND41 U1279 ( .A(n1085), .B(n1084), .C(n1083), .D(n1082), .Q(n1086) );
  AOI221 U1280 ( .A(n10), .B(regs[361]), .C(n33), .D(regs[297]), .Q(n1083) );
  NAND41 U1281 ( .A(n1081), .B(n1080), .C(n1079), .D(n1078), .Q(n1087) );
  AOI221 U1282 ( .A(n55), .B(regs[841]), .C(n1584), .D(regs[777]), .Q(n1078)
         );
  AOI221 U1283 ( .A(n10), .B(regs[873]), .C(n33), .D(regs[809]), .Q(n1079) );
  AOI221 U1284 ( .A(n82), .B(regs[969]), .C(n2), .D(regs[905]), .Q(n1080) );
  NAND22 U1285 ( .A(n1121), .B(n1120), .Q(o_data_Rt[10]) );
  NAND41 U1286 ( .A(n1117), .B(n1116), .C(n1115), .D(n1114), .Q(n1118) );
  AOI221 U1287 ( .A(n55), .B(regs[74]), .C(n4), .D(regs[10]), .Q(n1114) );
  AOI221 U1288 ( .A(n10), .B(regs[106]), .C(n33), .D(regs[42]), .Q(n1115) );
  NAND41 U1289 ( .A(n1113), .B(n1112), .C(n1111), .D(n1110), .Q(n1119) );
  AOI221 U1290 ( .A(n55), .B(regs[586]), .C(n4), .D(regs[522]), .Q(n1110) );
  AOI221 U1291 ( .A(n10), .B(regs[618]), .C(n33), .D(regs[554]), .Q(n1111) );
  NAND41 U1292 ( .A(n1107), .B(n1106), .C(n1105), .D(n1104), .Q(n1108) );
  AOI221 U1293 ( .A(n10), .B(regs[362]), .C(n33), .D(regs[298]), .Q(n1105) );
  NAND41 U1294 ( .A(n1103), .B(n1102), .C(n1101), .D(n1100), .Q(n1109) );
  AOI221 U1295 ( .A(n55), .B(regs[842]), .C(n1584), .D(regs[778]), .Q(n1100)
         );
  AOI221 U1296 ( .A(n10), .B(regs[874]), .C(n33), .D(regs[810]), .Q(n1101) );
  AOI221 U1297 ( .A(n48), .B(regs[970]), .C(n2), .D(regs[906]), .Q(n1102) );
  NAND22 U1298 ( .A(n1143), .B(n1142), .Q(o_data_Rt[11]) );
  NAND41 U1299 ( .A(n1139), .B(n1138), .C(n1137), .D(n1136), .Q(n1140) );
  AOI221 U1300 ( .A(n10), .B(regs[107]), .C(n33), .D(regs[43]), .Q(n1137) );
  NAND41 U1301 ( .A(n1135), .B(n1134), .C(n1133), .D(n1132), .Q(n1141) );
  AOI221 U1302 ( .A(n55), .B(regs[587]), .C(n4), .D(regs[523]), .Q(n1132) );
  AOI221 U1303 ( .A(n10), .B(regs[619]), .C(n33), .D(regs[555]), .Q(n1133) );
  NAND41 U1304 ( .A(n1129), .B(n1128), .C(n1127), .D(n1126), .Q(n1130) );
  AOI221 U1305 ( .A(n10), .B(regs[363]), .C(n33), .D(regs[299]), .Q(n1127) );
  NAND41 U1306 ( .A(n1125), .B(n1124), .C(n1123), .D(n1122), .Q(n1131) );
  AOI221 U1307 ( .A(n10), .B(regs[875]), .C(n33), .D(regs[811]), .Q(n1123) );
  NAND22 U1308 ( .A(n1429), .B(n1428), .Q(o_data_Rt[24]) );
  AOI221 U1309 ( .A(n1593), .B(n1427), .C(n1591), .D(n1426), .Q(n1428) );
  NAND41 U1310 ( .A(n1425), .B(n1424), .C(n1423), .D(n1422), .Q(n1426) );
  AOI221 U1311 ( .A(n1583), .B(regs[120]), .C(n8), .D(regs[56]), .Q(n1423) );
  NAND41 U1312 ( .A(n1421), .B(n1420), .C(n1419), .D(n1418), .Q(n1427) );
  AOI221 U1313 ( .A(n1583), .B(regs[632]), .C(n8), .D(regs[568]), .Q(n1419) );
  AOI221 U1314 ( .A(n1573), .B(n1417), .C(n1571), .D(n1416), .Q(n1429) );
  NAND41 U1315 ( .A(n1415), .B(n1414), .C(n1413), .D(n1412), .Q(n1416) );
  AOI221 U1316 ( .A(n10), .B(regs[376]), .C(n8), .D(regs[312]), .Q(n1413) );
  NAND41 U1317 ( .A(n1411), .B(n1410), .C(n1409), .D(n1408), .Q(n1417) );
  AOI221 U1318 ( .A(n7), .B(regs[856]), .C(n1584), .D(regs[792]), .Q(n1408) );
  AOI221 U1319 ( .A(n10), .B(regs[888]), .C(n8), .D(regs[824]), .Q(n1409) );
  NAND22 U1320 ( .A(n1517), .B(n1516), .Q(o_data_Rt[28]) );
  AOI221 U1321 ( .A(n1593), .B(n1515), .C(n1591), .D(n1514), .Q(n1516) );
  NAND41 U1322 ( .A(n1513), .B(n1512), .C(n1511), .D(n1510), .Q(n1514) );
  AOI221 U1323 ( .A(n55), .B(regs[92]), .C(n45), .D(regs[28]), .Q(n1510) );
  AOI221 U1324 ( .A(n1583), .B(regs[124]), .C(n8), .D(regs[60]), .Q(n1511) );
  NAND41 U1325 ( .A(n1509), .B(n1508), .C(n1507), .D(n1506), .Q(n1515) );
  AOI221 U1326 ( .A(n55), .B(regs[604]), .C(n45), .D(regs[540]), .Q(n1506) );
  AOI221 U1327 ( .A(n1583), .B(regs[636]), .C(n8), .D(regs[572]), .Q(n1507) );
  AOI221 U1328 ( .A(n1573), .B(n1505), .C(n1571), .D(n1504), .Q(n1517) );
  NAND41 U1329 ( .A(n1503), .B(n1502), .C(n1501), .D(n1500), .Q(n1504) );
  AOI221 U1330 ( .A(n10), .B(regs[380]), .C(n8), .D(regs[316]), .Q(n1501) );
  NAND41 U1331 ( .A(n1499), .B(n1498), .C(n1497), .D(n1496), .Q(n1505) );
  AOI221 U1332 ( .A(n1583), .B(regs[892]), .C(n8), .D(regs[828]), .Q(n1497) );
  AOI221 U1333 ( .A(n48), .B(regs[988]), .C(n2), .D(regs[924]), .Q(n1498) );
  NAND22 U1334 ( .A(n1539), .B(n1538), .Q(o_data_Rt[29]) );
  AOI221 U1335 ( .A(n1593), .B(n1537), .C(n1591), .D(n1536), .Q(n1538) );
  NAND41 U1336 ( .A(n1535), .B(n1534), .C(n1533), .D(n1532), .Q(n1536) );
  AOI221 U1337 ( .A(n1583), .B(regs[125]), .C(n8), .D(regs[61]), .Q(n1533) );
  NAND41 U1338 ( .A(n1531), .B(n1530), .C(n1529), .D(n1528), .Q(n1537) );
  AOI221 U1339 ( .A(n55), .B(regs[605]), .C(n45), .D(regs[541]), .Q(n1528) );
  AOI221 U1340 ( .A(n1583), .B(regs[637]), .C(n8), .D(regs[573]), .Q(n1529) );
  AOI221 U1341 ( .A(n1573), .B(n1527), .C(n1571), .D(n1526), .Q(n1539) );
  NAND41 U1342 ( .A(n1525), .B(n1524), .C(n1523), .D(n1522), .Q(n1526) );
  AOI221 U1343 ( .A(n10), .B(regs[381]), .C(n8), .D(regs[317]), .Q(n1523) );
  NAND41 U1344 ( .A(n1521), .B(n1520), .C(n1519), .D(n1518), .Q(n1527) );
  AOI221 U1345 ( .A(n1583), .B(regs[893]), .C(n8), .D(regs[829]), .Q(n1519) );
  NAND22 U1346 ( .A(n1451), .B(n1450), .Q(o_data_Rt[25]) );
  AOI221 U1347 ( .A(n1593), .B(n1449), .C(n1591), .D(n1448), .Q(n1450) );
  NAND41 U1348 ( .A(n1447), .B(n1446), .C(n1445), .D(n1444), .Q(n1448) );
  AOI221 U1349 ( .A(n1583), .B(regs[121]), .C(n8), .D(regs[57]), .Q(n1445) );
  NAND41 U1350 ( .A(n1443), .B(n1442), .C(n1441), .D(n1440), .Q(n1449) );
  AOI221 U1351 ( .A(n1583), .B(regs[633]), .C(n8), .D(regs[569]), .Q(n1441) );
  AOI221 U1352 ( .A(n1573), .B(n1439), .C(n1571), .D(n1438), .Q(n1451) );
  NAND41 U1353 ( .A(n1437), .B(n1436), .C(n1435), .D(n1434), .Q(n1438) );
  AOI221 U1354 ( .A(n10), .B(regs[377]), .C(n8), .D(regs[313]), .Q(n1435) );
  AOI221 U1355 ( .A(n55), .B(regs[857]), .C(n45), .D(regs[793]), .Q(n1430) );
  AOI221 U1356 ( .A(n1583), .B(regs[889]), .C(n8), .D(regs[825]), .Q(n1431) );
  NAND22 U1357 ( .A(n1495), .B(n1494), .Q(o_data_Rt[27]) );
  AOI221 U1358 ( .A(n1593), .B(n1493), .C(n1591), .D(n1492), .Q(n1494) );
  AOI221 U1359 ( .A(n1583), .B(regs[123]), .C(n8), .D(regs[59]), .Q(n1489) );
  AOI221 U1360 ( .A(n48), .B(regs[219]), .C(n2), .D(regs[155]), .Q(n1490) );
  NAND41 U1361 ( .A(n1487), .B(n1486), .C(n1485), .D(n1484), .Q(n1493) );
  AOI221 U1362 ( .A(n1583), .B(regs[635]), .C(n8), .D(regs[571]), .Q(n1485) );
  AOI221 U1363 ( .A(n1573), .B(n1483), .C(n1571), .D(n1482), .Q(n1495) );
  NAND41 U1364 ( .A(n1481), .B(n1480), .C(n1479), .D(n1478), .Q(n1482) );
  AOI221 U1365 ( .A(n10), .B(regs[379]), .C(n8), .D(regs[315]), .Q(n1479) );
  AOI221 U1366 ( .A(n48), .B(regs[475]), .C(n2), .D(regs[411]), .Q(n1480) );
  NAND41 U1367 ( .A(n1477), .B(n1476), .C(n1475), .D(n1474), .Q(n1483) );
  AOI221 U1368 ( .A(n1583), .B(regs[891]), .C(n8), .D(regs[827]), .Q(n1475) );
  AOI221 U1369 ( .A(n48), .B(regs[987]), .C(n2), .D(regs[923]), .Q(n1476) );
  NAND22 U1370 ( .A(n1473), .B(n1472), .Q(o_data_Rt[26]) );
  AOI221 U1371 ( .A(n1593), .B(n1471), .C(n1591), .D(n1470), .Q(n1472) );
  AOI221 U1372 ( .A(n1583), .B(regs[122]), .C(n8), .D(regs[58]), .Q(n1467) );
  AOI221 U1373 ( .A(n48), .B(regs[218]), .C(n2), .D(regs[154]), .Q(n1468) );
  NAND41 U1374 ( .A(n1465), .B(n1464), .C(n1463), .D(n1462), .Q(n1471) );
  AOI221 U1375 ( .A(n1583), .B(regs[634]), .C(n8), .D(regs[570]), .Q(n1463) );
  AOI221 U1376 ( .A(n1573), .B(n1461), .C(n1571), .D(n1460), .Q(n1473) );
  NAND41 U1377 ( .A(n1459), .B(n1458), .C(n1457), .D(n1456), .Q(n1460) );
  AOI221 U1378 ( .A(n10), .B(regs[378]), .C(n8), .D(regs[314]), .Q(n1457) );
  AOI221 U1379 ( .A(n48), .B(regs[474]), .C(n2), .D(regs[410]), .Q(n1458) );
  AOI221 U1380 ( .A(n1583), .B(regs[890]), .C(n8), .D(regs[826]), .Q(n1453) );
  NAND22 U1381 ( .A(n179), .B(n178), .Q(o_data_Rs[0]) );
  NAND41 U1382 ( .A(n175), .B(n174), .C(n173), .D(n172), .Q(n176) );
  AOI221 U1383 ( .A(n71), .B(regs[672]), .C(n65), .D(regs[640]), .Q(n172) );
  NAND41 U1384 ( .A(n170), .B(n169), .C(n168), .D(n167), .Q(n177) );
  NAND41 U1385 ( .A(n164), .B(n163), .C(n162), .D(n161), .Q(n165) );
  AOI221 U1386 ( .A(n71), .B(regs[416]), .C(n80), .D(regs[384]), .Q(n155) );
  NAND22 U1387 ( .A(n663), .B(n662), .Q(o_data_Rs[22]) );
  NAND41 U1388 ( .A(n659), .B(n658), .C(n657), .D(n656), .Q(n660) );
  AOI221 U1389 ( .A(n71), .B(regs[694]), .C(n65), .D(regs[662]), .Q(n656) );
  AOI221 U1390 ( .A(n46), .B(regs[598]), .C(n63), .D(regs[534]), .Q(n657) );
  AOI221 U1391 ( .A(n61), .B(regs[630]), .C(n12), .D(regs[566]), .Q(n658) );
  NAND41 U1392 ( .A(n655), .B(n654), .C(n653), .D(n652), .Q(n661) );
  AOI221 U1393 ( .A(n71), .B(regs[182]), .C(n65), .D(regs[150]), .Q(n652) );
  AOI221 U1394 ( .A(n46), .B(regs[86]), .C(n51), .D(regs[22]), .Q(n653) );
  NAND41 U1395 ( .A(n649), .B(n648), .C(n647), .D(n646), .Q(n650) );
  AOI221 U1396 ( .A(n861), .B(regs[854]), .C(n51), .D(regs[790]), .Q(n647) );
  NAND41 U1397 ( .A(n645), .B(n644), .C(n643), .D(n642), .Q(n651) );
  AOI221 U1398 ( .A(n861), .B(regs[342]), .C(n51), .D(regs[278]), .Q(n643) );
  AOI221 U1399 ( .A(n221), .B(n870), .C(n869), .D(n220), .Q(n222) );
  NAND41 U1400 ( .A(n219), .B(n218), .C(n217), .D(n216), .Q(n220) );
  NAND41 U1401 ( .A(n215), .B(n214), .C(n213), .D(n212), .Q(n221) );
  AOI221 U1402 ( .A(n72), .B(regs[162]), .C(n80), .D(regs[130]), .Q(n212) );
  AOI221 U1403 ( .A(n211), .B(n850), .C(n849), .D(n210), .Q(n223) );
  NAND41 U1404 ( .A(n209), .B(n208), .C(n207), .D(n206), .Q(n210) );
  NAND41 U1405 ( .A(n205), .B(n204), .C(n203), .D(n202), .Q(n211) );
  NAND22 U1406 ( .A(n201), .B(n200), .Q(o_data_Rs[1]) );
  AOI221 U1407 ( .A(n71), .B(regs[673]), .C(n80), .D(regs[641]), .Q(n194) );
  NAND41 U1408 ( .A(n193), .B(n192), .C(n191), .D(n190), .Q(n199) );
  NAND41 U1409 ( .A(n187), .B(n186), .C(n185), .D(n184), .Q(n188) );
  NAND41 U1410 ( .A(n183), .B(n182), .C(n181), .D(n180), .Q(n189) );
  AOI221 U1411 ( .A(n71), .B(regs[417]), .C(n65), .D(regs[385]), .Q(n180) );
  NAND22 U1412 ( .A(n641), .B(n640), .Q(o_data_Rs[21]) );
  NAND41 U1413 ( .A(n637), .B(n636), .C(n635), .D(n634), .Q(n638) );
  AOI221 U1414 ( .A(n46), .B(regs[597]), .C(n51), .D(regs[533]), .Q(n635) );
  AOI221 U1415 ( .A(n78), .B(regs[629]), .C(n12), .D(regs[565]), .Q(n636) );
  NAND41 U1416 ( .A(n633), .B(n632), .C(n631), .D(n630), .Q(n639) );
  AOI221 U1417 ( .A(n46), .B(regs[85]), .C(n51), .D(regs[21]), .Q(n631) );
  AOI221 U1418 ( .A(n78), .B(regs[117]), .C(n12), .D(regs[53]), .Q(n632) );
  NAND41 U1419 ( .A(n627), .B(n626), .C(n625), .D(n624), .Q(n628) );
  AOI221 U1420 ( .A(n861), .B(regs[853]), .C(n51), .D(regs[789]), .Q(n625) );
  AOI221 U1421 ( .A(n78), .B(regs[885]), .C(n12), .D(regs[821]), .Q(n626) );
  NAND41 U1422 ( .A(n623), .B(n622), .C(n621), .D(n620), .Q(n629) );
  AOI221 U1423 ( .A(n3), .B(regs[341]), .C(n51), .D(regs[277]), .Q(n621) );
  AOI221 U1424 ( .A(n78), .B(regs[373]), .C(n12), .D(regs[309]), .Q(n622) );
  NAND22 U1425 ( .A(n839), .B(n838), .Q(o_data_Rs[30]) );
  AOI221 U1426 ( .A(n72), .B(regs[702]), .C(n65), .D(regs[670]), .Q(n832) );
  NAND41 U1427 ( .A(n831), .B(n830), .C(n829), .D(n828), .Q(n837) );
  AOI221 U1428 ( .A(n72), .B(regs[958]), .C(n65), .D(regs[926]), .Q(n822) );
  AOI221 U1429 ( .A(n72), .B(regs[446]), .C(n65), .D(regs[414]), .Q(n818) );
  NAND41 U1430 ( .A(n791), .B(n790), .C(n789), .D(n788), .Q(n792) );
  AOI221 U1431 ( .A(n71), .B(regs[700]), .C(n65), .D(regs[668]), .Q(n788) );
  AOI221 U1432 ( .A(n56), .B(regs[604]), .C(n51), .D(regs[540]), .Q(n789) );
  AOI221 U1433 ( .A(n54), .B(regs[636]), .C(n12), .D(regs[572]), .Q(n790) );
  NAND41 U1434 ( .A(n787), .B(n786), .C(n785), .D(n784), .Q(n793) );
  AOI221 U1435 ( .A(n71), .B(regs[188]), .C(n65), .D(regs[156]), .Q(n784) );
  AOI221 U1436 ( .A(n56), .B(regs[92]), .C(n63), .D(regs[28]), .Q(n785) );
  AOI221 U1437 ( .A(n54), .B(regs[124]), .C(n12), .D(regs[60]), .Q(n786) );
  NAND41 U1438 ( .A(n781), .B(n780), .C(n779), .D(n778), .Q(n782) );
  AOI221 U1439 ( .A(n56), .B(regs[860]), .C(n79), .D(regs[796]), .Q(n779) );
  AOI221 U1440 ( .A(n54), .B(regs[892]), .C(n12), .D(regs[828]), .Q(n780) );
  NAND41 U1441 ( .A(n777), .B(n776), .C(n775), .D(n774), .Q(n783) );
  AOI221 U1442 ( .A(n71), .B(regs[444]), .C(n80), .D(regs[412]), .Q(n774) );
  AOI221 U1443 ( .A(n56), .B(regs[348]), .C(n51), .D(regs[284]), .Q(n775) );
  AOI221 U1444 ( .A(n54), .B(regs[380]), .C(n12), .D(regs[316]), .Q(n776) );
  NAND22 U1445 ( .A(n751), .B(n750), .Q(o_data_Rs[26]) );
  NAND41 U1446 ( .A(n747), .B(n746), .C(n745), .D(n744), .Q(n748) );
  AOI221 U1447 ( .A(n72), .B(regs[698]), .C(n80), .D(regs[666]), .Q(n744) );
  AOI221 U1448 ( .A(n3), .B(regs[602]), .C(n14), .D(regs[538]), .Q(n745) );
  AOI221 U1449 ( .A(n61), .B(regs[634]), .C(n12), .D(regs[570]), .Q(n746) );
  NAND41 U1450 ( .A(n743), .B(n742), .C(n741), .D(n740), .Q(n749) );
  AOI221 U1451 ( .A(n72), .B(regs[186]), .C(n80), .D(regs[154]), .Q(n740) );
  AOI221 U1452 ( .A(n3), .B(regs[90]), .C(n14), .D(regs[26]), .Q(n741) );
  AOI221 U1453 ( .A(n61), .B(regs[122]), .C(n12), .D(regs[58]), .Q(n742) );
  NAND41 U1454 ( .A(n737), .B(n736), .C(n735), .D(n734), .Q(n738) );
  AOI221 U1455 ( .A(n72), .B(regs[954]), .C(n65), .D(regs[922]), .Q(n734) );
  AOI221 U1456 ( .A(n3), .B(regs[858]), .C(n14), .D(regs[794]), .Q(n735) );
  AOI221 U1457 ( .A(n61), .B(regs[890]), .C(n12), .D(regs[826]), .Q(n736) );
  NAND41 U1458 ( .A(n733), .B(n732), .C(n731), .D(n730), .Q(n739) );
  AOI221 U1459 ( .A(n72), .B(regs[442]), .C(n80), .D(regs[410]), .Q(n730) );
  AOI221 U1460 ( .A(n3), .B(regs[346]), .C(n14), .D(regs[282]), .Q(n731) );
  AOI221 U1461 ( .A(n61), .B(regs[378]), .C(n12), .D(regs[314]), .Q(n732) );
  AOI221 U1462 ( .A(n71), .B(regs[703]), .C(n80), .D(regs[671]), .Q(n864) );
  AOI221 U1463 ( .A(n50), .B(regs[767]), .C(n76), .D(regs[735]), .Q(n867) );
  NAND41 U1464 ( .A(n855), .B(n854), .C(n853), .D(n852), .Q(n871) );
  NAND41 U1465 ( .A(n847), .B(n846), .C(n845), .D(n844), .Q(n848) );
  AOI221 U1466 ( .A(n72), .B(regs[447]), .C(n65), .D(regs[415]), .Q(n840) );
  NAND22 U1467 ( .A(n773), .B(n772), .Q(o_data_Rs[27]) );
  NAND41 U1468 ( .A(n769), .B(n768), .C(n767), .D(n766), .Q(n770) );
  AOI221 U1469 ( .A(n56), .B(regs[603]), .C(n14), .D(regs[539]), .Q(n767) );
  AOI221 U1470 ( .A(n54), .B(regs[635]), .C(n12), .D(regs[571]), .Q(n768) );
  NAND41 U1471 ( .A(n765), .B(n764), .C(n763), .D(n762), .Q(n771) );
  AOI221 U1472 ( .A(n71), .B(regs[187]), .C(n80), .D(regs[155]), .Q(n762) );
  AOI221 U1473 ( .A(n56), .B(regs[91]), .C(n63), .D(regs[27]), .Q(n763) );
  AOI221 U1474 ( .A(n54), .B(regs[123]), .C(n12), .D(regs[59]), .Q(n764) );
  NAND41 U1475 ( .A(n759), .B(n758), .C(n757), .D(n756), .Q(n760) );
  AOI221 U1476 ( .A(n71), .B(regs[955]), .C(n65), .D(regs[923]), .Q(n756) );
  AOI221 U1477 ( .A(n56), .B(regs[859]), .C(n79), .D(regs[795]), .Q(n757) );
  AOI221 U1478 ( .A(n54), .B(regs[891]), .C(n12), .D(regs[827]), .Q(n758) );
  NAND41 U1479 ( .A(n755), .B(n754), .C(n753), .D(n752), .Q(n761) );
  AOI221 U1480 ( .A(n71), .B(regs[443]), .C(n80), .D(regs[411]), .Q(n752) );
  AOI221 U1481 ( .A(n56), .B(regs[347]), .C(n63), .D(regs[283]), .Q(n753) );
  AOI221 U1482 ( .A(n54), .B(regs[379]), .C(n12), .D(regs[315]), .Q(n754) );
  NAND22 U1483 ( .A(n729), .B(n728), .Q(o_data_Rs[25]) );
  NAND41 U1484 ( .A(n725), .B(n724), .C(n723), .D(n722), .Q(n726) );
  AOI221 U1485 ( .A(n3), .B(regs[601]), .C(n14), .D(regs[537]), .Q(n723) );
  AOI221 U1486 ( .A(n61), .B(regs[633]), .C(n12), .D(regs[569]), .Q(n724) );
  NAND41 U1487 ( .A(n721), .B(n720), .C(n719), .D(n718), .Q(n727) );
  AOI221 U1488 ( .A(n72), .B(regs[185]), .C(n65), .D(regs[153]), .Q(n718) );
  AOI221 U1489 ( .A(n3), .B(regs[89]), .C(n14), .D(regs[25]), .Q(n719) );
  AOI221 U1490 ( .A(n61), .B(regs[121]), .C(n12), .D(regs[57]), .Q(n720) );
  NAND41 U1491 ( .A(n715), .B(n714), .C(n713), .D(n712), .Q(n716) );
  AOI221 U1492 ( .A(n3), .B(regs[857]), .C(n14), .D(regs[793]), .Q(n713) );
  AOI221 U1493 ( .A(n61), .B(regs[889]), .C(n12), .D(regs[825]), .Q(n714) );
  NAND41 U1494 ( .A(n711), .B(n710), .C(n709), .D(n708), .Q(n717) );
  AOI221 U1495 ( .A(n3), .B(regs[345]), .C(n14), .D(regs[281]), .Q(n709) );
  AOI221 U1496 ( .A(n61), .B(regs[377]), .C(n12), .D(regs[313]), .Q(n710) );
  NAND22 U1497 ( .A(n707), .B(n706), .Q(o_data_Rs[24]) );
  NAND41 U1498 ( .A(n703), .B(n702), .C(n701), .D(n700), .Q(n704) );
  AOI221 U1499 ( .A(n72), .B(regs[696]), .C(n65), .D(regs[664]), .Q(n700) );
  AOI221 U1500 ( .A(n3), .B(regs[600]), .C(n14), .D(regs[536]), .Q(n701) );
  AOI221 U1501 ( .A(n61), .B(regs[632]), .C(n12), .D(regs[568]), .Q(n702) );
  NAND41 U1502 ( .A(n699), .B(n698), .C(n697), .D(n696), .Q(n705) );
  AOI221 U1503 ( .A(n71), .B(regs[184]), .C(n80), .D(regs[152]), .Q(n696) );
  AOI221 U1504 ( .A(n46), .B(regs[88]), .C(n14), .D(regs[24]), .Q(n697) );
  AOI221 U1505 ( .A(n54), .B(regs[120]), .C(n12), .D(regs[56]), .Q(n698) );
  NAND41 U1506 ( .A(n693), .B(n692), .C(n691), .D(n690), .Q(n694) );
  AOI221 U1507 ( .A(n46), .B(regs[856]), .C(n14), .D(regs[792]), .Q(n691) );
  AOI221 U1508 ( .A(n61), .B(regs[888]), .C(n12), .D(regs[824]), .Q(n692) );
  NAND41 U1509 ( .A(n689), .B(n688), .C(n687), .D(n686), .Q(n695) );
  AOI221 U1510 ( .A(n71), .B(regs[440]), .C(n80), .D(regs[408]), .Q(n686) );
  AOI221 U1511 ( .A(n46), .B(regs[344]), .C(n14), .D(regs[280]), .Q(n687) );
  AOI221 U1512 ( .A(n54), .B(regs[376]), .C(n12), .D(regs[312]), .Q(n688) );
  NAND41 U1513 ( .A(n681), .B(n680), .C(n679), .D(n678), .Q(n682) );
  AOI221 U1514 ( .A(n46), .B(regs[599]), .C(n63), .D(regs[535]), .Q(n679) );
  AOI221 U1515 ( .A(n61), .B(regs[631]), .C(n12), .D(regs[567]), .Q(n680) );
  NAND41 U1516 ( .A(n677), .B(n676), .C(n675), .D(n674), .Q(n683) );
  AOI221 U1517 ( .A(n71), .B(regs[183]), .C(n80), .D(regs[151]), .Q(n674) );
  AOI221 U1518 ( .A(n46), .B(regs[87]), .C(n51), .D(regs[23]), .Q(n675) );
  AOI221 U1519 ( .A(n54), .B(regs[119]), .C(n12), .D(regs[55]), .Q(n676) );
  NAND41 U1520 ( .A(n671), .B(n670), .C(n669), .D(n668), .Q(n672) );
  AOI221 U1521 ( .A(n46), .B(regs[855]), .C(n79), .D(regs[791]), .Q(n669) );
  AOI221 U1522 ( .A(n61), .B(regs[887]), .C(n12), .D(regs[823]), .Q(n670) );
  NAND41 U1523 ( .A(n667), .B(n666), .C(n665), .D(n664), .Q(n673) );
  AOI221 U1524 ( .A(n71), .B(regs[439]), .C(n80), .D(regs[407]), .Q(n664) );
  AOI221 U1525 ( .A(n46), .B(regs[343]), .C(n63), .D(regs[279]), .Q(n665) );
  NAND41 U1526 ( .A(n813), .B(n812), .C(n811), .D(n810), .Q(n814) );
  AOI221 U1527 ( .A(n56), .B(regs[605]), .C(n63), .D(regs[541]), .Q(n811) );
  AOI221 U1528 ( .A(n66), .B(regs[637]), .C(n12), .D(regs[573]), .Q(n812) );
  NAND41 U1529 ( .A(n809), .B(n808), .C(n807), .D(n806), .Q(n815) );
  AOI221 U1530 ( .A(n72), .B(regs[189]), .C(n80), .D(regs[157]), .Q(n806) );
  AOI221 U1531 ( .A(n56), .B(regs[93]), .C(n51), .D(regs[29]), .Q(n807) );
  AOI221 U1532 ( .A(n66), .B(regs[125]), .C(n12), .D(regs[61]), .Q(n808) );
  NAND41 U1533 ( .A(n803), .B(n802), .C(n801), .D(n800), .Q(n804) );
  AOI221 U1534 ( .A(n72), .B(regs[957]), .C(n80), .D(regs[925]), .Q(n800) );
  AOI221 U1535 ( .A(n56), .B(regs[861]), .C(n79), .D(regs[797]), .Q(n801) );
  NAND41 U1536 ( .A(n799), .B(n798), .C(n797), .D(n796), .Q(n805) );
  AOI221 U1537 ( .A(n71), .B(regs[445]), .C(n65), .D(regs[413]), .Q(n796) );
  AOI221 U1538 ( .A(n56), .B(regs[349]), .C(n51), .D(regs[285]), .Q(n797) );
  AOI221 U1539 ( .A(n54), .B(regs[381]), .C(n12), .D(regs[317]), .Q(n798) );
  NAND22 U1540 ( .A(n245), .B(n244), .Q(o_data_Rs[3]) );
  NAND41 U1541 ( .A(n241), .B(n240), .C(n239), .D(n238), .Q(n242) );
  NAND41 U1542 ( .A(n237), .B(n236), .C(n235), .D(n234), .Q(n243) );
  NAND41 U1543 ( .A(n231), .B(n230), .C(n229), .D(n228), .Q(n232) );
  NAND41 U1544 ( .A(n227), .B(n226), .C(n225), .D(n224), .Q(n233) );
  NAND22 U1545 ( .A(n619), .B(n618), .Q(o_data_Rs[20]) );
  NAND41 U1546 ( .A(n615), .B(n614), .C(n613), .D(n612), .Q(n616) );
  NAND41 U1547 ( .A(n611), .B(n610), .C(n609), .D(n608), .Q(n617) );
  NAND41 U1548 ( .A(n605), .B(n604), .C(n603), .D(n602), .Q(n606) );
  NAND41 U1549 ( .A(n601), .B(n600), .C(n599), .D(n598), .Q(n607) );
  NAND22 U1550 ( .A(n465), .B(n464), .Q(o_data_Rs[13]) );
  NAND41 U1551 ( .A(n461), .B(n460), .C(n459), .D(n458), .Q(n462) );
  AOI221 U1552 ( .A(n71), .B(regs[685]), .C(n80), .D(regs[653]), .Q(n458) );
  NAND41 U1553 ( .A(n457), .B(n456), .C(n455), .D(n454), .Q(n463) );
  AOI221 U1554 ( .A(n71), .B(regs[173]), .C(n80), .D(regs[141]), .Q(n454) );
  NAND41 U1555 ( .A(n451), .B(n450), .C(n449), .D(n448), .Q(n452) );
  NAND41 U1556 ( .A(n447), .B(n446), .C(n445), .D(n444), .Q(n453) );
  NAND22 U1557 ( .A(n509), .B(n508), .Q(o_data_Rs[15]) );
  NAND41 U1558 ( .A(n505), .B(n504), .C(n503), .D(n502), .Q(n506) );
  AOI221 U1559 ( .A(n72), .B(regs[687]), .C(n65), .D(regs[655]), .Q(n502) );
  NAND41 U1560 ( .A(n501), .B(n500), .C(n499), .D(n498), .Q(n507) );
  AOI221 U1561 ( .A(n71), .B(regs[175]), .C(n65), .D(regs[143]), .Q(n498) );
  NAND41 U1562 ( .A(n495), .B(n494), .C(n493), .D(n492), .Q(n496) );
  NAND41 U1563 ( .A(n491), .B(n490), .C(n489), .D(n488), .Q(n497) );
  AOI221 U1564 ( .A(n71), .B(regs[431]), .C(n65), .D(regs[399]), .Q(n488) );
  NAND22 U1565 ( .A(n377), .B(n376), .Q(o_data_Rs[9]) );
  NAND41 U1566 ( .A(n373), .B(n372), .C(n371), .D(n370), .Q(n374) );
  AOI221 U1567 ( .A(n71), .B(regs[681]), .C(n65), .D(regs[649]), .Q(n370) );
  NAND41 U1568 ( .A(n369), .B(n368), .C(n367), .D(n366), .Q(n375) );
  AOI221 U1569 ( .A(n71), .B(regs[169]), .C(n65), .D(regs[137]), .Q(n366) );
  NAND41 U1570 ( .A(n363), .B(n362), .C(n361), .D(n360), .Q(n364) );
  NAND41 U1571 ( .A(n359), .B(n358), .C(n357), .D(n356), .Q(n365) );
  NAND22 U1572 ( .A(n289), .B(n288), .Q(o_data_Rs[5]) );
  NAND41 U1573 ( .A(n285), .B(n284), .C(n283), .D(n282), .Q(n286) );
  NAND41 U1574 ( .A(n281), .B(n280), .C(n279), .D(n278), .Q(n287) );
  NAND41 U1575 ( .A(n275), .B(n274), .C(n273), .D(n272), .Q(n276) );
  NAND41 U1576 ( .A(n271), .B(n270), .C(n269), .D(n268), .Q(n277) );
  NAND22 U1577 ( .A(n311), .B(n310), .Q(o_data_Rs[6]) );
  NAND41 U1578 ( .A(n307), .B(n306), .C(n305), .D(n304), .Q(n308) );
  AOI221 U1579 ( .A(n72), .B(regs[678]), .C(n80), .D(regs[646]), .Q(n304) );
  NAND41 U1580 ( .A(n303), .B(n302), .C(n301), .D(n300), .Q(n309) );
  AOI221 U1581 ( .A(n71), .B(regs[166]), .C(n80), .D(regs[134]), .Q(n300) );
  NAND41 U1582 ( .A(n297), .B(n296), .C(n295), .D(n294), .Q(n298) );
  NAND41 U1583 ( .A(n293), .B(n292), .C(n291), .D(n290), .Q(n299) );
  NAND22 U1584 ( .A(n399), .B(n398), .Q(o_data_Rs[10]) );
  NAND41 U1585 ( .A(n395), .B(n394), .C(n393), .D(n392), .Q(n396) );
  AOI221 U1586 ( .A(n71), .B(regs[682]), .C(n65), .D(regs[650]), .Q(n392) );
  NAND41 U1587 ( .A(n391), .B(n390), .C(n389), .D(n388), .Q(n397) );
  AOI221 U1588 ( .A(n71), .B(regs[170]), .C(n65), .D(regs[138]), .Q(n388) );
  NAND41 U1589 ( .A(n385), .B(n384), .C(n383), .D(n382), .Q(n386) );
  NAND41 U1590 ( .A(n381), .B(n380), .C(n379), .D(n378), .Q(n387) );
  NAND22 U1591 ( .A(n267), .B(n266), .Q(o_data_Rs[4]) );
  NAND41 U1592 ( .A(n263), .B(n262), .C(n261), .D(n260), .Q(n264) );
  NAND41 U1593 ( .A(n259), .B(n258), .C(n257), .D(n256), .Q(n265) );
  NAND41 U1594 ( .A(n253), .B(n252), .C(n251), .D(n250), .Q(n254) );
  NAND41 U1595 ( .A(n249), .B(n248), .C(n247), .D(n246), .Q(n255) );
  NAND22 U1596 ( .A(n597), .B(n596), .Q(o_data_Rs[19]) );
  NAND41 U1597 ( .A(n593), .B(n592), .C(n591), .D(n590), .Q(n594) );
  NAND41 U1598 ( .A(n589), .B(n588), .C(n587), .D(n586), .Q(n595) );
  NAND41 U1599 ( .A(n583), .B(n582), .C(n581), .D(n580), .Q(n584) );
  NAND41 U1600 ( .A(n579), .B(n578), .C(n577), .D(n576), .Q(n585) );
  NAND22 U1601 ( .A(n487), .B(n486), .Q(o_data_Rs[14]) );
  NAND41 U1602 ( .A(n483), .B(n482), .C(n481), .D(n480), .Q(n484) );
  AOI221 U1603 ( .A(n71), .B(regs[686]), .C(n80), .D(regs[654]), .Q(n480) );
  NAND41 U1604 ( .A(n479), .B(n478), .C(n477), .D(n476), .Q(n485) );
  AOI221 U1605 ( .A(n71), .B(regs[174]), .C(n80), .D(regs[142]), .Q(n476) );
  NAND41 U1606 ( .A(n473), .B(n472), .C(n471), .D(n470), .Q(n474) );
  NAND41 U1607 ( .A(n469), .B(n468), .C(n467), .D(n466), .Q(n475) );
  NAND22 U1608 ( .A(n575), .B(n574), .Q(o_data_Rs[18]) );
  NAND41 U1609 ( .A(n571), .B(n570), .C(n569), .D(n568), .Q(n572) );
  NAND41 U1610 ( .A(n567), .B(n566), .C(n565), .D(n564), .Q(n573) );
  NAND41 U1611 ( .A(n561), .B(n560), .C(n559), .D(n558), .Q(n562) );
  NAND41 U1612 ( .A(n557), .B(n556), .C(n555), .D(n554), .Q(n563) );
  NAND22 U1613 ( .A(n553), .B(n552), .Q(o_data_Rs[17]) );
  NAND41 U1614 ( .A(n549), .B(n548), .C(n547), .D(n546), .Q(n550) );
  AOI221 U1615 ( .A(n72), .B(regs[689]), .C(n80), .D(regs[657]), .Q(n546) );
  NAND41 U1616 ( .A(n545), .B(n544), .C(n543), .D(n542), .Q(n551) );
  AOI221 U1617 ( .A(n72), .B(regs[177]), .C(n80), .D(regs[145]), .Q(n542) );
  NAND41 U1618 ( .A(n539), .B(n538), .C(n537), .D(n536), .Q(n540) );
  NAND41 U1619 ( .A(n535), .B(n534), .C(n533), .D(n532), .Q(n541) );
  NAND22 U1620 ( .A(n333), .B(n332), .Q(o_data_Rs[7]) );
  NAND41 U1621 ( .A(n329), .B(n328), .C(n327), .D(n326), .Q(n330) );
  NAND41 U1622 ( .A(n325), .B(n324), .C(n323), .D(n322), .Q(n331) );
  NAND41 U1623 ( .A(n319), .B(n318), .C(n317), .D(n316), .Q(n320) );
  NAND41 U1624 ( .A(n315), .B(n314), .C(n313), .D(n312), .Q(n321) );
  NAND22 U1625 ( .A(n421), .B(n420), .Q(o_data_Rs[11]) );
  NAND41 U1626 ( .A(n417), .B(n416), .C(n415), .D(n414), .Q(n418) );
  AOI221 U1627 ( .A(n72), .B(regs[683]), .C(n65), .D(regs[651]), .Q(n414) );
  NAND41 U1628 ( .A(n413), .B(n412), .C(n411), .D(n410), .Q(n419) );
  AOI221 U1629 ( .A(n72), .B(regs[171]), .C(n65), .D(regs[139]), .Q(n410) );
  NAND41 U1630 ( .A(n407), .B(n406), .C(n405), .D(n404), .Q(n408) );
  NAND41 U1631 ( .A(n403), .B(n402), .C(n401), .D(n400), .Q(n409) );
  NAND22 U1632 ( .A(n443), .B(n442), .Q(o_data_Rs[12]) );
  NAND41 U1633 ( .A(n439), .B(n438), .C(n437), .D(n436), .Q(n440) );
  NAND41 U1634 ( .A(n435), .B(n434), .C(n433), .D(n432), .Q(n441) );
  NAND41 U1635 ( .A(n429), .B(n428), .C(n427), .D(n426), .Q(n430) );
  NAND41 U1636 ( .A(n425), .B(n424), .C(n423), .D(n422), .Q(n431) );
  NAND22 U1637 ( .A(n355), .B(n354), .Q(o_data_Rs[8]) );
  NAND41 U1638 ( .A(n351), .B(n350), .C(n349), .D(n348), .Q(n352) );
  NAND41 U1639 ( .A(n347), .B(n346), .C(n345), .D(n344), .Q(n353) );
  NAND41 U1640 ( .A(n341), .B(n340), .C(n339), .D(n338), .Q(n342) );
  NAND41 U1641 ( .A(n337), .B(n336), .C(n335), .D(n334), .Q(n343) );
  NAND22 U1642 ( .A(n531), .B(n530), .Q(o_data_Rs[16]) );
  NAND41 U1643 ( .A(n527), .B(n526), .C(n525), .D(n524), .Q(n528) );
  AOI221 U1644 ( .A(n72), .B(regs[688]), .C(n80), .D(regs[656]), .Q(n524) );
  NAND41 U1645 ( .A(n523), .B(n522), .C(n521), .D(n520), .Q(n529) );
  AOI221 U1646 ( .A(n72), .B(regs[176]), .C(n80), .D(regs[144]), .Q(n520) );
  NAND41 U1647 ( .A(n517), .B(n516), .C(n515), .D(n514), .Q(n518) );
  NAND41 U1648 ( .A(n513), .B(n512), .C(n511), .D(n510), .Q(n519) );
  AOI221 U1649 ( .A(n72), .B(regs[432]), .C(n65), .D(regs[400]), .Q(n510) );
  INV3 U1650 ( .A(i_addr_Rs[2]), .Q(n154) );
  NAND22 U1651 ( .A(n151), .B(i_addr_Rs[0]), .Q(n152) );
  INV6 U1652 ( .A(i_addr_Rs[1]), .Q(n151) );
  NAND22 U1653 ( .A(i_addr_Rs[2]), .B(i_addr_Rs[1]), .Q(n149) );
  NOR31 U1654 ( .A(i_addr_Rs[2]), .B(n150), .C(n151), .Q(n859) );
  AOI220 U1655 ( .A(n69), .B(regs[1014]), .C(n76), .D(regs[982]), .Q(n649) );
  AOI220 U1656 ( .A(n69), .B(regs[502]), .C(n76), .D(regs[470]), .Q(n645) );
  AOI220 U1657 ( .A(n66), .B(regs[610]), .C(n858), .D(regs[546]), .Q(n218) );
  AOI220 U1658 ( .A(n66), .B(regs[98]), .C(n858), .D(regs[34]), .Q(n214) );
  AOI220 U1659 ( .A(n66), .B(regs[866]), .C(n858), .D(regs[802]), .Q(n208) );
  AOI220 U1660 ( .A(n66), .B(regs[638]), .C(n858), .D(regs[574]), .Q(n834) );
  AOI220 U1661 ( .A(n66), .B(regs[126]), .C(n858), .D(regs[62]), .Q(n830) );
  AOI220 U1662 ( .A(n66), .B(regs[894]), .C(n858), .D(regs[830]), .Q(n824) );
  AOI220 U1663 ( .A(n66), .B(regs[382]), .C(n858), .D(regs[318]), .Q(n820) );
  AOI220 U1664 ( .A(n66), .B(regs[127]), .C(n858), .D(regs[63]), .Q(n854) );
  AOI220 U1665 ( .A(n72), .B(regs[959]), .C(n862), .D(regs[927]), .Q(n844) );
  AOI220 U1666 ( .A(n66), .B(regs[895]), .C(n858), .D(regs[831]), .Q(n846) );
  AOI220 U1667 ( .A(n66), .B(regs[383]), .C(n858), .D(regs[319]), .Q(n842) );
  AOI220 U1668 ( .A(n72), .B(regs[697]), .C(n862), .D(regs[665]), .Q(n722) );
  AOI220 U1669 ( .A(n71), .B(regs[695]), .C(n862), .D(regs[663]), .Q(n678) );
  AOI220 U1670 ( .A(n72), .B(regs[948]), .C(n862), .D(regs[916]), .Q(n602) );
  AOI220 U1671 ( .A(n55), .B(regs[89]), .C(n1584), .D(regs[25]), .Q(n1444) );
  AOI220 U1672 ( .A(n55), .B(regs[90]), .C(n1584), .D(regs[26]), .Q(n1466) );
  AOI220 U1673 ( .A(n55), .B(regs[91]), .C(n1584), .D(regs[27]), .Q(n1488) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, id_con_Wregwrite, ex_con_Wregwrite, mem_con_Wregwrite,
         for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst, ex_con_Mmemread,
         ex_con_Mmemwrite, ex_con_Malupc8, ex_con_Wmemtoreg, mem_con_Malupc8,
         mem_con_Wmemtoreg, wb_con_Wmemtoreg, u_fetch_jmux_i_addr_pc4_3_,
         u_fetch_jmux_i_addr_pc4_4_, u_fetch_jmux_i_addr_pc4_5_,
         u_fetch_jmux_i_addr_pc4_6_, u_fetch_jmux_i_addr_pc4_7_,
         u_fetch_jmux_i_addr_pc4_8_, u_fetch_jmux_i_addr_pc4_9_,
         u_fetch_jmux_i_addr_pc4_10_, u_fetch_jmux_i_addr_pc4_11_,
         u_fetch_jmux_i_addr_pc4_12_, u_fetch_jmux_i_addr_pc4_13_,
         u_fetch_jmux_i_addr_pc4_14_, u_fetch_jmux_i_addr_pc4_15_,
         u_fetch_jmux_i_addr_pc4_16_, u_fetch_jmux_i_addr_pc4_17_,
         u_fetch_jmux_i_addr_pc4_18_, u_fetch_jmux_i_addr_pc4_19_,
         u_fetch_jmux_i_addr_pc4_20_, u_fetch_jmux_i_addr_pc4_21_,
         u_fetch_jmux_i_addr_pc4_22_, u_fetch_jmux_i_addr_pc4_23_,
         u_fetch_jmux_i_addr_pc4_24_, u_fetch_jmux_i_addr_pc4_25_,
         u_fetch_jmux_i_addr_pc4_26_, u_fetch_jmux_i_addr_pc4_27_,
         u_fetch_jmux_i_addr_pc4_28_, u_fetch_jmux_i_addr_pc4_29_,
         u_fetch_jmux_i_addr_pc4_30_, u_fetch_jmux_i_addr_pc4_31_, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, u_decode_n23,
         u_decode_n17, u_decode_n6, u_decode_n4, u_decode_n3,
         u_decode_for_o_con_fb_0_, u_decode_for_o_con_fa_0_,
         u_decode_control_o_con_memtoreg, u_decode_control_o_con_memread,
         u_decode_jbcon_o_con_aluPC4, u_decode_control_o_con_regdst,
         u_decode_control_o_con_aluop_0_, u_decode_control_o_con_aluop_1_,
         u_decode_control_o_con_aluop_2_, u_decode_control_o_con_aluop_3_,
         u_decode_control_o_con_aluop_4_, u_decode_control_o_con_aluop_5_,
         u_decode_add_x_16_n209, u_decode_add_x_16_n208,
         u_decode_add_x_16_n205, u_decode_add_x_16_n203,
         u_decode_add_x_16_n202, u_decode_add_x_16_n199,
         u_decode_add_x_16_n197, u_decode_add_x_16_n193,
         u_decode_add_x_16_n191, u_decode_add_x_16_n189,
         u_decode_add_x_16_n186, u_decode_add_x_16_n183,
         u_decode_add_x_16_n182, u_decode_add_x_16_n180,
         u_decode_add_x_16_n179, u_decode_add_x_16_n178,
         u_decode_add_x_16_n177, u_decode_add_x_16_n176,
         u_decode_add_x_16_n175, u_decode_add_x_16_n174,
         u_decode_add_x_16_n173, u_decode_add_x_16_n172,
         u_decode_add_x_16_n171, u_decode_add_x_16_n170,
         u_decode_add_x_16_n169, u_decode_add_x_16_n168,
         u_decode_add_x_16_n167, u_decode_add_x_16_n166,
         u_decode_add_x_16_n162, u_decode_add_x_16_n161,
         u_decode_add_x_16_n160, u_decode_add_x_16_n159,
         u_decode_add_x_16_n158, u_decode_add_x_16_n157,
         u_decode_add_x_16_n156, u_decode_add_x_16_n155,
         u_decode_add_x_16_n154, u_decode_add_x_16_n153,
         u_decode_add_x_16_n152, u_decode_add_x_16_n151,
         u_decode_add_x_16_n150, u_decode_add_x_16_n149,
         u_decode_add_x_16_n148, u_decode_add_x_16_n147,
         u_decode_add_x_16_n146, u_decode_add_x_16_n145,
         u_decode_add_x_16_n144, u_decode_add_x_16_n143,
         u_decode_add_x_16_n142, u_decode_add_x_16_n141,
         u_decode_add_x_16_n140, u_decode_add_x_16_n139,
         u_decode_add_x_16_n138, u_decode_add_x_16_n137,
         u_decode_add_x_16_n136, u_decode_add_x_16_n135,
         u_decode_add_x_16_n131, u_decode_add_x_16_n130,
         u_decode_add_x_16_n129, u_decode_add_x_16_n128,
         u_decode_add_x_16_n127, u_decode_add_x_16_n126,
         u_decode_add_x_16_n125, u_decode_add_x_16_n124,
         u_decode_add_x_16_n123, u_decode_add_x_16_n122,
         u_decode_add_x_16_n121, u_decode_add_x_16_n120,
         u_decode_add_x_16_n119, u_decode_add_x_16_n118,
         u_decode_add_x_16_n117, u_decode_add_x_16_n116,
         u_decode_add_x_16_n115, u_decode_add_x_16_n114,
         u_decode_add_x_16_n113, u_decode_add_x_16_n112,
         u_decode_add_x_16_n111, u_decode_add_x_16_n110,
         u_decode_add_x_16_n109, u_decode_add_x_16_n108,
         u_decode_add_x_16_n107, u_decode_add_x_16_n106,
         u_decode_add_x_16_n105, u_decode_add_x_16_n104,
         u_decode_add_x_16_n103, u_decode_add_x_16_n102,
         u_decode_add_x_16_n101, u_decode_add_x_16_n99, u_decode_add_x_16_n97,
         u_decode_add_x_16_n96, u_decode_add_x_16_n95, u_decode_add_x_16_n94,
         u_decode_add_x_16_n93, u_decode_add_x_16_n92, u_decode_add_x_16_n91,
         u_decode_add_x_16_n90, u_decode_add_x_16_n89, u_decode_add_x_16_n88,
         u_decode_add_x_16_n87, u_decode_add_x_16_n86, u_decode_add_x_16_n85,
         u_decode_add_x_16_n84, u_decode_add_x_16_n83, u_decode_add_x_16_n82,
         u_decode_add_x_16_n81, u_decode_add_x_16_n80, u_decode_add_x_16_n79,
         u_decode_add_x_16_n78, u_decode_add_x_16_n77, u_decode_add_x_16_n76,
         u_decode_add_x_16_n75, u_decode_add_x_16_n74, u_decode_add_x_16_n73,
         u_decode_add_x_16_n72, u_decode_add_x_16_n71, u_decode_add_x_16_n70,
         u_decode_add_x_16_n69, u_decode_add_x_16_n68, u_decode_add_x_16_n67,
         u_decode_add_x_16_n66, u_decode_add_x_16_n65, u_decode_add_x_16_n64,
         u_decode_add_x_16_n63, u_decode_add_x_16_n62, u_decode_add_x_16_n59,
         u_decode_add_x_16_n58, u_decode_add_x_16_n57, u_decode_add_x_16_n56,
         u_decode_add_x_16_n55, u_decode_add_x_16_n54, u_decode_add_x_16_n53,
         u_decode_add_x_16_n52, u_decode_add_x_16_n51, u_decode_add_x_16_n50,
         u_decode_add_x_16_n49, u_decode_add_x_16_n48, u_decode_add_x_16_n47,
         u_decode_add_x_16_n46, u_decode_add_x_16_n45, u_decode_add_x_16_n44,
         u_decode_add_x_16_n43, u_decode_add_x_16_n42, u_decode_add_x_16_n41,
         u_decode_add_x_16_n40, u_decode_add_x_16_n39, u_decode_add_x_16_n37,
         u_decode_add_x_16_n36, u_decode_add_x_16_n35, u_decode_add_x_16_n34,
         u_decode_add_x_16_n33, u_decode_add_x_16_n32, u_decode_add_x_16_n31,
         u_decode_add_x_16_n30, u_decode_add_x_16_n27, u_decode_add_x_16_n26,
         u_decode_add_x_16_n23, u_decode_add_x_16_n21, u_decode_add_x_16_n20,
         u_decode_add_x_16_n17, u_decode_add_x_16_n15, u_decode_add_x_16_n14,
         u_decode_add_x_16_n11, u_decode_add_x_16_n9, u_decode_add_x_16_n7,
         u_decode_add_x_16_n6, u_decode_add_x_16_n5, u_decode_add_x_16_n4,
         u_decode_add_x_16_n3, u_decode_add_x_16_n1, add_x_4_n116,
         add_x_4_n111, add_x_4_n110, add_x_4_n107, add_x_4_n104, add_x_4_n103,
         add_x_4_n102, add_x_4_n98, add_x_4_n95, add_x_4_n94, add_x_4_n91,
         add_x_4_n88, add_x_4_n87, add_x_4_n86, add_x_4_n85, add_x_4_n82,
         add_x_4_n79, add_x_4_n78, add_x_4_n77, add_x_4_n73, add_x_4_n70,
         add_x_4_n69, add_x_4_n68, add_x_4_n67, add_x_4_n64, add_x_4_n61,
         add_x_4_n60, add_x_4_n57, add_x_4_n54, add_x_4_n53, add_x_4_n52,
         add_x_4_n51, add_x_4_n50, add_x_4_n46, add_x_4_n43, add_x_4_n42,
         add_x_4_n39, add_x_4_n36, add_x_4_n35, add_x_4_n34, add_x_4_n33,
         add_x_4_n30, add_x_4_n27, add_x_4_n26, add_x_4_n23, add_x_4_n18,
         add_x_4_n17, add_x_4_n14, add_x_4_n12, add_x_4_n11, add_x_4_n8,
         add_x_4_n7, add_x_4_n6, add_x_4_n4, add_x_4_n1, add_x_1_n118,
         add_x_1_n117, add_x_1_n111, add_x_1_n110, add_x_1_n109, add_x_1_n108,
         add_x_1_n102, add_x_1_n101, add_x_1_n95, add_x_1_n94, add_x_1_n93,
         add_x_1_n92, add_x_1_n86, add_x_1_n85, add_x_1_n84, add_x_1_n83,
         add_x_1_n77, add_x_1_n76, add_x_1_n75, add_x_1_n74, add_x_1_n73,
         add_x_1_n67, add_x_1_n66, add_x_1_n65, add_x_1_n64, add_x_1_n58,
         add_x_1_n57, add_x_1_n56, add_x_1_n55, add_x_1_n54, add_x_1_n53,
         add_x_1_n47, add_x_1_n46, add_x_1_n40, add_x_1_n39, add_x_1_n38,
         add_x_1_n37, add_x_1_n36, add_x_1_n35, add_x_1_n29, add_x_1_n28,
         add_x_1_n27, add_x_1_n26, add_x_1_n18, add_x_1_n17, add_x_1_n11,
         add_x_1_n10, add_x_1_n9, add_x_1_n7, add_x_1_n4, add_x_1_n2, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599;
  wire   [22:3] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [27:2] id_addr_pc4;
  wire   [31:26] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] wb_data_memout;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [1:0] for_o_con_Efamux;
  wire   [1:0] for_o_con_Efbmux;
  wire   [31:0] for_famemout;
  wire   [31:0] for_fbmemout;
  wire   [31:0] mem_data_alures;
  wire   [31:2] mem_data_pc4;
  wire   [31:0] u_mem_resmux_o_data_alu;
  wire   [31:0] u_mem_pc8;
  wire   [2:0] u_decode_jbcon_o_con_bop;
  wire   [31:0] u_decode_pcadd_o_addr_pcbranchE;
  wire   [31:0] u_decode_fbmemmux_o_data_fmem;
  wire   [31:0] u_decode_famemmux_o_data_fmem;
  wire   [31:0] u_decode_regbank_o_data_Rt;

  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext({n308, 
        n308, n308, n308, n308, n308, n308, n308, n308, n308, n308, n308, n308, 
        n308, n308, ex_data_immext[31], ex_addr_rd, ex_data_immext[10:0]}), 
        .i_addr_rt(ex_addr_rt), .i_addr_rd({n308, n308, n308, n308, n308}), 
        .i_data_FEalures(data_address), .i_data_FMalures(mem_data_alures), 
        .i_data_famemout(for_famemout), .i_data_fbmemout(for_fbmemout), 
        .i_con_Efamux(for_o_con_Efamux), .i_con_Efbmux(for_o_con_Efbmux), 
        .i_con_Ealuop(ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), 
        .i_con_Mmemwrite(ex_con_Mmemwrite), .i_con_Malupc8(ex_con_Malupc8), 
        .i_con_Wmemtoreg(ex_con_Wmemtoreg), .i_con_Wregwrite(ex_con_Wregwrite), 
        .i_con_bop(ex_con_bop), .o_data_alures(data_address), .o_data_rt(
        write_data), .o_addr_regdst(mem_addr_regdst), .o_con_Mmemread(mem_read), .o_con_Mmemwrite(mem_write), .o_con_Malupc8(mem_con_Malupc8), 
        .o_con_Wmemtoreg(mem_con_Wmemtoreg), .o_con_Wregwrite(
        mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), .o_addr_Mrt(
        for_addr_rtM), .o_con_ifbranch(if_con_b), .o_data_pc4_31__BAR(
        mem_data_pc4[31]), .o_data_pc4_29_(mem_data_pc4[29]), .o_data_pc4_27_(
        mem_data_pc4[27]), .o_data_pc4_26_(mem_data_pc4[26]), .o_data_pc4_25_(
        mem_data_pc4[25]), .o_data_pc4_24_(mem_data_pc4[24]), .o_data_pc4_23_(
        mem_data_pc4[23]), .o_data_pc4_22_(mem_data_pc4[22]), .o_data_pc4_21_(
        mem_data_pc4[21]), .o_data_pc4_20_(mem_data_pc4[20]), .o_data_pc4_19_(
        mem_data_pc4[19]), .o_data_pc4_18_(mem_data_pc4[18]), .o_data_pc4_17_(
        mem_data_pc4[17]), .o_data_pc4_16_(mem_data_pc4[16]), .o_data_pc4_15_(
        mem_data_pc4[15]), .o_data_pc4_14_(mem_data_pc4[14]), .o_data_pc4_13_(
        mem_data_pc4[13]), .o_data_pc4_12_(mem_data_pc4[12]), .o_data_pc4_11_(
        mem_data_pc4[11]), .o_data_pc4_10_(mem_data_pc4[10]), .o_data_pc4_9_(
        mem_data_pc4[9]), .o_data_pc4_8_(mem_data_pc4[8]), .o_data_pc4_7_(
        mem_data_pc4[7]), .o_data_pc4_6_(mem_data_pc4[6]), .o_data_pc4_5_(
        mem_data_pc4[5]), .o_data_pc4_4_(mem_data_pc4[4]), .o_data_pc4_3_(
        mem_data_pc4[3]), .o_data_pc4_2_(mem_data_pc4[2]), .o_data_pc4_1_(
        u_mem_pc8[1]), .o_data_pc4_0_(u_mem_pc8[0]), .o_data_pc4_30__BAR(
        mem_data_pc4[30]), .o_data_pc4_28__BAR(mem_data_pc4[28]) );
  DFC1 u_fetch_pipe_pc4_reg_0_ ( .D(instruction_address[0]), .C(clk), .RN(
        rst_n), .Q(u_decode_pcadd_o_addr_pcbranchE[0]) );
  DFC1 u_fetch_pipe_pc4_reg_1_ ( .D(instruction_address[1]), .C(clk), .RN(
        rst_n), .Q(u_decode_pcadd_o_addr_pcbranchE[1]) );
  DFC1 u_fetch_pipe_pc4_reg_2_ ( .D(n283), .C(clk), .RN(rst_n), .Q(
        id_addr_pc4[2]) );
  DFC1 u_fetch_pipe_pc4_reg_3_ ( .D(u_fetch_jmux_i_addr_pc4_3_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[3]) );
  DFC1 u_fetch_pipe_pc4_reg_4_ ( .D(u_fetch_jmux_i_addr_pc4_4_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[4]) );
  DFC1 u_fetch_pipe_pc4_reg_5_ ( .D(u_fetch_jmux_i_addr_pc4_5_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[5]) );
  DFC1 u_fetch_pipe_pc4_reg_6_ ( .D(u_fetch_jmux_i_addr_pc4_6_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[6]) );
  DFC1 u_fetch_pipe_pc4_reg_7_ ( .D(u_fetch_jmux_i_addr_pc4_7_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[7]) );
  DFC1 u_fetch_pipe_pc4_reg_8_ ( .D(u_fetch_jmux_i_addr_pc4_8_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[8]) );
  DFC1 u_fetch_pipe_pc4_reg_9_ ( .D(u_fetch_jmux_i_addr_pc4_9_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[9]) );
  DFC1 u_fetch_pipe_pc4_reg_10_ ( .D(u_fetch_jmux_i_addr_pc4_10_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[10]) );
  DFC1 u_fetch_pipe_pc4_reg_11_ ( .D(u_fetch_jmux_i_addr_pc4_11_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[11]) );
  DFC1 u_fetch_pipe_pc4_reg_12_ ( .D(u_fetch_jmux_i_addr_pc4_12_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[12]) );
  DFC1 u_fetch_pipe_pc4_reg_13_ ( .D(u_fetch_jmux_i_addr_pc4_13_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[13]) );
  DFC1 u_fetch_pipe_pc4_reg_14_ ( .D(u_fetch_jmux_i_addr_pc4_14_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[14]) );
  DFC1 u_fetch_pipe_pc4_reg_15_ ( .D(u_fetch_jmux_i_addr_pc4_15_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[15]) );
  DFC1 u_fetch_pipe_pc4_reg_16_ ( .D(u_fetch_jmux_i_addr_pc4_16_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[16]) );
  DFC1 u_fetch_pipe_pc4_reg_17_ ( .D(u_fetch_jmux_i_addr_pc4_17_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[17]) );
  DFC1 u_fetch_pipe_pc4_reg_18_ ( .D(u_fetch_jmux_i_addr_pc4_18_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[18]) );
  DFC1 u_fetch_pipe_pc4_reg_19_ ( .D(u_fetch_jmux_i_addr_pc4_19_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[19]) );
  DFC1 u_fetch_pipe_pc4_reg_20_ ( .D(u_fetch_jmux_i_addr_pc4_20_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[20]) );
  DFC1 u_fetch_pipe_pc4_reg_21_ ( .D(u_fetch_jmux_i_addr_pc4_21_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[21]) );
  DFC1 u_fetch_pipe_pc4_reg_22_ ( .D(u_fetch_jmux_i_addr_pc4_22_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[22]) );
  DFC1 u_fetch_pipe_pc4_reg_23_ ( .D(u_fetch_jmux_i_addr_pc4_23_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[23]) );
  DFC1 u_fetch_pipe_pc4_reg_24_ ( .D(u_fetch_jmux_i_addr_pc4_24_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[24]) );
  DFC1 u_fetch_pipe_pc4_reg_25_ ( .D(u_fetch_jmux_i_addr_pc4_25_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[25]) );
  DFC1 u_fetch_pipe_pc4_reg_26_ ( .D(u_fetch_jmux_i_addr_pc4_26_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[26]) );
  DFC1 u_fetch_pipe_pc4_reg_27_ ( .D(u_fetch_jmux_i_addr_pc4_27_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[27]) );
  DFC1 u_fetch_pipe_pc4_reg_28_ ( .D(u_fetch_jmux_i_addr_pc4_28_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[28]) );
  DFC1 u_fetch_pipe_pc4_reg_29_ ( .D(u_fetch_jmux_i_addr_pc4_29_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[29]) );
  DFC1 u_fetch_pipe_pc4_reg_30_ ( .D(u_fetch_jmux_i_addr_pc4_30_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[30]) );
  DFC1 u_fetch_pipe_pc4_reg_31_ ( .D(u_fetch_jmux_i_addr_pc4_31_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[31]) );
  DFC1 u_fetch_pipe_instr_reg_0_ ( .D(read_instruction[0]), .C(clk), .RN(rst_n), .Q(if_addr_j[2]), .QN(n259) );
  DFC1 u_fetch_pipe_instr_reg_6_ ( .D(read_instruction[6]), .C(clk), .RN(rst_n), .Q(if_addr_j[8]) );
  DFC1 u_fetch_pipe_instr_reg_8_ ( .D(read_instruction[8]), .C(clk), .RN(rst_n), .Q(if_addr_j[10]) );
  DFC1 u_fetch_pipe_instr_reg_9_ ( .D(read_instruction[9]), .C(clk), .RN(rst_n), .Q(if_addr_j[11]) );
  DFC1 u_fetch_pipe_instr_reg_10_ ( .D(read_instruction[10]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[12]) );
  DFC1 u_fetch_pipe_instr_reg_11_ ( .D(read_instruction[11]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[13]) );
  DFC1 u_fetch_pipe_instr_reg_12_ ( .D(read_instruction[12]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[14]) );
  DFC1 u_fetch_pipe_instr_reg_13_ ( .D(read_instruction[13]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[15]) );
  DFC1 u_fetch_pipe_instr_reg_14_ ( .D(read_instruction[14]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[16]) );
  DFC1 u_fetch_pipe_instr_reg_26_ ( .D(read_instruction[26]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[26]), .QN(n257) );
  DFC1 u_fetch_pipe_instr_reg_27_ ( .D(read_instruction[27]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[27]), .QN(n251) );
  DFC1 u_fetch_pipe_instr_reg_28_ ( .D(read_instruction[28]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[28]), .QN(n253) );
  DFC1 u_fetch_pipe_instr_reg_30_ ( .D(read_instruction[30]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[30]), .QN(n255) );
  DFC1 u_fetch_pipe_instr_reg_31_ ( .D(read_instruction[31]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[31]), .QN(n262) );
  DFC1 u_mem_pipe_data_memout_reg_0_ ( .D(read_data[0]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[0]) );
  DFC1 u_mem_pipe_data_memout_reg_1_ ( .D(read_data[1]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[1]) );
  DFC1 u_mem_pipe_data_memout_reg_2_ ( .D(read_data[2]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[2]) );
  DFC1 u_mem_pipe_data_memout_reg_3_ ( .D(read_data[3]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[3]) );
  DFC1 u_mem_pipe_data_memout_reg_4_ ( .D(read_data[4]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[4]) );
  DFC1 u_mem_pipe_data_memout_reg_5_ ( .D(read_data[5]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[5]) );
  DFC1 u_mem_pipe_data_memout_reg_6_ ( .D(read_data[6]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[6]) );
  DFC1 u_mem_pipe_data_memout_reg_7_ ( .D(read_data[7]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[7]) );
  DFC1 u_mem_pipe_data_memout_reg_8_ ( .D(read_data[8]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[8]) );
  DFC1 u_mem_pipe_data_memout_reg_9_ ( .D(read_data[9]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[9]) );
  DFC1 u_mem_pipe_data_memout_reg_10_ ( .D(read_data[10]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[10]) );
  DFC1 u_mem_pipe_data_memout_reg_11_ ( .D(read_data[11]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[11]) );
  DFC1 u_mem_pipe_data_memout_reg_12_ ( .D(read_data[12]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[12]) );
  DFC1 u_mem_pipe_data_memout_reg_13_ ( .D(read_data[13]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[13]) );
  DFC1 u_mem_pipe_data_memout_reg_14_ ( .D(read_data[14]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[14]) );
  DFC1 u_mem_pipe_data_memout_reg_15_ ( .D(read_data[15]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[15]) );
  DFC1 u_mem_pipe_data_memout_reg_16_ ( .D(read_data[16]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[16]) );
  DFC1 u_mem_pipe_data_memout_reg_17_ ( .D(read_data[17]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[17]) );
  DFC1 u_mem_pipe_data_memout_reg_18_ ( .D(read_data[18]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[18]) );
  DFC1 u_mem_pipe_data_memout_reg_19_ ( .D(read_data[19]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[19]) );
  DFC1 u_mem_pipe_data_memout_reg_20_ ( .D(read_data[20]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[20]) );
  DFC1 u_mem_pipe_data_memout_reg_21_ ( .D(read_data[21]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[21]) );
  DFC1 u_mem_pipe_data_memout_reg_22_ ( .D(read_data[22]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[22]) );
  DFC1 u_mem_pipe_data_memout_reg_23_ ( .D(read_data[23]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[23]) );
  DFC1 u_mem_pipe_data_memout_reg_24_ ( .D(read_data[24]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[24]) );
  DFC1 u_mem_pipe_data_memout_reg_25_ ( .D(read_data[25]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[25]) );
  DFC1 u_mem_pipe_data_memout_reg_26_ ( .D(read_data[26]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[26]) );
  DFC1 u_mem_pipe_data_memout_reg_27_ ( .D(read_data[27]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[27]) );
  DFC1 u_mem_pipe_data_memout_reg_28_ ( .D(read_data[28]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[28]) );
  DFC1 u_mem_pipe_data_memout_reg_29_ ( .D(read_data[29]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[29]) );
  DFC1 u_mem_pipe_data_memout_reg_30_ ( .D(read_data[30]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[30]) );
  DFC1 u_mem_pipe_data_memout_reg_31_ ( .D(read_data[31]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[31]) );
  DFC1 u_mem_pipe_rt_reg_4_ ( .D(for_addr_rtM[4]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[4]) );
  DFC1 u_mem_pipe_con_FWmemread_reg ( .D(ex_con_Mmemread), .C(clk), .RN(rst_n), 
        .Q(for_FWmemread) );
  DFC1 u_mem_pipe_rt_reg_0_ ( .D(for_addr_rtM[0]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[0]) );
  DFC1 u_mem_pipe_rt_reg_1_ ( .D(for_addr_rtM[1]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[1]) );
  DFC1 u_mem_pipe_rt_reg_2_ ( .D(for_addr_rtM[2]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[2]) );
  DFC1 u_mem_pipe_rt_reg_3_ ( .D(for_addr_rtM[3]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[3]) );
  DFC1 u_mem_pipe_con_Wregwrite_reg ( .D(mem_con_Wregwrite), .C(clk), .RN(
        rst_n), .Q(id_con_Wregwrite) );
  DFC1 u_mem_pipe_addr_regdst_reg_0_ ( .D(mem_addr_regdst[0]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[0]) );
  DFC1 u_mem_pipe_addr_regdst_reg_1_ ( .D(mem_addr_regdst[1]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[1]) );
  DFC1 u_mem_pipe_addr_regdst_reg_2_ ( .D(mem_addr_regdst[2]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[2]) );
  DFC1 u_mem_pipe_addr_regdst_reg_4_ ( .D(mem_addr_regdst[4]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[4]) );
  DFC1 u_mem_pipe_data_alures_reg_0_ ( .D(u_mem_resmux_o_data_alu[0]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[0]) );
  DFC1 u_mem_pipe_data_alures_reg_1_ ( .D(u_mem_resmux_o_data_alu[1]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[1]) );
  DFC1 u_mem_pipe_data_alures_reg_2_ ( .D(u_mem_resmux_o_data_alu[2]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[2]) );
  DFC1 u_mem_pipe_data_alures_reg_3_ ( .D(u_mem_resmux_o_data_alu[3]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[3]) );
  DFC1 u_mem_pipe_data_alures_reg_4_ ( .D(u_mem_resmux_o_data_alu[4]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[4]) );
  DFC1 u_mem_pipe_data_alures_reg_5_ ( .D(u_mem_resmux_o_data_alu[5]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[5]) );
  DFC1 u_mem_pipe_data_alures_reg_7_ ( .D(u_mem_resmux_o_data_alu[7]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[7]) );
  DFC1 u_mem_pipe_data_alures_reg_8_ ( .D(u_mem_resmux_o_data_alu[8]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[8]) );
  DFC1 u_mem_pipe_data_alures_reg_9_ ( .D(u_mem_resmux_o_data_alu[9]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[9]) );
  DFC1 u_mem_pipe_data_alures_reg_10_ ( .D(u_mem_resmux_o_data_alu[10]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[10]) );
  DFC1 u_mem_pipe_data_alures_reg_11_ ( .D(u_mem_resmux_o_data_alu[11]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[11]) );
  DFC1 u_mem_pipe_data_alures_reg_12_ ( .D(u_mem_resmux_o_data_alu[12]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[12]) );
  DFC1 u_mem_pipe_data_alures_reg_15_ ( .D(u_mem_resmux_o_data_alu[15]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[15]) );
  DFC1 u_mem_pipe_data_alures_reg_16_ ( .D(u_mem_resmux_o_data_alu[16]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[16]) );
  DFC1 u_mem_pipe_data_alures_reg_17_ ( .D(u_mem_resmux_o_data_alu[17]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[17]) );
  DFC1 u_mem_pipe_data_alures_reg_18_ ( .D(u_mem_resmux_o_data_alu[18]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[18]) );
  DFC1 u_mem_pipe_data_alures_reg_20_ ( .D(u_mem_resmux_o_data_alu[20]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[20]) );
  DFC1 u_mem_pipe_data_alures_reg_21_ ( .D(u_mem_resmux_o_data_alu[21]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[21]) );
  DFC1 u_mem_pipe_data_alures_reg_22_ ( .D(u_mem_resmux_o_data_alu[22]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[22]) );
  DFC1 u_mem_pipe_data_alures_reg_23_ ( .D(u_mem_resmux_o_data_alu[23]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[23]) );
  DFC1 u_mem_pipe_data_alures_reg_24_ ( .D(u_mem_resmux_o_data_alu[24]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[24]) );
  DFC1 u_mem_pipe_data_alures_reg_25_ ( .D(u_mem_resmux_o_data_alu[25]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[25]) );
  DFC1 u_mem_pipe_data_alures_reg_26_ ( .D(u_mem_resmux_o_data_alu[26]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[26]) );
  DFC1 u_mem_pipe_data_alures_reg_27_ ( .D(u_mem_resmux_o_data_alu[27]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[27]) );
  DFC1 u_mem_pipe_data_alures_reg_28_ ( .D(u_mem_resmux_o_data_alu[28]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[28]) );
  DFC1 u_mem_pipe_data_alures_reg_29_ ( .D(u_mem_resmux_o_data_alu[29]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[29]) );
  DFC1 u_mem_pipe_data_alures_reg_31_ ( .D(u_mem_resmux_o_data_alu[31]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[31]) );
  DFC1 u_fetch_u_pc_program_counter_reg_0_ ( .D(n137), .C(clk), .RN(rst_n), 
        .Q(instruction_address[0]) );
  DFC1 u_fetch_u_pc_program_counter_reg_1_ ( .D(n136), .C(clk), .RN(rst_n), 
        .Q(instruction_address[1]) );
  DFC1 u_fetch_u_pc_program_counter_reg_2_ ( .D(n135), .C(clk), .RN(rst_n), 
        .Q(instruction_address[2]), .QN(n283) );
  DFC1 u_fetch_u_pc_program_counter_reg_3_ ( .D(n134), .C(clk), .RN(rst_n), 
        .Q(instruction_address[3]), .QN(n296) );
  DFC1 u_fetch_u_pc_program_counter_reg_4_ ( .D(n133), .C(clk), .RN(rst_n), 
        .Q(instruction_address[4]), .QN(n274) );
  DFC1 u_fetch_u_pc_program_counter_reg_5_ ( .D(n132), .C(clk), .RN(rst_n), 
        .Q(instruction_address[5]), .QN(n292) );
  DFC1 u_fetch_u_pc_program_counter_reg_6_ ( .D(n131), .C(clk), .RN(rst_n), 
        .Q(instruction_address[6]), .QN(n295) );
  DFC1 u_fetch_u_pc_program_counter_reg_7_ ( .D(n130), .C(clk), .RN(rst_n), 
        .Q(instruction_address[7]), .QN(n291) );
  DFC1 u_fetch_u_pc_program_counter_reg_8_ ( .D(n129), .C(clk), .RN(rst_n), 
        .Q(instruction_address[8]), .QN(n273) );
  DFC1 u_fetch_u_pc_program_counter_reg_9_ ( .D(n128), .C(clk), .RN(rst_n), 
        .Q(instruction_address[9]), .QN(n290) );
  DFC1 u_fetch_u_pc_program_counter_reg_10_ ( .D(n127), .C(clk), .RN(rst_n), 
        .Q(instruction_address[10]), .QN(n272) );
  DFC1 u_fetch_u_pc_program_counter_reg_11_ ( .D(n126), .C(clk), .RN(rst_n), 
        .Q(instruction_address[11]), .QN(n289) );
  DFC1 u_fetch_u_pc_program_counter_reg_12_ ( .D(n125), .C(clk), .RN(rst_n), 
        .Q(instruction_address[12]), .QN(n294) );
  DFC1 u_fetch_u_pc_program_counter_reg_13_ ( .D(n124), .C(clk), .RN(rst_n), 
        .Q(instruction_address[13]), .QN(n288) );
  DFC1 u_fetch_u_pc_program_counter_reg_14_ ( .D(n123), .C(clk), .RN(rst_n), 
        .Q(instruction_address[14]), .QN(n271) );
  DFC1 u_fetch_u_pc_program_counter_reg_15_ ( .D(n122), .C(clk), .RN(rst_n), 
        .Q(instruction_address[15]), .QN(n287) );
  DFC1 u_fetch_u_pc_program_counter_reg_16_ ( .D(n121), .C(clk), .RN(rst_n), 
        .Q(instruction_address[16]), .QN(n270) );
  DFC1 u_fetch_u_pc_program_counter_reg_17_ ( .D(n120), .C(clk), .RN(rst_n), 
        .Q(instruction_address[17]), .QN(n286) );
  DFC1 u_fetch_u_pc_program_counter_reg_18_ ( .D(n119), .C(clk), .RN(rst_n), 
        .Q(instruction_address[18]), .QN(n293) );
  DFC1 u_fetch_u_pc_program_counter_reg_19_ ( .D(n118), .C(clk), .RN(rst_n), 
        .Q(instruction_address[19]), .QN(n285) );
  DFC1 u_fetch_u_pc_program_counter_reg_20_ ( .D(n117), .C(clk), .RN(rst_n), 
        .Q(instruction_address[20]), .QN(n269) );
  DFC1 u_fetch_u_pc_program_counter_reg_21_ ( .D(n116), .C(clk), .RN(rst_n), 
        .Q(instruction_address[21]), .QN(n284) );
  DFC1 u_fetch_u_pc_program_counter_reg_22_ ( .D(n115), .C(clk), .RN(rst_n), 
        .Q(instruction_address[22]), .QN(n268) );
  DFC1 u_fetch_u_pc_program_counter_reg_23_ ( .D(n114), .C(clk), .RN(rst_n), 
        .Q(instruction_address[23]), .QN(n267) );
  DFC1 u_fetch_u_pc_program_counter_reg_24_ ( .D(n113), .C(clk), .RN(rst_n), 
        .Q(instruction_address[24]), .QN(n263) );
  DFC1 u_fetch_u_pc_program_counter_reg_25_ ( .D(n112), .C(clk), .RN(rst_n), 
        .Q(instruction_address[25]), .QN(n266) );
  DFC1 u_fetch_u_pc_program_counter_reg_26_ ( .D(n111), .C(clk), .RN(rst_n), 
        .Q(instruction_address[26]), .QN(n252) );
  DFC1 u_fetch_u_pc_program_counter_reg_27_ ( .D(n110), .C(clk), .RN(rst_n), 
        .Q(instruction_address[27]), .QN(n276) );
  DFC1 u_fetch_u_pc_program_counter_reg_28_ ( .D(n109), .C(clk), .RN(rst_n), 
        .Q(instruction_address[28]), .QN(n265) );
  DFC1 u_fetch_u_pc_program_counter_reg_29_ ( .D(n108), .C(clk), .RN(rst_n), 
        .Q(instruction_address[29]), .QN(n275) );
  DFC1 u_fetch_u_pc_program_counter_reg_30_ ( .D(n107), .C(clk), .RN(rst_n), 
        .Q(instruction_address[30]), .QN(n264) );
  DFC1 u_fetch_u_pc_program_counter_reg_31_ ( .D(n138), .C(clk), .RN(rst_n), 
        .Q(instruction_address[31]) );
  DFC1 u_decode_pipe_addr_branch_reg_0_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[0]), .C(clk), .RN(rst_n), .Q(
        ex_data_pc4[0]) );
  DFC1 u_decode_pipe_addr_branch_reg_1_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[1]), .C(clk), .RN(rst_n), .Q(
        ex_data_pc4[1]) );
  DFC1 u_decode_pipe_addr_branch_reg_3_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[3]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[3]) );
  DFC1 u_decode_pipe_addr_branch_reg_4_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[4]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[4]) );
  DFC1 u_decode_pipe_addr_branch_reg_5_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[5]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[5]) );
  DFC1 u_decode_pipe_addr_branch_reg_6_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[6]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[6]) );
  DFC1 u_decode_pipe_addr_branch_reg_7_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[7]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[7]) );
  DFC1 u_decode_pipe_addr_branch_reg_8_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[8]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[8]) );
  DFC1 u_decode_pipe_addr_branch_reg_9_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[9]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[9]) );
  DFC1 u_decode_pipe_addr_branch_reg_10_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[10]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[10]) );
  DFC1 u_decode_pipe_addr_branch_reg_11_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[11]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[11]) );
  DFC1 u_decode_pipe_addr_branch_reg_12_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[12]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[12]) );
  DFC1 u_decode_pipe_addr_branch_reg_13_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[13]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[13]) );
  DFC1 u_decode_pipe_addr_branch_reg_14_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[14]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[14]) );
  DFC1 u_decode_pipe_addr_branch_reg_15_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[15]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[15]) );
  DFC1 u_decode_pipe_addr_branch_reg_16_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[16]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[16]) );
  DFC1 u_decode_pipe_addr_branch_reg_17_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[17]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[17]) );
  DFC1 u_decode_pipe_addr_branch_reg_18_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[18]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[18]) );
  DFC1 u_decode_pipe_addr_branch_reg_19_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[19]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[19]) );
  DFC1 u_decode_pipe_addr_branch_reg_20_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[20]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[20]) );
  DFC1 u_decode_pipe_addr_branch_reg_21_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[21]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[21]) );
  DFC1 u_decode_pipe_addr_branch_reg_22_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[22]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[22]) );
  DFC1 u_decode_pipe_addr_branch_reg_23_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[23]), .C(clk), .RN(rst_n), .QN(n306)
         );
  DFC1 u_decode_pipe_addr_branch_reg_24_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[24]), .C(clk), .RN(rst_n), .QN(n305)
         );
  DFC1 u_decode_pipe_addr_branch_reg_25_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[25]), .C(clk), .RN(rst_n), .QN(n304)
         );
  DFC1 u_decode_pipe_addr_branch_reg_26_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[26]), .C(clk), .RN(rst_n), .QN(n303)
         );
  DFC1 u_decode_pipe_addr_branch_reg_27_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[27]), .C(clk), .RN(rst_n), .QN(n302)
         );
  DFC1 u_decode_pipe_addr_branch_reg_28_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[28]), .C(clk), .RN(rst_n), .QN(n301)
         );
  DFC1 u_decode_pipe_addr_branch_reg_29_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[29]), .C(clk), .RN(rst_n), .QN(n300)
         );
  DFC1 u_decode_pipe_addr_branch_reg_30_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[30]), .C(clk), .RN(rst_n), .QN(n299)
         );
  DFC1 u_decode_pipe_addr_branch_reg_31_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[31]), .C(clk), .RN(rst_n), .QN(n298)
         );
  DFC1 u_decode_pipe_Fbmemout_reg_0_ ( .D(u_decode_fbmemmux_o_data_fmem[0]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[0]) );
  DFC1 u_decode_pipe_Fbmemout_reg_1_ ( .D(u_decode_fbmemmux_o_data_fmem[1]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[1]) );
  DFC1 u_decode_pipe_Fbmemout_reg_2_ ( .D(u_decode_fbmemmux_o_data_fmem[2]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[2]) );
  DFC1 u_decode_pipe_Fbmemout_reg_3_ ( .D(u_decode_fbmemmux_o_data_fmem[3]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[3]) );
  DFC1 u_decode_pipe_Fbmemout_reg_4_ ( .D(u_decode_fbmemmux_o_data_fmem[4]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[4]) );
  DFC1 u_decode_pipe_Fbmemout_reg_5_ ( .D(u_decode_fbmemmux_o_data_fmem[5]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[5]) );
  DFC1 u_decode_pipe_Fbmemout_reg_6_ ( .D(u_decode_fbmemmux_o_data_fmem[6]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[6]) );
  DFC1 u_decode_pipe_Fbmemout_reg_7_ ( .D(u_decode_fbmemmux_o_data_fmem[7]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[7]) );
  DFC1 u_decode_pipe_Fbmemout_reg_8_ ( .D(u_decode_fbmemmux_o_data_fmem[8]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[8]) );
  DFC1 u_decode_pipe_Fbmemout_reg_9_ ( .D(u_decode_fbmemmux_o_data_fmem[9]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[9]) );
  DFC1 u_decode_pipe_Fbmemout_reg_10_ ( .D(u_decode_fbmemmux_o_data_fmem[10]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[10]) );
  DFC1 u_decode_pipe_Fbmemout_reg_12_ ( .D(u_decode_fbmemmux_o_data_fmem[12]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[12]) );
  DFC1 u_decode_pipe_Fbmemout_reg_13_ ( .D(u_decode_fbmemmux_o_data_fmem[13]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[13]) );
  DFC1 u_decode_pipe_Fbmemout_reg_14_ ( .D(u_decode_fbmemmux_o_data_fmem[14]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[14]) );
  DFC1 u_decode_pipe_Fbmemout_reg_15_ ( .D(u_decode_fbmemmux_o_data_fmem[15]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[15]) );
  DFC1 u_decode_pipe_Fbmemout_reg_16_ ( .D(u_decode_fbmemmux_o_data_fmem[16]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[16]) );
  DFC1 u_decode_pipe_Fbmemout_reg_17_ ( .D(u_decode_fbmemmux_o_data_fmem[17]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[17]) );
  DFC1 u_decode_pipe_Fbmemout_reg_18_ ( .D(u_decode_fbmemmux_o_data_fmem[18]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[18]) );
  DFC1 u_decode_pipe_Fbmemout_reg_19_ ( .D(u_decode_fbmemmux_o_data_fmem[19]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[19]) );
  DFC1 u_decode_pipe_Fbmemout_reg_20_ ( .D(u_decode_fbmemmux_o_data_fmem[20]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[20]) );
  DFC1 u_decode_pipe_Fbmemout_reg_21_ ( .D(u_decode_fbmemmux_o_data_fmem[21]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[21]) );
  DFC1 u_decode_pipe_Fbmemout_reg_22_ ( .D(u_decode_fbmemmux_o_data_fmem[22]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[22]) );
  DFC1 u_decode_pipe_Fbmemout_reg_23_ ( .D(u_decode_fbmemmux_o_data_fmem[23]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[23]) );
  DFC1 u_decode_pipe_Fbmemout_reg_24_ ( .D(u_decode_fbmemmux_o_data_fmem[24]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[24]) );
  DFC1 u_decode_pipe_Fbmemout_reg_25_ ( .D(u_decode_fbmemmux_o_data_fmem[25]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[25]) );
  DFC1 u_decode_pipe_Fbmemout_reg_26_ ( .D(u_decode_fbmemmux_o_data_fmem[26]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[26]) );
  DFC1 u_decode_pipe_Fbmemout_reg_27_ ( .D(u_decode_fbmemmux_o_data_fmem[27]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[27]) );
  DFC1 u_decode_pipe_Fbmemout_reg_28_ ( .D(u_decode_fbmemmux_o_data_fmem[28]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[28]) );
  DFC1 u_decode_pipe_Fbmemout_reg_29_ ( .D(u_decode_fbmemmux_o_data_fmem[29]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[29]) );
  DFC1 u_decode_pipe_Fbmemout_reg_30_ ( .D(u_decode_fbmemmux_o_data_fmem[30]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[30]) );
  DFC1 u_decode_pipe_Fbmemout_reg_31_ ( .D(u_decode_fbmemmux_o_data_fmem[31]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[31]) );
  DFC1 u_decode_pipe_Famemout_reg_0_ ( .D(u_decode_famemmux_o_data_fmem[0]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[0]) );
  DFC1 u_decode_pipe_Famemout_reg_1_ ( .D(u_decode_famemmux_o_data_fmem[1]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[1]) );
  DFC1 u_decode_pipe_Famemout_reg_2_ ( .D(u_decode_famemmux_o_data_fmem[2]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[2]) );
  DFC1 u_decode_pipe_Famemout_reg_3_ ( .D(u_decode_famemmux_o_data_fmem[3]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[3]) );
  DFC1 u_decode_pipe_Famemout_reg_4_ ( .D(u_decode_famemmux_o_data_fmem[4]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[4]) );
  DFC1 u_decode_pipe_Famemout_reg_5_ ( .D(u_decode_famemmux_o_data_fmem[5]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[5]) );
  DFC1 u_decode_pipe_Famemout_reg_6_ ( .D(u_decode_famemmux_o_data_fmem[6]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[6]) );
  DFC1 u_decode_pipe_Famemout_reg_7_ ( .D(u_decode_famemmux_o_data_fmem[7]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[7]) );
  DFC1 u_decode_pipe_Famemout_reg_8_ ( .D(u_decode_famemmux_o_data_fmem[8]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[8]) );
  DFC1 u_decode_pipe_Famemout_reg_9_ ( .D(u_decode_famemmux_o_data_fmem[9]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[9]) );
  DFC1 u_decode_pipe_Famemout_reg_10_ ( .D(u_decode_famemmux_o_data_fmem[10]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[10]) );
  DFC1 u_decode_pipe_Famemout_reg_11_ ( .D(u_decode_famemmux_o_data_fmem[11]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[11]) );
  DFC1 u_decode_pipe_Famemout_reg_12_ ( .D(u_decode_famemmux_o_data_fmem[12]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[12]) );
  DFC1 u_decode_pipe_Famemout_reg_13_ ( .D(u_decode_famemmux_o_data_fmem[13]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[13]) );
  DFC1 u_decode_pipe_Famemout_reg_14_ ( .D(u_decode_famemmux_o_data_fmem[14]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[14]) );
  DFC1 u_decode_pipe_Famemout_reg_15_ ( .D(u_decode_famemmux_o_data_fmem[15]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[15]) );
  DFC1 u_decode_pipe_Famemout_reg_16_ ( .D(u_decode_famemmux_o_data_fmem[16]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[16]) );
  DFC1 u_decode_pipe_Famemout_reg_17_ ( .D(u_decode_famemmux_o_data_fmem[17]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[17]) );
  DFC1 u_decode_pipe_Famemout_reg_18_ ( .D(u_decode_famemmux_o_data_fmem[18]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[18]) );
  DFC1 u_decode_pipe_Famemout_reg_19_ ( .D(u_decode_famemmux_o_data_fmem[19]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[19]) );
  DFC1 u_decode_pipe_Famemout_reg_20_ ( .D(u_decode_famemmux_o_data_fmem[20]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[20]) );
  DFC1 u_decode_pipe_Famemout_reg_21_ ( .D(u_decode_famemmux_o_data_fmem[21]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[21]) );
  DFC1 u_decode_pipe_Famemout_reg_22_ ( .D(u_decode_famemmux_o_data_fmem[22]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[22]) );
  DFC1 u_decode_pipe_Famemout_reg_23_ ( .D(u_decode_famemmux_o_data_fmem[23]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[23]) );
  DFC1 u_decode_pipe_Famemout_reg_24_ ( .D(u_decode_famemmux_o_data_fmem[24]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[24]) );
  DFC1 u_decode_pipe_Famemout_reg_25_ ( .D(u_decode_famemmux_o_data_fmem[25]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[25]) );
  DFC1 u_decode_pipe_Famemout_reg_26_ ( .D(u_decode_famemmux_o_data_fmem[26]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[26]) );
  DFC1 u_decode_pipe_Famemout_reg_27_ ( .D(u_decode_famemmux_o_data_fmem[27]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[27]) );
  DFC1 u_decode_pipe_Famemout_reg_28_ ( .D(u_decode_famemmux_o_data_fmem[28]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[28]) );
  DFC1 u_decode_pipe_Famemout_reg_29_ ( .D(u_decode_famemmux_o_data_fmem[29]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[29]) );
  DFC1 u_decode_pipe_Famemout_reg_30_ ( .D(u_decode_famemmux_o_data_fmem[30]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[30]) );
  DFC1 u_decode_pipe_Famemout_reg_31_ ( .D(u_decode_famemmux_o_data_fmem[31]), 
        .C(clk), .RN(rst_n), .Q(for_famemout[31]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_4_ ( .D(if_addr_j[6]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[4]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_11_ ( .D(if_addr_j[13]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[0]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_12_ ( .D(if_addr_j[14]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[1]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_13_ ( .D(if_addr_j[15]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[2]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_14_ ( .D(if_addr_j[16]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[3]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_15_ ( .D(if_addr_j[17]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[4]) );
  DFC1 u_decode_pipe_con_Wmemtoreg_reg ( .D(u_decode_control_o_con_memtoreg), 
        .C(clk), .RN(rst_n), .Q(ex_con_Wmemtoreg) );
  DFC1 u_decode_pipe_con_Mmemwrite_reg ( .D(u_decode_n4), .C(clk), .RN(rst_n), 
        .Q(ex_con_Mmemwrite) );
  DFC1 u_decode_pipe_con_Mmemread_reg ( .D(u_decode_control_o_con_memread), 
        .C(clk), .RN(rst_n), .Q(ex_con_Mmemread) );
  DFC1 u_decode_pipe_con_MaluPC4_reg ( .D(u_decode_jbcon_o_con_aluPC4), .C(clk), .RN(rst_n), .Q(ex_con_Malupc8) );
  DFC1 u_decode_pipe_con_Ealuop_reg_5_ ( .D(u_decode_control_o_con_aluop_5_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[5]) );
  DFC1 u_decode_pipe_addr_pc4_reg_2_ ( .D(id_addr_pc4[2]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[2]) );
  DFC1 u_decode_pipe_addr_pc4_reg_3_ ( .D(id_addr_pc4[3]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[3]) );
  DFC1 u_decode_pipe_addr_pc4_reg_4_ ( .D(id_addr_pc4[4]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[4]) );
  DFC1 u_decode_pipe_addr_pc4_reg_5_ ( .D(id_addr_pc4[5]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[5]) );
  DFC1 u_decode_pipe_addr_pc4_reg_6_ ( .D(id_addr_pc4[6]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[6]) );
  DFC1 u_decode_pipe_addr_pc4_reg_7_ ( .D(id_addr_pc4[7]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[7]) );
  DFC1 u_decode_pipe_addr_pc4_reg_8_ ( .D(id_addr_pc4[8]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[8]) );
  DFC1 u_decode_pipe_addr_pc4_reg_9_ ( .D(id_addr_pc4[9]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[9]) );
  DFC1 u_decode_pipe_addr_pc4_reg_10_ ( .D(id_addr_pc4[10]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[10]) );
  DFC1 u_decode_pipe_addr_pc4_reg_11_ ( .D(id_addr_pc4[11]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[11]) );
  DFC1 u_decode_pipe_addr_pc4_reg_12_ ( .D(id_addr_pc4[12]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[12]) );
  DFC1 u_decode_pipe_addr_pc4_reg_13_ ( .D(id_addr_pc4[13]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[13]) );
  DFC1 u_decode_pipe_addr_pc4_reg_14_ ( .D(id_addr_pc4[14]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[14]) );
  DFC1 u_decode_pipe_addr_pc4_reg_15_ ( .D(id_addr_pc4[15]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[15]) );
  DFC1 u_decode_pipe_addr_pc4_reg_16_ ( .D(id_addr_pc4[16]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[16]) );
  DFC1 u_decode_pipe_addr_pc4_reg_17_ ( .D(id_addr_pc4[17]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[17]) );
  DFC1 u_decode_pipe_addr_pc4_reg_18_ ( .D(id_addr_pc4[18]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[18]) );
  DFC1 u_decode_pipe_addr_pc4_reg_19_ ( .D(id_addr_pc4[19]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[19]) );
  DFC1 u_decode_pipe_addr_pc4_reg_20_ ( .D(id_addr_pc4[20]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[20]) );
  DFC1 u_decode_pipe_addr_pc4_reg_21_ ( .D(id_addr_pc4[21]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[21]) );
  DFC1 u_decode_pipe_addr_pc4_reg_22_ ( .D(id_addr_pc4[22]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[22]) );
  DFC1 u_decode_pipe_addr_pc4_reg_23_ ( .D(id_addr_pc4[23]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[23]) );
  DFC1 u_decode_pipe_addr_pc4_reg_24_ ( .D(id_addr_pc4[24]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[24]) );
  DFC1 u_decode_pipe_addr_pc4_reg_25_ ( .D(id_addr_pc4[25]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[25]) );
  DFC1 u_decode_pipe_addr_pc4_reg_26_ ( .D(id_addr_pc4[26]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[26]) );
  DFC1 u_decode_pipe_addr_pc4_reg_27_ ( .D(id_addr_pc4[27]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[27]) );
  DFC1 u_decode_pipe_addr_pc4_reg_28_ ( .D(if_addr_j[28]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[28]) );
  DFC1 u_decode_pipe_addr_pc4_reg_29_ ( .D(if_addr_j[29]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[29]) );
  DFC1 u_decode_pipe_addr_pc4_reg_30_ ( .D(if_addr_j[30]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[30]) );
  DFC1 u_decode_pipe_addr_pc4_reg_31_ ( .D(if_addr_j[31]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[31]) );
  DFC1 u_decode_pipe_addr_rt_reg_0_ ( .D(n323), .C(clk), .RN(rst_n), .Q(
        ex_addr_rt[0]) );
  DFC1 u_decode_pipe_addr_rt_reg_1_ ( .D(n238), .C(clk), .RN(rst_n), .Q(
        ex_addr_rt[1]) );
  DFC1 u_decode_pipe_addr_rt_reg_2_ ( .D(n237), .C(clk), .RN(rst_n), .Q(
        ex_addr_rt[2]) );
  DFC1 u_decode_pipe_addr_rt_reg_3_ ( .D(if_addr_j[21]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[3]) );
  DFC1 u_decode_pipe_addr_rt_reg_4_ ( .D(if_addr_j[22]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[4]) );
  DFC1 u_decode_pipe_data_rt_reg_0_ ( .D(u_decode_regbank_o_data_Rt[0]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[0]) );
  DFC1 u_decode_pipe_data_rt_reg_1_ ( .D(u_decode_regbank_o_data_Rt[1]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[1]) );
  DFC1 u_decode_pipe_data_rt_reg_2_ ( .D(u_decode_regbank_o_data_Rt[2]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[2]) );
  DFC1 u_decode_pipe_data_rt_reg_3_ ( .D(u_decode_regbank_o_data_Rt[3]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[3]) );
  DFC1 u_decode_pipe_data_rt_reg_4_ ( .D(u_decode_regbank_o_data_Rt[4]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[4]) );
  DFC1 u_decode_pipe_data_rt_reg_5_ ( .D(u_decode_regbank_o_data_Rt[5]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[5]) );
  DFC1 u_decode_pipe_data_rt_reg_6_ ( .D(u_decode_regbank_o_data_Rt[6]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[6]) );
  DFC1 u_decode_pipe_data_rt_reg_7_ ( .D(u_decode_regbank_o_data_Rt[7]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[7]) );
  DFC1 u_decode_pipe_data_rt_reg_8_ ( .D(u_decode_regbank_o_data_Rt[8]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[8]) );
  DFC1 u_decode_pipe_data_rt_reg_9_ ( .D(u_decode_regbank_o_data_Rt[9]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[9]) );
  DFC1 u_decode_pipe_data_rt_reg_10_ ( .D(u_decode_regbank_o_data_Rt[10]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[10]) );
  DFC1 u_decode_pipe_data_rt_reg_11_ ( .D(u_decode_regbank_o_data_Rt[11]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[11]) );
  DFC1 u_decode_pipe_data_rt_reg_12_ ( .D(u_decode_regbank_o_data_Rt[12]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[12]) );
  DFC1 u_decode_pipe_data_rt_reg_13_ ( .D(u_decode_regbank_o_data_Rt[13]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[13]) );
  DFC1 u_decode_pipe_data_rt_reg_14_ ( .D(u_decode_regbank_o_data_Rt[14]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[14]) );
  DFC1 u_decode_pipe_data_rt_reg_15_ ( .D(u_decode_regbank_o_data_Rt[15]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[15]) );
  DFC1 u_decode_pipe_data_rt_reg_16_ ( .D(u_decode_regbank_o_data_Rt[16]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[16]) );
  DFC1 u_decode_pipe_data_rt_reg_17_ ( .D(u_decode_regbank_o_data_Rt[17]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[17]) );
  DFC1 u_decode_pipe_data_rt_reg_18_ ( .D(u_decode_regbank_o_data_Rt[18]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[18]) );
  DFC1 u_decode_pipe_data_rt_reg_19_ ( .D(u_decode_regbank_o_data_Rt[19]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[19]) );
  DFC1 u_decode_pipe_data_rt_reg_20_ ( .D(u_decode_regbank_o_data_Rt[20]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[20]) );
  DFC1 u_decode_pipe_data_rt_reg_21_ ( .D(u_decode_regbank_o_data_Rt[21]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[21]) );
  DFC1 u_decode_pipe_data_rt_reg_22_ ( .D(u_decode_regbank_o_data_Rt[22]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[22]) );
  DFC1 u_decode_pipe_data_rt_reg_23_ ( .D(u_decode_regbank_o_data_Rt[23]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[23]) );
  DFC1 u_decode_pipe_data_rt_reg_24_ ( .D(u_decode_regbank_o_data_Rt[24]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[24]) );
  DFC1 u_decode_pipe_data_rt_reg_25_ ( .D(u_decode_regbank_o_data_Rt[25]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[25]) );
  DFC1 u_decode_pipe_data_rt_reg_26_ ( .D(u_decode_regbank_o_data_Rt[26]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[26]) );
  DFC1 u_decode_pipe_data_rt_reg_27_ ( .D(u_decode_regbank_o_data_Rt[27]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[27]) );
  DFC1 u_decode_pipe_data_rt_reg_28_ ( .D(u_decode_regbank_o_data_Rt[28]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[28]) );
  DFC1 u_decode_pipe_data_rt_reg_29_ ( .D(u_decode_regbank_o_data_Rt[29]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[29]) );
  DFC1 u_decode_pipe_data_rt_reg_30_ ( .D(u_decode_regbank_o_data_Rt[30]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[30]) );
  DFC1 u_decode_pipe_data_rt_reg_31_ ( .D(u_decode_regbank_o_data_Rt[31]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[31]) );
  DFC1 u_decode_pipe_data_rs_reg_0_ ( .D(id_data_jr[0]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[0]) );
  DFC1 u_decode_pipe_data_rs_reg_1_ ( .D(id_data_jr[1]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[1]) );
  DFC1 u_decode_pipe_data_rs_reg_2_ ( .D(id_data_jr[2]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[2]) );
  DFC1 u_decode_pipe_data_rs_reg_3_ ( .D(id_data_jr[3]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[3]) );
  DFC1 u_decode_pipe_data_rs_reg_4_ ( .D(id_data_jr[4]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[4]) );
  DFC1 u_decode_pipe_data_rs_reg_5_ ( .D(id_data_jr[5]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[5]) );
  DFC1 u_decode_pipe_data_rs_reg_6_ ( .D(id_data_jr[6]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[6]) );
  DFC1 u_decode_pipe_data_rs_reg_7_ ( .D(id_data_jr[7]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[7]) );
  DFC1 u_decode_pipe_data_rs_reg_8_ ( .D(id_data_jr[8]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[8]) );
  DFC1 u_decode_pipe_data_rs_reg_9_ ( .D(id_data_jr[9]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[9]) );
  DFC1 u_decode_pipe_data_rs_reg_10_ ( .D(id_data_jr[10]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[10]) );
  DFC1 u_decode_pipe_data_rs_reg_11_ ( .D(id_data_jr[11]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[11]) );
  DFC1 u_decode_pipe_data_rs_reg_12_ ( .D(id_data_jr[12]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[12]) );
  DFC1 u_decode_pipe_data_rs_reg_13_ ( .D(id_data_jr[13]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[13]) );
  DFC1 u_decode_pipe_data_rs_reg_14_ ( .D(id_data_jr[14]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[14]) );
  DFC1 u_decode_pipe_data_rs_reg_16_ ( .D(id_data_jr[16]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[16]) );
  DFC1 u_decode_pipe_data_rs_reg_17_ ( .D(id_data_jr[17]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[17]) );
  DFC1 u_decode_pipe_data_rs_reg_18_ ( .D(id_data_jr[18]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[18]) );
  DFC1 u_decode_pipe_data_rs_reg_19_ ( .D(id_data_jr[19]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[19]) );
  DFC1 u_decode_pipe_data_rs_reg_20_ ( .D(id_data_jr[20]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[20]) );
  DFC1 u_decode_pipe_data_rs_reg_21_ ( .D(id_data_jr[21]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[21]) );
  DFC1 u_decode_pipe_data_rs_reg_22_ ( .D(id_data_jr[22]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[22]) );
  DFC1 u_decode_pipe_data_rs_reg_23_ ( .D(id_data_jr[23]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[23]) );
  DFC1 u_decode_pipe_data_rs_reg_24_ ( .D(id_data_jr[24]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[24]) );
  DFC1 u_decode_pipe_data_rs_reg_25_ ( .D(id_data_jr[25]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[25]) );
  DFC1 u_decode_pipe_data_rs_reg_26_ ( .D(id_data_jr[26]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[26]) );
  DFC1 u_decode_pipe_data_rs_reg_27_ ( .D(id_data_jr[27]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[27]) );
  DFC1 u_decode_pipe_data_rs_reg_28_ ( .D(id_data_jr[28]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[28]) );
  DFC1 u_decode_pipe_data_rs_reg_29_ ( .D(id_data_jr[29]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[29]) );
  DFC1 u_decode_pipe_data_rs_reg_30_ ( .D(id_data_jr[30]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[30]) );
  DFC1 u_decode_pipe_data_rs_reg_31_ ( .D(id_data_jr[31]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[31]) );
  DFC1 u_decode_pipe_bop_reg_0_ ( .D(u_decode_jbcon_o_con_bop[0]), .C(clk), 
        .RN(rst_n), .Q(ex_con_bop[0]) );
  DFC1 u_decode_pipe_bop_reg_1_ ( .D(u_decode_jbcon_o_con_bop[1]), .C(clk), 
        .RN(rst_n), .Q(ex_con_bop[1]) );
  DFC1 u_decode_pipe_bop_reg_2_ ( .D(u_decode_jbcon_o_con_bop[2]), .C(clk), 
        .RN(rst_n), .Q(ex_con_bop[2]) );
  D_register_bank u_decode_u_regbank ( .i_clk(clk), .i_rst_n(rst_n), 
        .i_addr_Rs(if_addr_j[27:23]), .i_addr_Rt({if_addr_j[22:19], n323}), 
        .i_con_RegWr(id_con_Wregwrite), .i_addr_Rd(id_addr_Wregwrite), 
        .i_data_Rd(id_data_Wregwrite), .o_data_Rs(id_data_jr), .o_data_Rt(
        u_decode_regbank_o_data_Rt) );
  OAI212 u_decode_add_x_16_U185 ( .A(u_decode_add_x_16_n149), .B(
        u_decode_add_x_16_n169), .C(u_decode_add_x_16_n150), .Q(
        u_decode_add_x_16_n148) );
  DFC3 u_fetch_pipe_instr_reg_16_ ( .D(read_instruction[16]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[18]) );
  DFC3 u_fetch_pipe_instr_reg_17_ ( .D(read_instruction[17]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[19]), .QN(n282) );
  DFC3 u_fetch_pipe_instr_reg_19_ ( .D(read_instruction[19]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[21]), .QN(n281) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_16_ ( .D(u_decode_n3), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[31]) );
  DFC3 u_fetch_pipe_instr_reg_23_ ( .D(read_instruction[23]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[25]), .QN(n277) );
  DFC3 u_decode_pipe_con_Ealusrc_reg ( .D(u_decode_n6), .C(clk), .RN(rst_n), 
        .Q(ex_con_Ealusrc) );
  DFC3 u_fetch_pipe_instr_reg_24_ ( .D(read_instruction[24]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[26]), .QN(n280) );
  DFC3 u_fetch_pipe_instr_reg_22_ ( .D(read_instruction[22]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[24]), .QN(n260) );
  DFC3 u_fetch_pipe_instr_reg_21_ ( .D(read_instruction[21]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[23]), .QN(n261) );
  DFC3 u_decode_pipe_con_Efamux_reg_1_ ( .D(u_decode_n17), .C(clk), .RN(rst_n), 
        .Q(for_o_con_Efamux[1]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_2_ ( .D(if_addr_j[4]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[2]) );
  DFC3 u_fetch_pipe_instr_reg_18_ ( .D(read_instruction[18]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[20]), .QN(n278) );
  DFC3 u_decode_pipe_con_Efbmux_reg_1_ ( .D(u_decode_n23), .C(clk), .RN(rst_n), 
        .Q(for_o_con_Efbmux[1]) );
  DFC3 u_decode_pipe_con_Efbmux_reg_0_ ( .D(u_decode_for_o_con_fb_0_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[0]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_3_ ( .D(if_addr_j[5]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[3]) );
  DFC3 u_fetch_pipe_instr_reg_29_ ( .D(read_instruction[29]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[29]), .QN(n312) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_5_ ( .D(if_addr_j[7]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[5]) );
  DFC3 u_decode_pipe_con_Efamux_reg_0_ ( .D(u_decode_for_o_con_fa_0_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[0]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_0_ ( .D(if_addr_j[2]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[0]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_1_ ( .D(if_addr_j[3]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[1]) );
  DFC3 u_decode_pipe_con_Eregdst_reg ( .D(u_decode_control_o_con_regdst), .C(
        clk), .RN(rst_n), .Q(ex_con_Eregdst) );
  DFC3 u_decode_pipe_con_Ealuop_reg_3_ ( .D(u_decode_control_o_con_aluop_3_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[3]) );
  DFC3 u_decode_pipe_con_Ealuop_reg_1_ ( .D(u_decode_control_o_con_aluop_1_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[1]) );
  DFC3 u_fetch_pipe_instr_reg_25_ ( .D(read_instruction[25]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[27]), .QN(n279) );
  DFC3 u_mem_pipe_addr_regdst_reg_3_ ( .D(mem_addr_regdst[3]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[3]) );
  DFC3 u_decode_pipe_con_Ealuop_reg_0_ ( .D(u_decode_control_o_con_aluop_0_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[0]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_7_ ( .D(if_addr_j[9]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[7]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_10_ ( .D(if_addr_j[12]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[10]) );
  DFC3 u_fetch_pipe_instr_reg_20_ ( .D(read_instruction[20]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[22]), .QN(n311) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_6_ ( .D(if_addr_j[8]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[6]) );
  DFC3 u_mem_pipe_con_Wmemtoreg_reg ( .D(mem_con_Wmemtoreg), .C(clk), .RN(
        rst_n), .Q(wb_con_Wmemtoreg) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_9_ ( .D(if_addr_j[11]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[9]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_8_ ( .D(if_addr_j[10]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[8]) );
  XNR21 add_x_4_U139 ( .A(instruction_address[2]), .B(n296), .Q(
        u_fetch_jmux_i_addr_pc4_3_) );
  OAI210 u_decode_add_x_16_U57 ( .A(u_decode_add_x_16_n73), .B(
        u_decode_add_x_16_n69), .C(u_decode_add_x_16_n70), .Q(
        u_decode_add_x_16_n68) );
  XNR21 u_decode_add_x_16_U134 ( .A(u_decode_add_x_16_n17), .B(
        u_decode_add_x_16_n121), .Q(u_decode_pcadd_o_addr_pcbranchE[15]) );
  XNR21 u_decode_add_x_16_U12 ( .A(u_decode_add_x_16_n3), .B(
        u_decode_add_x_16_n41), .Q(u_decode_pcadd_o_addr_pcbranchE[29]) );
  XNR21 u_decode_add_x_16_U159 ( .A(u_decode_add_x_16_n20), .B(
        u_decode_add_x_16_n137), .Q(u_decode_pcadd_o_addr_pcbranchE[12]) );
  XNR21 u_decode_add_x_16_U167 ( .A(u_decode_add_x_16_n21), .B(
        u_decode_add_x_16_n144), .Q(u_decode_pcadd_o_addr_pcbranchE[11]) );
  XNR21 add_x_1_U1 ( .A(mem_data_pc4[31]), .B(add_x_1_n2), .Q(u_mem_pc8[31])
         );
  XNR21 add_x_1_U87 ( .A(add_x_1_n73), .B(add_x_1_n74), .Q(u_mem_pc8[14]) );
  XNR21 u_decode_add_x_16_U183 ( .A(u_decode_add_x_16_n23), .B(
        u_decode_add_x_16_n155), .Q(u_decode_pcadd_o_addr_pcbranchE[9]) );
  NAND22 add_x_4_U141 ( .A(instruction_address[3]), .B(instruction_address[2]), 
        .Q(add_x_4_n111) );
  NAND22 add_x_4_U74 ( .A(add_x_4_n60), .B(instruction_address[16]), .Q(
        add_x_4_n57) );
  NAND22 add_x_4_U32 ( .A(add_x_4_n26), .B(instruction_address[24]), .Q(
        add_x_4_n23) );
  NAND22 add_x_4_U4 ( .A(add_x_4_n4), .B(instruction_address[30]), .Q(
        add_x_4_n1) );
  NAND22 add_x_4_U17 ( .A(add_x_4_n17), .B(add_x_4_n12), .Q(add_x_4_n11) );
  NAND22 add_x_4_U52 ( .A(add_x_4_n42), .B(instruction_address[20]), .Q(
        add_x_4_n39) );
  NAND22 u_decode_add_x_16_U2 ( .A(u_decode_add_x_16_n183), .B(
        u_decode_add_x_16_n32), .Q(u_decode_add_x_16_n1) );
  NOR21 u_decode_add_x_16_U38 ( .A(id_addr_pc4[27]), .B(n324), .Q(
        u_decode_add_x_16_n53) );
  NAND22 u_decode_add_x_16_U32 ( .A(u_decode_add_x_16_n58), .B(
        u_decode_add_x_16_n51), .Q(u_decode_add_x_16_n49) );
  NAND22 u_decode_add_x_16_U22 ( .A(u_decode_add_x_16_n63), .B(
        u_decode_add_x_16_n44), .Q(u_decode_add_x_16_n42) );
  NAND22 u_decode_add_x_16_U186 ( .A(u_decode_add_x_16_n159), .B(
        u_decode_add_x_16_n151), .Q(u_decode_add_x_16_n149) );
  OAI212 u_decode_add_x_16_U233 ( .A(u_decode_add_x_16_n182), .B(
        u_decode_add_x_16_n179), .C(u_decode_add_x_16_n180), .Q(
        u_decode_add_x_16_n178) );
  OAI212 u_decode_add_x_16_U203 ( .A(u_decode_add_x_16_n167), .B(
        u_decode_add_x_16_n161), .C(u_decode_add_x_16_n162), .Q(
        u_decode_add_x_16_n160) );
  OAI212 u_decode_add_x_16_U172 ( .A(u_decode_add_x_16_n146), .B(
        u_decode_add_x_16_n142), .C(u_decode_add_x_16_n143), .Q(
        u_decode_add_x_16_n141) );
  OAI212 u_decode_add_x_16_U137 ( .A(u_decode_add_x_16_n123), .B(
        u_decode_add_x_16_n119), .C(u_decode_add_x_16_n120), .Q(
        u_decode_add_x_16_n118) );
  AOI211 u_decode_add_x_16_U121 ( .A(u_decode_add_x_16_n109), .B(
        u_decode_add_x_16_n118), .C(u_decode_add_x_16_n110), .Q(
        u_decode_add_x_16_n108) );
  OAI212 u_decode_add_x_16_U119 ( .A(u_decode_add_x_16_n127), .B(
        u_decode_add_x_16_n107), .C(u_decode_add_x_16_n108), .Q(
        u_decode_add_x_16_n106) );
  AOI212 u_decode_add_x_16_U117 ( .A(u_decode_add_x_16_n148), .B(
        u_decode_add_x_16_n105), .C(u_decode_add_x_16_n106), .Q(
        u_decode_add_x_16_n104) );
  OAI212 u_decode_add_x_16_U102 ( .A(u_decode_add_x_16_n102), .B(
        u_decode_add_x_16_n96), .C(u_decode_add_x_16_n97), .Q(
        u_decode_add_x_16_n95) );
  OAI212 u_decode_add_x_16_U71 ( .A(u_decode_add_x_16_n81), .B(
        u_decode_add_x_16_n77), .C(u_decode_add_x_16_n78), .Q(
        u_decode_add_x_16_n76) );
  AOI211 u_decode_add_x_16_U55 ( .A(u_decode_add_x_16_n76), .B(
        u_decode_add_x_16_n67), .C(u_decode_add_x_16_n68), .Q(
        u_decode_add_x_16_n66) );
  OAI212 u_decode_add_x_16_U53 ( .A(u_decode_add_x_16_n65), .B(
        u_decode_add_x_16_n85), .C(u_decode_add_x_16_n66), .Q(
        u_decode_add_x_16_n64) );
  OAI212 u_decode_add_x_16_U21 ( .A(u_decode_add_x_16_n42), .B(
        u_decode_add_x_16_n104), .C(u_decode_add_x_16_n43), .Q(
        u_decode_add_x_16_n41) );
  OAI212 u_decode_add_x_16_U7 ( .A(u_decode_add_x_16_n34), .B(
        u_decode_add_x_16_n36), .C(u_decode_add_x_16_n35), .Q(
        u_decode_add_x_16_n33) );
  OAI212 u_decode_add_x_16_U41 ( .A(u_decode_add_x_16_n56), .B(
        u_decode_add_x_16_n62), .C(u_decode_add_x_16_n57), .Q(
        u_decode_add_x_16_n55) );
  NAND22 u_decode_add_x_16_U26 ( .A(u_decode_add_x_16_n186), .B(
        u_decode_add_x_16_n47), .Q(u_decode_add_x_16_n4) );
  OAI212 u_decode_add_x_16_U31 ( .A(u_decode_add_x_16_n49), .B(
        u_decode_add_x_16_n62), .C(u_decode_add_x_16_n50), .Q(
        u_decode_add_x_16_n48) );
  OAI212 u_decode_add_x_16_U150 ( .A(u_decode_add_x_16_n126), .B(
        u_decode_add_x_16_n147), .C(u_decode_add_x_16_n127), .Q(
        u_decode_add_x_16_n125) );
  OAI212 u_decode_add_x_16_U129 ( .A(u_decode_add_x_16_n114), .B(
        u_decode_add_x_16_n116), .C(u_decode_add_x_16_n115), .Q(
        u_decode_add_x_16_n113) );
  OAI212 u_decode_add_x_16_U143 ( .A(u_decode_add_x_16_n122), .B(
        u_decode_add_x_16_n124), .C(u_decode_add_x_16_n123), .Q(
        u_decode_add_x_16_n121) );
  OAI212 u_decode_add_x_16_U94 ( .A(u_decode_add_x_16_n91), .B(
        u_decode_add_x_16_n93), .C(u_decode_add_x_16_n92), .Q(
        u_decode_add_x_16_n90) );
  OAI212 u_decode_add_x_16_U84 ( .A(u_decode_add_x_16_n84), .B(
        u_decode_add_x_16_n104), .C(u_decode_add_x_16_n85), .Q(
        u_decode_add_x_16_n83) );
  OAI212 u_decode_add_x_16_U63 ( .A(u_decode_add_x_16_n72), .B(
        u_decode_add_x_16_n74), .C(u_decode_add_x_16_n73), .Q(
        u_decode_add_x_16_n71) );
  OAI212 u_decode_add_x_16_U77 ( .A(u_decode_add_x_16_n80), .B(
        u_decode_add_x_16_n82), .C(u_decode_add_x_16_n81), .Q(
        u_decode_add_x_16_n79) );
  XOR21 u_decode_add_x_16_U40 ( .A(u_decode_add_x_16_n6), .B(
        u_decode_add_x_16_n62), .Q(u_decode_pcadd_o_addr_pcbranchE[26]) );
  OAI212 u_decode_add_x_16_U168 ( .A(u_decode_add_x_16_n138), .B(
        u_decode_add_x_16_n147), .C(u_decode_add_x_16_n139), .Q(
        u_decode_add_x_16_n137) );
  NAND22 u_decode_add_x_16_U16 ( .A(u_decode_add_x_16_n37), .B(
        u_decode_add_x_16_n40), .Q(u_decode_add_x_16_n3) );
  NAND22 add_x_1_U118 ( .A(mem_data_pc4[8]), .B(mem_data_pc4[9]), .Q(
        add_x_1_n95) );
  NAND22 add_x_1_U127 ( .A(mem_data_pc4[6]), .B(mem_data_pc4[7]), .Q(
        add_x_1_n102) );
  NAND22 add_x_1_U147 ( .A(mem_data_pc4[2]), .B(mem_data_pc4[3]), .Q(
        add_x_1_n118) );
  NAND22 add_x_1_U138 ( .A(mem_data_pc4[4]), .B(mem_data_pc4[5]), .Q(
        add_x_1_n111) );
  NAND22 add_x_1_U107 ( .A(mem_data_pc4[10]), .B(mem_data_pc4[11]), .Q(
        add_x_1_n86) );
  NAND22 add_x_1_U84 ( .A(mem_data_pc4[14]), .B(mem_data_pc4[15]), .Q(
        add_x_1_n67) );
  XOR21 add_x_1_U41 ( .A(add_x_1_n35), .B(add_x_1_n36), .Q(u_mem_pc8[22]) );
  NAND22 add_x_1_U38 ( .A(mem_data_pc4[22]), .B(mem_data_pc4[23]), .Q(
        add_x_1_n29) );
  NAND22 add_x_1_U36 ( .A(add_x_1_n37), .B(add_x_1_n28), .Q(add_x_1_n27) );
  XOR21 add_x_1_U30 ( .A(add_x_1_n26), .B(add_x_1_n27), .Q(u_mem_pc8[24]) );
  NOR21 add_x_1_U15 ( .A(add_x_1_n11), .B(add_x_1_n18), .Q(add_x_1_n10) );
  NAND22 add_x_1_U14 ( .A(add_x_1_n10), .B(add_x_1_n55), .Q(add_x_1_n9) );
  XOR21 add_x_1_U3 ( .A(mem_data_pc4[30]), .B(add_x_1_n4), .Q(u_mem_pc8[30])
         );
  XOR21 add_x_1_U130 ( .A(add_x_1_n108), .B(add_x_1_n109), .Q(u_mem_pc8[6]) );
  XOR21 add_x_1_U76 ( .A(add_x_1_n64), .B(add_x_1_n65), .Q(u_mem_pc8[16]) );
  NAND22 add_x_1_U105 ( .A(add_x_1_n92), .B(add_x_1_n85), .Q(add_x_1_n84) );
  XOR21 add_x_1_U99 ( .A(add_x_1_n83), .B(add_x_1_n84), .Q(u_mem_pc8[12]) );
  OAI212 u_decode_add_x_16_U220 ( .A(u_decode_add_x_16_n176), .B(
        u_decode_add_x_16_n172), .C(u_decode_add_x_16_n173), .Q(
        u_decode_add_x_16_n171) );
  NAND22 u_decode_add_x_16_U127 ( .A(n324), .B(id_addr_pc4[17]), .Q(
        u_decode_add_x_16_n112) );
  NAND22 u_decode_add_x_16_U242 ( .A(if_addr_j[2]), .B(id_addr_pc4[2]), .Q(
        u_decode_add_x_16_n182) );
  NAND22 u_decode_add_x_16_U182 ( .A(if_addr_j[10]), .B(id_addr_pc4[10]), .Q(
        u_decode_add_x_16_n146) );
  NAND22 u_decode_add_x_16_U98 ( .A(n324), .B(id_addr_pc4[20]), .Q(
        u_decode_add_x_16_n92) );
  NAND22 u_decode_add_x_16_U49 ( .A(if_addr_j[17]), .B(id_addr_pc4[26]), .Q(
        u_decode_add_x_16_n57) );
  NAND22 add_x_4_U112 ( .A(instruction_address[8]), .B(instruction_address[9]), 
        .Q(add_x_4_n88) );
  NAND22 add_x_4_U121 ( .A(instruction_address[6]), .B(instruction_address[7]), 
        .Q(add_x_4_n95) );
  NAND22 add_x_4_U90 ( .A(instruction_address[12]), .B(instruction_address[13]), .Q(add_x_4_n70) );
  NAND22 add_x_4_U105 ( .A(add_x_4_n85), .B(instruction_address[10]), .Q(
        add_x_4_n82) );
  NAND22 add_x_4_U70 ( .A(instruction_address[16]), .B(instruction_address[17]), .Q(add_x_4_n54) );
  NAND22 add_x_4_U116 ( .A(add_x_4_n94), .B(instruction_address[8]), .Q(
        add_x_4_n91) );
  NAND22 add_x_4_U83 ( .A(add_x_4_n67), .B(instruction_address[14]), .Q(
        add_x_4_n64) );
  NAND22 add_x_4_U57 ( .A(instruction_address[18]), .B(instruction_address[19]), .Q(add_x_4_n43) );
  NOR21 add_x_4_U18 ( .A(n276), .B(n252), .Q(add_x_4_n12) );
  NAND22 add_x_4_U13 ( .A(add_x_4_n12), .B(instruction_address[28]), .Q(
        add_x_4_n8) );
  NAND22 add_x_4_U48 ( .A(instruction_address[20]), .B(instruction_address[21]), .Q(add_x_4_n36) );
  NAND22 add_x_4_U37 ( .A(instruction_address[22]), .B(instruction_address[23]), .Q(add_x_4_n27) );
  NAND22 add_x_4_U41 ( .A(add_x_4_n33), .B(instruction_address[22]), .Q(
        add_x_4_n30) );
  NAND22 u_decode_add_x_16_U237 ( .A(if_addr_j[3]), .B(id_addr_pc4[3]), .Q(
        u_decode_add_x_16_n180) );
  NAND22 u_decode_add_x_16_U230 ( .A(if_addr_j[4]), .B(id_addr_pc4[4]), .Q(
        u_decode_add_x_16_n176) );
  NAND22 u_decode_add_x_16_U215 ( .A(if_addr_j[6]), .B(id_addr_pc4[6]), .Q(
        u_decode_add_x_16_n167) );
  NAND22 u_decode_add_x_16_U199 ( .A(if_addr_j[8]), .B(id_addr_pc4[8]), .Q(
        u_decode_add_x_16_n157) );
  NAND22 u_decode_add_x_16_U166 ( .A(if_addr_j[12]), .B(id_addr_pc4[12]), .Q(
        u_decode_add_x_16_n136) );
  NAND22 u_decode_add_x_16_U147 ( .A(if_addr_j[14]), .B(id_addr_pc4[14]), .Q(
        u_decode_add_x_16_n123) );
  NAND22 u_decode_add_x_16_U114 ( .A(n324), .B(id_addr_pc4[18]), .Q(
        u_decode_add_x_16_n102) );
  NAND22 u_decode_add_x_16_U106 ( .A(n324), .B(id_addr_pc4[19]), .Q(
        u_decode_add_x_16_n97) );
  NAND22 u_decode_add_x_16_U92 ( .A(n324), .B(id_addr_pc4[21]), .Q(
        u_decode_add_x_16_n89) );
  NAND22 u_decode_add_x_16_U81 ( .A(n324), .B(id_addr_pc4[22]), .Q(
        u_decode_add_x_16_n81) );
  NAND22 u_decode_add_x_16_U75 ( .A(if_addr_j[17]), .B(id_addr_pc4[23]), .Q(
        u_decode_add_x_16_n78) );
  NAND22 u_decode_add_x_16_U67 ( .A(n324), .B(id_addr_pc4[24]), .Q(
        u_decode_add_x_16_n73) );
  NAND22 u_decode_add_x_16_U39 ( .A(if_addr_j[17]), .B(id_addr_pc4[27]), .Q(
        u_decode_add_x_16_n54) );
  NOR21 u_decode_add_x_16_U18 ( .A(if_addr_j[29]), .B(n324), .Q(
        u_decode_add_x_16_n39) );
  NAND22 u_decode_add_x_16_U19 ( .A(if_addr_j[17]), .B(if_addr_j[29]), .Q(
        u_decode_add_x_16_n40) );
  NAND22 u_decode_add_x_16_U11 ( .A(n324), .B(if_addr_j[30]), .Q(
        u_decode_add_x_16_n35) );
  NAND22 u_decode_add_x_16_U36 ( .A(u_decode_add_x_16_n51), .B(
        u_decode_add_x_16_n54), .Q(u_decode_add_x_16_n5) );
  NAND22 u_decode_add_x_16_U124 ( .A(u_decode_add_x_16_n197), .B(
        u_decode_add_x_16_n112), .Q(u_decode_add_x_16_n15) );
  NAND22 u_decode_add_x_16_U138 ( .A(u_decode_add_x_16_n199), .B(
        u_decode_add_x_16_n120), .Q(u_decode_add_x_16_n17) );
  NAND22 u_decode_add_x_16_U89 ( .A(u_decode_add_x_16_n193), .B(
        u_decode_add_x_16_n89), .Q(u_decode_add_x_16_n11) );
  NAND22 u_decode_add_x_16_U58 ( .A(u_decode_add_x_16_n189), .B(
        u_decode_add_x_16_n70), .Q(u_decode_add_x_16_n7) );
  NAND22 u_decode_add_x_16_U72 ( .A(u_decode_add_x_16_n191), .B(
        u_decode_add_x_16_n78), .Q(u_decode_add_x_16_n9) );
  NAND22 u_decode_add_x_16_U46 ( .A(u_decode_add_x_16_n58), .B(
        u_decode_add_x_16_n57), .Q(u_decode_add_x_16_n6) );
  NAND22 add_x_1_U51 ( .A(mem_data_pc4[20]), .B(mem_data_pc4[21]), .Q(
        add_x_1_n40) );
  NAND22 add_x_1_U60 ( .A(mem_data_pc4[18]), .B(mem_data_pc4[19]), .Q(
        add_x_1_n47) );
  NAND22 add_x_1_U96 ( .A(mem_data_pc4[12]), .B(mem_data_pc4[13]), .Q(
        add_x_1_n77) );
  NAND22 u_decode_add_x_16_U163 ( .A(u_decode_add_x_16_n202), .B(
        u_decode_add_x_16_n136), .Q(u_decode_add_x_16_n20) );
  NAND22 u_decode_add_x_16_U173 ( .A(u_decode_add_x_16_n203), .B(
        u_decode_add_x_16_n143), .Q(u_decode_add_x_16_n21) );
  NAND22 u_decode_add_x_16_U111 ( .A(u_decode_add_x_16_n99), .B(
        u_decode_add_x_16_n102), .Q(u_decode_add_x_16_n14) );
  XOR21 add_x_1_U63 ( .A(add_x_1_n53), .B(add_x_1_n54), .Q(u_mem_pc8[18]) );
  XOR21 add_x_1_U10 ( .A(mem_data_pc4[28]), .B(add_x_1_n9), .Q(u_mem_pc8[28])
         );
  NAND22 u_decode_add_x_16_U190 ( .A(u_decode_add_x_16_n205), .B(
        u_decode_add_x_16_n154), .Q(u_decode_add_x_16_n23) );
  NAND22 u_decode_add_x_16_U212 ( .A(u_decode_add_x_16_n208), .B(
        u_decode_add_x_16_n167), .Q(u_decode_add_x_16_n26) );
  NAND22 u_decode_add_x_16_U221 ( .A(u_decode_add_x_16_n209), .B(
        u_decode_add_x_16_n173), .Q(u_decode_add_x_16_n27) );
  DFC3 u_decode_pipe_con_Ealuop_reg_4_ ( .D(u_decode_control_o_con_aluop_4_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[4]) );
  DFC3 u_mem_pipe_data_alures_reg_30_ ( .D(u_mem_resmux_o_data_alu[30]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[30]) );
  DFC3 u_decode_pipe_Fbmemout_reg_11_ ( .D(u_decode_fbmemmux_o_data_fmem[11]), 
        .C(clk), .RN(rst_n), .Q(for_fbmemout[11]) );
  DFC3 u_mem_pipe_data_alures_reg_13_ ( .D(u_mem_resmux_o_data_alu[13]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[13]) );
  DFC3 u_fetch_pipe_instr_reg_2_ ( .D(read_instruction[2]), .C(clk), .RN(rst_n), .Q(if_addr_j[4]) );
  DFC3 u_fetch_pipe_instr_reg_4_ ( .D(read_instruction[4]), .C(clk), .RN(rst_n), .Q(if_addr_j[6]) );
  DFC3 u_fetch_pipe_instr_reg_5_ ( .D(read_instruction[5]), .C(clk), .RN(rst_n), .Q(if_addr_j[7]) );
  DFC3 u_fetch_pipe_instr_reg_3_ ( .D(read_instruction[3]), .C(clk), .RN(rst_n), .Q(if_addr_j[5]), .QN(n258) );
  DFC3 u_fetch_pipe_instr_reg_1_ ( .D(read_instruction[1]), .C(clk), .RN(rst_n), .Q(if_addr_j[3]), .QN(n254) );
  DFC3 u_fetch_pipe_instr_reg_7_ ( .D(read_instruction[7]), .C(clk), .RN(rst_n), .Q(if_addr_j[9]) );
  DFC3 u_mem_pipe_data_alures_reg_14_ ( .D(u_mem_resmux_o_data_alu[14]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[14]) );
  DFC3 u_mem_pipe_data_alures_reg_19_ ( .D(u_mem_resmux_o_data_alu[19]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[19]) );
  DFC3 u_decode_pipe_data_rs_reg_15_ ( .D(id_data_jr[15]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[15]) );
  DFC3 u_mem_pipe_data_alures_reg_6_ ( .D(u_mem_resmux_o_data_alu[6]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[6]) );
  NAND21 u_decode_add_x_16_U193 ( .A(if_addr_j[9]), .B(id_addr_pc4[9]), .Q(
        u_decode_add_x_16_n154) );
  NAND21 u_decode_add_x_16_U158 ( .A(if_addr_j[13]), .B(id_addr_pc4[13]), .Q(
        u_decode_add_x_16_n131) );
  NAND22 u_decode_add_x_16_U133 ( .A(if_addr_j[16]), .B(id_addr_pc4[16]), .Q(
        u_decode_add_x_16_n115) );
  NOR22 u_decode_add_x_16_U91 ( .A(id_addr_pc4[21]), .B(n324), .Q(
        u_decode_add_x_16_n88) );
  NOR22 u_decode_add_x_16_U60 ( .A(id_addr_pc4[25]), .B(n324), .Q(
        u_decode_add_x_16_n69) );
  OAI211 u_decode_add_x_16_U189 ( .A(u_decode_add_x_16_n157), .B(
        u_decode_add_x_16_n153), .C(u_decode_add_x_16_n154), .Q(
        u_decode_add_x_16_n152) );
  NOR22 u_decode_add_x_16_U66 ( .A(id_addr_pc4[24]), .B(n324), .Q(
        u_decode_add_x_16_n72) );
  NOR22 u_decode_add_x_16_U74 ( .A(id_addr_pc4[23]), .B(n324), .Q(
        u_decode_add_x_16_n77) );
  NOR22 u_decode_add_x_16_U80 ( .A(id_addr_pc4[22]), .B(n324), .Q(
        u_decode_add_x_16_n80) );
  NOR21 u_decode_add_x_16_U4 ( .A(if_addr_j[31]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n31) );
  NAND21 u_decode_add_x_16_U5 ( .A(n324), .B(if_addr_j[31]), .Q(
        u_decode_add_x_16_n32) );
  OAI211 u_decode_add_x_16_U154 ( .A(u_decode_add_x_16_n136), .B(
        u_decode_add_x_16_n130), .C(u_decode_add_x_16_n131), .Q(
        u_decode_add_x_16_n129) );
  OAI211 u_decode_add_x_16_U88 ( .A(u_decode_add_x_16_n92), .B(
        u_decode_add_x_16_n88), .C(u_decode_add_x_16_n89), .Q(
        u_decode_add_x_16_n87) );
  OAI211 u_decode_add_x_16_U25 ( .A(u_decode_add_x_16_n46), .B(
        u_decode_add_x_16_n50), .C(u_decode_add_x_16_n47), .Q(
        u_decode_add_x_16_n45) );
  OAI211 u_decode_add_x_16_U195 ( .A(u_decode_add_x_16_n156), .B(
        u_decode_add_x_16_n158), .C(u_decode_add_x_16_n157), .Q(
        u_decode_add_x_16_n155) );
  XOR22 add_x_4_U1 ( .A(instruction_address[31]), .B(add_x_4_n116), .Q(
        u_fetch_jmux_i_addr_pc4_31_) );
  NAND22 u_decode_add_x_16_U224 ( .A(if_addr_j[5]), .B(id_addr_pc4[5]), .Q(
        u_decode_add_x_16_n173) );
  OAI211 u_decode_add_x_16_U123 ( .A(u_decode_add_x_16_n115), .B(
        u_decode_add_x_16_n111), .C(u_decode_add_x_16_n112), .Q(
        u_decode_add_x_16_n110) );
  NAND22 u_decode_add_x_16_U54 ( .A(u_decode_add_x_16_n75), .B(
        u_decode_add_x_16_n67), .Q(u_decode_add_x_16_n65) );
  NAND22 add_x_1_U94 ( .A(add_x_1_n92), .B(add_x_1_n76), .Q(add_x_1_n75) );
  XNR21 u_decode_add_x_16_U216 ( .A(u_decode_add_x_16_n27), .B(
        u_decode_add_x_16_n174), .Q(u_decode_pcadd_o_addr_pcbranchE[5]) );
  XNR21 u_decode_add_x_16_U208 ( .A(u_decode_add_x_16_n26), .B(
        u_decode_add_x_16_n168), .Q(u_decode_pcadd_o_addr_pcbranchE[6]) );
  NAND22 add_x_1_U82 ( .A(add_x_1_n74), .B(add_x_1_n66), .Q(add_x_1_n65) );
  XNR21 u_decode_add_x_16_U107 ( .A(u_decode_add_x_16_n14), .B(
        u_decode_add_x_16_n103), .Q(u_decode_pcadd_o_addr_pcbranchE[18]) );
  XNR21 u_decode_add_x_16_U115 ( .A(u_decode_add_x_16_n15), .B(
        u_decode_add_x_16_n113), .Q(u_decode_pcadd_o_addr_pcbranchE[17]) );
  XNR21 u_decode_add_x_16_U50 ( .A(u_decode_add_x_16_n7), .B(
        u_decode_add_x_16_n71), .Q(u_decode_pcadd_o_addr_pcbranchE[25]) );
  XNR21 u_decode_add_x_16_U20 ( .A(u_decode_add_x_16_n4), .B(
        u_decode_add_x_16_n48), .Q(u_decode_pcadd_o_addr_pcbranchE[28]) );
  XNR21 u_decode_add_x_16_U1 ( .A(u_decode_add_x_16_n1), .B(
        u_decode_add_x_16_n33), .Q(u_decode_pcadd_o_addr_pcbranchE[31]) );
  XNR21 u_decode_add_x_16_U30 ( .A(u_decode_add_x_16_n5), .B(
        u_decode_add_x_16_n55), .Q(u_decode_pcadd_o_addr_pcbranchE[27]) );
  XNR21 u_decode_add_x_16_U68 ( .A(u_decode_add_x_16_n9), .B(
        u_decode_add_x_16_n79), .Q(u_decode_pcadd_o_addr_pcbranchE[23]) );
  XNR21 u_decode_add_x_16_U82 ( .A(u_decode_add_x_16_n11), .B(
        u_decode_add_x_16_n90), .Q(u_decode_pcadd_o_addr_pcbranchE[21]) );
  NAND22 add_x_4_U132 ( .A(instruction_address[4]), .B(instruction_address[5]), 
        .Q(add_x_4_n104) );
  NAND22 u_decode_add_x_16_U176 ( .A(if_addr_j[11]), .B(id_addr_pc4[11]), .Q(
        u_decode_add_x_16_n143) );
  NAND22 u_decode_add_x_16_U207 ( .A(if_addr_j[7]), .B(id_addr_pc4[7]), .Q(
        u_decode_add_x_16_n162) );
  NOR21 u_decode_add_x_16_U10 ( .A(if_addr_j[30]), .B(n324), .Q(
        u_decode_add_x_16_n34) );
  NOR21 add_x_1_U117 ( .A(add_x_1_n95), .B(add_x_1_n102), .Q(add_x_1_n94) );
  NOR21 add_x_1_U50 ( .A(add_x_1_n40), .B(add_x_1_n47), .Q(add_x_1_n39) );
  NOR21 add_x_1_U72 ( .A(add_x_1_n58), .B(add_x_1_n67), .Q(add_x_1_n57) );
  NOR22 u_decode_add_x_16_U105 ( .A(id_addr_pc4[19]), .B(n324), .Q(
        u_decode_add_x_16_n96) );
  NOR22 u_decode_add_x_16_U97 ( .A(id_addr_pc4[20]), .B(n324), .Q(
        u_decode_add_x_16_n91) );
  NOR21 u_decode_add_x_16_U219 ( .A(u_decode_add_x_16_n172), .B(
        u_decode_add_x_16_n175), .Q(u_decode_add_x_16_n170) );
  NAND22 add_x_1_U71 ( .A(add_x_1_n76), .B(add_x_1_n57), .Q(add_x_1_n56) );
  NOR22 u_decode_add_x_16_U87 ( .A(u_decode_add_x_16_n88), .B(
        u_decode_add_x_16_n91), .Q(u_decode_add_x_16_n86) );
  NAND22 u_decode_add_x_16_U151 ( .A(u_decode_add_x_16_n140), .B(
        u_decode_add_x_16_n128), .Q(u_decode_add_x_16_n126) );
  AOI211 u_decode_add_x_16_U187 ( .A(u_decode_add_x_16_n160), .B(
        u_decode_add_x_16_n151), .C(u_decode_add_x_16_n152), .Q(
        u_decode_add_x_16_n150) );
  XNR21 add_x_4_U135 ( .A(n274), .B(add_x_4_n110), .Q(
        u_fetch_jmux_i_addr_pc4_4_) );
  NAND22 add_x_4_U68 ( .A(add_x_4_n69), .B(add_x_4_n53), .Q(add_x_4_n52) );
  NAND22 add_x_1_U116 ( .A(add_x_1_n94), .B(add_x_1_n110), .Q(add_x_1_n93) );
  XOR21 add_x_4_U129 ( .A(n292), .B(add_x_4_n107), .Q(
        u_fetch_jmux_i_addr_pc4_5_) );
  XOR21 add_x_4_U124 ( .A(n295), .B(add_x_4_n102), .Q(
        u_fetch_jmux_i_addr_pc4_6_) );
  NOR21 add_x_4_U125 ( .A(n295), .B(add_x_4_n102), .Q(add_x_4_n98) );
  OAI211 u_decode_add_x_16_U226 ( .A(u_decode_add_x_16_n175), .B(
        u_decode_add_x_16_n177), .C(u_decode_add_x_16_n176), .Q(
        u_decode_add_x_16_n174) );
  AOI211 u_decode_add_x_16_U33 ( .A(u_decode_add_x_16_n51), .B(
        u_decode_add_x_16_n59), .C(u_decode_add_x_16_n52), .Q(
        u_decode_add_x_16_n50) );
  NAND22 u_decode_add_x_16_U85 ( .A(u_decode_add_x_16_n94), .B(
        u_decode_add_x_16_n86), .Q(u_decode_add_x_16_n84) );
  NOR21 add_x_4_U12 ( .A(add_x_4_n8), .B(add_x_4_n18), .Q(add_x_4_n7) );
  NOR21 add_x_1_U126 ( .A(add_x_1_n102), .B(add_x_1_n109), .Q(add_x_1_n101) );
  XNR21 add_x_4_U104 ( .A(n272), .B(add_x_4_n85), .Q(
        u_fetch_jmux_i_addr_pc4_10_) );
  XNR21 add_x_4_U119 ( .A(n291), .B(add_x_4_n98), .Q(
        u_fetch_jmux_i_addr_pc4_7_) );
  XNR21 add_x_4_U115 ( .A(n273), .B(add_x_4_n94), .Q(
        u_fetch_jmux_i_addr_pc4_8_) );
  XOR21 add_x_4_U98 ( .A(n289), .B(add_x_4_n82), .Q(
        u_fetch_jmux_i_addr_pc4_11_) );
  NOR21 add_x_4_U61 ( .A(n293), .B(add_x_4_n50), .Q(add_x_4_n46) );
  OAI211 u_decode_add_x_16_U178 ( .A(u_decode_add_x_16_n145), .B(
        u_decode_add_x_16_n147), .C(u_decode_add_x_16_n146), .Q(
        u_decode_add_x_16_n144) );
  AOI211 u_decode_add_x_16_U23 ( .A(u_decode_add_x_16_n64), .B(
        u_decode_add_x_16_n44), .C(u_decode_add_x_16_n45), .Q(
        u_decode_add_x_16_n43) );
  XOR21 add_x_4_U108 ( .A(n290), .B(add_x_4_n91), .Q(
        u_fetch_jmux_i_addr_pc4_9_) );
  XOR21 add_x_4_U93 ( .A(n294), .B(add_x_4_n77), .Q(
        u_fetch_jmux_i_addr_pc4_12_) );
  NOR21 add_x_1_U59 ( .A(add_x_1_n47), .B(add_x_1_n54), .Q(add_x_1_n46) );
  XOR21 add_x_4_U7 ( .A(n275), .B(add_x_4_n6), .Q(u_fetch_jmux_i_addr_pc4_29_)
         );
  XOR21 add_x_4_U60 ( .A(n293), .B(add_x_4_n50), .Q(
        u_fetch_jmux_i_addr_pc4_18_) );
  NOR21 add_x_4_U94 ( .A(n294), .B(add_x_4_n77), .Q(add_x_4_n73) );
  XNR21 add_x_4_U55 ( .A(n285), .B(add_x_4_n46), .Q(
        u_fetch_jmux_i_addr_pc4_19_) );
  XNR21 add_x_4_U86 ( .A(n288), .B(add_x_4_n73), .Q(
        u_fetch_jmux_i_addr_pc4_13_) );
  XNR21 add_x_4_U82 ( .A(n271), .B(add_x_4_n67), .Q(
        u_fetch_jmux_i_addr_pc4_14_) );
  XOR21 add_x_4_U44 ( .A(n284), .B(add_x_4_n39), .Q(
        u_fetch_jmux_i_addr_pc4_21_) );
  XOR21 add_x_4_U77 ( .A(n287), .B(add_x_4_n64), .Q(
        u_fetch_jmux_i_addr_pc4_15_) );
  XOR21 add_x_4_U65 ( .A(n286), .B(add_x_4_n57), .Q(
        u_fetch_jmux_i_addr_pc4_17_) );
  XOR21 add_x_4_U35 ( .A(n267), .B(add_x_4_n30), .Q(
        u_fetch_jmux_i_addr_pc4_23_) );
  XOR21 add_x_4_U24 ( .A(n266), .B(add_x_4_n23), .Q(
        u_fetch_jmux_i_addr_pc4_25_) );
  XOR21 add_x_4_U10 ( .A(n265), .B(add_x_4_n11), .Q(
        u_fetch_jmux_i_addr_pc4_28_) );
  NOR21 add_x_1_U4 ( .A(mem_data_pc4[30]), .B(add_x_1_n4), .Q(add_x_1_n2) );
  NOR21 u_decode_add_x_16_U236 ( .A(id_addr_pc4[3]), .B(if_addr_j[3]), .Q(
        u_decode_add_x_16_n179) );
  NOR21 u_decode_add_x_16_U214 ( .A(id_addr_pc4[6]), .B(if_addr_j[6]), .Q(
        u_decode_add_x_16_n166) );
  NAND22 add_x_4_U101 ( .A(instruction_address[10]), .B(
        instruction_address[11]), .Q(add_x_4_n79) );
  NAND22 add_x_4_U79 ( .A(instruction_address[14]), .B(instruction_address[15]), .Q(add_x_4_n61) );
  NAND22 u_decode_add_x_16_U141 ( .A(if_addr_j[15]), .B(id_addr_pc4[15]), .Q(
        u_decode_add_x_16_n120) );
  NOR21 add_x_1_U95 ( .A(add_x_1_n77), .B(add_x_1_n86), .Q(add_x_1_n76) );
  NOR21 add_x_4_U47 ( .A(add_x_4_n36), .B(add_x_4_n43), .Q(add_x_4_n35) );
  NAND22 u_decode_add_x_16_U61 ( .A(n324), .B(id_addr_pc4[25]), .Q(
        u_decode_add_x_16_n70) );
  NOR21 u_decode_add_x_16_U202 ( .A(u_decode_add_x_16_n161), .B(
        u_decode_add_x_16_n166), .Q(u_decode_add_x_16_n159) );
  NOR21 add_x_4_U69 ( .A(add_x_4_n54), .B(add_x_4_n61), .Q(add_x_4_n53) );
  NOR21 u_decode_add_x_16_U188 ( .A(u_decode_add_x_16_n153), .B(
        u_decode_add_x_16_n156), .Q(u_decode_add_x_16_n151) );
  NOR21 u_decode_add_x_16_U171 ( .A(u_decode_add_x_16_n142), .B(
        u_decode_add_x_16_n145), .Q(u_decode_add_x_16_n140) );
  NOR22 add_x_4_U131 ( .A(add_x_4_n111), .B(add_x_4_n104), .Q(add_x_4_n103) );
  NOR21 add_x_4_U111 ( .A(add_x_4_n88), .B(add_x_4_n95), .Q(add_x_4_n87) );
  NAND21 add_x_4_U136 ( .A(add_x_4_n110), .B(instruction_address[4]), .Q(
        add_x_4_n107) );
  NAND22 u_decode_add_x_16_U120 ( .A(u_decode_add_x_16_n109), .B(
        u_decode_add_x_16_n117), .Q(u_decode_add_x_16_n107) );
  NOR21 add_x_4_U120 ( .A(add_x_4_n95), .B(add_x_4_n102), .Q(add_x_4_n94) );
  NOR21 u_decode_add_x_16_U118 ( .A(u_decode_add_x_16_n126), .B(
        u_decode_add_x_16_n107), .Q(u_decode_add_x_16_n105) );
  NAND22 add_x_4_U46 ( .A(add_x_4_n51), .B(add_x_4_n35), .Q(add_x_4_n34) );
  AOI211 u_decode_add_x_16_U201 ( .A(u_decode_add_x_16_n168), .B(
        u_decode_add_x_16_n159), .C(u_decode_add_x_16_n160), .Q(
        u_decode_add_x_16_n158) );
  NAND22 add_x_4_U11 ( .A(add_x_4_n7), .B(add_x_4_n51), .Q(add_x_4_n6) );
  NAND22 add_x_4_U88 ( .A(add_x_4_n85), .B(add_x_4_n69), .Q(add_x_4_n68) );
  NAND22 add_x_4_U99 ( .A(add_x_4_n85), .B(add_x_4_n78), .Q(add_x_4_n77) );
  NOR21 add_x_1_U24 ( .A(add_x_1_n18), .B(add_x_1_n54), .Q(add_x_1_n17) );
  NAND22 add_x_1_U7 ( .A(add_x_1_n7), .B(mem_data_pc4[29]), .Q(add_x_1_n4) );
  XNR21 add_x_4_U73 ( .A(n270), .B(add_x_4_n60), .Q(
        u_fetch_jmux_i_addr_pc4_16_) );
  XNR21 add_x_4_U51 ( .A(n269), .B(add_x_4_n42), .Q(
        u_fetch_jmux_i_addr_pc4_20_) );
  XNR21 add_x_4_U40 ( .A(n268), .B(add_x_4_n33), .Q(
        u_fetch_jmux_i_addr_pc4_22_) );
  XOR21 add_x_4_U16 ( .A(n276), .B(add_x_4_n14), .Q(
        u_fetch_jmux_i_addr_pc4_27_) );
  NAND22 add_x_1_U73 ( .A(mem_data_pc4[16]), .B(mem_data_pc4[17]), .Q(
        add_x_1_n58) );
  NOR21 u_decode_add_x_16_U165 ( .A(id_addr_pc4[12]), .B(if_addr_j[12]), .Q(
        u_decode_add_x_16_n135) );
  NOR21 u_decode_add_x_16_U153 ( .A(u_decode_add_x_16_n130), .B(
        u_decode_add_x_16_n135), .Q(u_decode_add_x_16_n128) );
  NAND22 u_decode_add_x_16_U29 ( .A(if_addr_j[17]), .B(if_addr_j[28]), .Q(
        u_decode_add_x_16_n47) );
  NOR21 add_x_4_U89 ( .A(add_x_4_n70), .B(add_x_4_n79), .Q(add_x_4_n69) );
  NOR21 add_x_1_U137 ( .A(add_x_1_n118), .B(add_x_1_n111), .Q(add_x_1_n110) );
  NOR21 u_decode_add_x_16_U122 ( .A(u_decode_add_x_16_n114), .B(
        u_decode_add_x_16_n111), .Q(u_decode_add_x_16_n109) );
  AOI211 u_decode_add_x_16_U152 ( .A(u_decode_add_x_16_n141), .B(
        u_decode_add_x_16_n128), .C(u_decode_add_x_16_n129), .Q(
        u_decode_add_x_16_n127) );
  NAND22 add_x_4_U110 ( .A(add_x_4_n87), .B(add_x_4_n103), .Q(add_x_4_n86) );
  NOR22 add_x_4_U67 ( .A(add_x_4_n86), .B(add_x_4_n52), .Q(add_x_4_n51) );
  NOR21 add_x_4_U78 ( .A(add_x_4_n61), .B(add_x_4_n68), .Q(add_x_4_n60) );
  NOR21 add_x_1_U48 ( .A(add_x_1_n38), .B(add_x_1_n54), .Q(add_x_1_n37) );
  NOR21 add_x_1_U11 ( .A(mem_data_pc4[28]), .B(add_x_1_n9), .Q(add_x_1_n7) );
  NOR21 add_x_4_U56 ( .A(add_x_4_n43), .B(add_x_4_n50), .Q(add_x_4_n42) );
  XNR21 add_x_4_U3 ( .A(n264), .B(add_x_4_n4), .Q(u_fetch_jmux_i_addr_pc4_30_)
         );
  NAND22 add_x_4_U21 ( .A(add_x_4_n17), .B(instruction_address[26]), .Q(
        add_x_4_n14) );
  XNR21 add_x_4_U20 ( .A(n252), .B(add_x_4_n17), .Q(
        u_fetch_jmux_i_addr_pc4_26_) );
  XNR21 add_x_4_U31 ( .A(n263), .B(add_x_4_n26), .Q(
        u_fetch_jmux_i_addr_pc4_24_) );
  NAND22 add_x_1_U16 ( .A(mem_data_pc4[26]), .B(mem_data_pc4[27]), .Q(
        add_x_1_n11) );
  NOR21 u_decode_add_x_16_U136 ( .A(u_decode_add_x_16_n119), .B(
        u_decode_add_x_16_n122), .Q(u_decode_add_x_16_n117) );
  NOR21 add_x_4_U8 ( .A(n275), .B(add_x_4_n6), .Q(add_x_4_n4) );
  NOR21 add_x_4_U36 ( .A(add_x_4_n27), .B(add_x_4_n34), .Q(add_x_4_n26) );
  NOR21 u_decode_add_x_16_U198 ( .A(id_addr_pc4[8]), .B(if_addr_j[8]), .Q(
        u_decode_add_x_16_n156) );
  NOR21 u_decode_add_x_16_U181 ( .A(id_addr_pc4[10]), .B(if_addr_j[10]), .Q(
        u_decode_add_x_16_n145) );
  AOI211 u_decode_add_x_16_U218 ( .A(u_decode_add_x_16_n178), .B(
        u_decode_add_x_16_n170), .C(u_decode_add_x_16_n171), .Q(
        u_decode_add_x_16_n169) );
  NOR21 u_decode_add_x_16_U24 ( .A(u_decode_add_x_16_n46), .B(
        u_decode_add_x_16_n49), .Q(u_decode_add_x_16_n44) );
  DFP1 u_decode_pipe_con_Wregwrite_reg ( .D(n336), .C(clk), .SN(rst_n), .Q(
        n297), .QN(ex_con_Wregwrite) );
  DFP1 u_decode_pipe_addr_branch_reg_2_ ( .D(u_decode_add_x_16_n30), .C(clk), 
        .SN(rst_n), .Q(n307) );
  DFC3 u_decode_pipe_con_Ealuop_reg_2_ ( .D(u_decode_control_o_con_aluop_2_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[2]) );
  DFC3 u_fetch_pipe_instr_reg_15_ ( .D(read_instruction[15]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[17]), .QN(n256) );
  INV3 U204 ( .A(n282), .Q(n238) );
  NOR21 U205 ( .A(n370), .B(n369), .Q(n373) );
  NOR40 U206 ( .A(if_addr_j[7]), .B(if_addr_j[6]), .C(if_addr_j[4]), .D(n258), 
        .Q(n368) );
  NOR21 U207 ( .A(u_decode_add_x_16_n69), .B(u_decode_add_x_16_n72), .Q(
        u_decode_add_x_16_n67) );
  AOI211 U208 ( .A(u_decode_add_x_16_n95), .B(u_decode_add_x_16_n86), .C(
        u_decode_add_x_16_n87), .Q(u_decode_add_x_16_n85) );
  NOR21 U209 ( .A(n374), .B(n373), .Q(n377) );
  NOR31 U210 ( .A(n348), .B(n347), .C(n346), .Q(n354) );
  NOR22 U211 ( .A(id_data_instr[29]), .B(n333), .Q(n366) );
  NOR21 U212 ( .A(u_decode_add_x_16_n65), .B(u_decode_add_x_16_n84), .Q(
        u_decode_add_x_16_n63) );
  NOR21 U213 ( .A(u_decode_add_x_16_n77), .B(u_decode_add_x_16_n80), .Q(
        u_decode_add_x_16_n75) );
  NOR21 U214 ( .A(u_decode_add_x_16_n96), .B(u_decode_add_x_16_n101), .Q(
        u_decode_add_x_16_n94) );
  NOR21 U215 ( .A(id_addr_pc4[18]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n101) );
  NOR21 U216 ( .A(add_x_1_n93), .B(add_x_1_n56), .Q(add_x_1_n55) );
  NAND31 U217 ( .A(n340), .B(n339), .C(n311), .Q(n358) );
  BUF6 U218 ( .A(n573), .Q(n240) );
  BUF6 U219 ( .A(n363), .Q(n239) );
  NOR21 U220 ( .A(if_addr_j[28]), .B(n324), .Q(u_decode_add_x_16_n46) );
  NOR21 U221 ( .A(id_addr_pc4[26]), .B(n324), .Q(u_decode_add_x_16_n56) );
  AOI211 U222 ( .A(u_decode_add_x_16_n103), .B(u_decode_add_x_16_n63), .C(
        u_decode_add_x_16_n64), .Q(u_decode_add_x_16_n62) );
  AOI211 U223 ( .A(u_decode_add_x_16_n83), .B(u_decode_add_x_16_n75), .C(
        u_decode_add_x_16_n76), .Q(u_decode_add_x_16_n74) );
  AOI211 U224 ( .A(u_decode_add_x_16_n103), .B(u_decode_add_x_16_n94), .C(
        u_decode_add_x_16_n95), .Q(u_decode_add_x_16_n93) );
  NOR21 U225 ( .A(id_addr_pc4[17]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n111) );
  NOR21 U226 ( .A(id_addr_pc4[16]), .B(if_addr_j[16]), .Q(
        u_decode_add_x_16_n114) );
  AOI211 U227 ( .A(u_decode_add_x_16_n125), .B(u_decode_add_x_16_n117), .C(
        u_decode_add_x_16_n118), .Q(u_decode_add_x_16_n116) );
  NOR21 U228 ( .A(id_addr_pc4[15]), .B(if_addr_j[15]), .Q(
        u_decode_add_x_16_n119) );
  NOR21 U229 ( .A(id_addr_pc4[14]), .B(if_addr_j[14]), .Q(
        u_decode_add_x_16_n122) );
  NOR21 U230 ( .A(id_addr_pc4[13]), .B(if_addr_j[13]), .Q(
        u_decode_add_x_16_n130) );
  NOR21 U231 ( .A(id_addr_pc4[11]), .B(if_addr_j[11]), .Q(
        u_decode_add_x_16_n142) );
  NOR21 U232 ( .A(id_addr_pc4[9]), .B(if_addr_j[9]), .Q(u_decode_add_x_16_n153) );
  NOR21 U233 ( .A(id_addr_pc4[7]), .B(if_addr_j[7]), .Q(u_decode_add_x_16_n161) );
  NOR21 U234 ( .A(id_addr_pc4[5]), .B(if_addr_j[5]), .Q(u_decode_add_x_16_n172) );
  NOR21 U235 ( .A(id_addr_pc4[4]), .B(if_addr_j[4]), .Q(u_decode_add_x_16_n175) );
  NOR21 U236 ( .A(add_x_4_n18), .B(add_x_4_n50), .Q(add_x_4_n17) );
  AOI211 U237 ( .A(n316), .B(id_data_jr[21]), .C(n425), .Q(n427) );
  NAND31 U238 ( .A(n440), .B(n438), .C(n439), .Q(n118) );
  NAND31 U239 ( .A(n446), .B(n445), .C(n444), .Q(n119) );
  AOI211 U240 ( .A(n318), .B(n323), .C(n442), .Q(n446) );
  AOI211 U241 ( .A(n316), .B(id_data_jr[17]), .C(n449), .Q(n451) );
  NAND31 U242 ( .A(n456), .B(n458), .C(n457), .Q(n121) );
  AOI211 U243 ( .A(n316), .B(id_data_jr[15]), .C(n461), .Q(n463) );
  NAND31 U244 ( .A(n482), .B(n481), .C(n480), .Q(n125) );
  AOI211 U245 ( .A(n319), .B(if_addr_j[12]), .C(n478), .Q(n482) );
  NAND31 U246 ( .A(n502), .B(n500), .C(n501), .Q(n128) );
  AOI211 U247 ( .A(n318), .B(if_addr_j[9]), .C(n498), .Q(n502) );
  NAND31 U248 ( .A(n520), .B(n519), .C(n518), .Q(n131) );
  NAND31 U249 ( .A(n538), .B(n536), .C(n537), .Q(n134) );
  AOI211 U250 ( .A(n318), .B(if_addr_j[3]), .C(n534), .Q(n538) );
  NOR40 U251 ( .A(if_addr_j[23]), .B(if_addr_j[25]), .C(if_addr_j[27]), .D(
        if_addr_j[24]), .Q(n590) );
  NOR40 U252 ( .A(n591), .B(n592), .C(n593), .D(n594), .Q(n582) );
  CLKIN0 U253 ( .A(add_x_1_n29), .Q(n140) );
  NAND40 U254 ( .A(mem_data_pc4[24]), .B(mem_data_pc4[25]), .C(add_x_1_n39), 
        .D(n140), .Q(add_x_1_n18) );
  CLKIN0 U255 ( .A(data_address[19]), .Q(n141) );
  NOR20 U256 ( .A(add_x_1_n54), .B(add_x_1_n53), .Q(n142) );
  XNR20 U257 ( .A(mem_data_pc4[19]), .B(n142), .Q(n143) );
  IMUX20 U258 ( .A(n141), .B(n143), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[19]) );
  CLKIN0 U259 ( .A(data_address[13]), .Q(n144) );
  NOR20 U260 ( .A(add_x_1_n84), .B(add_x_1_n83), .Q(n145) );
  XNR20 U261 ( .A(mem_data_pc4[13]), .B(n145), .Q(n146) );
  IMUX20 U262 ( .A(n144), .B(n146), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[13]) );
  NAND20 U263 ( .A(add_x_1_n17), .B(mem_data_pc4[26]), .Q(n147) );
  XNR20 U264 ( .A(mem_data_pc4[27]), .B(n147), .Q(n148) );
  MUX21 U265 ( .A(data_address[27]), .B(n148), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[27]) );
  CLKIN0 U266 ( .A(data_address[26]), .Q(n149) );
  XNR20 U267 ( .A(add_x_1_n17), .B(mem_data_pc4[26]), .Q(n150) );
  IMUX20 U268 ( .A(n149), .B(n150), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[26]) );
  CLKIN0 U269 ( .A(data_address[15]), .Q(n151) );
  NOR20 U270 ( .A(add_x_1_n75), .B(add_x_1_n73), .Q(n152) );
  XNR20 U271 ( .A(mem_data_pc4[15]), .B(n152), .Q(n153) );
  IMUX20 U272 ( .A(n151), .B(n153), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[15]) );
  NAND20 U273 ( .A(add_x_1_n101), .B(mem_data_pc4[8]), .Q(n154) );
  XNR20 U274 ( .A(mem_data_pc4[9]), .B(n154), .Q(n155) );
  MUX21 U275 ( .A(data_address[9]), .B(n155), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[9]) );
  XNR20 U276 ( .A(n323), .B(for_o_addr_Erd[0]), .Q(n156) );
  IMUX20 U277 ( .A(n282), .B(n238), .S(for_o_addr_Erd[1]), .Q(n157) );
  IMUX20 U278 ( .A(n281), .B(if_addr_j[21]), .S(for_o_addr_Erd[3]), .Q(n158)
         );
  XNR20 U279 ( .A(n311), .B(for_o_addr_Erd[4]), .Q(n159) );
  NOR40 U280 ( .A(n297), .B(n157), .C(n158), .D(n159), .Q(n160) );
  OAI2110 U281 ( .A(n278), .B(for_o_addr_Erd[2]), .C(n160), .D(n156), .Q(n161)
         );
  AOI210 U282 ( .A(n278), .B(for_o_addr_Erd[2]), .C(n161), .Q(n360) );
  CLKIN0 U283 ( .A(u_decode_add_x_16_n40), .Q(n162) );
  AOI211 U284 ( .A(u_decode_add_x_16_n41), .B(u_decode_add_x_16_n37), .C(n162), 
        .Q(u_decode_add_x_16_n36) );
  OAI210 U285 ( .A(id_addr_pc4[2]), .B(if_addr_j[2]), .C(
        u_decode_add_x_16_n182), .Q(u_decode_add_x_16_n30) );
  CLKIN0 U286 ( .A(u_decode_add_x_16_n73), .Q(n163) );
  NOR20 U287 ( .A(u_decode_add_x_16_n72), .B(n163), .Q(n164) );
  XNR20 U288 ( .A(u_decode_add_x_16_n74), .B(n164), .Q(
        u_decode_pcadd_o_addr_pcbranchE[24]) );
  CLKIN0 U289 ( .A(u_decode_add_x_16_n92), .Q(n165) );
  NOR20 U290 ( .A(u_decode_add_x_16_n91), .B(n165), .Q(n166) );
  XNR20 U291 ( .A(u_decode_add_x_16_n93), .B(n166), .Q(
        u_decode_pcadd_o_addr_pcbranchE[20]) );
  CLKIN0 U292 ( .A(u_decode_add_x_16_n115), .Q(n167) );
  NOR20 U293 ( .A(u_decode_add_x_16_n114), .B(n167), .Q(n168) );
  XNR20 U294 ( .A(u_decode_add_x_16_n116), .B(n168), .Q(
        u_decode_pcadd_o_addr_pcbranchE[16]) );
  CLKIN0 U295 ( .A(u_decode_add_x_16_n136), .Q(n169) );
  AOI210 U296 ( .A(u_decode_add_x_16_n137), .B(u_decode_add_x_16_n202), .C(
        n169), .Q(n170) );
  CLKIN0 U297 ( .A(u_decode_add_x_16_n131), .Q(n171) );
  NOR20 U298 ( .A(u_decode_add_x_16_n130), .B(n171), .Q(n172) );
  XNR20 U299 ( .A(n170), .B(n172), .Q(u_decode_pcadd_o_addr_pcbranchE[13]) );
  CLKIN0 U300 ( .A(u_decode_add_x_16_n157), .Q(n173) );
  NOR20 U301 ( .A(u_decode_add_x_16_n156), .B(n173), .Q(n174) );
  XNR20 U302 ( .A(u_decode_add_x_16_n158), .B(n174), .Q(
        u_decode_pcadd_o_addr_pcbranchE[8]) );
  CLKIN0 U303 ( .A(data_address[25]), .Q(n175) );
  NOR20 U304 ( .A(add_x_1_n27), .B(add_x_1_n26), .Q(n176) );
  XNR20 U305 ( .A(mem_data_pc4[25]), .B(n176), .Q(n177) );
  IMUX20 U306 ( .A(n175), .B(n177), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[25]) );
  NAND20 U307 ( .A(add_x_1_n46), .B(mem_data_pc4[20]), .Q(n178) );
  XNR20 U308 ( .A(mem_data_pc4[21]), .B(n178), .Q(n179) );
  MUX21 U309 ( .A(data_address[21]), .B(n179), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[21]) );
  NAND20 U310 ( .A(add_x_1_n92), .B(mem_data_pc4[10]), .Q(n180) );
  XNR20 U311 ( .A(mem_data_pc4[11]), .B(n180), .Q(n181) );
  MUX21 U312 ( .A(data_address[11]), .B(n181), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[11]) );
  CLKIN0 U313 ( .A(data_address[8]), .Q(n182) );
  XNR20 U314 ( .A(add_x_1_n101), .B(mem_data_pc4[8]), .Q(n183) );
  IMUX20 U315 ( .A(n182), .B(n183), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[8]) );
  NAND20 U316 ( .A(add_x_1_n117), .B(mem_data_pc4[4]), .Q(n184) );
  XNR20 U317 ( .A(mem_data_pc4[5]), .B(n184), .Q(n185) );
  MUX21 U318 ( .A(data_address[5]), .B(n185), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[5]) );
  CLKIN0 U319 ( .A(data_address[3]), .Q(n186) );
  XNR20 U320 ( .A(mem_data_pc4[3]), .B(mem_data_pc4[2]), .Q(n187) );
  IMUX20 U321 ( .A(n186), .B(n187), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[3]) );
  CLKIN0 U322 ( .A(add_x_4_n27), .Q(n188) );
  NAND40 U323 ( .A(instruction_address[24]), .B(instruction_address[25]), .C(
        add_x_4_n35), .D(n188), .Q(add_x_4_n18) );
  IMUX20 U324 ( .A(n261), .B(if_addr_j[23]), .S(for_o_addr_Erd[0]), .Q(n189)
         );
  IMUX20 U325 ( .A(n260), .B(if_addr_j[24]), .S(for_o_addr_Erd[1]), .Q(n190)
         );
  NOR40 U326 ( .A(if_addr_j[27]), .B(for_o_addr_Erd[1]), .C(for_o_addr_Erd[3]), 
        .D(for_o_addr_Erd[0]), .Q(n191) );
  IMUX20 U327 ( .A(if_addr_j[26]), .B(n280), .S(for_o_addr_Erd[3]), .Q(n192)
         );
  OAI210 U328 ( .A(for_o_addr_Erd[2]), .B(n191), .C(n277), .Q(n193) );
  OAI2110 U329 ( .A(for_o_addr_Erd[2]), .B(n277), .C(n192), .D(n193), .Q(n194)
         );
  NAND20 U330 ( .A(n279), .B(for_o_addr_Erd[4]), .Q(n195) );
  OAI2110 U331 ( .A(n279), .B(for_o_addr_Erd[4]), .C(ex_con_Wregwrite), .D(
        n195), .Q(n196) );
  NOR40 U332 ( .A(n189), .B(n190), .C(n194), .D(n196), .Q(n565) );
  NAND20 U333 ( .A(u_decode_control_o_con_aluop_0_), .B(n364), .Q(n197) );
  AOI210 U334 ( .A(n197), .B(n598), .C(n251), .Q(
        u_decode_control_o_con_aluop_4_) );
  NAND20 U335 ( .A(n358), .B(n360), .Q(n198) );
  NAND20 U336 ( .A(n359), .B(n198), .Q(u_decode_n23) );
  CLKIN0 U337 ( .A(u_decode_add_x_16_n35), .Q(n199) );
  NOR20 U338 ( .A(u_decode_add_x_16_n34), .B(n199), .Q(n200) );
  XNR20 U339 ( .A(u_decode_add_x_16_n36), .B(n200), .Q(
        u_decode_pcadd_o_addr_pcbranchE[30]) );
  CLKIN0 U340 ( .A(u_decode_add_x_16_n81), .Q(n201) );
  NOR20 U341 ( .A(u_decode_add_x_16_n80), .B(n201), .Q(n202) );
  XNR20 U342 ( .A(u_decode_add_x_16_n82), .B(n202), .Q(
        u_decode_pcadd_o_addr_pcbranchE[22]) );
  CLKIN0 U343 ( .A(u_decode_add_x_16_n102), .Q(n203) );
  AOI210 U344 ( .A(u_decode_add_x_16_n103), .B(u_decode_add_x_16_n99), .C(n203), .Q(n204) );
  CLKIN0 U345 ( .A(u_decode_add_x_16_n97), .Q(n205) );
  NOR20 U346 ( .A(u_decode_add_x_16_n96), .B(n205), .Q(n206) );
  XNR20 U347 ( .A(n204), .B(n206), .Q(u_decode_pcadd_o_addr_pcbranchE[19]) );
  CLKIN0 U348 ( .A(u_decode_add_x_16_n123), .Q(n207) );
  NOR20 U349 ( .A(u_decode_add_x_16_n122), .B(n207), .Q(n208) );
  XNR20 U350 ( .A(u_decode_add_x_16_n124), .B(n208), .Q(
        u_decode_pcadd_o_addr_pcbranchE[14]) );
  CLKIN0 U351 ( .A(u_decode_add_x_16_n146), .Q(n209) );
  NOR20 U352 ( .A(u_decode_add_x_16_n145), .B(n209), .Q(n210) );
  XNR20 U353 ( .A(u_decode_add_x_16_n147), .B(n210), .Q(
        u_decode_pcadd_o_addr_pcbranchE[10]) );
  CLKIN0 U354 ( .A(u_decode_add_x_16_n167), .Q(n211) );
  AOI210 U355 ( .A(u_decode_add_x_16_n168), .B(u_decode_add_x_16_n208), .C(
        n211), .Q(n212) );
  CLKIN0 U356 ( .A(u_decode_add_x_16_n162), .Q(n213) );
  NOR20 U357 ( .A(u_decode_add_x_16_n161), .B(n213), .Q(n214) );
  XNR20 U358 ( .A(n212), .B(n214), .Q(u_decode_pcadd_o_addr_pcbranchE[7]) );
  CLKIN0 U359 ( .A(u_decode_add_x_16_n176), .Q(n215) );
  NOR20 U360 ( .A(u_decode_add_x_16_n175), .B(n215), .Q(n216) );
  XNR20 U361 ( .A(u_decode_add_x_16_n177), .B(n216), .Q(
        u_decode_pcadd_o_addr_pcbranchE[4]) );
  CLKIN0 U362 ( .A(u_decode_add_x_16_n180), .Q(n217) );
  NOR20 U363 ( .A(u_decode_add_x_16_n179), .B(n217), .Q(n218) );
  XNR20 U364 ( .A(u_decode_add_x_16_n182), .B(n218), .Q(
        u_decode_pcadd_o_addr_pcbranchE[3]) );
  CLKIN0 U365 ( .A(data_address[29]), .Q(n219) );
  XNR20 U366 ( .A(add_x_1_n7), .B(mem_data_pc4[29]), .Q(n220) );
  IMUX20 U367 ( .A(n219), .B(n220), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[29]) );
  CLKIN0 U368 ( .A(data_address[23]), .Q(n221) );
  NOR20 U369 ( .A(add_x_1_n36), .B(add_x_1_n35), .Q(n222) );
  XNR20 U370 ( .A(mem_data_pc4[23]), .B(n222), .Q(n223) );
  IMUX20 U371 ( .A(n221), .B(n223), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[23]) );
  CLKIN0 U372 ( .A(data_address[20]), .Q(n224) );
  XNR20 U373 ( .A(add_x_1_n46), .B(mem_data_pc4[20]), .Q(n225) );
  IMUX20 U374 ( .A(n224), .B(n225), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[20]) );
  CLKIN0 U375 ( .A(data_address[17]), .Q(n226) );
  NOR20 U376 ( .A(add_x_1_n65), .B(add_x_1_n64), .Q(n227) );
  XNR20 U377 ( .A(mem_data_pc4[17]), .B(n227), .Q(n228) );
  IMUX20 U378 ( .A(n226), .B(n228), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[17]) );
  CLKIN0 U379 ( .A(data_address[10]), .Q(n229) );
  XNR20 U380 ( .A(add_x_1_n92), .B(mem_data_pc4[10]), .Q(n230) );
  IMUX20 U381 ( .A(n229), .B(n230), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[10]) );
  CLKIN0 U382 ( .A(data_address[7]), .Q(n231) );
  NOR20 U383 ( .A(add_x_1_n109), .B(add_x_1_n108), .Q(n232) );
  XNR20 U384 ( .A(mem_data_pc4[7]), .B(n232), .Q(n233) );
  IMUX20 U385 ( .A(n231), .B(n233), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[7]) );
  CLKIN0 U386 ( .A(data_address[4]), .Q(n234) );
  XNR20 U387 ( .A(add_x_1_n117), .B(mem_data_pc4[4]), .Q(n235) );
  IMUX20 U388 ( .A(n234), .B(n235), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[4]) );
  CLKIN0 U389 ( .A(data_address[2]), .Q(n236) );
  IMUX20 U390 ( .A(n236), .B(mem_data_pc4[2]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[2]) );
  NAND23 U391 ( .A(n320), .B(if_addr_b[10]), .Q(n494) );
  NAND23 U392 ( .A(n320), .B(if_addr_b[4]), .Q(n530) );
  NAND24 U393 ( .A(n406), .B(n407), .Q(n241) );
  NOR22 U394 ( .A(n533), .B(n322), .Q(n534) );
  NOR22 U395 ( .A(n497), .B(n322), .Q(n498) );
  AOI212 U396 ( .A(n319), .B(if_addr_j[16]), .C(n454), .Q(n458) );
  NOR22 U397 ( .A(n483), .B(n322), .Q(n484) );
  NOR22 U398 ( .A(n503), .B(n322), .Q(n504) );
  NAND33 U399 ( .A(n428), .B(n427), .C(n426), .Q(n116) );
  NAND33 U400 ( .A(n550), .B(n549), .C(n548), .Q(n136) );
  NAND33 U401 ( .A(n434), .B(n433), .C(n432), .Q(n117) );
  NOR21 U402 ( .A(n423), .B(n546), .Q(n424) );
  AOI211 U403 ( .A(n319), .B(if_addr_j[10]), .C(n492), .Q(n496) );
  INV15 U404 ( .A(if_con_b), .Q(n490) );
  NAND33 U405 ( .A(n545), .B(n544), .C(n543), .Q(n135) );
  NOR23 U406 ( .A(n515), .B(n309), .Q(n516) );
  NOR22 U407 ( .A(n441), .B(n309), .Q(n442) );
  NOR22 U408 ( .A(n477), .B(n309), .Q(n478) );
  NOR22 U409 ( .A(n465), .B(n309), .Q(n466) );
  AOI212 U410 ( .A(n244), .B(u_fetch_jmux_i_addr_pc4_26_), .C(n400), .Q(n403)
         );
  AOI212 U411 ( .A(n244), .B(u_fetch_jmux_i_addr_pc4_24_), .C(n410), .Q(n413)
         );
  AOI212 U412 ( .A(n244), .B(u_fetch_jmux_i_addr_pc4_30_), .C(n380), .Q(n383)
         );
  INV3 U413 ( .A(n278), .Q(n237) );
  NAND33 U414 ( .A(n464), .B(n463), .C(n462), .Q(n122) );
  AOI212 U415 ( .A(n542), .B(u_fetch_jmux_i_addr_pc4_28_), .C(n390), .Q(n393)
         );
  NAND33 U416 ( .A(n246), .B(n249), .C(n250), .Q(n138) );
  NOR24 U417 ( .A(n378), .B(if_con_b), .Q(n540) );
  NOR22 U418 ( .A(n298), .B(n554), .Q(n247) );
  NOR31 U419 ( .A(n353), .B(n352), .C(n354), .Q(n363) );
  NAND31 U420 ( .A(n582), .B(n583), .C(n572), .Q(n573) );
  NOR23 U421 ( .A(n364), .B(n369), .Q(n541) );
  AOI212 U422 ( .A(n244), .B(u_fetch_jmux_i_addr_pc4_23_), .C(n415), .Q(n418)
         );
  NAND33 U423 ( .A(n452), .B(n451), .C(n450), .Q(n120) );
  AOI212 U424 ( .A(n318), .B(if_addr_j[13]), .C(n472), .Q(n476) );
  NAND33 U425 ( .A(n508), .B(n507), .C(n506), .Q(n129) );
  AOI212 U426 ( .A(n319), .B(if_addr_j[8]), .C(n504), .Q(n508) );
  NAND22 U427 ( .A(n408), .B(n242), .Q(n112) );
  CLKIN6 U428 ( .A(n241), .Q(n242) );
  NAND23 U429 ( .A(n315), .B(id_data_jr[25]), .Q(n407) );
  NAND23 U430 ( .A(n319), .B(if_addr_j[25]), .Q(n406) );
  NAND33 U431 ( .A(n470), .B(n469), .C(n468), .Q(n123) );
  AOI212 U432 ( .A(n319), .B(if_addr_j[14]), .C(n466), .Q(n470) );
  NAND33 U433 ( .A(n488), .B(n487), .C(n486), .Q(n126) );
  AOI212 U434 ( .A(n318), .B(if_addr_j[11]), .C(n484), .Q(n488) );
  AOI212 U435 ( .A(n244), .B(u_fetch_jmux_i_addr_pc4_27_), .C(n395), .Q(n398)
         );
  AOI212 U436 ( .A(n244), .B(u_fetch_jmux_i_addr_pc4_29_), .C(n385), .Q(n388)
         );
  IMUX23 U437 ( .A(n244), .B(n541), .S(instruction_address[2]), .Q(n544) );
  NAND26 U438 ( .A(n490), .B(n489), .Q(n243) );
  INV15 U439 ( .A(n317), .Q(n319) );
  INV12 U440 ( .A(n540), .Q(n317) );
  NOR22 U441 ( .A(n453), .B(n546), .Q(n454) );
  NOR22 U442 ( .A(n471), .B(n322), .Q(n472) );
  CLKBU15 U443 ( .A(n542), .Q(n244) );
  NAND33 U444 ( .A(n393), .B(n392), .C(n391), .Q(n109) );
  AOI211 U445 ( .A(n244), .B(u_fetch_jmux_i_addr_pc4_25_), .C(n405), .Q(n408)
         );
  NAND33 U446 ( .A(n532), .B(n531), .C(n530), .Q(n133) );
  NAND33 U447 ( .A(n496), .B(n495), .C(n494), .Q(n127) );
  NAND33 U448 ( .A(n474), .B(n476), .C(n475), .Q(n124) );
  NAND28 U449 ( .A(n490), .B(n489), .Q(n546) );
  NAND28 U450 ( .A(n490), .B(n489), .Q(n322) );
  NAND26 U451 ( .A(n490), .B(n489), .Q(n309) );
  NOR22 U452 ( .A(n554), .B(n307), .Q(n539) );
  NAND28 U453 ( .A(if_con_b), .B(n313), .Q(n554) );
  INV3 U454 ( .A(add_x_4_n51), .Q(add_x_4_n50) );
  INV3 U455 ( .A(add_x_1_n55), .Q(add_x_1_n54) );
  INV1 U456 ( .A(u_decode_add_x_16_n111), .Q(u_decode_add_x_16_n197) );
  INV1 U457 ( .A(u_decode_add_x_16_n142), .Q(u_decode_add_x_16_n203) );
  INV1 U458 ( .A(u_decode_add_x_16_n153), .Q(u_decode_add_x_16_n205) );
  INV1 U459 ( .A(u_decode_add_x_16_n119), .Q(u_decode_add_x_16_n199) );
  INV3 U460 ( .A(n541), .Q(n313) );
  NOR20 U461 ( .A(n335), .B(n334), .Q(u_decode_jbcon_o_con_aluPC4) );
  AOI311 U462 ( .A(n254), .B(n259), .C(n368), .D(n367), .Q(n370) );
  INV1 U463 ( .A(add_x_1_n118), .Q(add_x_1_n117) );
  IMUX20 U464 ( .A(n260), .B(if_addr_j[24]), .S(for_addr_rtM[1]), .Q(n588) );
  INV1 U465 ( .A(u_fetch_jmux_i_addr_pc4_16_), .Q(n453) );
  INV3 U466 ( .A(n377), .Q(n378) );
  NAND41 U467 ( .A(for_FWmemread), .B(n358), .C(n351), .D(n580), .Q(n352) );
  NOR20 U468 ( .A(n365), .B(n334), .Q(u_decode_control_o_con_regdst) );
  INV2 U469 ( .A(add_x_1_n39), .Q(add_x_1_n38) );
  INV2 U470 ( .A(u_decode_add_x_16_n69), .Q(u_decode_add_x_16_n189) );
  INV2 U471 ( .A(n560), .Q(u_decode_n4) );
  INV1 U472 ( .A(n366), .Q(n334) );
  NAND22 U473 ( .A(n366), .B(n325), .Q(n369) );
  INV2 U474 ( .A(add_x_1_n110), .Q(add_x_1_n109) );
  NAND41 U475 ( .A(mem_read), .B(n584), .C(n583), .D(n585), .Q(n572) );
  INV2 U476 ( .A(u_decode_add_x_16_n46), .Q(u_decode_add_x_16_n186) );
  NAND31 U477 ( .A(n581), .B(n350), .C(n349), .Q(n353) );
  MUX21 U478 ( .A(data_address[0]), .B(u_mem_pc8[0]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[0]) );
  INV3 U479 ( .A(n367), .Q(n364) );
  NOR40 U480 ( .A(n586), .B(n587), .C(n588), .D(n589), .Q(n584) );
  INV2 U481 ( .A(u_decode_add_x_16_n135), .Q(u_decode_add_x_16_n202) );
  MUX21 U482 ( .A(mem_data_alures[16]), .B(wb_data_memout[16]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[16]) );
  MUX21 U483 ( .A(mem_data_alures[23]), .B(wb_data_memout[23]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[23]) );
  MUX21 U484 ( .A(mem_data_alures[18]), .B(wb_data_memout[18]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[18]) );
  MUX21 U485 ( .A(mem_data_alures[8]), .B(wb_data_memout[8]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[8]) );
  MUX21 U486 ( .A(mem_data_alures[6]), .B(wb_data_memout[6]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[6]) );
  MUX21 U487 ( .A(mem_data_alures[3]), .B(wb_data_memout[3]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[3]) );
  MUX21 U488 ( .A(mem_data_alures[2]), .B(wb_data_memout[2]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[2]) );
  MUX21 U489 ( .A(mem_data_alures[17]), .B(wb_data_memout[17]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[17]) );
  MUX21 U490 ( .A(mem_data_alures[31]), .B(wb_data_memout[31]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[31]) );
  BUF6 U491 ( .A(if_addr_j[17]), .Q(n324) );
  MUX21 U492 ( .A(mem_data_alures[19]), .B(wb_data_memout[19]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[19]) );
  MUX21 U493 ( .A(mem_data_alures[21]), .B(wb_data_memout[21]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[21]) );
  MUX21 U494 ( .A(mem_data_alures[0]), .B(wb_data_memout[0]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[0]) );
  MUX21 U495 ( .A(mem_data_alures[12]), .B(wb_data_memout[12]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[12]) );
  MUX21 U496 ( .A(mem_data_alures[13]), .B(wb_data_memout[13]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[13]) );
  MUX21 U497 ( .A(mem_data_alures[11]), .B(wb_data_memout[11]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[11]) );
  INV2 U498 ( .A(mem_data_pc4[12]), .Q(add_x_1_n83) );
  INV2 U499 ( .A(mem_data_pc4[14]), .Q(add_x_1_n73) );
  INV1 U500 ( .A(u_fetch_jmux_i_addr_pc4_15_), .Q(n459) );
  INV1 U501 ( .A(u_fetch_jmux_i_addr_pc4_17_), .Q(n447) );
  INV1 U502 ( .A(u_fetch_jmux_i_addr_pc4_19_), .Q(n435) );
  INV1 U503 ( .A(u_fetch_jmux_i_addr_pc4_14_), .Q(n465) );
  INV1 U504 ( .A(u_fetch_jmux_i_addr_pc4_20_), .Q(n429) );
  INV1 U505 ( .A(u_fetch_jmux_i_addr_pc4_12_), .Q(n477) );
  INV1 U506 ( .A(u_fetch_jmux_i_addr_pc4_9_), .Q(n497) );
  INV3 U507 ( .A(u_decode_add_x_16_n104), .Q(u_decode_add_x_16_n103) );
  INV1 U508 ( .A(u_fetch_jmux_i_addr_pc4_11_), .Q(n483) );
  INV1 U509 ( .A(u_fetch_jmux_i_addr_pc4_18_), .Q(n441) );
  INV3 U510 ( .A(add_x_1_n75), .Q(add_x_1_n74) );
  NOR23 U511 ( .A(n372), .B(n371), .Q(n376) );
  INV1 U512 ( .A(u_fetch_jmux_i_addr_pc4_7_), .Q(n509) );
  INV1 U513 ( .A(u_fetch_jmux_i_addr_pc4_8_), .Q(n503) );
  INV2 U514 ( .A(u_decode_control_o_con_aluop_5_), .Q(n330) );
  INV1 U515 ( .A(u_fetch_jmux_i_addr_pc4_5_), .Q(n521) );
  INV3 U516 ( .A(n373), .Q(n371) );
  INV1 U517 ( .A(u_fetch_jmux_i_addr_pc4_6_), .Q(n515) );
  NAND31 U518 ( .A(n358), .B(mem_read), .C(n345), .Q(n346) );
  INV3 U519 ( .A(add_x_4_n86), .Q(add_x_4_n85) );
  NAND22 U520 ( .A(n366), .B(n365), .Q(n374) );
  INV3 U521 ( .A(add_x_1_n93), .Q(add_x_1_n92) );
  INV1 U522 ( .A(u_fetch_jmux_i_addr_pc4_4_), .Q(n527) );
  INV2 U523 ( .A(u_decode_add_x_16_n141), .Q(u_decode_add_x_16_n139) );
  NOR21 U524 ( .A(id_data_instr[31]), .B(n562), .Q(
        u_decode_control_o_con_aluop_0_) );
  NAND22 U525 ( .A(n590), .B(n280), .Q(n583) );
  MUX21 U526 ( .A(data_address[1]), .B(u_mem_pc8[1]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[1]) );
  INV2 U527 ( .A(u_decode_add_x_16_n166), .Q(u_decode_add_x_16_n208) );
  INV2 U528 ( .A(add_x_4_n79), .Q(add_x_4_n78) );
  INV2 U529 ( .A(add_x_4_n111), .Q(add_x_4_n110) );
  NOR21 U530 ( .A(n312), .B(id_data_instr[30]), .Q(n558) );
  BUF12 U531 ( .A(if_addr_j[18]), .Q(n323) );
  INV2 U532 ( .A(mem_data_pc4[18]), .Q(add_x_1_n53) );
  NAND31 U533 ( .A(n526), .B(n524), .C(n525), .Q(n132) );
  INV12 U534 ( .A(n314), .Q(n316) );
  INV12 U535 ( .A(n317), .Q(n318) );
  INV12 U536 ( .A(n314), .Q(n315) );
  INV1 U537 ( .A(u_fetch_jmux_i_addr_pc4_21_), .Q(n423) );
  OAI311 U538 ( .A(n362), .B(n361), .C(n360), .D(n359), .Q(
        u_decode_for_o_con_fb_0_) );
  INV2 U539 ( .A(n563), .Q(u_decode_n17) );
  INV3 U540 ( .A(u_decode_add_x_16_n83), .Q(u_decode_add_x_16_n82) );
  INV3 U541 ( .A(n489), .Q(n552) );
  INV3 U542 ( .A(n375), .Q(n248) );
  INV1 U543 ( .A(u_fetch_jmux_i_addr_pc4_13_), .Q(n471) );
  OAI311 U544 ( .A(n565), .B(n569), .C(n570), .D(n571), .Q(
        u_decode_for_o_con_fa_0_) );
  INV3 U545 ( .A(u_decode_add_x_16_n125), .Q(u_decode_add_x_16_n124) );
  NAND21 U546 ( .A(n541), .B(instruction_address[31]), .Q(n375) );
  INV3 U547 ( .A(add_x_1_n37), .Q(add_x_1_n36) );
  NAND21 U548 ( .A(n541), .B(instruction_address[29]), .Q(n384) );
  NAND21 U549 ( .A(n541), .B(instruction_address[27]), .Q(n394) );
  NOR21 U550 ( .A(n564), .B(n565), .Q(n563) );
  INV3 U551 ( .A(add_x_4_n68), .Q(add_x_4_n67) );
  INV1 U552 ( .A(u_fetch_jmux_i_addr_pc4_10_), .Q(n491) );
  INV3 U553 ( .A(add_x_4_n34), .Q(add_x_4_n33) );
  NOR21 U554 ( .A(n599), .B(n335), .Q(u_decode_control_o_con_aluop_5_) );
  INV3 U555 ( .A(u_decode_add_x_16_n148), .Q(u_decode_add_x_16_n147) );
  INV3 U556 ( .A(n374), .Q(n372) );
  INV3 U557 ( .A(u_decode_add_x_16_n169), .Q(u_decode_add_x_16_n168) );
  INV2 U558 ( .A(n329), .Q(n331) );
  NAND22 U559 ( .A(n364), .B(n251), .Q(n365) );
  NAND22 U560 ( .A(n344), .B(n343), .Q(n347) );
  INV3 U561 ( .A(add_x_4_n103), .Q(add_x_4_n102) );
  NAND22 U562 ( .A(n342), .B(n341), .Q(n348) );
  NOR21 U563 ( .A(n328), .B(n333), .Q(n329) );
  NOR21 U564 ( .A(n238), .B(n323), .Q(n339) );
  INV3 U565 ( .A(n558), .Q(n562) );
  XNR21 U566 ( .A(for_addr_rtW[0]), .B(n323), .Q(n351) );
  XNR21 U567 ( .A(for_addr_rtW[1]), .B(n238), .Q(n350) );
  INV2 U568 ( .A(add_x_1_n67), .Q(add_x_1_n66) );
  NAND22 U569 ( .A(n262), .B(n255), .Q(n333) );
  NOR21 U570 ( .A(n435), .B(n546), .Q(n436) );
  NOR21 U571 ( .A(n521), .B(n243), .Q(n522) );
  NOR21 U572 ( .A(n459), .B(n243), .Q(n460) );
  NOR21 U573 ( .A(n447), .B(n546), .Q(n448) );
  NOR21 U574 ( .A(n491), .B(n243), .Q(n492) );
  NOR22 U575 ( .A(n429), .B(n322), .Q(n430) );
  NAND21 U576 ( .A(n541), .B(instruction_address[25]), .Q(n404) );
  NAND21 U577 ( .A(n541), .B(instruction_address[28]), .Q(n389) );
  XNR21 U578 ( .A(n238), .B(for_addr_rtM[1]), .Q(n341) );
  NAND31 U579 ( .A(n514), .B(n512), .C(n513), .Q(n130) );
  AOI211 U580 ( .A(n319), .B(if_addr_j[2]), .C(n539), .Q(n545) );
  AOI211 U581 ( .A(n318), .B(if_addr_j[15]), .C(n460), .Q(n464) );
  NAND22 U582 ( .A(n318), .B(if_addr_j[31]), .Q(n250) );
  NAND22 U583 ( .A(n315), .B(id_data_jr[31]), .Q(n249) );
  AOI211 U584 ( .A(n319), .B(n237), .C(n430), .Q(n434) );
  AOI211 U585 ( .A(n319), .B(if_addr_j[17]), .C(n448), .Q(n452) );
  AOI211 U586 ( .A(id_data_jr[22]), .B(n316), .C(n310), .Q(n422) );
  AOI211 U587 ( .A(n318), .B(n238), .C(n436), .Q(n440) );
  AOI211 U588 ( .A(n318), .B(if_addr_j[21]), .C(n424), .Q(n428) );
  NAND22 U589 ( .A(n547), .B(instruction_address[1]), .Q(n550) );
  AOI212 U590 ( .A(n315), .B(id_data_jr[16]), .C(n455), .Q(n457) );
  NAND22 U591 ( .A(n309), .B(n313), .Q(n547) );
  NOR21 U592 ( .A(n317), .B(n311), .Q(n310) );
  INV6 U593 ( .A(if_con_b), .Q(n245) );
  MUX22 U594 ( .A(data_address[31]), .B(u_mem_pc8[31]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[31]) );
  MUX22 U595 ( .A(data_address[16]), .B(u_mem_pc8[16]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[16]) );
  MUX22 U596 ( .A(data_address[24]), .B(u_mem_pc8[24]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[24]) );
  MUX22 U597 ( .A(data_address[30]), .B(u_mem_pc8[30]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[30]) );
  NAND21 U598 ( .A(n552), .B(n313), .Q(n553) );
  OAI2111 U599 ( .A(n331), .B(n251), .C(n338), .D(n598), .Q(
        u_decode_control_o_con_aluop_3_) );
  MUX22 U600 ( .A(data_address[14]), .B(u_mem_pc8[14]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[14]) );
  NOR21 U601 ( .A(n292), .B(n313), .Q(n523) );
  INV2 U602 ( .A(u_decode_control_o_con_aluop_4_), .Q(n338) );
  NOR21 U603 ( .A(n287), .B(n313), .Q(n461) );
  NOR21 U604 ( .A(n296), .B(n313), .Q(n535) );
  MUX22 U605 ( .A(data_address[28]), .B(u_mem_pc8[28]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[28]) );
  NOR21 U606 ( .A(n284), .B(n313), .Q(n425) );
  NOR21 U607 ( .A(n291), .B(n313), .Q(n511) );
  MUX22 U608 ( .A(data_address[18]), .B(u_mem_pc8[18]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[18]) );
  NOR21 U609 ( .A(n274), .B(n313), .Q(n529) );
  NOR21 U610 ( .A(n286), .B(n313), .Q(n449) );
  NOR33 U611 ( .A(n541), .B(n376), .C(n377), .Q(n489) );
  NOR21 U612 ( .A(n285), .B(n313), .Q(n437) );
  MUX22 U613 ( .A(data_address[12]), .B(u_mem_pc8[12]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[12]) );
  INV2 U614 ( .A(n564), .Q(n571) );
  NOR21 U615 ( .A(n268), .B(n313), .Q(n419) );
  NOR21 U616 ( .A(n269), .B(n313), .Q(n431) );
  NOR21 U617 ( .A(n270), .B(n313), .Q(n455) );
  OAI211 U618 ( .A(n332), .B(n331), .C(n330), .Q(
        u_decode_control_o_con_aluop_2_) );
  NOR21 U619 ( .A(n288), .B(n313), .Q(n473) );
  NOR21 U620 ( .A(n290), .B(n313), .Q(n499) );
  NOR21 U621 ( .A(n289), .B(n313), .Q(n485) );
  NOR21 U622 ( .A(n273), .B(n313), .Q(n505) );
  NOR21 U623 ( .A(n271), .B(n313), .Q(n467) );
  NOR21 U624 ( .A(n272), .B(n313), .Q(n493) );
  NAND21 U625 ( .A(n572), .B(n240), .Q(n564) );
  MUX22 U626 ( .A(data_address[6]), .B(u_mem_pc8[6]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[6]) );
  AOI211 U627 ( .A(n365), .B(n312), .C(n333), .Q(
        u_decode_control_o_con_aluop_1_) );
  INV2 U628 ( .A(u_decode_control_o_con_aluop_0_), .Q(n599) );
  INV2 U629 ( .A(u_decode_add_x_16_n31), .Q(u_decode_add_x_16_n183) );
  INV2 U630 ( .A(u_decode_add_x_16_n54), .Q(u_decode_add_x_16_n52) );
  INV2 U631 ( .A(u_decode_add_x_16_n57), .Q(u_decode_add_x_16_n59) );
  NAND21 U632 ( .A(n366), .B(n332), .Q(n327) );
  INV2 U633 ( .A(u_decode_add_x_16_n88), .Q(u_decode_add_x_16_n193) );
  INV2 U634 ( .A(u_decode_add_x_16_n77), .Q(u_decode_add_x_16_n191) );
  INV2 U635 ( .A(u_decode_add_x_16_n140), .Q(u_decode_add_x_16_n138) );
  INV2 U636 ( .A(add_x_1_n86), .Q(add_x_1_n85) );
  INV2 U637 ( .A(u_decode_add_x_16_n172), .Q(u_decode_add_x_16_n209) );
  NAND22 U638 ( .A(id_data_instr[31]), .B(n558), .Q(n560) );
  INV1 U639 ( .A(u_fetch_jmux_i_addr_pc4_3_), .Q(n533) );
  NAND21 U640 ( .A(id_data_instr[28]), .B(id_data_instr[29]), .Q(n328) );
  INV2 U641 ( .A(mem_data_pc4[6]), .Q(add_x_1_n108) );
  IMUX21 U642 ( .A(n277), .B(if_addr_j[25]), .S(for_addr_rtW[2]), .Q(n591) );
  IMUX21 U643 ( .A(n280), .B(if_addr_j[26]), .S(for_addr_rtW[3]), .Q(n592) );
  IMUX21 U644 ( .A(n261), .B(if_addr_j[23]), .S(for_addr_rtW[0]), .Q(n593) );
  IMUX21 U645 ( .A(if_addr_j[21]), .B(n281), .S(for_addr_rtW[3]), .Q(n580) );
  IMUX21 U646 ( .A(if_addr_j[22]), .B(n311), .S(for_addr_rtW[4]), .Q(n581) );
  IMUX21 U647 ( .A(if_addr_j[23]), .B(n261), .S(for_addr_rtM[0]), .Q(n585) );
  NAND28 U648 ( .A(n245), .B(n376), .Q(n314) );
  AOI212 U649 ( .A(n315), .B(id_data_jr[20]), .C(n431), .Q(n433) );
  NOR23 U650 ( .A(n552), .B(if_con_b), .Q(n542) );
  AOI2112 U651 ( .A(n244), .B(u_fetch_jmux_i_addr_pc4_31_), .C(n247), .D(n248), 
        .Q(n246) );
  NOR24 U652 ( .A(n541), .B(n490), .Q(n551) );
  NOR24 U653 ( .A(n541), .B(n490), .Q(n321) );
  AOI212 U654 ( .A(n551), .B(if_addr_b[22]), .C(n419), .Q(n421) );
  AOI212 U655 ( .A(n316), .B(id_data_jr[13]), .C(n473), .Q(n475) );
  AOI212 U656 ( .A(n316), .B(id_data_jr[9]), .C(n499), .Q(n501) );
  AOI212 U657 ( .A(n316), .B(id_data_jr[5]), .C(n523), .Q(n525) );
  AOI212 U658 ( .A(n316), .B(id_data_jr[7]), .C(n511), .Q(n513) );
  AOI212 U659 ( .A(n316), .B(id_data_jr[11]), .C(n485), .Q(n487) );
  AOI212 U660 ( .A(n316), .B(id_data_jr[3]), .C(n535), .Q(n537) );
  AOI212 U661 ( .A(n316), .B(id_data_jr[19]), .C(n437), .Q(n439) );
  NAND33 U662 ( .A(n422), .B(n421), .C(n420), .Q(n115) );
  NAND33 U663 ( .A(n403), .B(n402), .C(n401), .Q(n111) );
  NAND22 U664 ( .A(n319), .B(if_addr_j[26]), .Q(n401) );
  OAI212 U665 ( .A(n299), .B(n554), .C(n379), .Q(n380) );
  OAI212 U666 ( .A(n302), .B(n554), .C(n394), .Q(n395) );
  OAI212 U667 ( .A(n304), .B(n554), .C(n404), .Q(n405) );
  OAI212 U668 ( .A(n305), .B(n554), .C(n409), .Q(n410) );
  OAI212 U669 ( .A(n306), .B(n554), .C(n414), .Q(n415) );
  NAND33 U670 ( .A(n418), .B(n417), .C(n416), .Q(n114) );
  NAND33 U671 ( .A(n413), .B(n412), .C(n411), .Q(n113) );
  NAND33 U672 ( .A(n398), .B(n397), .C(n396), .Q(n110) );
  NAND22 U673 ( .A(n318), .B(if_addr_j[27]), .Q(n396) );
  OAI212 U674 ( .A(n301), .B(n554), .C(n389), .Q(n390) );
  OAI212 U675 ( .A(n303), .B(n554), .C(n399), .Q(n400) );
  NAND33 U676 ( .A(n388), .B(n387), .C(n386), .Q(n108) );
  OAI212 U677 ( .A(n300), .B(n554), .C(n384), .Q(n385) );
  NAND33 U678 ( .A(n383), .B(n382), .C(n381), .Q(n107) );
  NOR21 U679 ( .A(n597), .B(u_decode_control_o_con_aluop_1_), .Q(n336) );
  INV3 U680 ( .A(u_decode_add_x_16_n178), .Q(u_decode_add_x_16_n177) );
  NAND22 U681 ( .A(n561), .B(n562), .Q(u_decode_n6) );
  INV3 U682 ( .A(mem_data_pc4[16]), .Q(add_x_1_n64) );
  INV3 U683 ( .A(add_x_1_n29), .Q(add_x_1_n28) );
  INV3 U684 ( .A(mem_data_pc4[24]), .Q(add_x_1_n26) );
  INV3 U685 ( .A(u_decode_add_x_16_n101), .Q(u_decode_add_x_16_n99) );
  INV3 U686 ( .A(mem_data_pc4[22]), .Q(add_x_1_n35) );
  NAND22 U687 ( .A(n597), .B(id_data_instr[31]), .Q(n561) );
  NOR31 U688 ( .A(id_data_instr[29]), .B(id_data_instr[30]), .C(n335), .Q(n597) );
  NAND22 U689 ( .A(n329), .B(id_data_instr[26]), .Q(n598) );
  NAND41 U690 ( .A(mem_con_Wregwrite), .B(n358), .C(n357), .D(n568), .Q(n361)
         );
  NAND31 U691 ( .A(n253), .B(id_data_instr[27]), .C(id_data_instr[26]), .Q(
        n335) );
  NOR21 U692 ( .A(if_addr_j[20]), .B(if_addr_j[21]), .Q(n340) );
  OAI2111 U693 ( .A(mem_addr_regdst[4]), .B(n279), .C(n574), .D(n575), .Q(n570) );
  NAND41 U694 ( .A(mem_con_Wregwrite), .B(n577), .C(n578), .D(n579), .Q(n569)
         );
  NAND22 U695 ( .A(n253), .B(id_data_instr[27]), .Q(n325) );
  NAND22 U696 ( .A(n257), .B(n253), .Q(n367) );
  NAND22 U697 ( .A(n318), .B(if_addr_j[23]), .Q(n416) );
  NOR20 U698 ( .A(n257), .B(id_data_instr[27]), .Q(n332) );
  NAND22 U699 ( .A(n315), .B(id_data_jr[0]), .Q(n556) );
  NAND22 U700 ( .A(n542), .B(u_fetch_jmux_i_addr_pc4_22_), .Q(n420) );
  NAND22 U701 ( .A(n316), .B(id_data_jr[1]), .Q(n549) );
  NAND22 U702 ( .A(n316), .B(id_data_jr[30]), .Q(n382) );
  NAND22 U703 ( .A(n316), .B(id_data_jr[28]), .Q(n392) );
  NAND22 U704 ( .A(n316), .B(id_data_jr[26]), .Q(n402) );
  NAND22 U705 ( .A(n315), .B(id_data_jr[27]), .Q(n397) );
  NAND22 U706 ( .A(n319), .B(if_addr_j[24]), .Q(n411) );
  NAND22 U707 ( .A(n316), .B(id_data_jr[24]), .Q(n412) );
  NAND22 U708 ( .A(n315), .B(id_data_jr[23]), .Q(n417) );
  NAND22 U709 ( .A(n315), .B(id_data_jr[29]), .Q(n387) );
  AOI211 U710 ( .A(n318), .B(if_addr_j[5]), .C(n522), .Q(n526) );
  AOI211 U711 ( .A(n315), .B(id_data_jr[6]), .C(n517), .Q(n519) );
  AOI211 U712 ( .A(n319), .B(if_addr_j[6]), .C(n516), .Q(n520) );
  AOI211 U713 ( .A(n315), .B(id_data_jr[10]), .C(n493), .Q(n495) );
  AOI211 U714 ( .A(n315), .B(id_data_jr[4]), .C(n529), .Q(n531) );
  AOI211 U715 ( .A(n319), .B(if_addr_j[4]), .C(n528), .Q(n532) );
  AOI211 U716 ( .A(n315), .B(id_data_jr[14]), .C(n467), .Q(n469) );
  AOI211 U717 ( .A(n315), .B(id_data_jr[18]), .C(n443), .Q(n445) );
  AOI211 U718 ( .A(n318), .B(if_addr_j[7]), .C(n510), .Q(n514) );
  AOI211 U719 ( .A(n315), .B(id_data_jr[12]), .C(n479), .Q(n481) );
  AOI211 U720 ( .A(n315), .B(id_data_jr[8]), .C(n505), .Q(n507) );
  NOR24 U721 ( .A(n541), .B(n490), .Q(n320) );
  OAI310 U722 ( .A(id_data_instr[28]), .B(n323), .C(n327), .D(n326), .Q(
        u_decode_jbcon_o_con_bop[0]) );
  NAND30 U723 ( .A(n366), .B(id_data_instr[28]), .C(n257), .Q(n326) );
  NAND22 U724 ( .A(n319), .B(if_addr_j[30]), .Q(n381) );
  NAND22 U725 ( .A(n319), .B(if_addr_j[28]), .Q(n391) );
  NAND22 U726 ( .A(n318), .B(if_addr_j[29]), .Q(n386) );
  AOI211 U727 ( .A(n338), .B(n337), .C(n256), .Q(u_decode_n3) );
  NAND22 U728 ( .A(n561), .B(n560), .Q(u_decode_control_o_con_memtoreg) );
  NOR21 U729 ( .A(n354), .B(n239), .Q(n359) );
  NAND31 U730 ( .A(n567), .B(n356), .C(n355), .Q(n362) );
  MUX21 U731 ( .A(mem_data_alures[4]), .B(wb_data_memout[4]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[4]) );
  MUX21 U732 ( .A(mem_data_alures[5]), .B(wb_data_memout[5]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[5]) );
  MUX21 U733 ( .A(mem_data_alures[10]), .B(wb_data_memout[10]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[10]) );
  MUX21 U734 ( .A(mem_data_alures[9]), .B(wb_data_memout[9]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[9]) );
  MUX21 U735 ( .A(mem_data_alures[20]), .B(wb_data_memout[20]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[20]) );
  MUX21 U736 ( .A(mem_data_alures[1]), .B(wb_data_memout[1]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[1]) );
  MUX21 U737 ( .A(mem_data_alures[15]), .B(wb_data_memout[15]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[15]) );
  MUX21 U738 ( .A(mem_data_alures[7]), .B(wb_data_memout[7]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[7]) );
  MUX22 U739 ( .A(mem_data_alures[27]), .B(wb_data_memout[27]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[27]) );
  MUX22 U740 ( .A(mem_data_alures[26]), .B(wb_data_memout[26]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[26]) );
  MUX22 U741 ( .A(mem_data_alures[14]), .B(wb_data_memout[14]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[14]) );
  MUX22 U742 ( .A(mem_data_alures[24]), .B(wb_data_memout[24]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[24]) );
  MUX22 U743 ( .A(mem_data_alures[28]), .B(wb_data_memout[28]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[28]) );
  MUX22 U744 ( .A(mem_data_alures[22]), .B(wb_data_memout[22]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[22]) );
  MUX22 U745 ( .A(mem_data_alures[29]), .B(wb_data_memout[29]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[29]) );
  MUX22 U746 ( .A(mem_data_alures[30]), .B(wb_data_memout[30]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[30]) );
  MUX22 U747 ( .A(mem_data_alures[25]), .B(wb_data_memout[25]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[25]) );
  OAI2111 U748 ( .A(for_addr_rtW[4]), .B(n279), .C(for_FWmemread), .D(n595), 
        .Q(n594) );
  AOI211 U749 ( .A(for_addr_rtW[4]), .B(n279), .C(n596), .Q(n595) );
  NAND31 U750 ( .A(n557), .B(n556), .C(n555), .Q(n137) );
  NAND31 U751 ( .A(n554), .B(instruction_address[0]), .C(n553), .Q(n555) );
  NAND22 U752 ( .A(n320), .B(ex_data_pc4[0]), .Q(n557) );
  NAND22 U753 ( .A(n315), .B(id_data_jr[2]), .Q(n543) );
  NAND22 U754 ( .A(n551), .B(ex_data_pc4[1]), .Q(n548) );
  NAND22 U755 ( .A(n321), .B(if_addr_b[21]), .Q(n426) );
  INV3 U756 ( .A(add_x_4_n1), .Q(add_x_4_n116) );
  NAND22 U757 ( .A(n321), .B(if_addr_b[3]), .Q(n536) );
  NAND22 U758 ( .A(n551), .B(if_addr_b[20]), .Q(n432) );
  NAND22 U759 ( .A(n320), .B(if_addr_b[13]), .Q(n474) );
  NAND22 U760 ( .A(n321), .B(if_addr_b[15]), .Q(n462) );
  NAND22 U761 ( .A(n321), .B(if_addr_b[9]), .Q(n500) );
  NAND22 U762 ( .A(n320), .B(if_addr_b[5]), .Q(n524) );
  NAND22 U763 ( .A(n321), .B(if_addr_b[6]), .Q(n518) );
  NOR21 U764 ( .A(n527), .B(n546), .Q(n528) );
  NAND22 U765 ( .A(n320), .B(if_addr_b[19]), .Q(n438) );
  NAND22 U766 ( .A(n551), .B(if_addr_b[14]), .Q(n468) );
  NAND22 U767 ( .A(n321), .B(if_addr_b[18]), .Q(n444) );
  NAND22 U768 ( .A(n551), .B(if_addr_b[17]), .Q(n450) );
  NAND22 U769 ( .A(n320), .B(if_addr_b[7]), .Q(n512) );
  NOR21 U770 ( .A(n509), .B(n243), .Q(n510) );
  NAND22 U771 ( .A(n551), .B(if_addr_b[11]), .Q(n486) );
  NAND22 U772 ( .A(n321), .B(if_addr_b[12]), .Q(n480) );
  NAND22 U773 ( .A(n551), .B(if_addr_b[8]), .Q(n506) );
  NAND22 U774 ( .A(n320), .B(if_addr_b[16]), .Q(n456) );
  MUX21 U775 ( .A(read_data[12]), .B(wb_data_memout[12]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[12]) );
  MUX21 U776 ( .A(read_data[4]), .B(wb_data_memout[4]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[4]) );
  MUX21 U777 ( .A(read_data[8]), .B(wb_data_memout[8]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[8]) );
  MUX21 U778 ( .A(read_data[30]), .B(wb_data_memout[30]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[30]) );
  MUX21 U779 ( .A(read_data[10]), .B(wb_data_memout[10]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[10]) );
  MUX21 U780 ( .A(read_data[9]), .B(wb_data_memout[9]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[9]) );
  MUX21 U781 ( .A(read_data[7]), .B(wb_data_memout[7]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[7]) );
  MUX21 U782 ( .A(read_data[26]), .B(wb_data_memout[26]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[26]) );
  MUX21 U783 ( .A(read_data[2]), .B(wb_data_memout[2]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[2]) );
  MUX21 U784 ( .A(read_data[1]), .B(wb_data_memout[1]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[1]) );
  MUX21 U785 ( .A(read_data[0]), .B(wb_data_memout[0]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[0]) );
  MUX21 U786 ( .A(read_data[28]), .B(wb_data_memout[28]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[28]) );
  MUX21 U787 ( .A(read_data[11]), .B(wb_data_memout[11]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[11]) );
  MUX21 U788 ( .A(read_data[6]), .B(wb_data_memout[6]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[6]) );
  MUX21 U789 ( .A(read_data[3]), .B(wb_data_memout[3]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[3]) );
  MUX21 U790 ( .A(read_data[5]), .B(wb_data_memout[5]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[5]) );
  MUX21 U791 ( .A(read_data[15]), .B(wb_data_memout[15]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[15]) );
  MUX21 U792 ( .A(read_data[14]), .B(wb_data_memout[14]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[14]) );
  MUX21 U793 ( .A(read_data[13]), .B(wb_data_memout[13]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[13]) );
  MUX21 U794 ( .A(read_data[20]), .B(wb_data_memout[20]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[20]) );
  MUX21 U795 ( .A(read_data[21]), .B(wb_data_memout[21]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[21]) );
  MUX21 U796 ( .A(read_data[22]), .B(wb_data_memout[22]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[22]) );
  MUX21 U797 ( .A(read_data[17]), .B(wb_data_memout[17]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[17]) );
  MUX21 U798 ( .A(read_data[24]), .B(wb_data_memout[24]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[24]) );
  MUX21 U799 ( .A(read_data[25]), .B(wb_data_memout[25]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[25]) );
  MUX21 U800 ( .A(read_data[27]), .B(wb_data_memout[27]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[27]) );
  MUX21 U801 ( .A(read_data[29]), .B(wb_data_memout[29]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[29]) );
  MUX21 U802 ( .A(read_data[31]), .B(wb_data_memout[31]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[31]) );
  MUX21 U803 ( .A(read_data[23]), .B(wb_data_memout[23]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[23]) );
  MUX21 U804 ( .A(read_data[16]), .B(wb_data_memout[16]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[16]) );
  MUX21 U805 ( .A(read_data[19]), .B(wb_data_memout[19]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[19]) );
  MUX21 U806 ( .A(read_data[18]), .B(wb_data_memout[18]), .S(n239), .Q(
        u_decode_fbmemmux_o_data_fmem[18]) );
  AOI2110 U807 ( .A(id_data_instr[28]), .B(n251), .C(n257), .D(n369), .Q(
        u_decode_jbcon_o_con_bop[2]) );
  OAI220 U808 ( .A(n326), .B(n251), .C(n327), .D(n566), .Q(
        u_decode_jbcon_o_con_bop[1]) );
  MUX21 U809 ( .A(data_address[22]), .B(u_mem_pc8[22]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[22]) );
  AOI310 U810 ( .A(n559), .B(n558), .C(n253), .D(
        u_decode_control_o_con_memtoreg), .Q(n337) );
  XNR21 U811 ( .A(n323), .B(mem_addr_regdst[0]), .Q(n357) );
  XNR21 U812 ( .A(if_addr_j[22]), .B(mem_addr_regdst[4]), .Q(n355) );
  XNR21 U813 ( .A(n237), .B(mem_addr_regdst[2]), .Q(n356) );
  XNR21 U814 ( .A(if_addr_j[22]), .B(for_addr_rtM[4]), .Q(n345) );
  XNR21 U815 ( .A(n323), .B(for_addr_rtM[0]), .Q(n343) );
  XNR21 U816 ( .A(if_addr_j[21]), .B(for_addr_rtM[3]), .Q(n344) );
  XNR21 U817 ( .A(if_addr_j[20]), .B(for_addr_rtM[2]), .Q(n342) );
  XNR21 U818 ( .A(for_addr_rtW[2]), .B(n237), .Q(n349) );
  INV3 U819 ( .A(u_decode_add_x_16_n39), .Q(u_decode_add_x_16_n37) );
  INV3 U820 ( .A(u_decode_add_x_16_n53), .Q(u_decode_add_x_16_n51) );
  INV3 U821 ( .A(u_decode_add_x_16_n56), .Q(u_decode_add_x_16_n58) );
  NAND20 U822 ( .A(n541), .B(instruction_address[30]), .Q(n379) );
  NAND20 U823 ( .A(n541), .B(instruction_address[26]), .Q(n399) );
  NAND20 U824 ( .A(n541), .B(instruction_address[24]), .Q(n409) );
  NAND20 U825 ( .A(n541), .B(instruction_address[23]), .Q(n414) );
  NOR20 U826 ( .A(n295), .B(n313), .Q(n517) );
  NOR20 U827 ( .A(n293), .B(n313), .Q(n443) );
  NOR20 U828 ( .A(n294), .B(n313), .Q(n479) );
  LOGIC0 U829 ( .Q(n308) );
  NAND20 U830 ( .A(id_data_instr[26]), .B(id_data_instr[27]), .Q(n559) );
  NOR20 U831 ( .A(id_data_instr[28]), .B(n323), .Q(n566) );
  IMUX20 U832 ( .A(n238), .B(n282), .S(mem_addr_regdst[1]), .Q(n568) );
  IMUX20 U833 ( .A(if_addr_j[21]), .B(n281), .S(mem_addr_regdst[3]), .Q(n567)
         );
  OAI210 U834 ( .A(mem_addr_regdst[4]), .B(n576), .C(n279), .Q(n575) );
  NOR40 U835 ( .A(if_addr_j[26]), .B(mem_addr_regdst[2]), .C(
        mem_addr_regdst[1]), .D(mem_addr_regdst[0]), .Q(n576) );
  IMUX20 U836 ( .A(if_addr_j[23]), .B(n261), .S(mem_addr_regdst[0]), .Q(n574)
         );
  IMUX20 U837 ( .A(if_addr_j[25]), .B(n277), .S(mem_addr_regdst[2]), .Q(n579)
         );
  IMUX20 U838 ( .A(if_addr_j[26]), .B(n280), .S(mem_addr_regdst[3]), .Q(n578)
         );
  IMUX20 U839 ( .A(if_addr_j[24]), .B(n260), .S(mem_addr_regdst[1]), .Q(n577)
         );
  MUX21 U840 ( .A(wb_data_memout[9]), .B(read_data[9]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[9]) );
  MUX21 U841 ( .A(wb_data_memout[8]), .B(read_data[8]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[8]) );
  MUX21 U842 ( .A(wb_data_memout[7]), .B(read_data[7]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[7]) );
  MUX21 U843 ( .A(wb_data_memout[6]), .B(read_data[6]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[6]) );
  MUX21 U844 ( .A(wb_data_memout[5]), .B(read_data[5]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[5]) );
  MUX21 U845 ( .A(wb_data_memout[4]), .B(read_data[4]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[4]) );
  MUX21 U846 ( .A(wb_data_memout[3]), .B(read_data[3]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[3]) );
  MUX21 U847 ( .A(wb_data_memout[31]), .B(read_data[31]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[31]) );
  MUX21 U848 ( .A(wb_data_memout[30]), .B(read_data[30]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[30]) );
  MUX21 U849 ( .A(wb_data_memout[2]), .B(read_data[2]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[2]) );
  MUX21 U850 ( .A(wb_data_memout[29]), .B(read_data[29]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[29]) );
  MUX21 U851 ( .A(wb_data_memout[28]), .B(read_data[28]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[28]) );
  MUX21 U852 ( .A(wb_data_memout[27]), .B(read_data[27]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[27]) );
  MUX21 U853 ( .A(wb_data_memout[26]), .B(read_data[26]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[26]) );
  MUX21 U854 ( .A(wb_data_memout[25]), .B(read_data[25]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[25]) );
  MUX21 U855 ( .A(wb_data_memout[24]), .B(read_data[24]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[24]) );
  MUX21 U856 ( .A(wb_data_memout[23]), .B(read_data[23]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[23]) );
  MUX21 U857 ( .A(wb_data_memout[22]), .B(read_data[22]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[22]) );
  MUX21 U858 ( .A(wb_data_memout[21]), .B(read_data[21]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[21]) );
  MUX21 U859 ( .A(wb_data_memout[20]), .B(read_data[20]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[20]) );
  MUX21 U860 ( .A(wb_data_memout[1]), .B(read_data[1]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[1]) );
  MUX21 U861 ( .A(wb_data_memout[19]), .B(read_data[19]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[19]) );
  MUX21 U862 ( .A(wb_data_memout[18]), .B(read_data[18]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[18]) );
  MUX21 U863 ( .A(wb_data_memout[17]), .B(read_data[17]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[17]) );
  MUX21 U864 ( .A(wb_data_memout[16]), .B(read_data[16]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[16]) );
  MUX21 U865 ( .A(wb_data_memout[15]), .B(read_data[15]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[15]) );
  MUX21 U866 ( .A(wb_data_memout[14]), .B(read_data[14]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[14]) );
  MUX21 U867 ( .A(wb_data_memout[13]), .B(read_data[13]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[13]) );
  MUX21 U868 ( .A(wb_data_memout[12]), .B(read_data[12]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[12]) );
  MUX21 U869 ( .A(wb_data_memout[11]), .B(read_data[11]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[11]) );
  MUX21 U870 ( .A(wb_data_memout[10]), .B(read_data[10]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[10]) );
  MUX21 U871 ( .A(wb_data_memout[0]), .B(read_data[0]), .S(n240), .Q(
        u_decode_famemmux_o_data_fmem[0]) );
  IMUX20 U872 ( .A(n277), .B(if_addr_j[25]), .S(for_addr_rtM[2]), .Q(n589) );
  IMUX20 U873 ( .A(n279), .B(if_addr_j[27]), .S(for_addr_rtM[4]), .Q(n587) );
  IMUX20 U874 ( .A(n280), .B(if_addr_j[26]), .S(for_addr_rtM[3]), .Q(n586) );
  IMUX20 U875 ( .A(n260), .B(if_addr_j[24]), .S(for_addr_rtW[1]), .Q(n596) );
  OAI210 U876 ( .A(n251), .B(n598), .C(n561), .Q(
        u_decode_control_o_con_memread) );
endmodule

