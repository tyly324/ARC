// Verilog simulation library for c35_IOLIB_ANA_3M
// Owner: austriamicrosystems AG  HIT-Kit: Digital
module APRIO500P (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module APRIO50P (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module APRIOWP (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module APRIO500SP (PAD,Z,Z0);
  inout PAD ;
  inout Z ;
  inout Z0 ;
endmodule
module AGNDALLP (VSSA);
  input VSSA ;
endmodule
module AVDDALLP (VDDA);
  input VDDA ;
endmodule
module APRIOP (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module APRIO1K5P (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
module APRIO200P (Z,PAD);
  inout Z ;
  inout PAD ;
endmodule
