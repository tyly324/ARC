module W_loadmux4