
module F_jumpmux ( i_addr_j, i_addr_jr, i_addr_pc4, i_con_jump, o_addr_jumpmux
 );
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [31:0] i_addr_pc4;
  input [1:0] i_con_jump;
  output [31:0] o_addr_jumpmux;
  wire   n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n24,
         n25, n46, n47, n68, n69, n1, n2, n3, n6, n7, n20, n21, n22, n23, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97;

  OAI2111 U1 ( .A(n1), .B(n58), .C(n57), .D(n56), .Q(o_addr_jumpmux[16]) );
  OAI2111 U2 ( .A(n1), .B(n52), .C(n51), .D(n50), .Q(o_addr_jumpmux[14]) );
  OAI2111 U3 ( .A(n1), .B(n31), .C(n78), .D(n77), .Q(o_addr_jumpmux[25]) );
  OAI2111 U4 ( .A(n1), .B(n55), .C(n54), .D(n53), .Q(o_addr_jumpmux[15]) );
  OAI2111 U5 ( .A(n1), .B(n85), .C(n84), .D(n83), .Q(o_addr_jumpmux[28]) );
  OAI2111 U6 ( .A(n95), .B(n88), .C(n87), .D(n86), .Q(o_addr_jumpmux[29]) );
  OAI2111 U7 ( .A(n1), .B(n29), .C(n74), .D(n73), .Q(o_addr_jumpmux[23]) );
  OAI2111 U8 ( .A(n1), .B(n33), .C(n82), .D(n81), .Q(o_addr_jumpmux[27]) );
  OAI2111 U9 ( .A(n1), .B(n94), .C(n93), .D(n92), .Q(o_addr_jumpmux[31]) );
  BUF2 U10 ( .A(n97), .Q(n7) );
  INV6 U11 ( .A(n37), .Q(n96) );
  NAND22 U12 ( .A(n95), .B(n36), .Q(n37) );
  OAI2111 U13 ( .A(n95), .B(n40), .C(n39), .D(n38), .Q(o_addr_jumpmux[10]) );
  OAI2111 U14 ( .A(n1), .B(n21), .C(n60), .D(n59), .Q(o_addr_jumpmux[17]) );
  OAI2111 U15 ( .A(n1), .B(n32), .C(n80), .D(n79), .Q(o_addr_jumpmux[26]) );
  INV3 U16 ( .A(n95), .Q(n2) );
  INV1 U17 ( .A(n95), .Q(n3) );
  NAND22 U18 ( .A(i_addr_pc4[15]), .B(n96), .Q(n53) );
  OAI2111 U19 ( .A(n1), .B(n43), .C(n42), .D(n41), .Q(o_addr_jumpmux[11]) );
  NAND22 U20 ( .A(i_addr_pc4[11]), .B(n96), .Q(n41) );
  NAND22 U21 ( .A(n35), .B(i_con_jump[1]), .Q(n36) );
  INV3 U22 ( .A(n36), .Q(n97) );
  AOI221 U23 ( .A(i_addr_pc4[7]), .B(n96), .C(i_addr_jr[7]), .D(n7), .Q(n10)
         );
  NAND20 U24 ( .A(i_addr_pc4[16]), .B(n96), .Q(n56) );
  NAND20 U25 ( .A(i_addr_pc4[19]), .B(n96), .Q(n63) );
  INV0 U26 ( .A(i_addr_j[26]), .Q(n32) );
  INV0 U27 ( .A(i_addr_j[12]), .Q(n45) );
  INV0 U28 ( .A(i_addr_j[27]), .Q(n33) );
  NAND20 U29 ( .A(i_addr_pc4[14]), .B(n96), .Q(n50) );
  NAND20 U30 ( .A(i_addr_pc4[17]), .B(n96), .Q(n59) );
  NAND20 U31 ( .A(i_addr_pc4[18]), .B(n96), .Q(n61) );
  AOI220 U32 ( .A(i_addr_pc4[5]), .B(n96), .C(i_addr_jr[5]), .D(n7), .Q(n14)
         );
  AOI220 U33 ( .A(i_addr_pc4[6]), .B(n96), .C(i_addr_jr[6]), .D(n7), .Q(n12)
         );
  AOI220 U34 ( .A(i_addr_pc4[8]), .B(n96), .C(i_addr_jr[8]), .D(n7), .Q(n8) );
  AOI220 U35 ( .A(i_addr_jr[12]), .B(n20), .C(i_addr_pc4[12]), .D(n96), .Q(n44) );
  AOI220 U36 ( .A(i_addr_jr[13]), .B(n20), .C(i_addr_pc4[13]), .D(n96), .Q(n48) );
  NAND20 U37 ( .A(i_addr_j[5]), .B(n3), .Q(n15) );
  NAND20 U38 ( .A(i_addr_j[6]), .B(n3), .Q(n13) );
  NAND20 U39 ( .A(i_addr_j[7]), .B(n3), .Q(n11) );
  NAND20 U40 ( .A(i_addr_j[8]), .B(n3), .Q(n9) );
  NAND20 U41 ( .A(i_addr_j[4]), .B(n3), .Q(n17) );
  NAND20 U42 ( .A(i_addr_j[3]), .B(n3), .Q(n19) );
  NAND20 U43 ( .A(i_addr_j[2]), .B(n2), .Q(n25) );
  INV0 U44 ( .A(i_addr_j[20]), .Q(n26) );
  INV0 U45 ( .A(i_addr_j[21]), .Q(n27) );
  INV0 U46 ( .A(i_addr_j[22]), .Q(n28) );
  INV0 U47 ( .A(i_addr_j[17]), .Q(n21) );
  BUF2 U48 ( .A(n97), .Q(n6) );
  BUF2 U49 ( .A(n97), .Q(n20) );
  INV3 U50 ( .A(n2), .Q(n1) );
  NAND22 U51 ( .A(i_addr_pc4[10]), .B(n96), .Q(n38) );
  NAND22 U52 ( .A(i_addr_pc4[21]), .B(n96), .Q(n67) );
  NAND22 U53 ( .A(i_addr_pc4[22]), .B(n96), .Q(n71) );
  NAND22 U54 ( .A(i_addr_pc4[25]), .B(n96), .Q(n77) );
  NAND22 U55 ( .A(i_addr_pc4[26]), .B(n96), .Q(n79) );
  NAND22 U56 ( .A(i_con_jump[0]), .B(n34), .Q(n95) );
  INV3 U57 ( .A(i_con_jump[1]), .Q(n34) );
  AOI221 U58 ( .A(i_addr_pc4[9]), .B(n96), .C(i_addr_jr[9]), .D(n7), .Q(n4) );
  AOI221 U59 ( .A(i_addr_pc4[4]), .B(n96), .C(i_addr_jr[4]), .D(n7), .Q(n16)
         );
  AOI221 U60 ( .A(i_addr_pc4[2]), .B(n96), .C(i_addr_jr[2]), .D(n20), .Q(n24)
         );
  AOI221 U61 ( .A(i_addr_pc4[3]), .B(n96), .C(i_addr_jr[3]), .D(n20), .Q(n18)
         );
  NAND22 U62 ( .A(i_addr_pc4[20]), .B(n96), .Q(n65) );
  NAND22 U63 ( .A(i_addr_pc4[23]), .B(n96), .Q(n73) );
  NAND22 U64 ( .A(i_addr_pc4[24]), .B(n96), .Q(n75) );
  NAND22 U65 ( .A(i_addr_pc4[27]), .B(n96), .Q(n81) );
  NAND22 U66 ( .A(i_addr_pc4[28]), .B(n96), .Q(n83) );
  NAND22 U67 ( .A(i_addr_pc4[29]), .B(n96), .Q(n86) );
  NAND22 U68 ( .A(i_addr_pc4[30]), .B(n96), .Q(n89) );
  NAND22 U69 ( .A(i_addr_pc4[31]), .B(n96), .Q(n92) );
  NAND22 U70 ( .A(i_addr_jr[10]), .B(n6), .Q(n39) );
  NAND22 U71 ( .A(i_addr_jr[20]), .B(n6), .Q(n66) );
  NAND22 U72 ( .A(i_addr_jr[21]), .B(n6), .Q(n70) );
  NAND22 U73 ( .A(i_addr_jr[22]), .B(n6), .Q(n72) );
  NAND22 U74 ( .A(i_addr_jr[23]), .B(n6), .Q(n74) );
  NAND22 U75 ( .A(i_addr_jr[24]), .B(n6), .Q(n76) );
  NAND22 U76 ( .A(i_addr_jr[25]), .B(n6), .Q(n78) );
  NAND22 U77 ( .A(i_addr_jr[26]), .B(n6), .Q(n80) );
  NAND22 U78 ( .A(i_addr_jr[27]), .B(n6), .Q(n82) );
  NAND22 U79 ( .A(i_addr_jr[28]), .B(n6), .Q(n84) );
  NAND22 U80 ( .A(i_addr_jr[29]), .B(n6), .Q(n87) );
  NAND22 U81 ( .A(i_addr_jr[30]), .B(n6), .Q(n90) );
  NAND22 U82 ( .A(i_addr_jr[31]), .B(n6), .Q(n93) );
  NAND22 U83 ( .A(i_addr_jr[11]), .B(n7), .Q(n42) );
  NAND22 U84 ( .A(i_addr_jr[14]), .B(n7), .Q(n51) );
  NAND22 U85 ( .A(i_addr_jr[15]), .B(n7), .Q(n54) );
  NAND22 U86 ( .A(i_addr_jr[16]), .B(n7), .Q(n57) );
  NAND22 U87 ( .A(i_addr_jr[17]), .B(n7), .Q(n60) );
  NAND22 U88 ( .A(i_addr_jr[18]), .B(n7), .Q(n62) );
  NAND22 U89 ( .A(i_addr_jr[19]), .B(n7), .Q(n64) );
  INV3 U90 ( .A(i_addr_j[18]), .Q(n22) );
  INV3 U91 ( .A(i_addr_j[23]), .Q(n29) );
  AOI221 U92 ( .A(i_addr_pc4[0]), .B(n96), .C(i_addr_jr[0]), .D(n7), .Q(n68)
         );
  AOI221 U93 ( .A(i_addr_pc4[1]), .B(n96), .C(i_addr_jr[1]), .D(n20), .Q(n46)
         );
  NAND22 U94 ( .A(n68), .B(n69), .Q(o_addr_jumpmux[0]) );
  NAND22 U95 ( .A(i_addr_j[0]), .B(n3), .Q(n69) );
  NAND22 U96 ( .A(n46), .B(n47), .Q(o_addr_jumpmux[1]) );
  NAND22 U97 ( .A(i_addr_j[1]), .B(n3), .Q(n47) );
  NAND22 U98 ( .A(n24), .B(n25), .Q(o_addr_jumpmux[2]) );
  NAND22 U99 ( .A(n18), .B(n19), .Q(o_addr_jumpmux[3]) );
  NAND22 U100 ( .A(n4), .B(n5), .Q(o_addr_jumpmux[9]) );
  NAND22 U101 ( .A(i_addr_j[9]), .B(n2), .Q(n5) );
  NAND22 U102 ( .A(n16), .B(n17), .Q(o_addr_jumpmux[4]) );
  NAND22 U103 ( .A(n14), .B(n15), .Q(o_addr_jumpmux[5]) );
  NAND22 U104 ( .A(n12), .B(n13), .Q(o_addr_jumpmux[6]) );
  NAND22 U105 ( .A(n10), .B(n11), .Q(o_addr_jumpmux[7]) );
  NAND22 U106 ( .A(n8), .B(n9), .Q(o_addr_jumpmux[8]) );
  INV3 U107 ( .A(i_addr_j[25]), .Q(n31) );
  INV3 U108 ( .A(i_addr_j[16]), .Q(n58) );
  INV3 U109 ( .A(i_addr_j[19]), .Q(n23) );
  INV3 U110 ( .A(i_addr_j[24]), .Q(n30) );
  INV3 U111 ( .A(i_addr_j[15]), .Q(n55) );
  INV3 U112 ( .A(i_addr_j[11]), .Q(n43) );
  INV3 U113 ( .A(i_addr_j[13]), .Q(n49) );
  INV3 U114 ( .A(i_addr_j[14]), .Q(n52) );
  INV3 U115 ( .A(i_addr_j[28]), .Q(n85) );
  INV3 U116 ( .A(i_addr_j[29]), .Q(n88) );
  INV3 U117 ( .A(i_addr_j[30]), .Q(n91) );
  INV3 U118 ( .A(i_addr_j[10]), .Q(n40) );
  INV3 U119 ( .A(i_addr_j[31]), .Q(n94) );
  CLKIN3 U120 ( .A(i_con_jump[0]), .Q(n35) );
  OAI212 U121 ( .A(n1), .B(n45), .C(n44), .Q(o_addr_jumpmux[12]) );
  OAI212 U122 ( .A(n1), .B(n49), .C(n48), .Q(o_addr_jumpmux[13]) );
  OAI2112 U123 ( .A(n1), .B(n22), .C(n62), .D(n61), .Q(o_addr_jumpmux[18]) );
  OAI2112 U124 ( .A(n1), .B(n23), .C(n64), .D(n63), .Q(o_addr_jumpmux[19]) );
  OAI2112 U125 ( .A(n1), .B(n26), .C(n66), .D(n65), .Q(o_addr_jumpmux[20]) );
  OAI2112 U126 ( .A(n1), .B(n27), .C(n70), .D(n67), .Q(o_addr_jumpmux[21]) );
  OAI2112 U127 ( .A(n1), .B(n28), .C(n72), .D(n71), .Q(o_addr_jumpmux[22]) );
  OAI2112 U128 ( .A(n1), .B(n30), .C(n76), .D(n75), .Q(o_addr_jumpmux[24]) );
  OAI2112 U129 ( .A(n95), .B(n91), .C(n90), .D(n89), .Q(o_addr_jumpmux[30]) );
endmodule


module F_branchmux ( i_addr_jumpmux, i_addr_b, i_con_ifbranch, o_addr_nextpc
 );
  input [31:0] i_addr_jumpmux;
  input [31:0] i_addr_b;
  output [31:0] o_addr_nextpc;
  input i_con_ifbranch;
  wire   n35, n36, n37, n38, n39, n40, n41, n44, n55, n66, n1, n2, n3;

  CLKIN3 U1 ( .A(n39), .Q(o_addr_nextpc[5]) );
  CLKIN3 U2 ( .A(n38), .Q(o_addr_nextpc[6]) );
  CLKIN3 U3 ( .A(n37), .Q(o_addr_nextpc[7]) );
  CLKIN3 U4 ( .A(n36), .Q(o_addr_nextpc[8]) );
  CLKIN3 U5 ( .A(n40), .Q(o_addr_nextpc[4]) );
  CLKIN3 U6 ( .A(n66), .Q(o_addr_nextpc[0]) );
  CLKIN3 U7 ( .A(n41), .Q(o_addr_nextpc[3]) );
  CLKIN3 U8 ( .A(n44), .Q(o_addr_nextpc[2]) );
  CLKIN3 U9 ( .A(n55), .Q(o_addr_nextpc[1]) );
  CLKIN3 U10 ( .A(n35), .Q(o_addr_nextpc[9]) );
  INV3 U11 ( .A(n3), .Q(n2) );
  INV3 U12 ( .A(n3), .Q(n1) );
  INV3 U13 ( .A(i_con_ifbranch), .Q(n3) );
  MUX22 U14 ( .A(i_addr_jumpmux[11]), .B(i_addr_b[11]), .S(n1), .Q(
        o_addr_nextpc[11]) );
  MUX22 U15 ( .A(i_addr_jumpmux[14]), .B(i_addr_b[14]), .S(n1), .Q(
        o_addr_nextpc[14]) );
  MUX22 U16 ( .A(i_addr_jumpmux[15]), .B(i_addr_b[15]), .S(n1), .Q(
        o_addr_nextpc[15]) );
  MUX22 U17 ( .A(i_addr_jumpmux[19]), .B(i_addr_b[19]), .S(n1), .Q(
        o_addr_nextpc[19]) );
  MUX22 U18 ( .A(i_addr_jumpmux[22]), .B(i_addr_b[22]), .S(n2), .Q(
        o_addr_nextpc[22]) );
  MUX22 U19 ( .A(i_addr_jumpmux[23]), .B(i_addr_b[23]), .S(n2), .Q(
        o_addr_nextpc[23]) );
  MUX22 U20 ( .A(i_addr_jumpmux[24]), .B(i_addr_b[24]), .S(n2), .Q(
        o_addr_nextpc[24]) );
  MUX22 U21 ( .A(i_addr_jumpmux[25]), .B(i_addr_b[25]), .S(n2), .Q(
        o_addr_nextpc[25]) );
  MUX22 U22 ( .A(i_addr_jumpmux[26]), .B(i_addr_b[26]), .S(n2), .Q(
        o_addr_nextpc[26]) );
  MUX22 U23 ( .A(i_addr_jumpmux[27]), .B(i_addr_b[27]), .S(n2), .Q(
        o_addr_nextpc[27]) );
  MUX22 U24 ( .A(i_addr_jumpmux[28]), .B(i_addr_b[28]), .S(n2), .Q(
        o_addr_nextpc[28]) );
  MUX22 U25 ( .A(i_addr_jumpmux[29]), .B(i_addr_b[29]), .S(n2), .Q(
        o_addr_nextpc[29]) );
  MUX22 U26 ( .A(i_addr_jumpmux[30]), .B(i_addr_b[30]), .S(n2), .Q(
        o_addr_nextpc[30]) );
  MUX22 U27 ( .A(i_addr_jumpmux[31]), .B(i_addr_b[31]), .S(n2), .Q(
        o_addr_nextpc[31]) );
  MUX22 U28 ( .A(i_addr_jumpmux[10]), .B(i_addr_b[10]), .S(n1), .Q(
        o_addr_nextpc[10]) );
  MUX22 U29 ( .A(i_addr_jumpmux[12]), .B(i_addr_b[12]), .S(n1), .Q(
        o_addr_nextpc[12]) );
  MUX22 U30 ( .A(i_addr_jumpmux[13]), .B(i_addr_b[13]), .S(n1), .Q(
        o_addr_nextpc[13]) );
  MUX22 U31 ( .A(i_addr_jumpmux[16]), .B(i_addr_b[16]), .S(n1), .Q(
        o_addr_nextpc[16]) );
  MUX22 U32 ( .A(i_addr_jumpmux[17]), .B(i_addr_b[17]), .S(n1), .Q(
        o_addr_nextpc[17]) );
  MUX22 U33 ( .A(i_addr_jumpmux[18]), .B(i_addr_b[18]), .S(n1), .Q(
        o_addr_nextpc[18]) );
  MUX22 U34 ( .A(i_addr_jumpmux[20]), .B(i_addr_b[20]), .S(n1), .Q(
        o_addr_nextpc[20]) );
  MUX22 U35 ( .A(i_addr_jumpmux[21]), .B(i_addr_b[21]), .S(n1), .Q(
        o_addr_nextpc[21]) );
  AOI221 U36 ( .A(i_addr_b[0]), .B(n2), .C(i_addr_jumpmux[0]), .D(n3), .Q(n66)
         );
  AOI221 U37 ( .A(i_addr_b[1]), .B(n2), .C(i_addr_jumpmux[1]), .D(n3), .Q(n55)
         );
  AOI221 U38 ( .A(i_addr_b[2]), .B(n2), .C(i_addr_jumpmux[2]), .D(n3), .Q(n44)
         );
  AOI221 U39 ( .A(i_addr_b[3]), .B(n2), .C(i_addr_jumpmux[3]), .D(n3), .Q(n41)
         );
  AOI221 U40 ( .A(i_con_ifbranch), .B(i_addr_b[9]), .C(i_addr_jumpmux[9]), .D(
        n3), .Q(n35) );
  AOI221 U41 ( .A(i_addr_b[4]), .B(n1), .C(i_addr_jumpmux[4]), .D(n3), .Q(n40)
         );
  AOI221 U42 ( .A(i_addr_b[5]), .B(n1), .C(i_addr_jumpmux[5]), .D(n3), .Q(n39)
         );
  AOI221 U43 ( .A(i_addr_b[6]), .B(n1), .C(i_addr_jumpmux[6]), .D(n3), .Q(n38)
         );
  AOI221 U44 ( .A(i_addr_b[7]), .B(n2), .C(i_addr_jumpmux[7]), .D(n3), .Q(n37)
         );
  AOI221 U45 ( .A(i_addr_b[8]), .B(n1), .C(i_addr_jumpmux[8]), .D(n3), .Q(n36)
         );
endmodule


module F_pc ( i_clk, i_rst_n, i_con_stall, i_addr_next_pc, o_addr_pc );
  input [31:0] i_addr_next_pc;
  output [31:0] o_addr_pc;
  input i_clk, i_rst_n, i_con_stall;


  DFEC1 program_counter_reg_31_ ( .D(i_addr_next_pc[31]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[31]) );
  DFEC1 program_counter_reg_1_ ( .D(i_addr_next_pc[1]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[1]) );
  DFEC1 program_counter_reg_0_ ( .D(i_addr_next_pc[0]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[0]) );
  DFEC1 program_counter_reg_27_ ( .D(i_addr_next_pc[27]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[27]) );
  DFEC1 program_counter_reg_23_ ( .D(i_addr_next_pc[23]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[23]) );
  DFEC1 program_counter_reg_30_ ( .D(i_addr_next_pc[30]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[30]) );
  DFEC1 program_counter_reg_29_ ( .D(i_addr_next_pc[29]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[29]) );
  DFEC1 program_counter_reg_28_ ( .D(i_addr_next_pc[28]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[28]) );
  DFEC1 program_counter_reg_19_ ( .D(i_addr_next_pc[19]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[19]) );
  DFEC1 program_counter_reg_2_ ( .D(i_addr_next_pc[2]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[2]) );
  DFEC1 program_counter_reg_15_ ( .D(i_addr_next_pc[15]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[15]) );
  DFEC1 program_counter_reg_11_ ( .D(i_addr_next_pc[11]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[11]) );
  DFEC1 program_counter_reg_9_ ( .D(i_addr_next_pc[9]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[9]) );
  DFEC1 program_counter_reg_7_ ( .D(i_addr_next_pc[7]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[7]) );
  DFEC1 program_counter_reg_5_ ( .D(i_addr_next_pc[5]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[5]) );
  DFEC1 program_counter_reg_4_ ( .D(i_addr_next_pc[4]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[4]) );
  DFEC1 program_counter_reg_8_ ( .D(i_addr_next_pc[8]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[8]) );
  DFEC1 program_counter_reg_3_ ( .D(i_addr_next_pc[3]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[3]) );
  DFEC1 program_counter_reg_12_ ( .D(i_addr_next_pc[12]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[12]) );
  DFEC1 program_counter_reg_26_ ( .D(i_addr_next_pc[26]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[26]) );
  DFEC1 program_counter_reg_25_ ( .D(i_addr_next_pc[25]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[25]) );
  DFEC1 program_counter_reg_22_ ( .D(i_addr_next_pc[22]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[22]) );
  DFEC1 program_counter_reg_21_ ( .D(i_addr_next_pc[21]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[21]) );
  DFEC1 program_counter_reg_18_ ( .D(i_addr_next_pc[18]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[18]) );
  DFEC1 program_counter_reg_17_ ( .D(i_addr_next_pc[17]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[17]) );
  DFEC1 program_counter_reg_13_ ( .D(i_addr_next_pc[13]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[13]) );
  DFEC1 program_counter_reg_10_ ( .D(i_addr_next_pc[10]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[10]) );
  DFEC1 program_counter_reg_6_ ( .D(i_addr_next_pc[6]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[6]) );
  DFEC1 program_counter_reg_14_ ( .D(i_addr_next_pc[14]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[14]) );
  DFEC1 program_counter_reg_16_ ( .D(i_addr_next_pc[16]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[16]) );
  DFEC1 program_counter_reg_24_ ( .D(i_addr_next_pc[24]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[24]) );
  DFEC1 program_counter_reg_20_ ( .D(i_addr_next_pc[20]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[20]) );
endmodule


module F_add4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   A_1_, A_0_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101;
  assign SUM[1] = A_1_;
  assign A_1_ = A[1];
  assign SUM[0] = A_0_;
  assign A_0_ = A[0];

  NAND22 U2 ( .A(n2), .B(n3), .Q(n1) );
  NAND22 U3 ( .A(n90), .B(n3), .Q(n89) );
  NAND22 U4 ( .A(n88), .B(n3), .Q(n87) );
  NAND22 U5 ( .A(A[16]), .B(n33), .Q(n73) );
  NAND22 U6 ( .A(n70), .B(n33), .Q(n71) );
  NAND22 U7 ( .A(n59), .B(n33), .Q(n60) );
  NAND22 U8 ( .A(n57), .B(n33), .Q(n58) );
  NAND31 U9 ( .A(n33), .B(A[21]), .C(n57), .Q(n56) );
  NAND22 U10 ( .A(n19), .B(n33), .Q(n46) );
  NAND31 U11 ( .A(n19), .B(n33), .C(A[24]), .Q(n45) );
  NAND31 U12 ( .A(n31), .B(n33), .C(n19), .Q(n32) );
  INV3 U13 ( .A(n34), .Q(n33) );
  CLKIN3 U14 ( .A(A[2]), .Q(SUM[2]) );
  NAND31 U15 ( .A(n43), .B(n19), .C(n33), .Q(n42) );
  CLKIN0 U16 ( .A(A[8]), .Q(n4) );
  INV0 U17 ( .A(A[13]), .Q(n86) );
  INV0 U18 ( .A(A[6]), .Q(n10) );
  INV0 U19 ( .A(A[10]), .Q(n95) );
  XOR21 U20 ( .A(n37), .B(n42), .Q(SUM[26]) );
  XOR21 U21 ( .A(n51), .B(n56), .Q(SUM[22]) );
  XOR21 U22 ( .A(n36), .B(n45), .Q(SUM[25]) );
  XOR21 U23 ( .A(n63), .B(n73), .Q(SUM[17]) );
  XOR21 U24 ( .A(n64), .B(n71), .Q(SUM[18]) );
  XOR21 U25 ( .A(n50), .B(n58), .Q(SUM[21]) );
  NOR20 U26 ( .A(n34), .B(n69), .Q(n68) );
  XOR20 U27 ( .A(n33), .B(A[16]), .Q(SUM[16]) );
  XNR20 U28 ( .A(A[11]), .B(n93), .Q(SUM[11]) );
  XNR20 U29 ( .A(A[15]), .B(n80), .Q(SUM[15]) );
  XNR20 U30 ( .A(A[7]), .B(n8), .Q(SUM[7]) );
  NAND20 U31 ( .A(A[4]), .B(n14), .Q(n13) );
  CLKIN3 U32 ( .A(n90), .Q(n79) );
  CLKIN3 U33 ( .A(n99), .Q(n78) );
  XNR20 U34 ( .A(A[12]), .B(n89), .Q(SUM[12]) );
  XOR20 U35 ( .A(A[4]), .B(n14), .Q(SUM[4]) );
  XNR20 U36 ( .A(A[3]), .B(SUM[2]), .Q(SUM[3]) );
  XNR20 U37 ( .A(A[8]), .B(n7), .Q(SUM[8]) );
  INV0 U38 ( .A(A[5]), .Q(n11) );
  INV0 U39 ( .A(A[9]), .Q(n6) );
  INV3 U40 ( .A(n7), .Q(n3) );
  INV3 U41 ( .A(n47), .Q(n19) );
  NAND22 U42 ( .A(n59), .B(n48), .Q(n47) );
  NOR31 U43 ( .A(n49), .B(n50), .C(n51), .Q(n48) );
  XNR21 U44 ( .A(n94), .B(n95), .Q(SUM[10]) );
  XNR21 U45 ( .A(n81), .B(n82), .Q(SUM[14]) );
  NOR21 U46 ( .A(n44), .B(n36), .Q(n43) );
  INV3 U47 ( .A(n98), .Q(n7) );
  NOR31 U48 ( .A(n78), .B(n16), .C(SUM[2]), .Q(n98) );
  INV3 U49 ( .A(n96), .Q(n94) );
  NAND22 U50 ( .A(n97), .B(n3), .Q(n96) );
  NOR21 U51 ( .A(n6), .B(n4), .Q(n97) );
  INV3 U52 ( .A(n83), .Q(n81) );
  NAND22 U53 ( .A(n84), .B(n3), .Q(n83) );
  NOR21 U54 ( .A(n85), .B(n86), .Q(n84) );
  XNR21 U55 ( .A(n12), .B(n11), .Q(SUM[5]) );
  XNR21 U56 ( .A(n9), .B(n10), .Q(SUM[6]) );
  NOR21 U57 ( .A(n63), .B(n72), .Q(n70) );
  NOR21 U58 ( .A(n11), .B(n13), .Q(n9) );
  NOR21 U59 ( .A(SUM[2]), .B(n16), .Q(n14) );
  XNR21 U60 ( .A(n5), .B(n1), .Q(SUM[9]) );
  INV3 U61 ( .A(n6), .Q(n5) );
  XNR21 U62 ( .A(A[13]), .B(n87), .Q(SUM[13]) );
  NOR21 U63 ( .A(n37), .B(n36), .Q(n41) );
  NOR21 U64 ( .A(n51), .B(n50), .Q(n54) );
  INV3 U65 ( .A(n52), .Q(n59) );
  INV3 U66 ( .A(n68), .Q(n67) );
  INV3 U67 ( .A(n70), .Q(n69) );
  INV3 U68 ( .A(n4), .Q(n2) );
  XNR21 U69 ( .A(A[20]), .B(n60), .Q(SUM[20]) );
  XNR21 U70 ( .A(A[24]), .B(n46), .Q(SUM[24]) );
  NAND22 U71 ( .A(n94), .B(A[10]), .Q(n93) );
  XOR21 U72 ( .A(n28), .B(n29), .Q(SUM[29]) );
  INV3 U73 ( .A(A[29]), .Q(n28) );
  NAND31 U74 ( .A(n19), .B(n33), .C(n30), .Q(n29) );
  NOR21 U75 ( .A(n27), .B(n22), .Q(n30) );
  NAND22 U76 ( .A(n81), .B(A[14]), .Q(n80) );
  NAND22 U77 ( .A(n74), .B(n75), .Q(n34) );
  NOR21 U78 ( .A(n78), .B(n79), .Q(n74) );
  NOR21 U79 ( .A(n76), .B(n77), .Q(n75) );
  NAND41 U80 ( .A(A[14]), .B(A[13]), .C(A[12]), .D(A[15]), .Q(n76) );
  XNR21 U81 ( .A(A[28]), .B(n32), .Q(SUM[28]) );
  XOR21 U82 ( .A(n23), .B(n24), .Q(SUM[30]) );
  INV3 U83 ( .A(A[30]), .Q(n23) );
  NAND31 U84 ( .A(n25), .B(n33), .C(n19), .Q(n24) );
  NOR21 U85 ( .A(n22), .B(n21), .Q(n25) );
  XOR21 U86 ( .A(n17), .B(n18), .Q(SUM[31]) );
  INV3 U87 ( .A(A[31]), .Q(n17) );
  NAND31 U88 ( .A(n20), .B(n33), .C(n19), .Q(n18) );
  NOR31 U89 ( .A(n21), .B(n23), .C(n22), .Q(n20) );
  XNR21 U90 ( .A(A[23]), .B(n53), .Q(SUM[23]) );
  NAND31 U91 ( .A(n54), .B(n57), .C(n33), .Q(n53) );
  NAND22 U92 ( .A(n61), .B(n62), .Q(n52) );
  NOR21 U93 ( .A(n72), .B(n65), .Q(n61) );
  NOR21 U94 ( .A(n63), .B(n64), .Q(n62) );
  INV3 U95 ( .A(A[19]), .Q(n65) );
  INV3 U96 ( .A(A[17]), .Q(n63) );
  INV3 U97 ( .A(A[18]), .Q(n64) );
  NAND22 U98 ( .A(A[23]), .B(A[20]), .Q(n49) );
  NOR21 U99 ( .A(n91), .B(n92), .Q(n90) );
  NAND22 U100 ( .A(A[10]), .B(A[11]), .Q(n92) );
  NAND22 U101 ( .A(A[8]), .B(A[9]), .Q(n91) );
  NAND22 U102 ( .A(A[3]), .B(A[2]), .Q(n77) );
  NOR21 U103 ( .A(n100), .B(n101), .Q(n99) );
  NAND22 U104 ( .A(A[6]), .B(A[7]), .Q(n101) );
  NAND22 U105 ( .A(A[4]), .B(A[5]), .Q(n100) );
  XNR21 U106 ( .A(n38), .B(n39), .Q(SUM[27]) );
  INV3 U107 ( .A(A[27]), .Q(n38) );
  NOR21 U108 ( .A(n40), .B(n34), .Q(n39) );
  NAND31 U109 ( .A(n41), .B(A[24]), .C(n19), .Q(n40) );
  NAND22 U110 ( .A(n9), .B(A[6]), .Q(n8) );
  INV3 U111 ( .A(A[25]), .Q(n36) );
  INV3 U112 ( .A(A[21]), .Q(n50) );
  NOR31 U113 ( .A(n37), .B(n35), .C(n36), .Q(n31) );
  NAND22 U114 ( .A(A[27]), .B(A[24]), .Q(n35) );
  NAND22 U115 ( .A(n90), .B(A[12]), .Q(n85) );
  INV3 U116 ( .A(A[26]), .Q(n37) );
  INV3 U117 ( .A(A[22]), .Q(n51) );
  NAND22 U118 ( .A(n59), .B(A[20]), .Q(n55) );
  INV3 U119 ( .A(A[3]), .Q(n16) );
  INV3 U120 ( .A(A[28]), .Q(n27) );
  INV3 U121 ( .A(A[24]), .Q(n44) );
  INV3 U122 ( .A(A[16]), .Q(n72) );
  INV3 U123 ( .A(A[14]), .Q(n82) );
  INV3 U124 ( .A(n26), .Q(n21) );
  NOR21 U125 ( .A(n27), .B(n28), .Q(n26) );
  INV3 U126 ( .A(n13), .Q(n12) );
  XOR21 U127 ( .A(A[19]), .B(n66), .Q(SUM[19]) );
  NOR21 U128 ( .A(n64), .B(n67), .Q(n66) );
  CLKIN3 U129 ( .A(n31), .Q(n22) );
  CLKIN3 U130 ( .A(n55), .Q(n57) );
  CLKIN3 U131 ( .A(n85), .Q(n88) );
endmodule


module F_add4 ( i_addr_pc, o_addr_pcadd4 );
  input [31:0] i_addr_pc;
  output [31:0] o_addr_pcadd4;
  wire   n2, n1;

  F_add4_DW01_add_1 add_5 ( .A(i_addr_pc), .B({n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n2, n1, n1}), .CI(n1), .SUM(o_addr_pcadd4) );
  LOGIC0 U3 ( .Q(n1) );
  LOGIC1 U4 ( .Q(n2) );
endmodule


module fetch ( i_clk, i_nrst, i_addr_b, i_addr_j, i_addr_jr, i_con_b, i_con_j, 
        i_data_instr, i_con_ifstall, o_addr_pc, o_addr_pc4, o_data_instr );
  input [31:0] i_addr_b;
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [1:0] i_con_j;
  input [31:0] i_data_instr;
  output [31:0] o_addr_pc;
  output [31:0] o_addr_pc4;
  output [31:0] o_data_instr;
  input i_clk, i_nrst, i_con_b, i_con_ifstall;

  wire   [31:0] jmux_i_addr_pc4;
  wire   [31:0] bmux_i_addr_jumpmux;
  wire   [31:0] pc_i_addr_next_pc;

  DFC3 pipe_instr_reg_31_ ( .D(i_data_instr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[31]) );
  DFC3 pipe_instr_reg_30_ ( .D(i_data_instr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[30]) );
  DFC3 pipe_instr_reg_29_ ( .D(i_data_instr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[29]) );
  DFC3 pipe_instr_reg_28_ ( .D(i_data_instr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[28]) );
  DFC3 pipe_instr_reg_27_ ( .D(i_data_instr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[27]) );
  DFC3 pipe_instr_reg_26_ ( .D(i_data_instr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[26]) );
  DFC3 pipe_instr_reg_25_ ( .D(i_data_instr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[25]) );
  DFC3 pipe_instr_reg_24_ ( .D(i_data_instr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[24]) );
  DFC3 pipe_instr_reg_23_ ( .D(i_data_instr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[23]) );
  DFC3 pipe_instr_reg_22_ ( .D(i_data_instr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[22]) );
  DFC3 pipe_instr_reg_21_ ( .D(i_data_instr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[21]) );
  DFC3 pipe_instr_reg_20_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[20]) );
  DFC3 pipe_instr_reg_19_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[19]) );
  DFC3 pipe_instr_reg_18_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[18]) );
  DFC3 pipe_instr_reg_17_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[17]) );
  DFC3 pipe_instr_reg_16_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[16]) );
  DFC3 pipe_instr_reg_15_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[15]) );
  DFC3 pipe_instr_reg_14_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[14]) );
  DFC3 pipe_instr_reg_13_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[13]) );
  DFC3 pipe_instr_reg_12_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[12]) );
  DFC3 pipe_instr_reg_11_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[11]) );
  DFC3 pipe_instr_reg_10_ ( .D(i_data_instr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[10]) );
  DFC3 pipe_instr_reg_9_ ( .D(i_data_instr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[9]) );
  DFC3 pipe_instr_reg_8_ ( .D(i_data_instr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[8]) );
  DFC3 pipe_instr_reg_7_ ( .D(i_data_instr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[7]) );
  DFC3 pipe_instr_reg_6_ ( .D(i_data_instr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[6]) );
  DFC3 pipe_instr_reg_5_ ( .D(i_data_instr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[5]) );
  DFC3 pipe_instr_reg_4_ ( .D(i_data_instr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[4]) );
  DFC3 pipe_instr_reg_3_ ( .D(i_data_instr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[3]) );
  DFC3 pipe_instr_reg_2_ ( .D(i_data_instr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[2]) );
  DFC3 pipe_instr_reg_1_ ( .D(i_data_instr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[1]) );
  DFC3 pipe_instr_reg_0_ ( .D(i_data_instr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(jmux_i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(jmux_i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(jmux_i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(jmux_i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(jmux_i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(jmux_i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(jmux_i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(jmux_i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_pc4_reg_22_ ( .D(jmux_i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(jmux_i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(jmux_i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(jmux_i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(jmux_i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(jmux_i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(jmux_i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(jmux_i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(jmux_i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(jmux_i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(jmux_i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(jmux_i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(jmux_i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(jmux_i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(jmux_i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(jmux_i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(jmux_i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(jmux_i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(jmux_i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(jmux_i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(jmux_i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(jmux_i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(jmux_i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  F_jumpmux u_jumpmux ( .i_addr_j(i_addr_j), .i_addr_jr(i_addr_jr), 
        .i_addr_pc4(jmux_i_addr_pc4), .i_con_jump(i_con_j), .o_addr_jumpmux(
        bmux_i_addr_jumpmux) );
  F_branchmux u_branchmux ( .i_addr_jumpmux(bmux_i_addr_jumpmux), .i_addr_b(
        i_addr_b), .i_con_ifbranch(i_con_b), .o_addr_nextpc(pc_i_addr_next_pc)
         );
  F_pc u_pc ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_con_stall(i_con_ifstall), 
        .i_addr_next_pc(pc_i_addr_next_pc), .o_addr_pc(o_addr_pc) );
  F_add4 u_add4 ( .i_addr_pc(o_addr_pc), .o_addr_pcadd4(jmux_i_addr_pc4) );
  DFC1 pipe_pc4_reg_23_ ( .D(jmux_i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
endmodule


module D_control ( o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite, 
        o_con_alusrc, o_con_regwrite, o_con_ifsign, o_con_loadsig, o_con_aluop, 
        i_con_instru );
  output [1:0] o_con_loadsig;
  output [5:0] o_con_aluop;
  input [5:0] i_con_instru;
  output o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite,
         o_con_alusrc, o_con_regwrite, o_con_ifsign;
  wire   n_Logic0_, o_con_alusrc, n9, n10, n11, n12, n13, n14, n15, n16, n1,
         n2, n3, n4, n5, n6, n7;
  assign o_con_loadsig[0] = n_Logic0_;
  assign o_con_loadsig[1] = n_Logic0_;
  assign o_con_memwrite = n_Logic0_;
  assign o_con_memtoreg = n_Logic0_;
  assign o_con_memread = n_Logic0_;
  assign o_con_aluop[0] = o_con_alusrc;

  OAI212 U2 ( .A(n6), .B(n2), .C(n9), .Q(o_con_regwrite) );
  OAI222 U9 ( .A(n10), .B(n11), .C(n4), .D(n14), .Q(o_con_aluop[2]) );
  OAI212 U11 ( .A(n6), .B(n9), .C(n1), .Q(o_con_aluop[1]) );
  OAI212 U15 ( .A(n6), .B(n2), .C(n10), .Q(o_con_alusrc) );
  OAI2110 U3 ( .A(i_con_instru[1]), .B(n7), .C(n12), .D(n16), .Q(n9) );
  NOR30 U4 ( .A(i_con_instru[2]), .B(i_con_instru[5]), .C(i_con_instru[4]), 
        .Q(n16) );
  NOR30 U5 ( .A(i_con_instru[4]), .B(i_con_instru[5]), .C(n3), .Q(n15) );
  INV0 U6 ( .A(i_con_instru[3]), .Q(n3) );
  NAND20 U7 ( .A(i_con_instru[1]), .B(i_con_instru[0]), .Q(n11) );
  NAND20 U8 ( .A(i_con_instru[1]), .B(n7), .Q(n12) );
  NOR30 U10 ( .A(n9), .B(i_con_instru[3]), .C(n6), .Q(o_con_regdst) );
  INV0 U12 ( .A(i_con_instru[0]), .Q(n7) );
  INV0 U13 ( .A(i_con_instru[2]), .Q(n4) );
  NAND30 U14 ( .A(i_con_instru[0]), .B(n5), .C(i_con_instru[2]), .Q(n13) );
  INV0 U16 ( .A(i_con_instru[1]), .Q(n5) );
  NAND22 U17 ( .A(n15), .B(n4), .Q(n10) );
  INV3 U18 ( .A(n11), .Q(n6) );
  NAND22 U19 ( .A(n15), .B(n7), .Q(n14) );
  INV3 U20 ( .A(o_con_alusrc), .Q(n1) );
  INV3 U21 ( .A(n15), .Q(n2) );
  NOR21 U22 ( .A(n10), .B(n12), .Q(o_con_aluop[4]) );
  NOR21 U23 ( .A(n10), .B(n11), .Q(o_con_aluop[5]) );
  NOR21 U24 ( .A(n6), .B(n10), .Q(o_con_ifsign) );
  AOI211 U25 ( .A(n12), .B(n13), .C(n2), .Q(o_con_aluop[3]) );
  LOGIC0 U26 ( .Q(n_Logic0_) );
endmodule


module D_jb_control ( o_con_jump, o_con_bop, o_con_aluPC4, o_con_ifstall, 
        i_con_instru, i_con_func, i_con_rt );
  output [1:0] o_con_jump;
  output [2:0] o_con_bop;
  input [5:0] i_con_instru;
  input [5:0] i_con_func;
  input i_con_rt;
  output o_con_aluPC4, o_con_ifstall;
  wire   n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n1, n3, n4,
         n5, n6;

  OAI222 U13 ( .A(n5), .B(n17), .C(n15), .D(n18), .Q(o_con_bop[1]) );
  NOR31 U3 ( .A(i_con_instru[3]), .B(i_con_instru[5]), .C(i_con_instru[4]), 
        .Q(n8) );
  NOR40 U4 ( .A(n12), .B(i_con_func[2]), .C(i_con_func[5]), .D(i_con_func[4]), 
        .Q(n10) );
  CLKIN3 U5 ( .A(i_con_instru[1]), .Q(n5) );
  CLKIN3 U6 ( .A(i_con_instru[0]), .Q(n6) );
  CLKIN3 U7 ( .A(i_con_instru[2]), .Q(n4) );
  NAND20 U8 ( .A(i_con_instru[0]), .B(n5), .Q(n15) );
  NAND30 U9 ( .A(n8), .B(n6), .C(i_con_instru[2]), .Q(n17) );
  NOR30 U10 ( .A(n16), .B(n3), .C(n6), .Q(o_con_bop[2]) );
  XNR20 U11 ( .A(n5), .B(i_con_instru[2]), .Q(n16) );
  NOR20 U12 ( .A(i_con_instru[2]), .B(i_con_rt), .Q(n19) );
  NAND31 U14 ( .A(n5), .B(n4), .C(n6), .Q(n9) );
  NAND22 U15 ( .A(n8), .B(n9), .Q(o_con_jump[1]) );
  INV3 U16 ( .A(n8), .Q(n3) );
  INV3 U17 ( .A(n14), .Q(o_con_ifstall) );
  AOI211 U18 ( .A(n4), .B(n15), .C(n3), .Q(n14) );
  OAI311 U19 ( .A(n1), .B(n3), .C(n15), .D(n17), .Q(o_con_bop[0]) );
  NAND22 U20 ( .A(n8), .B(n1), .Q(n18) );
  OAI2111 U21 ( .A(n10), .B(n9), .C(n11), .D(n8), .Q(o_con_jump[0]) );
  NAND22 U22 ( .A(i_con_instru[1]), .B(n4), .Q(n11) );
  NAND22 U23 ( .A(n13), .B(i_con_func[3]), .Q(n12) );
  NOR21 U24 ( .A(i_con_func[1]), .B(i_con_func[0]), .Q(n13) );
  NOR40 U25 ( .A(i_con_instru[2]), .B(n3), .C(n5), .D(n6), .Q(o_con_aluPC4) );
  INV3 U26 ( .A(n19), .Q(n1) );
endmodule


module D_pcadd_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318;

  INV3 U2 ( .A(n41), .Q(n36) );
  NAND31 U3 ( .A(n290), .B(n291), .C(n292), .Q(n41) );
  NAND22 U4 ( .A(n254), .B(n220), .Q(n256) );
  NAND22 U5 ( .A(n184), .B(n195), .Q(n196) );
  NAND22 U6 ( .A(n25), .B(n27), .Q(n28) );
  NAND22 U7 ( .A(n14), .B(n15), .Q(n12) );
  NAND22 U8 ( .A(n259), .B(n219), .Q(n260) );
  OAI312 U9 ( .A(n123), .B(n124), .C(n125), .D(n126), .Q(n122) );
  NAND42 U10 ( .A(n208), .B(n209), .C(n210), .D(n41), .Q(n132) );
  OAI210 U11 ( .A(n29), .B(n30), .C(n31), .Q(n24) );
  NAND20 U12 ( .A(B[6]), .B(A[6]), .Q(n27) );
  INV0 U13 ( .A(B[22]), .Q(n9) );
  AOI211 U14 ( .A(n253), .B(n254), .C(n255), .Q(n252) );
  AOI211 U15 ( .A(n154), .B(n148), .C(n159), .Q(n158) );
  NAND20 U16 ( .A(n142), .B(n144), .Q(n157) );
  XOR20 U17 ( .A(n32), .B(n34), .Q(SUM[5]) );
  NOR20 U18 ( .A(n29), .B(n35), .Q(n34) );
  XNR20 U19 ( .A(n260), .B(n258), .Q(SUM[13]) );
  XNR20 U20 ( .A(n28), .B(n24), .Q(SUM[6]) );
  XNR20 U21 ( .A(n12), .B(n13), .Q(SUM[9]) );
  INV3 U22 ( .A(n195), .Q(n177) );
  NAND20 U23 ( .A(n129), .B(n130), .Q(n125) );
  CLKIN3 U24 ( .A(n185), .Q(n183) );
  NAND21 U25 ( .A(n133), .B(n134), .Q(n123) );
  INV3 U26 ( .A(n237), .Q(n209) );
  INV0 U27 ( .A(n142), .Q(n156) );
  INV1 U28 ( .A(n128), .Q(n135) );
  INV1 U29 ( .A(n33), .Q(n25) );
  NOR21 U30 ( .A(A[2]), .B(B[2]), .Q(n49) );
  NAND22 U31 ( .A(B[26]), .B(A[26]), .Q(n96) );
  NAND20 U32 ( .A(A[12]), .B(B[12]), .Q(n218) );
  CLKIN2 U33 ( .A(B[18]), .Q(n7) );
  XOR20 U34 ( .A(B[23]), .B(A[23]), .Q(n3) );
  NOR20 U35 ( .A(A[20]), .B(B[20]), .Q(n168) );
  AOI210 U36 ( .A(n82), .B(n53), .C(n79), .Q(n85) );
  AOI210 U37 ( .A(n66), .B(n53), .C(n63), .Q(n76) );
  AOI210 U38 ( .A(n52), .B(n53), .C(n57), .Q(n60) );
  CLKIN3 U39 ( .A(B[17]), .Q(n6) );
  NOR20 U40 ( .A(B[24]), .B(A[24]), .Q(n99) );
  NAND21 U41 ( .A(B[20]), .B(A[20]), .Q(n146) );
  INV0 U42 ( .A(A[3]), .Q(n298) );
  NAND20 U43 ( .A(B[24]), .B(A[24]), .Q(n108) );
  IMUX20 U44 ( .A(n16), .B(n17), .S(n18), .Q(SUM[8]) );
  XNR20 U45 ( .A(B[12]), .B(A[12]), .Q(n268) );
  AOI210 U46 ( .A(n208), .B(n270), .C(n264), .Q(n269) );
  NOR20 U47 ( .A(n236), .B(n237), .Q(n226) );
  NAND20 U48 ( .A(B[24]), .B(A[24]), .Q(n92) );
  NAND20 U49 ( .A(n283), .B(n284), .Q(n282) );
  NOR20 U50 ( .A(A[24]), .B(B[24]), .Q(n116) );
  NOR20 U51 ( .A(B[20]), .B(A[20]), .Q(n189) );
  NOR20 U52 ( .A(B[24]), .B(A[24]), .Q(n152) );
  NOR20 U53 ( .A(A[12]), .B(B[12]), .Q(n266) );
  NAND20 U54 ( .A(B[12]), .B(A[12]), .Q(n263) );
  NOR20 U55 ( .A(B[12]), .B(A[12]), .Q(n278) );
  XOR20 U56 ( .A(n154), .B(n161), .Q(SUM[21]) );
  AOI210 U57 ( .A(n111), .B(n53), .C(n115), .Q(n114) );
  AOI210 U58 ( .A(n102), .B(n53), .C(n105), .Q(n107) );
  NAND20 U59 ( .A(n210), .B(n41), .Q(n289) );
  AOI210 U60 ( .A(n198), .B(n165), .C(n199), .Q(n202) );
  NOR20 U61 ( .A(n127), .B(n168), .Q(n164) );
  XNR20 U62 ( .A(n196), .B(n194), .Q(SUM[18]) );
  INV3 U63 ( .A(n148), .Q(n145) );
  INV0 U64 ( .A(n127), .Q(n173) );
  NAND20 U65 ( .A(B[3]), .B(A[3]), .Q(n292) );
  NOR20 U66 ( .A(A[5]), .B(B[5]), .Q(n29) );
  INV0 U67 ( .A(B[25]), .Q(n10) );
  INV0 U68 ( .A(B[26]), .Q(n11) );
  NOR20 U69 ( .A(A[6]), .B(B[6]), .Q(n33) );
  OAI2110 U70 ( .A(A[6]), .B(B[6]), .C(A[5]), .D(B[5]), .Q(n314) );
  NOR20 U71 ( .A(A[3]), .B(B[3]), .Q(n301) );
  NAND21 U72 ( .A(B[25]), .B(A[25]), .Q(n93) );
  NAND21 U73 ( .A(B[22]), .B(A[22]), .Q(n144) );
  XNR20 U74 ( .A(B[28]), .B(A[28]), .Q(n84) );
  XNR20 U75 ( .A(B[29]), .B(A[29]), .Q(n75) );
  XNR20 U76 ( .A(B[30]), .B(A[30]), .Q(n59) );
  NAND21 U77 ( .A(B[18]), .B(A[18]), .Q(n195) );
  NOR20 U78 ( .A(A[4]), .B(B[4]), .Q(n37) );
  NOR20 U79 ( .A(A[19]), .B(B[19]), .Q(n179) );
  NOR20 U80 ( .A(A[7]), .B(B[7]), .Q(n315) );
  NOR20 U81 ( .A(B[7]), .B(A[7]), .Q(n307) );
  OAI220 U82 ( .A(A[5]), .B(B[5]), .C(A[6]), .D(B[6]), .Q(n312) );
  INV0 U83 ( .A(B[3]), .Q(n297) );
  XNR21 U84 ( .A(n1), .B(n101), .Q(SUM[27]) );
  XOR20 U85 ( .A(B[27]), .B(A[27]), .Q(n1) );
  XNR21 U86 ( .A(n2), .B(n193), .Q(SUM[19]) );
  XOR20 U87 ( .A(B[19]), .B(A[19]), .Q(n2) );
  XNR21 U88 ( .A(n3), .B(n153), .Q(SUM[23]) );
  XNR21 U89 ( .A(n4), .B(n50), .Q(SUM[31]) );
  XOR20 U90 ( .A(B[31]), .B(A[31]), .Q(n4) );
  XNR20 U91 ( .A(B[7]), .B(A[7]), .Q(n22) );
  AOI210 U92 ( .A(n173), .B(n165), .C(n136), .Q(n172) );
  IMUX20 U93 ( .A(n205), .B(n206), .S(n165), .Q(SUM[16]) );
  NOR20 U94 ( .A(B[4]), .B(A[4]), .Q(n306) );
  NAND20 U95 ( .A(A[2]), .B(B[2]), .Q(n302) );
  NAND20 U96 ( .A(B[19]), .B(A[19]), .Q(n174) );
  NAND20 U97 ( .A(B[28]), .B(A[28]), .Q(n78) );
  NAND20 U98 ( .A(B[29]), .B(A[29]), .Q(n62) );
  AOI210 U99 ( .A(A[27]), .B(B[27]), .C(n95), .Q(n86) );
  NOR20 U100 ( .A(A[28]), .B(B[28]), .Q(n83) );
  NOR20 U101 ( .A(A[29]), .B(B[29]), .Q(n67) );
  NAND20 U102 ( .A(B[7]), .B(A[7]), .Q(n308) );
  NAND20 U103 ( .A(B[4]), .B(A[4]), .Q(n313) );
  NOR20 U104 ( .A(B[27]), .B(A[27]), .Q(n100) );
  NAND20 U105 ( .A(B[4]), .B(A[4]), .Q(n38) );
  XNR21 U106 ( .A(n44), .B(n5), .Q(SUM[3]) );
  XNR20 U107 ( .A(B[3]), .B(A[3]), .Q(n5) );
  XNR20 U108 ( .A(B[4]), .B(A[4]), .Q(n40) );
  NOR20 U109 ( .A(B[4]), .B(A[4]), .Q(n42) );
  NAND20 U110 ( .A(B[30]), .B(A[30]), .Q(n56) );
  NOR20 U111 ( .A(A[30]), .B(B[30]), .Q(n58) );
  NAND20 U112 ( .A(B[5]), .B(A[5]), .Q(n31) );
  NAND20 U113 ( .A(B[2]), .B(A[2]), .Q(n45) );
  NAND22 U114 ( .A(n242), .B(n225), .Q(n133) );
  NOR21 U115 ( .A(n159), .B(n145), .Q(n161) );
  NAND41 U116 ( .A(n133), .B(n134), .C(n207), .D(n132), .Q(n165) );
  NOR21 U117 ( .A(n212), .B(n131), .Q(n207) );
  OAI2111 U118 ( .A(n18), .B(n261), .C(n262), .D(n263), .Q(n258) );
  NAND22 U119 ( .A(n265), .B(n208), .Q(n261) );
  NAND22 U120 ( .A(n264), .B(n265), .Q(n262) );
  INV3 U121 ( .A(n266), .Q(n265) );
  INV3 U122 ( .A(n211), .Q(n210) );
  AOI211 U123 ( .A(n198), .B(n165), .C(n199), .Q(n197) );
  XOR21 U124 ( .A(n113), .B(n114), .Q(SUM[25]) );
  NAND22 U125 ( .A(n90), .B(n93), .Q(n113) );
  XOR21 U126 ( .A(n106), .B(n107), .Q(SUM[26]) );
  NAND22 U127 ( .A(n88), .B(n96), .Q(n106) );
  AOI2111 U128 ( .A(n180), .B(n181), .C(n182), .D(n183), .Q(n176) );
  NAND22 U129 ( .A(n208), .B(n209), .Q(n243) );
  NAND22 U130 ( .A(n310), .B(n311), .Q(n309) );
  INV3 U131 ( .A(n315), .Q(n310) );
  OAI2111 U132 ( .A(n312), .B(n313), .C(n314), .D(n27), .Q(n311) );
  NAND22 U133 ( .A(n121), .B(n122), .Q(n53) );
  AOI211 U134 ( .A(n135), .B(n136), .C(n137), .Q(n121) );
  NAND22 U135 ( .A(n286), .B(n15), .Q(n283) );
  NAND22 U136 ( .A(n14), .B(n13), .Q(n286) );
  NAND22 U137 ( .A(n224), .B(n225), .Q(n130) );
  XOR21 U138 ( .A(n201), .B(n202), .Q(SUM[17]) );
  NAND22 U139 ( .A(n185), .B(n181), .Q(n201) );
  XOR21 U140 ( .A(n157), .B(n158), .Q(SUM[22]) );
  NAND22 U141 ( .A(n82), .B(n80), .Q(n81) );
  INV3 U142 ( .A(n163), .Q(n154) );
  AOI2111 U143 ( .A(n164), .B(n165), .C(n166), .D(n167), .Q(n163) );
  NOR21 U144 ( .A(n168), .B(n169), .Q(n167) );
  NAND22 U145 ( .A(n66), .B(n64), .Q(n65) );
  NAND22 U146 ( .A(n219), .B(n257), .Q(n253) );
  NAND22 U147 ( .A(n258), .B(n259), .Q(n257) );
  NAND22 U148 ( .A(n288), .B(n289), .Q(n270) );
  NOR21 U149 ( .A(n242), .B(n224), .Q(n288) );
  NOR21 U150 ( .A(n127), .B(n128), .Q(n126) );
  NAND22 U151 ( .A(n57), .B(n51), .Q(n55) );
  INV3 U152 ( .A(n136), .Q(n169) );
  INV3 U153 ( .A(n94), .Q(n89) );
  NAND22 U154 ( .A(n229), .B(n271), .Q(n264) );
  NAND22 U155 ( .A(n272), .B(n273), .Q(n271) );
  AOI211 U156 ( .A(n275), .B(n233), .C(n241), .Q(n272) );
  AOI311 U157 ( .A(n274), .B(n15), .C(n233), .D(n240), .Q(n273) );
  INV3 U158 ( .A(n31), .Q(n35) );
  XOR21 U159 ( .A(n283), .B(n285), .Q(SUM[10]) );
  NOR21 U160 ( .A(n235), .B(n240), .Q(n285) );
  NAND22 U161 ( .A(n111), .B(n90), .Q(n110) );
  INV3 U162 ( .A(n275), .Q(n14) );
  NOR21 U163 ( .A(n238), .B(n239), .Q(n236) );
  INV3 U164 ( .A(n229), .Q(n239) );
  NOR21 U165 ( .A(n240), .B(n241), .Q(n238) );
  XNR21 U166 ( .A(n256), .B(n253), .Q(SUM[14]) );
  NAND22 U167 ( .A(n105), .B(n88), .Q(n104) );
  NOR21 U168 ( .A(n14), .B(n232), .Q(n231) );
  NAND22 U169 ( .A(n229), .B(n233), .Q(n232) );
  NOR21 U170 ( .A(n234), .B(n235), .Q(n230) );
  INV3 U171 ( .A(n15), .Q(n234) );
  INV3 U172 ( .A(n233), .Q(n235) );
  AOI211 U173 ( .A(n108), .B(n93), .C(n109), .Q(n105) );
  INV3 U174 ( .A(n90), .Q(n109) );
  NAND22 U175 ( .A(n70), .B(n71), .Q(n47) );
  NAND22 U176 ( .A(n72), .B(n73), .Q(n71) );
  INV3 U177 ( .A(n74), .Q(n73) );
  XOR21 U178 ( .A(n47), .B(n68), .Q(SUM[2]) );
  NOR21 U179 ( .A(n69), .B(n49), .Q(n68) );
  XOR21 U180 ( .A(n72), .B(n190), .Q(SUM[1]) );
  NOR21 U181 ( .A(n191), .B(n74), .Q(n190) );
  INV3 U182 ( .A(n217), .Q(n259) );
  INV3 U183 ( .A(n223), .Q(n254) );
  INV3 U184 ( .A(n49), .Q(n48) );
  INV3 U185 ( .A(n240), .Q(n284) );
  NAND22 U186 ( .A(n11), .B(n112), .Q(n88) );
  INV3 U187 ( .A(A[26]), .Q(n112) );
  NAND22 U188 ( .A(n294), .B(n295), .Q(n291) );
  NOR21 U189 ( .A(n299), .B(n300), .Q(n290) );
  NOR21 U190 ( .A(A[8]), .B(B[8]), .Q(n287) );
  NAND31 U191 ( .A(n142), .B(n148), .C(n149), .Q(n128) );
  NOR21 U192 ( .A(n150), .B(n151), .Q(n149) );
  NOR21 U193 ( .A(B[23]), .B(A[23]), .Q(n151) );
  NOR21 U194 ( .A(B[20]), .B(A[20]), .Q(n150) );
  NOR21 U195 ( .A(n276), .B(n277), .Q(n208) );
  XOR21 U196 ( .A(n84), .B(n85), .Q(SUM[28]) );
  XOR21 U197 ( .A(n75), .B(n76), .Q(SUM[29]) );
  XOR21 U198 ( .A(n59), .B(n60), .Q(SUM[30]) );
  NAND22 U199 ( .A(B[17]), .B(A[17]), .Q(n181) );
  NAND22 U200 ( .A(n174), .B(n175), .Q(n136) );
  INV3 U201 ( .A(n179), .Q(n178) );
  NAND22 U202 ( .A(B[23]), .B(A[23]), .Q(n140) );
  NOR21 U203 ( .A(A[23]), .B(B[23]), .Q(n139) );
  AOI211 U204 ( .A(n141), .B(n142), .C(n143), .Q(n138) );
  NOR21 U205 ( .A(B[12]), .B(A[12]), .Q(n246) );
  NOR31 U206 ( .A(n303), .B(n49), .C(n301), .Q(n299) );
  NAND22 U207 ( .A(B[1]), .B(A[1]), .Q(n303) );
  NAND22 U208 ( .A(n6), .B(n204), .Q(n185) );
  INV3 U209 ( .A(A[17]), .Q(n204) );
  NOR21 U210 ( .A(A[27]), .B(B[27]), .Q(n94) );
  NAND22 U211 ( .A(B[21]), .B(A[21]), .Q(n147) );
  NAND22 U212 ( .A(n244), .B(n245), .Q(n237) );
  NOR21 U213 ( .A(n248), .B(n249), .Q(n244) );
  NOR21 U214 ( .A(n246), .B(n247), .Q(n245) );
  NOR21 U215 ( .A(A[14]), .B(B[14]), .Q(n249) );
  NOR21 U216 ( .A(B[15]), .B(A[15]), .Q(n247) );
  NAND22 U217 ( .A(n304), .B(n305), .Q(n211) );
  NOR21 U218 ( .A(n306), .B(n307), .Q(n304) );
  NOR21 U219 ( .A(n29), .B(n33), .Q(n305) );
  NAND22 U220 ( .A(n86), .B(n87), .Q(n79) );
  NAND41 U221 ( .A(n88), .B(n89), .C(n90), .D(n91), .Q(n87) );
  NOR21 U222 ( .A(n94), .B(n96), .Q(n95) );
  NAND22 U223 ( .A(n77), .B(n78), .Q(n63) );
  NAND22 U224 ( .A(n79), .B(n80), .Q(n77) );
  NAND22 U225 ( .A(n61), .B(n62), .Q(n57) );
  NAND22 U226 ( .A(n63), .B(n64), .Q(n61) );
  NOR21 U227 ( .A(n49), .B(n296), .Q(n295) );
  NAND22 U228 ( .A(B[0]), .B(A[0]), .Q(n296) );
  NAND31 U229 ( .A(n88), .B(n90), .C(n98), .Q(n97) );
  NOR21 U230 ( .A(n99), .B(n100), .Q(n98) );
  XOR21 U231 ( .A(n251), .B(n252), .Q(SUM[15]) );
  XNR21 U232 ( .A(B[15]), .B(A[15]), .Q(n251) );
  AOI211 U233 ( .A(n194), .B(n184), .C(n177), .Q(n193) );
  AOI311 U234 ( .A(n142), .B(n148), .C(n154), .D(n155), .Q(n153) );
  AOI311 U235 ( .A(n88), .B(n102), .C(n53), .D(n103), .Q(n101) );
  NAND22 U236 ( .A(n104), .B(n96), .Q(n103) );
  AOI311 U237 ( .A(n51), .B(n52), .C(n53), .D(n54), .Q(n50) );
  NAND22 U238 ( .A(n55), .B(n56), .Q(n54) );
  XOR21 U239 ( .A(n280), .B(n281), .Q(SUM[11]) );
  XOR21 U240 ( .A(B[11]), .B(A[11]), .Q(n281) );
  NAND22 U241 ( .A(n282), .B(n233), .Q(n280) );
  NOR21 U242 ( .A(A[13]), .B(B[13]), .Q(n248) );
  NAND31 U243 ( .A(n184), .B(n185), .C(n186), .Q(n127) );
  NOR21 U244 ( .A(n187), .B(n188), .Q(n186) );
  NOR21 U245 ( .A(B[16]), .B(A[16]), .Q(n187) );
  NOR21 U246 ( .A(B[19]), .B(A[19]), .Q(n188) );
  XNR21 U247 ( .A(B[16]), .B(A[16]), .Q(n205) );
  NOR21 U248 ( .A(n250), .B(n199), .Q(n206) );
  NOR21 U249 ( .A(B[16]), .B(A[16]), .Q(n250) );
  IMUX21 U250 ( .A(n118), .B(n119), .S(n120), .Q(SUM[24]) );
  XNR21 U251 ( .A(B[24]), .B(A[24]), .Q(n119) );
  NOR21 U252 ( .A(n152), .B(n115), .Q(n118) );
  IMUX21 U253 ( .A(n170), .B(n171), .S(n172), .Q(SUM[20]) );
  XNR21 U254 ( .A(B[20]), .B(A[20]), .Q(n171) );
  NOR21 U255 ( .A(n189), .B(n166), .Q(n170) );
  NAND22 U256 ( .A(n92), .B(n93), .Q(n91) );
  NAND22 U257 ( .A(n8), .B(n162), .Q(n148) );
  INV3 U258 ( .A(A[21]), .Q(n162) );
  INV3 U259 ( .A(B[21]), .Q(n8) );
  NAND22 U260 ( .A(n10), .B(n117), .Q(n90) );
  INV3 U261 ( .A(A[25]), .Q(n117) );
  NAND22 U262 ( .A(n7), .B(n200), .Q(n184) );
  INV3 U263 ( .A(A[18]), .Q(n200) );
  NAND22 U264 ( .A(n9), .B(n160), .Q(n142) );
  INV3 U265 ( .A(A[22]), .Q(n160) );
  NAND22 U266 ( .A(B[10]), .B(A[10]), .Q(n233) );
  OAI2111 U267 ( .A(n217), .B(n218), .C(n219), .D(n220), .Q(n216) );
  NAND22 U268 ( .A(B[9]), .B(A[9]), .Q(n15) );
  NOR21 U269 ( .A(A[10]), .B(B[10]), .Q(n240) );
  NAND22 U270 ( .A(B[11]), .B(A[11]), .Q(n229) );
  IMUX21 U271 ( .A(n267), .B(n268), .S(n269), .Q(SUM[12]) );
  NOR21 U272 ( .A(n278), .B(n279), .Q(n267) );
  NAND22 U273 ( .A(B[14]), .B(A[14]), .Q(n220) );
  NAND22 U274 ( .A(B[13]), .B(A[13]), .Q(n219) );
  NOR21 U275 ( .A(A[1]), .B(B[1]), .Q(n74) );
  AOI211 U276 ( .A(n297), .B(n298), .C(n74), .Q(n294) );
  NOR21 U277 ( .A(A[11]), .B(B[11]), .Q(n241) );
  NOR21 U278 ( .A(A[14]), .B(B[14]), .Q(n223) );
  NOR21 U279 ( .A(A[13]), .B(B[13]), .Q(n217) );
  NAND22 U280 ( .A(B[16]), .B(A[16]), .Q(n180) );
  NAND22 U281 ( .A(n213), .B(n214), .Q(n131) );
  NAND22 U282 ( .A(B[15]), .B(A[15]), .Q(n213) );
  NAND22 U283 ( .A(n215), .B(n216), .Q(n214) );
  AOI211 U284 ( .A(n221), .B(n222), .C(n223), .Q(n215) );
  NAND22 U285 ( .A(B[8]), .B(A[8]), .Q(n21) );
  NOR21 U286 ( .A(A[9]), .B(B[9]), .Q(n275) );
  NOR21 U287 ( .A(n301), .B(n302), .Q(n300) );
  NAND22 U288 ( .A(B[8]), .B(A[8]), .Q(n274) );
  XOR21 U289 ( .A(n22), .B(n23), .Q(SUM[7]) );
  AOI211 U290 ( .A(n24), .B(n25), .C(n26), .Q(n23) );
  NOR21 U291 ( .A(n19), .B(n20), .Q(n16) );
  XNR21 U292 ( .A(B[8]), .B(A[8]), .Q(n17) );
  NOR21 U293 ( .A(B[8]), .B(A[8]), .Q(n19) );
  IMUX21 U294 ( .A(n39), .B(n40), .S(n36), .Q(SUM[4]) );
  NOR21 U295 ( .A(n42), .B(n43), .Q(n39) );
  INV3 U296 ( .A(n83), .Q(n80) );
  INV3 U297 ( .A(n67), .Q(n64) );
  INV3 U298 ( .A(n58), .Q(n51) );
  INV3 U299 ( .A(B[15]), .Q(n221) );
  NAND22 U300 ( .A(n226), .B(n227), .Q(n134) );
  AOI311 U301 ( .A(n228), .B(n229), .C(n230), .D(n231), .Q(n227) );
  NAND22 U302 ( .A(B[8]), .B(A[8]), .Q(n228) );
  INV3 U303 ( .A(n116), .Q(n111) );
  INV3 U304 ( .A(A[15]), .Q(n222) );
  INV3 U305 ( .A(n203), .Q(n198) );
  NOR21 U306 ( .A(A[16]), .B(B[16]), .Q(n203) );
  INV3 U307 ( .A(B[0]), .Q(n316) );
  INV3 U308 ( .A(n318), .Q(n317) );
  NOR21 U309 ( .A(B[0]), .B(n293), .Q(n318) );
  NAND22 U310 ( .A(B[1]), .B(A[1]), .Q(n70) );
  NAND22 U311 ( .A(n45), .B(n46), .Q(n44) );
  NAND22 U312 ( .A(n47), .B(n48), .Q(n46) );
  INV3 U313 ( .A(n192), .Q(n72) );
  NAND22 U314 ( .A(B[0]), .B(A[0]), .Q(n192) );
  INV3 U315 ( .A(A[0]), .Q(n293) );
  CLKIN3 U316 ( .A(n21), .Q(n20) );
  CLKIN3 U317 ( .A(n27), .Q(n26) );
  CLKIN3 U318 ( .A(n32), .Q(n30) );
  OAI212 U319 ( .A(n36), .B(n37), .C(n38), .Q(n32) );
  CLKIN3 U320 ( .A(n38), .Q(n43) );
  CLKIN3 U321 ( .A(n65), .Q(n52) );
  CLKIN3 U322 ( .A(n45), .Q(n69) );
  CLKIN3 U323 ( .A(n81), .Q(n66) );
  CLKIN3 U324 ( .A(n97), .Q(n82) );
  CLKIN3 U325 ( .A(n110), .Q(n102) );
  CLKIN3 U326 ( .A(n53), .Q(n120) );
  CLKIN3 U327 ( .A(n131), .Q(n129) );
  CLKIN3 U328 ( .A(n132), .Q(n124) );
  OAI212 U329 ( .A(n138), .B(n139), .C(n140), .Q(n137) );
  CLKIN3 U330 ( .A(n144), .Q(n143) );
  OAI212 U331 ( .A(n145), .B(n146), .C(n147), .Q(n141) );
  CLKIN3 U332 ( .A(n108), .Q(n115) );
  OAI212 U333 ( .A(n156), .B(n147), .C(n144), .Q(n155) );
  CLKIN3 U334 ( .A(n147), .Q(n159) );
  OAI212 U335 ( .A(n176), .B(n177), .C(n178), .Q(n175) );
  CLKIN3 U336 ( .A(n184), .Q(n182) );
  CLKIN3 U337 ( .A(n146), .Q(n166) );
  CLKIN3 U338 ( .A(n70), .Q(n191) );
  OAI212 U339 ( .A(n183), .B(n197), .C(n181), .Q(n194) );
  CLKIN3 U340 ( .A(n130), .Q(n212) );
  CLKIN3 U341 ( .A(n243), .Q(n225) );
  CLKIN3 U342 ( .A(n180), .Q(n199) );
  CLKIN3 U343 ( .A(n220), .Q(n255) );
  OAI222 U344 ( .A(A[9]), .B(B[9]), .C(A[10]), .D(B[10]), .Q(n277) );
  OAI222 U345 ( .A(B[8]), .B(A[8]), .C(B[11]), .D(A[11]), .Q(n276) );
  CLKIN3 U346 ( .A(n263), .Q(n279) );
  OAI212 U347 ( .A(n18), .B(n287), .C(n21), .Q(n13) );
  CLKIN3 U348 ( .A(n270), .Q(n18) );
  CLKIN3 U349 ( .A(n308), .Q(n224) );
  CLKIN3 U350 ( .A(n309), .Q(n242) );
  OAI212 U351 ( .A(A[0]), .B(n316), .C(n317), .Q(SUM[0]) );
endmodule


module D_pcadd ( i_addr_pcadd4E, i_data_immshiftl, o_addr_pcbranchE );
  input [31:0] i_addr_pcadd4E;
  input [31:0] i_data_immshiftl;
  output [31:0] o_addr_pcbranchE;
  wire   n1;

  D_pcadd_DW01_add_1 add_5 ( .A(i_addr_pcadd4E), .B(i_data_immshiftl), .CI(n1), 
        .SUM(o_addr_pcbranchE) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_addr_Rt, i_con_RegWr, 
        i_addr_Rd, i_data_Rd, o_data_Rs, o_data_Rt );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rt;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr;
  wire   n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1, n2, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987;
  wire   [1023:0] regs;

  DFEC1 regs_reg_30__31_ ( .D(i_data_Rd[31]), .E(n1960), .C(i_clk), .RN(n1934), 
        .Q(regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(n1926), .E(n1960), .C(i_clk), .RN(n1934), .Q(
        regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(i_data_Rd[29]), .E(n1960), .C(i_clk), .RN(n1934), 
        .Q(regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(i_data_Rd[28]), .E(n1960), .C(i_clk), .RN(n1934), 
        .Q(regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(i_data_Rd[27]), .E(n1960), .C(i_clk), .RN(n1935), 
        .Q(regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(i_data_Rd[26]), .E(n1960), .C(i_clk), .RN(n1935), 
        .Q(regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(i_data_Rd[25]), .E(n1960), .C(i_clk), .RN(n1935), 
        .Q(regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(i_data_Rd[24]), .E(n1960), .C(i_clk), .RN(n1935), 
        .Q(regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(i_data_Rd[23]), .E(n1960), .C(i_clk), .RN(n1935), 
        .Q(regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(i_data_Rd[22]), .E(n1960), .C(i_clk), .RN(n1935), 
        .Q(regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(i_data_Rd[21]), .E(n1960), .C(i_clk), .RN(n1935), 
        .Q(regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(i_data_Rd[20]), .E(n1960), .C(i_clk), .RN(n1935), 
        .Q(regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n1960), .C(i_clk), .RN(n1935), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(i_data_Rd[18]), .E(n1960), .C(i_clk), .RN(n1936), 
        .Q(regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(i_data_Rd[17]), .E(n1960), .C(i_clk), .RN(n1936), 
        .Q(regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(i_data_Rd[16]), .E(n1960), .C(i_clk), .RN(n1936), 
        .Q(regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(n1881), .E(n1960), .C(i_clk), .RN(n1936), .Q(
        regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(n1877), .E(n1960), .C(i_clk), .RN(n1936), .Q(
        regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(n1873), .E(n1960), .C(i_clk), .RN(n1936), .Q(
        regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(n1869), .E(n1960), .C(i_clk), .RN(n1936), .Q(
        regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(n1865), .E(n1960), .C(i_clk), .RN(n1936), .Q(
        regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(n1861), .E(n1960), .C(i_clk), .RN(n1936), .Q(
        regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(n1857), .E(n1960), .C(i_clk), .RN(n1937), .Q(
        regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(n1853), .E(n1960), .C(i_clk), .RN(n1937), .Q(
        regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(n1849), .E(n1960), .C(i_clk), .RN(n1937), .Q(
        regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n1960), .C(i_clk), .RN(n1937), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(i_data_Rd[5]), .E(n1960), .C(i_clk), .RN(n1937), 
        .Q(regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(n1839), .E(n1960), .C(i_clk), .RN(n1937), .Q(
        regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(i_data_Rd[3]), .E(n1960), .C(i_clk), .RN(n1937), 
        .Q(regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(i_data_Rd[2]), .E(n1960), .C(i_clk), .RN(n1937), 
        .Q(regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n1960), .C(i_clk), .RN(n1937), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(i_data_Rd[0]), .E(n1960), .C(i_clk), .RN(n1938), 
        .Q(regs[960]) );
  DFEC1 regs_reg_26__31_ ( .D(i_data_Rd[31]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(n1926), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(i_data_Rd[29]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(i_data_Rd[28]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(i_data_Rd[27]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(i_data_Rd[26]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(i_data_Rd[25]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(i_data_Rd[24]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(i_data_Rd[23]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(i_data_Rd[22]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(i_data_Rd[21]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(i_data_Rd[20]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(i_data_Rd[18]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(i_data_Rd[17]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(i_data_Rd[16]), .E(n1964), .C(i_clk), .RN(
        i_rst_n), .Q(regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(n1881), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(n1877), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(n1873), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(n1869), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(n1865), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(n1861), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(n1857), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(n1853), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(n1849), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n1964), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(i_data_Rd[5]), .E(n1964), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(n1839), .E(n1964), .C(i_clk), .RN(i_rst_n), .Q(
        regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(i_data_Rd[3]), .E(n1964), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(i_data_Rd[2]), .E(n1964), .C(i_clk), .RN(n1938), 
        .Q(regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n1964), .C(i_clk), .RN(n1939), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(i_data_Rd[0]), .E(n1964), .C(i_clk), .RN(n1931), 
        .Q(regs[832]) );
  DFEC1 regs_reg_22__31_ ( .D(n1929), .E(n1952), .C(i_clk), .RN(n1945), .Q(
        regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(i_data_Rd[30]), .E(n1952), .C(i_clk), .RN(n1931), 
        .Q(regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(n1923), .E(n1952), .C(i_clk), .RN(n1932), .Q(
        regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(n1920), .E(n1952), .C(i_clk), .RN(n1933), .Q(
        regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(n1917), .E(n1952), .C(i_clk), .RN(n1934), .Q(
        regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(n1914), .E(n1952), .C(i_clk), .RN(n1935), .Q(
        regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(n1911), .E(n1952), .C(i_clk), .RN(n1936), .Q(
        regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(n1908), .E(n1952), .C(i_clk), .RN(n1937), .Q(
        regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(n1905), .E(n1952), .C(i_clk), .RN(n1938), .Q(
        regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(n1902), .E(n1952), .C(i_clk), .RN(n1942), .Q(
        regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(n1899), .E(n1952), .C(i_clk), .RN(n1943), .Q(
        regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(n1896), .E(n1952), .C(i_clk), .RN(n1944), .Q(
        regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(n1893), .E(n1952), .C(i_clk), .RN(n1945), .Q(
        regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(n1890), .E(n1952), .C(i_clk), .RN(n1931), .Q(
        regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(n1887), .E(n1952), .C(i_clk), .RN(n1932), .Q(
        regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(n1884), .E(n1952), .C(i_clk), .RN(n1933), .Q(
        regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(n1880), .E(n1952), .C(i_clk), .RN(n1934), .Q(
        regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(n1876), .E(n1952), .C(i_clk), .RN(n1935), .Q(
        regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(n1872), .E(n1952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(n1868), .E(n1952), .C(i_clk), .RN(n1950), .Q(
        regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(n1864), .E(n1952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(n1860), .E(n1952), .C(i_clk), .RN(n1947), .Q(
        regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(n1856), .E(n1952), .C(i_clk), .RN(n1937), .Q(
        regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(n1852), .E(n1952), .C(i_clk), .RN(n1949), .Q(
        regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(n1848), .E(n1952), .C(i_clk), .RN(n1948), .Q(
        regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(n1845), .E(n1952), .C(i_clk), .RN(n1947), .Q(
        regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(n1842), .E(n1952), .C(i_clk), .RN(i_rst_n), .Q(
        regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(i_data_Rd[4]), .E(n1952), .C(i_clk), .RN(n1936), 
        .Q(regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(n1836), .E(n1952), .C(i_clk), .RN(n1937), .Q(
        regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(n1833), .E(n1952), .C(i_clk), .RN(n1938), .Q(
        regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(n1830), .E(n1952), .C(i_clk), .RN(n1939), .Q(
        regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(n1827), .E(n1952), .C(i_clk), .RN(n1940), .Q(
        regs[704]) );
  DFEC1 regs_reg_18__31_ ( .D(n1929), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(i_data_Rd[30]), .E(n1956), .C(i_clk), .RN(
        i_rst_n), .Q(regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(n1923), .E(n1956), .C(i_clk), .RN(n1945), .Q(
        regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(n1920), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(n1917), .E(n1956), .C(i_clk), .RN(n1934), .Q(
        regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(n1914), .E(n1956), .C(i_clk), .RN(n1935), .Q(
        regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(n1911), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(n1908), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(n1905), .E(n1956), .C(i_clk), .RN(n1942), .Q(
        regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(n1902), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(n1899), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(n1896), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(n1893), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(n1890), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(n1887), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(n1884), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(n1880), .E(n1956), .C(i_clk), .RN(n1941), .Q(
        regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(n1876), .E(n1956), .C(i_clk), .RN(n1939), .Q(
        regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(n1872), .E(n1956), .C(i_clk), .RN(n1947), .Q(
        regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(n1868), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(n1864), .E(n1956), .C(i_clk), .RN(n1949), .Q(
        regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(n1860), .E(n1956), .C(i_clk), .RN(n1948), .Q(
        regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(n1856), .E(n1956), .C(i_clk), .RN(n1947), .Q(
        regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(n1852), .E(n1956), .C(i_clk), .RN(n1950), .Q(
        regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(n1848), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(n1845), .E(n1956), .C(i_clk), .RN(n1942), .Q(
        regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(n1842), .E(n1956), .C(i_clk), .RN(n1932), .Q(
        regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(i_data_Rd[4]), .E(n1956), .C(i_clk), .RN(n1933), 
        .Q(regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(n1836), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(n1833), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(n1830), .E(n1956), .C(i_clk), .RN(i_rst_n), .Q(
        regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(n1827), .E(n1956), .C(i_clk), .RN(n1939), .Q(
        regs[576]) );
  DFEC1 regs_reg_14__31_ ( .D(n1928), .E(n1969), .C(i_clk), .RN(n1942), .Q(
        regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(n1925), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(n1922), .E(n1969), .C(i_clk), .RN(n1950), .Q(
        regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(n1919), .E(n1969), .C(i_clk), .RN(n1950), .Q(
        regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(n1916), .E(n1969), .C(i_clk), .RN(n1938), .Q(
        regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(n1913), .E(n1969), .C(i_clk), .RN(n1947), .Q(
        regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(n1910), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(n1907), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(n1904), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(n1901), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(n1898), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(n1895), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(n1892), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(n1889), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(n1886), .E(n1969), .C(i_clk), .RN(n1930), .Q(
        regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(n1883), .E(n1969), .C(i_clk), .RN(n1946), .Q(
        regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(n1879), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(n1875), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(n1871), .E(n1969), .C(i_clk), .RN(n1946), .Q(
        regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(n1867), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(n1863), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(n1859), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(n1855), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(n1851), .E(n1969), .C(i_clk), .RN(n1948), .Q(
        regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(n1847), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(n1844), .E(n1969), .C(i_clk), .RN(n1938), .Q(
        regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(n1841), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(n1838), .E(n1969), .C(i_clk), .RN(n1948), .Q(
        regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(n1835), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(n1832), .E(n1969), .C(i_clk), .RN(i_rst_n), .Q(
        regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(n1829), .E(n1969), .C(i_clk), .RN(n1936), .Q(
        regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(n1826), .E(n1969), .C(i_clk), .RN(n1934), .Q(
        regs[448]) );
  DFEC1 regs_reg_10__31_ ( .D(n1928), .E(n1973), .C(i_clk), .RN(n1940), .Q(
        regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(n1925), .E(n1973), .C(i_clk), .RN(n1950), .Q(
        regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(n1922), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(n1919), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(n1916), .E(n1973), .C(i_clk), .RN(n1939), .Q(
        regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(n1913), .E(n1973), .C(i_clk), .RN(n1930), .Q(
        regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(n1910), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(n1907), .E(n1973), .C(i_clk), .RN(n1950), .Q(
        regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(n1904), .E(n1973), .C(i_clk), .RN(n1949), .Q(
        regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(n1901), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(n1898), .E(n1973), .C(i_clk), .RN(n1937), .Q(
        regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(n1895), .E(n1973), .C(i_clk), .RN(n1949), .Q(
        regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(n1892), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(n1889), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(n1886), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(n1883), .E(n1973), .C(i_clk), .RN(n1950), .Q(
        regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(n1879), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(n1875), .E(n1973), .C(i_clk), .RN(n1930), .Q(
        regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(n1871), .E(n1973), .C(i_clk), .RN(n1941), .Q(
        regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(n1867), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(n1863), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(n1859), .E(n1973), .C(i_clk), .RN(n1949), .Q(
        regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(n1855), .E(n1973), .C(i_clk), .RN(n1944), .Q(
        regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(n1851), .E(n1973), .C(i_clk), .RN(n1942), .Q(
        regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(n1847), .E(n1973), .C(i_clk), .RN(n1940), .Q(
        regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(n1844), .E(n1973), .C(i_clk), .RN(n1930), .Q(
        regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(n1841), .E(n1973), .C(i_clk), .RN(n1944), .Q(
        regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(n1838), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(n1835), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(n1832), .E(n1973), .C(i_clk), .RN(n1935), .Q(
        regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(n1829), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(n1826), .E(n1973), .C(i_clk), .RN(i_rst_n), .Q(
        regs[320]) );
  DFEC1 regs_reg_6__31_ ( .D(n1927), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(n1924), .E(n1977), .C(i_clk), .RN(n1950), .Q(
        regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(n1921), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(n1918), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(n1915), .E(n1977), .C(i_clk), .RN(n1943), .Q(
        regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(n1912), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(n1909), .E(n1977), .C(i_clk), .RN(n1936), .Q(
        regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(n1906), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(n1903), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(n1900), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(n1897), .E(n1977), .C(i_clk), .RN(n1947), .Q(
        regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(n1894), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(n1891), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(n1888), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(n1885), .E(n1977), .C(i_clk), .RN(n1939), .Q(
        regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(n1882), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(n1878), .E(n1977), .C(i_clk), .RN(n1942), .Q(
        regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(n1874), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(n1870), .E(n1977), .C(i_clk), .RN(n1950), .Q(
        regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(n1866), .E(n1977), .C(i_clk), .RN(n1948), .Q(
        regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(n1862), .E(n1977), .C(i_clk), .RN(n1944), .Q(
        regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(n1858), .E(n1977), .C(i_clk), .RN(n1945), .Q(
        regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(n1854), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(n1850), .E(n1977), .C(i_clk), .RN(n1949), .Q(
        regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(n1846), .E(n1977), .C(i_clk), .RN(n1948), .Q(
        regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(n1843), .E(n1977), .C(i_clk), .RN(n1947), .Q(
        regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(n1840), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(n1837), .E(n1977), .C(i_clk), .RN(i_rst_n), .Q(
        regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(n1834), .E(n1977), .C(i_clk), .RN(n1942), .Q(
        regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(n1831), .E(n1977), .C(i_clk), .RN(n1933), .Q(
        regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(n1828), .E(n1977), .C(i_clk), .RN(n1931), .Q(
        regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(n1825), .E(n1977), .C(i_clk), .RN(n1932), .Q(
        regs[192]) );
  DFEC1 regs_reg_2__31_ ( .D(n1927), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(n1924), .E(n1981), .C(i_clk), .RN(n1932), .Q(
        regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(n1921), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(n1918), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(n1915), .E(n1981), .C(i_clk), .RN(n1932), .Q(
        regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(n1912), .E(n1981), .C(i_clk), .RN(n1945), .Q(
        regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(n1909), .E(n1981), .C(i_clk), .RN(n1933), .Q(
        regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(n1906), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(n1903), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(n1900), .E(n1981), .C(i_clk), .RN(n1941), .Q(
        regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(n1897), .E(n1981), .C(i_clk), .RN(n1946), .Q(
        regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(n1894), .E(n1981), .C(i_clk), .RN(n1944), .Q(
        regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(n1891), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(n1888), .E(n1981), .C(i_clk), .RN(n1930), .Q(
        regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(n1885), .E(n1981), .C(i_clk), .RN(n1946), .Q(
        regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(n1882), .E(n1981), .C(i_clk), .RN(n1946), .Q(
        regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(n1878), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(n1874), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(n1870), .E(n1981), .C(i_clk), .RN(n1941), .Q(
        regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(n1866), .E(n1981), .C(i_clk), .RN(n1940), .Q(
        regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(n1862), .E(n1981), .C(i_clk), .RN(n1948), .Q(
        regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(n1858), .E(n1981), .C(i_clk), .RN(n1930), .Q(
        regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(n1854), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(n1850), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(n1846), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(n1843), .E(n1981), .C(i_clk), .RN(n1947), .Q(
        regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(n1840), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(n1837), .E(n1981), .C(i_clk), .RN(n1930), .Q(
        regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(n1834), .E(n1981), .C(i_clk), .RN(n1947), .Q(
        regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(n1831), .E(n1981), .C(i_clk), .RN(n1940), .Q(
        regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(n1828), .E(n1981), .C(i_clk), .RN(i_rst_n), .Q(
        regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(n1825), .E(n1981), .C(i_clk), .RN(n1939), .Q(
        regs[64]) );
  DFEC1 regs_reg_31__31_ ( .D(i_data_Rd[31]), .E(n1959), .C(i_clk), .RN(n1931), 
        .Q(regs[1023]) );
  DFEC1 regs_reg_31__30_ ( .D(n1926), .E(n1959), .C(i_clk), .RN(n1931), .Q(
        regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(i_data_Rd[29]), .E(n1959), .C(i_clk), .RN(n1931), 
        .Q(regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(i_data_Rd[28]), .E(n1959), .C(i_clk), .RN(n1931), 
        .Q(regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(i_data_Rd[27]), .E(n1959), .C(i_clk), .RN(n1931), 
        .Q(regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(i_data_Rd[26]), .E(n1959), .C(i_clk), .RN(n1931), 
        .Q(regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(i_data_Rd[25]), .E(n1959), .C(i_clk), .RN(n1931), 
        .Q(regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(i_data_Rd[24]), .E(n1959), .C(i_clk), .RN(n1931), 
        .Q(regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(i_data_Rd[23]), .E(n1959), .C(i_clk), .RN(n1931), 
        .Q(regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(i_data_Rd[22]), .E(n1959), .C(i_clk), .RN(n1932), 
        .Q(regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(i_data_Rd[21]), .E(n1959), .C(i_clk), .RN(n1932), 
        .Q(regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(i_data_Rd[20]), .E(n1959), .C(i_clk), .RN(n1932), 
        .Q(regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n1959), .C(i_clk), .RN(n1932), 
        .Q(regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(i_data_Rd[18]), .E(n1959), .C(i_clk), .RN(n1932), 
        .Q(regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(i_data_Rd[17]), .E(n1959), .C(i_clk), .RN(n1932), 
        .Q(regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(i_data_Rd[16]), .E(n1959), .C(i_clk), .RN(n1932), 
        .Q(regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(n1881), .E(n1959), .C(i_clk), .RN(n1932), .Q(
        regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(n1877), .E(n1959), .C(i_clk), .RN(n1932), .Q(
        regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(n1873), .E(n1959), .C(i_clk), .RN(n1933), .Q(
        regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(n1869), .E(n1959), .C(i_clk), .RN(n1933), .Q(
        regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(n1865), .E(n1959), .C(i_clk), .RN(n1933), .Q(
        regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(n1861), .E(n1959), .C(i_clk), .RN(n1933), .Q(
        regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(n1857), .E(n1959), .C(i_clk), .RN(n1933), .Q(
        regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(n1853), .E(n1959), .C(i_clk), .RN(n1933), .Q(
        regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(n1849), .E(n1959), .C(i_clk), .RN(n1933), .Q(
        regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n1959), .C(i_clk), .RN(n1933), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(i_data_Rd[5]), .E(n1959), .C(i_clk), .RN(n1933), 
        .Q(regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(n1839), .E(n1959), .C(i_clk), .RN(n1934), .Q(
        regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(i_data_Rd[3]), .E(n1959), .C(i_clk), .RN(n1934), 
        .Q(regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(i_data_Rd[2]), .E(n1959), .C(i_clk), .RN(n1934), 
        .Q(regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n1959), .C(i_clk), .RN(n1934), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(i_data_Rd[0]), .E(n1959), .C(i_clk), .RN(n1934), 
        .Q(regs[992]) );
  DFEC1 regs_reg_29__31_ ( .D(i_data_Rd[31]), .E(n1961), .C(i_clk), .RN(n1938), 
        .Q(regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(n1926), .E(n1961), .C(i_clk), .RN(n1938), .Q(
        regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(i_data_Rd[29]), .E(n1961), .C(i_clk), .RN(n1938), 
        .Q(regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(i_data_Rd[28]), .E(n1961), .C(i_clk), .RN(n1938), 
        .Q(regs[956]) );
  DFEC1 regs_reg_29__27_ ( .D(i_data_Rd[27]), .E(n1961), .C(i_clk), .RN(n1938), 
        .Q(regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(i_data_Rd[26]), .E(n1961), .C(i_clk), .RN(n1938), 
        .Q(regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(i_data_Rd[25]), .E(n1961), .C(i_clk), .RN(n1938), 
        .Q(regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(i_data_Rd[24]), .E(n1961), .C(i_clk), .RN(n1938), 
        .Q(regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(i_data_Rd[23]), .E(n1961), .C(i_clk), .RN(n1939), 
        .Q(regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(i_data_Rd[22]), .E(n1961), .C(i_clk), .RN(n1939), 
        .Q(regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(i_data_Rd[21]), .E(n1961), .C(i_clk), .RN(n1939), 
        .Q(regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(i_data_Rd[20]), .E(n1961), .C(i_clk), .RN(n1939), 
        .Q(regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n1961), .C(i_clk), .RN(n1939), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(i_data_Rd[18]), .E(n1961), .C(i_clk), .RN(n1939), 
        .Q(regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(i_data_Rd[17]), .E(n1961), .C(i_clk), .RN(n1939), 
        .Q(regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(i_data_Rd[16]), .E(n1961), .C(i_clk), .RN(n1939), 
        .Q(regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(n1881), .E(n1961), .C(i_clk), .RN(n1939), .Q(
        regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(n1877), .E(n1961), .C(i_clk), .RN(n1940), .Q(
        regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(n1873), .E(n1961), .C(i_clk), .RN(n1940), .Q(
        regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(n1869), .E(n1961), .C(i_clk), .RN(n1940), .Q(
        regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(n1865), .E(n1961), .C(i_clk), .RN(n1940), .Q(
        regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(n1861), .E(n1961), .C(i_clk), .RN(n1940), .Q(
        regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(n1857), .E(n1961), .C(i_clk), .RN(n1940), .Q(
        regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(n1853), .E(n1961), .C(i_clk), .RN(n1940), .Q(
        regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(n1849), .E(n1961), .C(i_clk), .RN(n1940), .Q(
        regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n1961), .C(i_clk), .RN(n1940), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(i_data_Rd[5]), .E(n1961), .C(i_clk), .RN(n1941), 
        .Q(regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(n1839), .E(n1961), .C(i_clk), .RN(n1941), .Q(
        regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(i_data_Rd[3]), .E(n1961), .C(i_clk), .RN(n1941), 
        .Q(regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(i_data_Rd[2]), .E(n1961), .C(i_clk), .RN(n1941), 
        .Q(regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n1961), .C(i_clk), .RN(n1941), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(i_data_Rd[0]), .E(n1961), .C(i_clk), .RN(n1941), 
        .Q(regs[928]) );
  DFEC1 regs_reg_28__31_ ( .D(i_data_Rd[31]), .E(n1962), .C(i_clk), .RN(n1941), 
        .Q(regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(n1926), .E(n1962), .C(i_clk), .RN(n1941), .Q(
        regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(i_data_Rd[29]), .E(n1962), .C(i_clk), .RN(n1941), 
        .Q(regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(i_data_Rd[28]), .E(n1962), .C(i_clk), .RN(
        i_rst_n), .Q(regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(i_data_Rd[27]), .E(n1962), .C(i_clk), .RN(
        i_rst_n), .Q(regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(i_data_Rd[26]), .E(n1962), .C(i_clk), .RN(
        i_rst_n), .Q(regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(i_data_Rd[25]), .E(n1962), .C(i_clk), .RN(
        i_rst_n), .Q(regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(i_data_Rd[24]), .E(n1962), .C(i_clk), .RN(
        i_rst_n), .Q(regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(i_data_Rd[23]), .E(n1962), .C(i_clk), .RN(
        i_rst_n), .Q(regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(i_data_Rd[22]), .E(n1962), .C(i_clk), .RN(
        i_rst_n), .Q(regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(i_data_Rd[21]), .E(n1962), .C(i_clk), .RN(
        i_rst_n), .Q(regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(i_data_Rd[20]), .E(n1962), .C(i_clk), .RN(
        i_rst_n), .Q(regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n1962), .C(i_clk), .RN(n1942), 
        .Q(regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(i_data_Rd[18]), .E(n1962), .C(i_clk), .RN(n1942), 
        .Q(regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(i_data_Rd[17]), .E(n1962), .C(i_clk), .RN(n1942), 
        .Q(regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(i_data_Rd[16]), .E(n1962), .C(i_clk), .RN(n1942), 
        .Q(regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(n1881), .E(n1962), .C(i_clk), .RN(n1942), .Q(
        regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(n1877), .E(n1962), .C(i_clk), .RN(n1942), .Q(
        regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(n1873), .E(n1962), .C(i_clk), .RN(n1942), .Q(
        regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(n1869), .E(n1962), .C(i_clk), .RN(n1942), .Q(
        regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(n1865), .E(n1962), .C(i_clk), .RN(n1942), .Q(
        regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(n1861), .E(n1962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(n1857), .E(n1962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(n1853), .E(n1962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(n1849), .E(n1962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n1962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(i_data_Rd[5]), .E(n1962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(n1839), .E(n1962), .C(i_clk), .RN(i_rst_n), .Q(
        regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(i_data_Rd[3]), .E(n1962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(i_data_Rd[2]), .E(n1962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n1962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(i_data_Rd[0]), .E(n1962), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(i_data_Rd[31]), .E(n1963), .C(i_clk), .RN(n1943), 
        .Q(regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(n1926), .E(n1963), .C(i_clk), .RN(n1942), .Q(
        regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(i_data_Rd[29]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(i_data_Rd[28]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(i_data_Rd[27]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(i_data_Rd[26]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(i_data_Rd[25]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(i_data_Rd[24]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(i_data_Rd[23]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(i_data_Rd[22]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(i_data_Rd[21]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(i_data_Rd[20]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(i_data_Rd[18]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(i_data_Rd[17]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(i_data_Rd[16]), .E(n1963), .C(i_clk), .RN(
        i_rst_n), .Q(regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(n1881), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(n1877), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(n1873), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(n1869), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(n1865), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(n1861), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(n1857), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(n1853), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(n1849), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n1963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(i_data_Rd[5]), .E(n1963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(n1839), .E(n1963), .C(i_clk), .RN(i_rst_n), .Q(
        regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(i_data_Rd[3]), .E(n1963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(i_data_Rd[2]), .E(n1963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(i_data_Rd[1]), .E(n1963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(i_data_Rd[0]), .E(n1963), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[864]) );
  DFEC1 regs_reg_25__31_ ( .D(i_data_Rd[31]), .E(n1965), .C(i_clk), .RN(n1932), 
        .Q(regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(n1926), .E(n1965), .C(i_clk), .RN(n1933), .Q(
        regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(i_data_Rd[29]), .E(n1965), .C(i_clk), .RN(n1934), 
        .Q(regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(i_data_Rd[28]), .E(n1965), .C(i_clk), .RN(n1935), 
        .Q(regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(i_data_Rd[27]), .E(n1965), .C(i_clk), .RN(n1936), 
        .Q(regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(i_data_Rd[26]), .E(n1965), .C(i_clk), .RN(n1940), 
        .Q(regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(i_data_Rd[25]), .E(n1965), .C(i_clk), .RN(
        i_rst_n), .Q(regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(i_data_Rd[24]), .E(n1965), .C(i_clk), .RN(
        i_rst_n), .Q(regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(i_data_Rd[23]), .E(n1965), .C(i_clk), .RN(
        i_rst_n), .Q(regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(i_data_Rd[22]), .E(n1965), .C(i_clk), .RN(
        i_rst_n), .Q(regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(i_data_Rd[21]), .E(n1965), .C(i_clk), .RN(
        i_rst_n), .Q(regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(i_data_Rd[20]), .E(n1965), .C(i_clk), .RN(n1949), 
        .Q(regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(i_data_Rd[19]), .E(n1965), .C(i_clk), .RN(
        i_rst_n), .Q(regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(i_data_Rd[18]), .E(n1965), .C(i_clk), .RN(
        i_rst_n), .Q(regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(i_data_Rd[17]), .E(n1965), .C(i_clk), .RN(n1950), 
        .Q(regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(i_data_Rd[16]), .E(n1965), .C(i_clk), .RN(
        i_rst_n), .Q(regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(n1881), .E(n1965), .C(i_clk), .RN(n1947), .Q(
        regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(n1877), .E(n1965), .C(i_clk), .RN(n1944), .Q(
        regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(n1873), .E(n1965), .C(i_clk), .RN(n1937), .Q(
        regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(n1869), .E(n1965), .C(i_clk), .RN(n1938), .Q(
        regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(n1865), .E(n1965), .C(i_clk), .RN(n1939), .Q(
        regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(n1861), .E(n1965), .C(i_clk), .RN(n1931), .Q(
        regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(n1857), .E(n1965), .C(i_clk), .RN(n1932), .Q(
        regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(n1853), .E(n1965), .C(i_clk), .RN(n1933), .Q(
        regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(n1849), .E(n1965), .C(i_clk), .RN(n1947), .Q(
        regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(i_data_Rd[6]), .E(n1965), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(i_data_Rd[5]), .E(n1965), .C(i_clk), .RN(n1931), 
        .Q(regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(n1839), .E(n1965), .C(i_clk), .RN(n1932), .Q(
        regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(i_data_Rd[3]), .E(n1965), .C(i_clk), .RN(n1943), 
        .Q(regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(i_data_Rd[2]), .E(n1965), .C(i_clk), .RN(n1944), 
        .Q(regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(i_data_Rd[1]), .E(n1965), .C(i_clk), .RN(n1945), 
        .Q(regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(i_data_Rd[0]), .E(n1965), .C(i_clk), .RN(n1942), 
        .Q(regs[800]) );
  DFEC1 regs_reg_24__31_ ( .D(i_data_Rd[31]), .E(n1966), .C(i_clk), .RN(
        i_rst_n), .Q(regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(n1926), .E(n1966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(i_data_Rd[29]), .E(n1966), .C(i_clk), .RN(
        i_rst_n), .Q(regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(i_data_Rd[28]), .E(n1966), .C(i_clk), .RN(n1937), 
        .Q(regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(i_data_Rd[27]), .E(n1966), .C(i_clk), .RN(n1930), 
        .Q(regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(i_data_Rd[26]), .E(n1966), .C(i_clk), .RN(n1938), 
        .Q(regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(i_data_Rd[25]), .E(n1966), .C(i_clk), .RN(
        i_rst_n), .Q(regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(i_data_Rd[24]), .E(n1966), .C(i_clk), .RN(n1950), 
        .Q(regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(i_data_Rd[23]), .E(n1966), .C(i_clk), .RN(n1949), 
        .Q(regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(i_data_Rd[22]), .E(n1966), .C(i_clk), .RN(n1948), 
        .Q(regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(i_data_Rd[21]), .E(n1966), .C(i_clk), .RN(n1939), 
        .Q(regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(i_data_Rd[20]), .E(n1966), .C(i_clk), .RN(n1931), 
        .Q(regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(i_data_Rd[19]), .E(n1966), .C(i_clk), .RN(n1932), 
        .Q(regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(i_data_Rd[18]), .E(n1966), .C(i_clk), .RN(n1933), 
        .Q(regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(i_data_Rd[17]), .E(n1966), .C(i_clk), .RN(n1934), 
        .Q(regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(i_data_Rd[16]), .E(n1966), .C(i_clk), .RN(n1935), 
        .Q(regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(n1881), .E(n1966), .C(i_clk), .RN(n1936), .Q(
        regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(n1877), .E(n1966), .C(i_clk), .RN(n1940), .Q(
        regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(n1873), .E(n1966), .C(i_clk), .RN(n1941), .Q(
        regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(n1869), .E(n1966), .C(i_clk), .RN(n1931), .Q(
        regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(n1865), .E(n1966), .C(i_clk), .RN(n1932), .Q(
        regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(n1861), .E(n1966), .C(i_clk), .RN(n1933), .Q(
        regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(n1857), .E(n1966), .C(i_clk), .RN(n1934), .Q(
        regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(n1853), .E(n1966), .C(i_clk), .RN(n1935), .Q(
        regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(n1849), .E(n1966), .C(i_clk), .RN(n1936), .Q(
        regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(i_data_Rd[6]), .E(n1966), .C(i_clk), .RN(n1940), 
        .Q(regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(i_data_Rd[5]), .E(n1966), .C(i_clk), .RN(n1941), 
        .Q(regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(n1839), .E(n1966), .C(i_clk), .RN(i_rst_n), .Q(
        regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(i_data_Rd[3]), .E(n1966), .C(i_clk), .RN(n1947), 
        .Q(regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(i_data_Rd[2]), .E(n1966), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(i_data_Rd[1]), .E(n1966), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(i_data_Rd[0]), .E(n1966), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(n1929), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(i_data_Rd[30]), .E(n1951), .C(i_clk), .RN(
        i_rst_n), .Q(regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(n1923), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(n1920), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(n1917), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(n1914), .E(n1951), .C(i_clk), .RN(n1931), .Q(
        regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(n1911), .E(n1951), .C(i_clk), .RN(n1932), .Q(
        regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(n1908), .E(n1951), .C(i_clk), .RN(n1933), .Q(
        regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(n1905), .E(n1951), .C(i_clk), .RN(n1934), .Q(
        regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(n1902), .E(n1951), .C(i_clk), .RN(n1935), .Q(
        regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(n1899), .E(n1951), .C(i_clk), .RN(n1936), .Q(
        regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(n1896), .E(n1951), .C(i_clk), .RN(n1937), .Q(
        regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(n1893), .E(n1951), .C(i_clk), .RN(n1938), .Q(
        regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(n1890), .E(n1951), .C(i_clk), .RN(n1939), .Q(
        regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(n1887), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(n1884), .E(n1951), .C(i_clk), .RN(n1944), .Q(
        regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(n1880), .E(n1951), .C(i_clk), .RN(n1946), .Q(
        regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(n1876), .E(n1951), .C(i_clk), .RN(n1944), .Q(
        regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(n1872), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(n1868), .E(n1951), .C(i_clk), .RN(n1942), .Q(
        regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(n1864), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(n1860), .E(n1951), .C(i_clk), .RN(n1947), .Q(
        regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(n1856), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(n1852), .E(n1951), .C(i_clk), .RN(n1946), .Q(
        regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(n1848), .E(n1951), .C(i_clk), .RN(n1949), .Q(
        regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(n1845), .E(n1951), .C(i_clk), .RN(n1948), .Q(
        regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(n1842), .E(n1951), .C(i_clk), .RN(n1947), .Q(
        regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(i_data_Rd[4]), .E(n1951), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(n1836), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(n1833), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(n1830), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(n1827), .E(n1951), .C(i_clk), .RN(i_rst_n), .Q(
        regs[736]) );
  DFEC1 regs_reg_21__31_ ( .D(n1929), .E(n1953), .C(i_clk), .RN(n1941), .Q(
        regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(i_data_Rd[30]), .E(n1953), .C(i_clk), .RN(
        i_rst_n), .Q(regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(n1923), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(n1920), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(n1917), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(n1914), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(n1911), .E(n1953), .C(i_clk), .RN(n1945), .Q(
        regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(n1908), .E(n1953), .C(i_clk), .RN(n1933), .Q(
        regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(n1905), .E(n1953), .C(i_clk), .RN(n1945), .Q(
        regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(n1902), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(n1899), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(n1896), .E(n1953), .C(i_clk), .RN(n1930), .Q(
        regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(n1893), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(n1890), .E(n1953), .C(i_clk), .RN(n1940), .Q(
        regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(n1887), .E(n1953), .C(i_clk), .RN(n1950), .Q(
        regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(n1884), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(n1880), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(n1876), .E(n1953), .C(i_clk), .RN(n1948), .Q(
        regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(n1872), .E(n1953), .C(i_clk), .RN(n1939), .Q(
        regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(n1868), .E(n1953), .C(i_clk), .RN(n1946), .Q(
        regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(n1864), .E(n1953), .C(i_clk), .RN(n1949), .Q(
        regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(n1860), .E(n1953), .C(i_clk), .RN(n1948), .Q(
        regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(n1856), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(n1852), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(n1848), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(n1845), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(n1842), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(i_data_Rd[4]), .E(n1953), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(n1836), .E(n1953), .C(i_clk), .RN(n1942), .Q(
        regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(n1833), .E(n1953), .C(i_clk), .RN(n1943), .Q(
        regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(n1830), .E(n1953), .C(i_clk), .RN(i_rst_n), .Q(
        regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(n1827), .E(n1953), .C(i_clk), .RN(n1942), .Q(
        regs[672]) );
  DFEC1 regs_reg_20__31_ ( .D(n1929), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(i_data_Rd[30]), .E(n1954), .C(i_clk), .RN(
        i_rst_n), .Q(regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(n1923), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(n1920), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(n1917), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(n1914), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(n1911), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(n1908), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(n1905), .E(n1954), .C(i_clk), .RN(n1943), .Q(
        regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(n1902), .E(n1954), .C(i_clk), .RN(n1944), .Q(
        regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(n1899), .E(n1954), .C(i_clk), .RN(n1945), .Q(
        regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(n1896), .E(n1954), .C(i_clk), .RN(n1931), .Q(
        regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(n1893), .E(n1954), .C(i_clk), .RN(n1932), .Q(
        regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(n1890), .E(n1954), .C(i_clk), .RN(n1933), .Q(
        regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(n1887), .E(n1954), .C(i_clk), .RN(n1934), .Q(
        regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(n1884), .E(n1954), .C(i_clk), .RN(n1935), .Q(
        regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(n1880), .E(n1954), .C(i_clk), .RN(n1936), .Q(
        regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(n1876), .E(n1954), .C(i_clk), .RN(n1941), .Q(
        regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(n1872), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(n1868), .E(n1954), .C(i_clk), .RN(n1942), .Q(
        regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(n1864), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(n1860), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(n1856), .E(n1954), .C(i_clk), .RN(n1930), .Q(
        regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(n1852), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(n1848), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(n1845), .E(n1954), .C(i_clk), .RN(n1946), .Q(
        regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(n1842), .E(n1954), .C(i_clk), .RN(i_rst_n), .Q(
        regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(i_data_Rd[4]), .E(n1954), .C(i_clk), .RN(n1931), 
        .Q(regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(n1836), .E(n1954), .C(i_clk), .RN(n1932), .Q(
        regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(n1833), .E(n1954), .C(i_clk), .RN(n1933), .Q(
        regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(n1830), .E(n1954), .C(i_clk), .RN(n1934), .Q(
        regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(n1827), .E(n1954), .C(i_clk), .RN(n1935), .Q(
        regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(n1929), .E(n1955), .C(i_clk), .RN(n1936), .Q(
        regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(i_data_Rd[30]), .E(n1955), .C(i_clk), .RN(n1937), 
        .Q(regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(n1923), .E(n1955), .C(i_clk), .RN(n1938), .Q(
        regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(n1920), .E(n1955), .C(i_clk), .RN(n1949), .Q(
        regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(n1917), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(n1914), .E(n1955), .C(i_clk), .RN(n1941), .Q(
        regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(n1911), .E(n1955), .C(i_clk), .RN(n1937), .Q(
        regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(n1908), .E(n1955), .C(i_clk), .RN(n1943), .Q(
        regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(n1905), .E(n1955), .C(i_clk), .RN(n1944), .Q(
        regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(n1902), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(n1899), .E(n1955), .C(i_clk), .RN(n1941), .Q(
        regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(n1896), .E(n1955), .C(i_clk), .RN(n1943), .Q(
        regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(n1893), .E(n1955), .C(i_clk), .RN(n1943), .Q(
        regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(n1890), .E(n1955), .C(i_clk), .RN(n1942), .Q(
        regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(n1887), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(n1884), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(n1880), .E(n1955), .C(i_clk), .RN(n1950), .Q(
        regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(n1876), .E(n1955), .C(i_clk), .RN(n1930), .Q(
        regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(n1872), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(n1868), .E(n1955), .C(i_clk), .RN(n1931), .Q(
        regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(n1864), .E(n1955), .C(i_clk), .RN(n1947), .Q(
        regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(n1860), .E(n1955), .C(i_clk), .RN(n1946), .Q(
        regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(n1856), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(n1852), .E(n1955), .C(i_clk), .RN(n1949), .Q(
        regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(n1848), .E(n1955), .C(i_clk), .RN(n1948), .Q(
        regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(n1845), .E(n1955), .C(i_clk), .RN(n1947), .Q(
        regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(n1842), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(i_data_Rd[4]), .E(n1955), .C(i_clk), .RN(n1931), 
        .Q(regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(n1836), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(n1833), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(n1830), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(n1827), .E(n1955), .C(i_clk), .RN(i_rst_n), .Q(
        regs[608]) );
  DFEC1 regs_reg_17__31_ ( .D(n1929), .E(n1957), .C(i_clk), .RN(n1944), .Q(
        regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(i_data_Rd[30]), .E(n1957), .C(i_clk), .RN(n1950), 
        .Q(regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(n1923), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(n1920), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(n1917), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(n1914), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(n1911), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(n1908), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(n1905), .E(n1957), .C(i_clk), .RN(n1946), .Q(
        regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(n1902), .E(n1957), .C(i_clk), .RN(n1940), .Q(
        regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(n1899), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(n1896), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(n1893), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(n1890), .E(n1957), .C(i_clk), .RN(n1943), .Q(
        regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(n1887), .E(n1957), .C(i_clk), .RN(n1944), .Q(
        regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(n1884), .E(n1957), .C(i_clk), .RN(n1945), .Q(
        regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(n1880), .E(n1957), .C(i_clk), .RN(n1950), .Q(
        regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(n1876), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(n1872), .E(n1957), .C(i_clk), .RN(n1936), .Q(
        regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(n1868), .E(n1957), .C(i_clk), .RN(n1946), .Q(
        regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(n1864), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(n1860), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(n1856), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(n1852), .E(n1957), .C(i_clk), .RN(n1943), .Q(
        regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(n1848), .E(n1957), .C(i_clk), .RN(n1947), .Q(
        regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(n1845), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(n1842), .E(n1957), .C(i_clk), .RN(n1944), .Q(
        regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(i_data_Rd[4]), .E(n1957), .C(i_clk), .RN(n1930), 
        .Q(regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(n1836), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(n1833), .E(n1957), .C(i_clk), .RN(n1946), .Q(
        regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(n1830), .E(n1957), .C(i_clk), .RN(i_rst_n), .Q(
        regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(n1827), .E(n1957), .C(i_clk), .RN(n1940), .Q(
        regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(n1929), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(i_data_Rd[30]), .E(n1958), .C(i_clk), .RN(n1949), 
        .Q(regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(n1923), .E(n1958), .C(i_clk), .RN(n1948), .Q(
        regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(n1920), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(n1917), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(n1914), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(n1911), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(n1908), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(n1905), .E(n1958), .C(i_clk), .RN(n1949), .Q(
        regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(n1902), .E(n1958), .C(i_clk), .RN(n1948), .Q(
        regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(n1899), .E(n1958), .C(i_clk), .RN(n1931), .Q(
        regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(n1896), .E(n1958), .C(i_clk), .RN(n1932), .Q(
        regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(n1893), .E(n1958), .C(i_clk), .RN(n1933), .Q(
        regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(n1890), .E(n1958), .C(i_clk), .RN(n1934), .Q(
        regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(n1887), .E(n1958), .C(i_clk), .RN(n1935), .Q(
        regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(n1884), .E(n1958), .C(i_clk), .RN(n1947), .Q(
        regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(n1880), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(n1876), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(n1872), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(n1868), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(n1864), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(n1860), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(n1856), .E(n1958), .C(i_clk), .RN(n1943), .Q(
        regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(n1852), .E(n1958), .C(i_clk), .RN(n1941), .Q(
        regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(n1848), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(n1845), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(n1842), .E(n1958), .C(i_clk), .RN(n1950), .Q(
        regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(i_data_Rd[4]), .E(n1958), .C(i_clk), .RN(n1946), 
        .Q(regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(n1836), .E(n1958), .C(i_clk), .RN(n1950), .Q(
        regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(n1833), .E(n1958), .C(i_clk), .RN(n1938), .Q(
        regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(n1830), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(n1827), .E(n1958), .C(i_clk), .RN(i_rst_n), .Q(
        regs[512]) );
  DFEC1 regs_reg_15__31_ ( .D(n1928), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(n1925), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(n1922), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(n1919), .E(n1968), .C(i_clk), .RN(n1936), .Q(
        regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(n1916), .E(n1968), .C(i_clk), .RN(n1950), .Q(
        regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(n1913), .E(n1968), .C(i_clk), .RN(n1938), .Q(
        regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(n1910), .E(n1968), .C(i_clk), .RN(n1939), .Q(
        regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(n1907), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(n1904), .E(n1968), .C(i_clk), .RN(n1948), .Q(
        regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(n1901), .E(n1968), .C(i_clk), .RN(n1937), .Q(
        regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(n1898), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(n1895), .E(n1968), .C(i_clk), .RN(n1942), .Q(
        regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(n1892), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(n1889), .E(n1968), .C(i_clk), .RN(n1949), .Q(
        regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(n1886), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(n1883), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(n1879), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(n1875), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(n1871), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(n1867), .E(n1968), .C(i_clk), .RN(n1931), .Q(
        regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(n1863), .E(n1968), .C(i_clk), .RN(n1932), .Q(
        regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(n1859), .E(n1968), .C(i_clk), .RN(n1933), .Q(
        regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(n1855), .E(n1968), .C(i_clk), .RN(n1934), .Q(
        regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(n1851), .E(n1968), .C(i_clk), .RN(n1935), .Q(
        regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(n1847), .E(n1968), .C(i_clk), .RN(n1936), .Q(
        regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(n1844), .E(n1968), .C(i_clk), .RN(n1937), .Q(
        regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(n1841), .E(n1968), .C(i_clk), .RN(n1938), .Q(
        regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(n1838), .E(n1968), .C(i_clk), .RN(n1939), .Q(
        regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(n1835), .E(n1968), .C(i_clk), .RN(n1930), .Q(
        regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(n1832), .E(n1968), .C(i_clk), .RN(i_rst_n), .Q(
        regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(n1829), .E(n1968), .C(i_clk), .RN(n1937), .Q(
        regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(n1826), .E(n1968), .C(i_clk), .RN(n1939), .Q(
        regs[480]) );
  DFEC1 regs_reg_13__31_ ( .D(n1928), .E(n1970), .C(i_clk), .RN(n1944), .Q(
        regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(n1925), .E(n1970), .C(i_clk), .RN(n1939), .Q(
        regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(n1922), .E(n1970), .C(i_clk), .RN(n1949), .Q(
        regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(n1919), .E(n1970), .C(i_clk), .RN(n1948), .Q(
        regs[444]) );
  DFEC1 regs_reg_13__27_ ( .D(n1916), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(n1913), .E(n1970), .C(i_clk), .RN(n1945), .Q(
        regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(n1910), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(n1907), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(n1904), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(n1901), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(n1898), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(n1895), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(n1892), .E(n1970), .C(i_clk), .RN(n1938), .Q(
        regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(n1889), .E(n1970), .C(i_clk), .RN(n1944), .Q(
        regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(n1886), .E(n1970), .C(i_clk), .RN(n1940), .Q(
        regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(n1883), .E(n1970), .C(i_clk), .RN(n1945), .Q(
        regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(n1879), .E(n1970), .C(i_clk), .RN(n1945), .Q(
        regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(n1875), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(n1871), .E(n1970), .C(i_clk), .RN(n1935), .Q(
        regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(n1867), .E(n1970), .C(i_clk), .RN(n1941), .Q(
        regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(n1863), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(n1859), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(n1855), .E(n1970), .C(i_clk), .RN(n1940), .Q(
        regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(n1851), .E(n1970), .C(i_clk), .RN(n1946), .Q(
        regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(n1847), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(n1844), .E(n1970), .C(i_clk), .RN(n1941), .Q(
        regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(n1841), .E(n1970), .C(i_clk), .RN(n1937), .Q(
        regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(n1838), .E(n1970), .C(i_clk), .RN(n1940), .Q(
        regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(n1835), .E(n1970), .C(i_clk), .RN(n1937), .Q(
        regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(n1832), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(n1829), .E(n1970), .C(i_clk), .RN(n1948), .Q(
        regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(n1826), .E(n1970), .C(i_clk), .RN(i_rst_n), .Q(
        regs[416]) );
  DFEC1 regs_reg_12__31_ ( .D(n1928), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(n1925), .E(n1971), .C(i_clk), .RN(n1941), .Q(
        regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(n1922), .E(n1971), .C(i_clk), .RN(n1946), .Q(
        regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(n1919), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(n1916), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(n1913), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(n1910), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(n1907), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(n1904), .E(n1971), .C(i_clk), .RN(n1948), .Q(
        regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(n1901), .E(n1971), .C(i_clk), .RN(n1935), .Q(
        regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(n1898), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(n1895), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(n1892), .E(n1971), .C(i_clk), .RN(n1943), .Q(
        regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(n1889), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(n1886), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(n1883), .E(n1971), .C(i_clk), .RN(n1937), .Q(
        regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(n1879), .E(n1971), .C(i_clk), .RN(n1938), .Q(
        regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(n1875), .E(n1971), .C(i_clk), .RN(n1931), .Q(
        regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(n1871), .E(n1971), .C(i_clk), .RN(n1932), .Q(
        regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(n1867), .E(n1971), .C(i_clk), .RN(n1933), .Q(
        regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(n1863), .E(n1971), .C(i_clk), .RN(n1934), .Q(
        regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(n1859), .E(n1971), .C(i_clk), .RN(n1935), .Q(
        regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(n1855), .E(n1971), .C(i_clk), .RN(n1945), .Q(
        regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(n1851), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(n1847), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(n1844), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(n1841), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(n1838), .E(n1971), .C(i_clk), .RN(n1947), .Q(
        regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(n1835), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(n1832), .E(n1971), .C(i_clk), .RN(n1945), .Q(
        regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(n1829), .E(n1971), .C(i_clk), .RN(n1937), .Q(
        regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(n1826), .E(n1971), .C(i_clk), .RN(i_rst_n), .Q(
        regs[384]) );
  DFEC1 regs_reg_11__31_ ( .D(n1928), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(n1925), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(n1922), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(n1919), .E(n1972), .C(i_clk), .RN(n1941), .Q(
        regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(n1916), .E(n1972), .C(i_clk), .RN(n1949), .Q(
        regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(n1913), .E(n1972), .C(i_clk), .RN(n1934), .Q(
        regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(n1910), .E(n1972), .C(i_clk), .RN(n1943), .Q(
        regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(n1907), .E(n1972), .C(i_clk), .RN(n1944), .Q(
        regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(n1904), .E(n1972), .C(i_clk), .RN(n1936), .Q(
        regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(n1901), .E(n1972), .C(i_clk), .RN(n1939), .Q(
        regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(n1898), .E(n1972), .C(i_clk), .RN(n1948), .Q(
        regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(n1895), .E(n1972), .C(i_clk), .RN(n1938), .Q(
        regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(n1892), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(n1889), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(n1886), .E(n1972), .C(i_clk), .RN(n1935), .Q(
        regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(n1883), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(n1879), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(n1875), .E(n1972), .C(i_clk), .RN(n1946), .Q(
        regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(n1871), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(n1867), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(n1863), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(n1859), .E(n1972), .C(i_clk), .RN(n1939), .Q(
        regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(n1855), .E(n1972), .C(i_clk), .RN(n1930), .Q(
        regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(n1851), .E(n1972), .C(i_clk), .RN(n1946), .Q(
        regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(n1847), .E(n1972), .C(i_clk), .RN(n1940), .Q(
        regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(n1844), .E(n1972), .C(i_clk), .RN(n1939), .Q(
        regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(n1841), .E(n1972), .C(i_clk), .RN(n1936), .Q(
        regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(n1838), .E(n1972), .C(i_clk), .RN(n1941), .Q(
        regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(n1835), .E(n1972), .C(i_clk), .RN(n1949), .Q(
        regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(n1832), .E(n1972), .C(i_clk), .RN(n1941), .Q(
        regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(n1829), .E(n1972), .C(i_clk), .RN(i_rst_n), .Q(
        regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(n1826), .E(n1972), .C(i_clk), .RN(n1940), .Q(
        regs[352]) );
  DFEC1 regs_reg_9__31_ ( .D(n1928), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(n1925), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(n1922), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(n1919), .E(n1974), .C(i_clk), .RN(n1949), .Q(
        regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(n1916), .E(n1974), .C(i_clk), .RN(n1948), .Q(
        regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(n1913), .E(n1974), .C(i_clk), .RN(n1947), .Q(
        regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(n1910), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(n1907), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(n1904), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(n1901), .E(n1974), .C(i_clk), .RN(n1950), .Q(
        regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(n1898), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(n1895), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(n1892), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(n1889), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(n1886), .E(n1974), .C(i_clk), .RN(n1937), .Q(
        regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(n1883), .E(n1974), .C(i_clk), .RN(n1947), .Q(
        regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(n1879), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(n1875), .E(n1974), .C(i_clk), .RN(n1947), .Q(
        regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(n1871), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(n1867), .E(n1974), .C(i_clk), .RN(n1950), .Q(
        regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(n1863), .E(n1974), .C(i_clk), .RN(n1936), .Q(
        regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(n1859), .E(n1974), .C(i_clk), .RN(n1930), .Q(
        regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(n1855), .E(n1974), .C(i_clk), .RN(n1939), .Q(
        regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(n1851), .E(n1974), .C(i_clk), .RN(n1930), .Q(
        regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(n1847), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(n1844), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(n1841), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(n1838), .E(n1974), .C(i_clk), .RN(n1934), .Q(
        regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(n1835), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(n1832), .E(n1974), .C(i_clk), .RN(i_rst_n), .Q(
        regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(n1829), .E(n1974), .C(i_clk), .RN(n1943), .Q(
        regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(n1826), .E(n1974), .C(i_clk), .RN(n1936), .Q(
        regs[288]) );
  DFEC1 regs_reg_8__31_ ( .D(n1928), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(n1925), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(n1922), .E(n1975), .C(i_clk), .RN(n1946), .Q(
        regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(n1919), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(n1916), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(n1913), .E(n1975), .C(i_clk), .RN(n1949), .Q(
        regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(n1910), .E(n1975), .C(i_clk), .RN(n1948), .Q(
        regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(n1907), .E(n1975), .C(i_clk), .RN(n1947), .Q(
        regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(n1904), .E(n1975), .C(i_clk), .RN(n1930), .Q(
        regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(n1901), .E(n1975), .C(i_clk), .RN(n1950), .Q(
        regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(n1898), .E(n1975), .C(i_clk), .RN(n1950), .Q(
        regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(n1895), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(n1892), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(n1889), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(n1886), .E(n1975), .C(i_clk), .RN(n1949), .Q(
        regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(n1883), .E(n1975), .C(i_clk), .RN(n1948), .Q(
        regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(n1879), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(n1875), .E(n1975), .C(i_clk), .RN(n1946), .Q(
        regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(n1871), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(n1867), .E(n1975), .C(i_clk), .RN(n1938), .Q(
        regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(n1863), .E(n1975), .C(i_clk), .RN(n1947), .Q(
        regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(n1859), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(n1855), .E(n1975), .C(i_clk), .RN(n1934), .Q(
        regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(n1851), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(n1847), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(n1844), .E(n1975), .C(i_clk), .RN(i_rst_n), .Q(
        regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(n1841), .E(n1975), .C(i_clk), .RN(n1935), .Q(
        regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(n1838), .E(n1975), .C(i_clk), .RN(n1950), .Q(
        regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(n1835), .E(n1975), .C(i_clk), .RN(n1941), .Q(
        regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(n1832), .E(n1975), .C(i_clk), .RN(n1946), .Q(
        regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(n1829), .E(n1975), .C(i_clk), .RN(n1940), .Q(
        regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(n1826), .E(n1975), .C(i_clk), .RN(n1938), .Q(
        regs[256]) );
  DFEC1 regs_reg_7__31_ ( .D(n1927), .E(n1976), .C(i_clk), .RN(n1933), .Q(
        regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(n1924), .E(n1976), .C(i_clk), .RN(n1930), .Q(
        regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(n1921), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(n1918), .E(n1976), .C(i_clk), .RN(n1930), .Q(
        regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(n1915), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(n1912), .E(n1976), .C(i_clk), .RN(n1940), .Q(
        regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(n1909), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(n1906), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(n1903), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(n1900), .E(n1976), .C(i_clk), .RN(n1937), .Q(
        regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(n1897), .E(n1976), .C(i_clk), .RN(n1933), .Q(
        regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(n1894), .E(n1976), .C(i_clk), .RN(n1947), .Q(
        regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(n1891), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(n1888), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(n1885), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(n1882), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(n1878), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(n1874), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(n1870), .E(n1976), .C(i_clk), .RN(n1930), .Q(
        regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(n1866), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(n1862), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(n1858), .E(n1976), .C(i_clk), .RN(n1934), .Q(
        regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(n1854), .E(n1976), .C(i_clk), .RN(n1935), .Q(
        regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(n1850), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(n1846), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(n1843), .E(n1976), .C(i_clk), .RN(n1946), .Q(
        regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(n1840), .E(n1976), .C(i_clk), .RN(n1936), .Q(
        regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(n1837), .E(n1976), .C(i_clk), .RN(n1930), .Q(
        regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(n1834), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(n1831), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(n1828), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(n1825), .E(n1976), .C(i_clk), .RN(i_rst_n), .Q(
        regs[224]) );
  DFEC1 regs_reg_5__31_ ( .D(n1927), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(n1924), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(n1921), .E(n1978), .C(i_clk), .RN(n1936), .Q(
        regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(n1918), .E(n1978), .C(i_clk), .RN(n1943), .Q(
        regs[188]) );
  DFEC1 regs_reg_5__27_ ( .D(n1915), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(n1912), .E(n1978), .C(i_clk), .RN(n1946), .Q(
        regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(n1909), .E(n1978), .C(i_clk), .RN(n1946), .Q(
        regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(n1906), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(n1903), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(n1900), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(n1897), .E(n1978), .C(i_clk), .RN(n1933), .Q(
        regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(n1894), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(n1891), .E(n1978), .C(i_clk), .RN(n1950), .Q(
        regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(n1888), .E(n1978), .C(i_clk), .RN(n1940), .Q(
        regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(n1885), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(n1882), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(n1878), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(n1874), .E(n1978), .C(i_clk), .RN(n1945), .Q(
        regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(n1870), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(n1866), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(n1862), .E(n1978), .C(i_clk), .RN(n1930), .Q(
        regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(n1858), .E(n1978), .C(i_clk), .RN(n1948), .Q(
        regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(n1854), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(n1850), .E(n1978), .C(i_clk), .RN(n1934), .Q(
        regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(n1846), .E(n1978), .C(i_clk), .RN(n1932), .Q(
        regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(n1843), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(n1840), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(n1837), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(n1834), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(n1831), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(n1828), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(n1825), .E(n1978), .C(i_clk), .RN(i_rst_n), .Q(
        regs[160]) );
  DFEC1 regs_reg_4__31_ ( .D(n1927), .E(n1979), .C(i_clk), .RN(n1942), .Q(
        regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(n1924), .E(n1979), .C(i_clk), .RN(n1945), .Q(
        regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(n1921), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(n1918), .E(n1979), .C(i_clk), .RN(n1931), .Q(
        regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(n1915), .E(n1979), .C(i_clk), .RN(n1938), .Q(
        regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(n1912), .E(n1979), .C(i_clk), .RN(n1949), .Q(
        regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(n1909), .E(n1979), .C(i_clk), .RN(n1948), .Q(
        regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(n1906), .E(n1979), .C(i_clk), .RN(n1947), .Q(
        regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(n1903), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(n1900), .E(n1979), .C(i_clk), .RN(n1949), .Q(
        regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(n1897), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(n1894), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(n1891), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(n1888), .E(n1979), .C(i_clk), .RN(n1935), .Q(
        regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(n1885), .E(n1979), .C(i_clk), .RN(n1938), .Q(
        regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(n1882), .E(n1979), .C(i_clk), .RN(n1931), .Q(
        regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(n1878), .E(n1979), .C(i_clk), .RN(n1943), .Q(
        regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(n1874), .E(n1979), .C(i_clk), .RN(n1942), .Q(
        regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(n1870), .E(n1979), .C(i_clk), .RN(n1941), .Q(
        regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(n1866), .E(n1979), .C(i_clk), .RN(n1930), .Q(
        regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(n1862), .E(n1979), .C(i_clk), .RN(n1943), .Q(
        regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(n1858), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(n1854), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(n1850), .E(n1979), .C(i_clk), .RN(n1948), .Q(
        regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(n1846), .E(n1979), .C(i_clk), .RN(n1946), .Q(
        regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(n1843), .E(n1979), .C(i_clk), .RN(n1943), .Q(
        regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(n1840), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(n1837), .E(n1979), .C(i_clk), .RN(n1947), .Q(
        regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(n1834), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(n1831), .E(n1979), .C(i_clk), .RN(n1948), .Q(
        regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(n1828), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(n1825), .E(n1979), .C(i_clk), .RN(i_rst_n), .Q(
        regs[128]) );
  DFEC1 regs_reg_3__31_ ( .D(n1927), .E(n1980), .C(i_clk), .RN(n1942), .Q(
        regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(n1924), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(n1921), .E(n1980), .C(i_clk), .RN(n1945), .Q(
        regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(n1918), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(n1915), .E(n1980), .C(i_clk), .RN(n1930), .Q(
        regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(n1912), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(n1909), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(n1906), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(n1903), .E(n1980), .C(i_clk), .RN(n1946), .Q(
        regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(n1900), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(n1897), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(n1894), .E(n1980), .C(i_clk), .RN(n1948), .Q(
        regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(n1891), .E(n1980), .C(i_clk), .RN(n1946), .Q(
        regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(n1888), .E(n1980), .C(i_clk), .RN(n1949), .Q(
        regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(n1885), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(n1882), .E(n1980), .C(i_clk), .RN(n1949), .Q(
        regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(n1878), .E(n1980), .C(i_clk), .RN(n1932), .Q(
        regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(n1874), .E(n1980), .C(i_clk), .RN(n1930), .Q(
        regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(n1870), .E(n1980), .C(i_clk), .RN(n1950), .Q(
        regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(n1866), .E(n1980), .C(i_clk), .RN(n1930), .Q(
        regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(n1862), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(n1858), .E(n1980), .C(i_clk), .RN(n1949), .Q(
        regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(n1854), .E(n1980), .C(i_clk), .RN(n1934), .Q(
        regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(n1850), .E(n1980), .C(i_clk), .RN(n1944), .Q(
        regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(n1846), .E(n1980), .C(i_clk), .RN(n1942), .Q(
        regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(n1843), .E(n1980), .C(i_clk), .RN(n1950), .Q(
        regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(n1840), .E(n1980), .C(i_clk), .RN(n1950), .Q(
        regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(n1837), .E(n1980), .C(i_clk), .RN(n1944), .Q(
        regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(n1834), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(n1831), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(n1828), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(n1825), .E(n1980), .C(i_clk), .RN(i_rst_n), .Q(
        regs[96]) );
  DFEC1 regs_reg_1__31_ ( .D(n1927), .E(n1982), .C(i_clk), .RN(i_rst_n), .Q(
        regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(n1924), .E(n1982), .C(i_clk), .RN(n1937), .Q(
        regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(n1921), .E(n1982), .C(i_clk), .RN(i_rst_n), .Q(
        regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(n1918), .E(n1982), .C(i_clk), .RN(n1949), .Q(
        regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(n1915), .E(n1982), .C(i_clk), .RN(i_rst_n), .Q(
        regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(n1912), .E(n1982), .C(i_clk), .RN(i_rst_n), .Q(
        regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(n1909), .E(n1982), .C(i_clk), .RN(n1945), .Q(
        regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(n1906), .E(n1982), .C(i_clk), .RN(n1930), .Q(
        regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(n1903), .E(n1982), .C(i_clk), .RN(i_rst_n), .Q(
        regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(n1900), .E(n1982), .C(i_clk), .RN(i_rst_n), .Q(
        regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(n1897), .E(n1982), .C(i_clk), .RN(i_rst_n), .Q(
        regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(n1894), .E(n1982), .C(i_clk), .RN(n1931), .Q(
        regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(n1891), .E(n1982), .C(i_clk), .RN(n1943), .Q(
        regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(n1888), .E(n1982), .C(i_clk), .RN(n1943), .Q(
        regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(n1885), .E(n1982), .C(i_clk), .RN(n1943), .Q(
        regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(n1882), .E(n1982), .C(i_clk), .RN(n1943), .Q(
        regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(n1878), .E(n1982), .C(i_clk), .RN(n1943), .Q(
        regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(n1874), .E(n1982), .C(i_clk), .RN(n1943), .Q(
        regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(n1870), .E(n1982), .C(i_clk), .RN(n1943), .Q(
        regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(n1866), .E(n1982), .C(i_clk), .RN(n1943), .Q(
        regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(n1862), .E(n1982), .C(i_clk), .RN(n1943), .Q(
        regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(n1858), .E(n1982), .C(i_clk), .RN(n1944), .Q(
        regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(n1854), .E(n1982), .C(i_clk), .RN(n1944), .Q(
        regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(n1850), .E(n1982), .C(i_clk), .RN(n1944), .Q(
        regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(n1846), .E(n1982), .C(i_clk), .RN(n1944), .Q(
        regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(n1843), .E(n1982), .C(i_clk), .RN(n1944), .Q(
        regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(n1840), .E(n1982), .C(i_clk), .RN(n1944), .Q(
        regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(n1837), .E(n1982), .C(i_clk), .RN(n1944), .Q(
        regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(n1834), .E(n1982), .C(i_clk), .RN(n1944), .Q(
        regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(n1831), .E(n1982), .C(i_clk), .RN(n1944), .Q(
        regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(n1828), .E(n1982), .C(i_clk), .RN(n1945), .Q(
        regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(n1825), .E(n1982), .C(i_clk), .RN(n1945), .Q(
        regs[32]) );
  DFEC1 regs_reg_0__31_ ( .D(n1927), .E(n1983), .C(i_clk), .RN(n1945), .Q(
        regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(n1924), .E(n1983), .C(i_clk), .RN(n1945), .Q(
        regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(n1921), .E(n1983), .C(i_clk), .RN(n1945), .Q(
        regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(n1918), .E(n1983), .C(i_clk), .RN(n1945), .Q(
        regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(n1915), .E(n1983), .C(i_clk), .RN(n1945), .Q(
        regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(n1912), .E(n1983), .C(i_clk), .RN(n1945), .Q(
        regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(n1909), .E(n1983), .C(i_clk), .RN(n1945), .Q(
        regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(n1906), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(n1903), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(n1900), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(n1897), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(n1894), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(n1891), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(n1888), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(n1885), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(n1882), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(n1878), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(n1874), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(n1870), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(n1866), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(n1862), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(n1858), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(n1854), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(n1850), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(n1846), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(n1843), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(n1840), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(n1837), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(n1834), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(n1831), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(n1828), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(n1825), .E(n1983), .C(i_clk), .RN(i_rst_n), .Q(
        regs[0]) );
  CLKBU12 U2 ( .A(i_addr_Rs[0]), .Q(n1818) );
  BUF6 U3 ( .A(n1824), .Q(n1819) );
  IMUX40 U4 ( .A(n1577), .B(n1578), .C(n1579), .D(n1580), .S0(n1774), .S1(
        n1777), .Q(n1576) );
  IMUX40 U5 ( .A(n1587), .B(n1588), .C(n1589), .D(n1590), .S0(n1774), .S1(
        n1777), .Q(n1586) );
  IMUX40 U6 ( .A(n1582), .B(n1583), .C(n1584), .D(n1585), .S0(n1774), .S1(
        n1777), .Q(n1581) );
  BUF4 U7 ( .A(i_addr_Rs[0]), .Q(n1823) );
  BUF6 U8 ( .A(i_addr_Rs[0]), .Q(n1817) );
  BUF6 U9 ( .A(i_addr_Rs[3]), .Q(n1774) );
  BUF8 U10 ( .A(n1824), .Q(n1820) );
  BUF6 U11 ( .A(i_addr_Rs[0]), .Q(n1) );
  BUF6 U12 ( .A(i_addr_Rs[0]), .Q(n2) );
  CLKBU4 U13 ( .A(n1823), .Q(n1816) );
  BUF2 U14 ( .A(i_addr_Rs[4]), .Q(n1772) );
  BUF2 U15 ( .A(i_addr_Rt[4]), .Q(n1392) );
  BUF2 U16 ( .A(n1945), .Q(n1942) );
  BUF2 U17 ( .A(n1930), .Q(n1941) );
  BUF2 U18 ( .A(n1950), .Q(n1940) );
  BUF2 U19 ( .A(n1947), .Q(n1939) );
  BUF2 U20 ( .A(n1947), .Q(n1938) );
  BUF2 U21 ( .A(n1947), .Q(n1937) );
  BUF2 U22 ( .A(n1948), .Q(n1936) );
  BUF2 U23 ( .A(n1948), .Q(n1935) );
  BUF2 U24 ( .A(n1948), .Q(n1934) );
  BUF2 U25 ( .A(n1949), .Q(n1933) );
  BUF2 U26 ( .A(n1949), .Q(n1932) );
  BUF2 U27 ( .A(n1949), .Q(n1931) );
  BUF2 U28 ( .A(n1946), .Q(n1945) );
  BUF2 U29 ( .A(n1946), .Q(n1944) );
  BUF2 U30 ( .A(n1946), .Q(n1943) );
  BUF2 U31 ( .A(n1950), .Q(n1947) );
  BUF2 U32 ( .A(n1940), .Q(n1948) );
  BUF2 U33 ( .A(n1941), .Q(n1949) );
  BUF2 U34 ( .A(n1950), .Q(n1946) );
  BUF2 U35 ( .A(n1823), .Q(n1815) );
  BUF2 U36 ( .A(i_addr_Rs[0]), .Q(n1821) );
  BUF2 U37 ( .A(n1787), .Q(n1789) );
  BUF2 U38 ( .A(n1787), .Q(n1790) );
  BUF2 U39 ( .A(n1786), .Q(n1791) );
  BUF2 U40 ( .A(n1786), .Q(n1792) );
  BUF2 U41 ( .A(n1786), .Q(n1793) );
  BUF2 U42 ( .A(n1813), .Q(n1794) );
  BUF2 U43 ( .A(n1813), .Q(n1795) );
  BUF2 U44 ( .A(n1811), .Q(n1796) );
  BUF2 U45 ( .A(n1811), .Q(n1797) );
  BUF2 U46 ( .A(n1781), .Q(n1798) );
  BUF2 U47 ( .A(n1784), .Q(n1799) );
  BUF2 U48 ( .A(n1784), .Q(n1800) );
  BUF2 U49 ( .A(n1784), .Q(n1801) );
  BUF2 U50 ( .A(n1783), .Q(n1802) );
  BUF2 U51 ( .A(n1783), .Q(n1803) );
  BUF2 U52 ( .A(n1783), .Q(n1804) );
  BUF2 U53 ( .A(n1782), .Q(n1805) );
  BUF2 U54 ( .A(n1782), .Q(n1806) );
  BUF2 U55 ( .A(n1782), .Q(n1807) );
  BUF2 U56 ( .A(n1781), .Q(n1808) );
  BUF2 U57 ( .A(n1781), .Q(n1809) );
  BUF2 U58 ( .A(n1781), .Q(n1810) );
  BUF2 U59 ( .A(n1787), .Q(n1788) );
  BUF2 U60 ( .A(i_addr_Rt[0]), .Q(n1430) );
  BUF2 U61 ( .A(i_addr_Rt[0]), .Q(n1431) );
  BUF2 U62 ( .A(i_addr_Rt[0]), .Q(n1432) );
  BUF2 U63 ( .A(i_addr_Rt[0]), .Q(n1433) );
  BUF2 U64 ( .A(i_addr_Rt[0]), .Q(n1434) );
  BUF2 U65 ( .A(i_addr_Rt[0]), .Q(n1435) );
  BUF2 U66 ( .A(i_addr_Rt[0]), .Q(n1436) );
  BUF2 U67 ( .A(i_addr_Rt[0]), .Q(n1437) );
  BUF2 U68 ( .A(i_addr_Rt[0]), .Q(n1438) );
  BUF2 U69 ( .A(n1449), .Q(n1439) );
  BUF2 U70 ( .A(n1450), .Q(n1440) );
  BUF2 U71 ( .A(n1449), .Q(n1441) );
  BUF2 U72 ( .A(i_addr_Rt[0]), .Q(n1442) );
  BUF2 U73 ( .A(n1449), .Q(n1443) );
  BUF2 U74 ( .A(n1449), .Q(n1444) );
  BUF2 U75 ( .A(n1449), .Q(n1445) );
  BUF2 U76 ( .A(n1450), .Q(n1446) );
  BUF2 U77 ( .A(n1450), .Q(n1447) );
  BUF2 U78 ( .A(n1450), .Q(n1448) );
  BUF2 U79 ( .A(n1429), .Q(n1409) );
  BUF2 U80 ( .A(n1408), .Q(n1410) );
  BUF2 U81 ( .A(n1408), .Q(n1411) );
  BUF2 U82 ( .A(n1407), .Q(n1412) );
  BUF2 U83 ( .A(n1407), .Q(n1413) );
  BUF2 U84 ( .A(n1407), .Q(n1414) );
  BUF2 U85 ( .A(n1407), .Q(n1415) );
  BUF2 U86 ( .A(n1406), .Q(n1416) );
  BUF2 U87 ( .A(n1406), .Q(n1417) );
  BUF2 U88 ( .A(n1406), .Q(n1418) );
  BUF2 U89 ( .A(n1405), .Q(n1419) );
  BUF2 U90 ( .A(n1405), .Q(n1420) );
  BUF2 U91 ( .A(n1405), .Q(n1421) );
  BUF2 U92 ( .A(n1404), .Q(n1422) );
  BUF2 U93 ( .A(n1404), .Q(n1423) );
  BUF2 U94 ( .A(n1404), .Q(n1424) );
  BUF2 U95 ( .A(i_data_Rd[0]), .Q(n1825) );
  BUF2 U96 ( .A(i_data_Rd[1]), .Q(n1828) );
  BUF2 U97 ( .A(i_data_Rd[2]), .Q(n1831) );
  BUF2 U98 ( .A(i_data_Rd[3]), .Q(n1834) );
  BUF2 U99 ( .A(i_data_Rd[4]), .Q(n1837) );
  BUF2 U100 ( .A(i_data_Rd[5]), .Q(n1840) );
  BUF2 U101 ( .A(i_data_Rd[6]), .Q(n1843) );
  BUF2 U102 ( .A(i_data_Rd[7]), .Q(n1846) );
  BUF2 U103 ( .A(i_data_Rd[8]), .Q(n1850) );
  BUF2 U104 ( .A(i_data_Rd[9]), .Q(n1854) );
  BUF2 U105 ( .A(i_data_Rd[10]), .Q(n1858) );
  BUF2 U106 ( .A(i_data_Rd[11]), .Q(n1862) );
  BUF2 U107 ( .A(i_data_Rd[12]), .Q(n1866) );
  BUF2 U108 ( .A(i_data_Rd[13]), .Q(n1870) );
  BUF2 U109 ( .A(i_data_Rd[14]), .Q(n1874) );
  BUF2 U110 ( .A(i_data_Rd[15]), .Q(n1878) );
  BUF2 U111 ( .A(i_data_Rd[16]), .Q(n1882) );
  BUF2 U112 ( .A(i_data_Rd[17]), .Q(n1885) );
  BUF2 U113 ( .A(i_data_Rd[18]), .Q(n1888) );
  BUF2 U114 ( .A(i_data_Rd[19]), .Q(n1891) );
  BUF2 U115 ( .A(i_data_Rd[20]), .Q(n1894) );
  BUF2 U116 ( .A(i_data_Rd[21]), .Q(n1897) );
  BUF2 U117 ( .A(i_data_Rd[22]), .Q(n1900) );
  BUF2 U118 ( .A(i_data_Rd[23]), .Q(n1903) );
  BUF2 U119 ( .A(i_data_Rd[24]), .Q(n1906) );
  BUF2 U120 ( .A(i_data_Rd[25]), .Q(n1909) );
  BUF2 U121 ( .A(i_data_Rd[26]), .Q(n1912) );
  BUF2 U122 ( .A(i_data_Rd[27]), .Q(n1915) );
  BUF2 U123 ( .A(i_data_Rd[28]), .Q(n1918) );
  BUF2 U124 ( .A(i_data_Rd[29]), .Q(n1921) );
  BUF2 U125 ( .A(i_data_Rd[30]), .Q(n1924) );
  BUF2 U126 ( .A(i_data_Rd[31]), .Q(n1927) );
  BUF2 U127 ( .A(i_data_Rd[0]), .Q(n1826) );
  BUF2 U128 ( .A(i_data_Rd[1]), .Q(n1829) );
  BUF2 U129 ( .A(i_data_Rd[2]), .Q(n1832) );
  BUF2 U130 ( .A(i_data_Rd[3]), .Q(n1835) );
  BUF2 U131 ( .A(i_data_Rd[4]), .Q(n1838) );
  BUF2 U132 ( .A(i_data_Rd[5]), .Q(n1841) );
  BUF2 U133 ( .A(i_data_Rd[6]), .Q(n1844) );
  BUF2 U134 ( .A(i_data_Rd[7]), .Q(n1847) );
  BUF2 U135 ( .A(i_data_Rd[8]), .Q(n1851) );
  BUF2 U136 ( .A(i_data_Rd[9]), .Q(n1855) );
  BUF2 U137 ( .A(i_data_Rd[10]), .Q(n1859) );
  BUF2 U138 ( .A(i_data_Rd[11]), .Q(n1863) );
  BUF2 U139 ( .A(i_data_Rd[12]), .Q(n1867) );
  BUF2 U140 ( .A(i_data_Rd[13]), .Q(n1871) );
  BUF2 U141 ( .A(i_data_Rd[14]), .Q(n1875) );
  BUF2 U142 ( .A(i_data_Rd[15]), .Q(n1879) );
  BUF2 U143 ( .A(i_data_Rd[16]), .Q(n1883) );
  BUF2 U144 ( .A(i_data_Rd[17]), .Q(n1886) );
  BUF2 U145 ( .A(i_data_Rd[18]), .Q(n1889) );
  BUF2 U146 ( .A(i_data_Rd[19]), .Q(n1892) );
  BUF2 U147 ( .A(i_data_Rd[20]), .Q(n1895) );
  BUF2 U148 ( .A(i_data_Rd[21]), .Q(n1898) );
  BUF2 U149 ( .A(i_data_Rd[22]), .Q(n1901) );
  BUF2 U150 ( .A(i_data_Rd[23]), .Q(n1904) );
  BUF2 U151 ( .A(i_data_Rd[24]), .Q(n1907) );
  BUF2 U152 ( .A(i_data_Rd[25]), .Q(n1910) );
  BUF2 U153 ( .A(i_data_Rd[26]), .Q(n1913) );
  BUF2 U154 ( .A(i_data_Rd[27]), .Q(n1916) );
  BUF2 U155 ( .A(i_data_Rd[28]), .Q(n1919) );
  BUF2 U156 ( .A(i_data_Rd[29]), .Q(n1922) );
  BUF2 U157 ( .A(i_data_Rd[30]), .Q(n1925) );
  BUF2 U158 ( .A(i_data_Rd[31]), .Q(n1928) );
  BUF2 U159 ( .A(i_data_Rd[0]), .Q(n1827) );
  BUF2 U160 ( .A(i_data_Rd[1]), .Q(n1830) );
  BUF2 U161 ( .A(i_data_Rd[2]), .Q(n1833) );
  BUF2 U162 ( .A(i_data_Rd[3]), .Q(n1836) );
  BUF2 U163 ( .A(i_data_Rd[5]), .Q(n1842) );
  BUF2 U164 ( .A(i_data_Rd[6]), .Q(n1845) );
  BUF2 U165 ( .A(i_data_Rd[7]), .Q(n1848) );
  BUF2 U166 ( .A(i_data_Rd[8]), .Q(n1852) );
  BUF2 U167 ( .A(i_data_Rd[9]), .Q(n1856) );
  BUF2 U168 ( .A(i_data_Rd[10]), .Q(n1860) );
  BUF2 U169 ( .A(i_data_Rd[11]), .Q(n1864) );
  BUF2 U170 ( .A(i_data_Rd[12]), .Q(n1868) );
  BUF2 U171 ( .A(i_data_Rd[13]), .Q(n1872) );
  BUF2 U172 ( .A(i_data_Rd[14]), .Q(n1876) );
  BUF2 U173 ( .A(i_data_Rd[15]), .Q(n1880) );
  BUF2 U174 ( .A(i_data_Rd[16]), .Q(n1884) );
  BUF2 U175 ( .A(i_data_Rd[17]), .Q(n1887) );
  BUF2 U176 ( .A(i_data_Rd[18]), .Q(n1890) );
  BUF2 U177 ( .A(i_data_Rd[19]), .Q(n1893) );
  BUF2 U178 ( .A(i_data_Rd[20]), .Q(n1896) );
  BUF2 U179 ( .A(i_data_Rd[21]), .Q(n1899) );
  BUF2 U180 ( .A(i_data_Rd[22]), .Q(n1902) );
  BUF2 U181 ( .A(i_data_Rd[23]), .Q(n1905) );
  BUF2 U182 ( .A(i_data_Rd[24]), .Q(n1908) );
  BUF2 U183 ( .A(i_data_Rd[25]), .Q(n1911) );
  BUF2 U184 ( .A(i_data_Rd[26]), .Q(n1914) );
  BUF2 U185 ( .A(i_data_Rd[27]), .Q(n1917) );
  BUF2 U186 ( .A(i_data_Rd[28]), .Q(n1920) );
  BUF2 U187 ( .A(i_data_Rd[29]), .Q(n1923) );
  BUF2 U188 ( .A(i_data_Rd[31]), .Q(n1929) );
  BUF2 U189 ( .A(i_data_Rd[4]), .Q(n1839) );
  BUF2 U190 ( .A(i_data_Rd[7]), .Q(n1849) );
  BUF2 U191 ( .A(i_data_Rd[8]), .Q(n1853) );
  BUF2 U192 ( .A(i_data_Rd[9]), .Q(n1857) );
  BUF2 U193 ( .A(i_data_Rd[10]), .Q(n1861) );
  BUF2 U194 ( .A(i_data_Rd[11]), .Q(n1865) );
  BUF2 U195 ( .A(i_data_Rd[12]), .Q(n1869) );
  BUF2 U196 ( .A(i_data_Rd[13]), .Q(n1873) );
  BUF2 U197 ( .A(i_data_Rd[14]), .Q(n1877) );
  BUF2 U198 ( .A(i_data_Rd[15]), .Q(n1881) );
  BUF2 U199 ( .A(i_data_Rd[30]), .Q(n1926) );
  BUF2 U200 ( .A(n1930), .Q(n1950) );
  BUF2 U201 ( .A(i_rst_n), .Q(n1930) );
  BUF2 U202 ( .A(i_addr_Rs[0]), .Q(n1824) );
  BUF2 U203 ( .A(n1814), .Q(n1787) );
  BUF2 U204 ( .A(n1814), .Q(n1786) );
  BUF2 U205 ( .A(n1814), .Q(n1785) );
  BUF2 U206 ( .A(n1813), .Q(n1784) );
  BUF2 U207 ( .A(n1812), .Q(n1783) );
  BUF2 U208 ( .A(n1812), .Q(n1782) );
  BUF2 U209 ( .A(n1812), .Q(n1781) );
  NOR21 U210 ( .A(n1967), .B(n1984), .Q(n1099) );
  NOR31 U211 ( .A(n1986), .B(n1987), .C(n1985), .Q(n1079) );
  INV3 U212 ( .A(n1063), .Q(n1983) );
  NAND31 U213 ( .A(n1064), .B(n1065), .C(i_con_RegWr), .Q(n1063) );
  INV3 U214 ( .A(n1080), .Q(n1975) );
  NAND31 U215 ( .A(i_con_RegWr), .B(n1064), .C(n1081), .Q(n1080) );
  INV3 U216 ( .A(n1082), .Q(n1974) );
  NAND31 U217 ( .A(n1067), .B(i_con_RegWr), .C(n1081), .Q(n1082) );
  INV3 U218 ( .A(n1083), .Q(n1973) );
  NAND31 U219 ( .A(n1069), .B(i_con_RegWr), .C(n1081), .Q(n1083) );
  INV3 U220 ( .A(n1084), .Q(n1972) );
  NAND31 U221 ( .A(n1071), .B(i_con_RegWr), .C(n1081), .Q(n1084) );
  INV3 U222 ( .A(n1085), .Q(n1971) );
  NAND31 U223 ( .A(n1073), .B(i_con_RegWr), .C(n1081), .Q(n1085) );
  INV3 U224 ( .A(n1086), .Q(n1970) );
  NAND31 U225 ( .A(n1075), .B(i_con_RegWr), .C(n1081), .Q(n1086) );
  INV3 U226 ( .A(n1087), .Q(n1969) );
  NAND31 U227 ( .A(n1077), .B(i_con_RegWr), .C(n1081), .Q(n1087) );
  INV3 U228 ( .A(n1088), .Q(n1968) );
  NAND31 U229 ( .A(n1079), .B(i_con_RegWr), .C(n1081), .Q(n1088) );
  INV3 U230 ( .A(n1089), .Q(n1958) );
  NAND31 U231 ( .A(i_con_RegWr), .B(n1064), .C(n1090), .Q(n1089) );
  INV3 U232 ( .A(n1091), .Q(n1957) );
  NAND31 U233 ( .A(n1067), .B(i_con_RegWr), .C(n1090), .Q(n1091) );
  INV3 U234 ( .A(n1092), .Q(n1956) );
  NAND31 U235 ( .A(n1069), .B(i_con_RegWr), .C(n1090), .Q(n1092) );
  INV3 U236 ( .A(n1093), .Q(n1955) );
  NAND31 U237 ( .A(n1071), .B(i_con_RegWr), .C(n1090), .Q(n1093) );
  INV3 U238 ( .A(n1094), .Q(n1954) );
  NAND31 U239 ( .A(n1073), .B(i_con_RegWr), .C(n1090), .Q(n1094) );
  INV3 U240 ( .A(n1095), .Q(n1953) );
  NAND31 U241 ( .A(n1075), .B(i_con_RegWr), .C(n1090), .Q(n1095) );
  INV3 U242 ( .A(n1096), .Q(n1952) );
  NAND31 U243 ( .A(n1077), .B(i_con_RegWr), .C(n1090), .Q(n1096) );
  INV3 U244 ( .A(n1097), .Q(n1951) );
  NAND31 U245 ( .A(n1079), .B(i_con_RegWr), .C(n1090), .Q(n1097) );
  INV3 U246 ( .A(n1098), .Q(n1966) );
  NAND31 U247 ( .A(i_con_RegWr), .B(n1064), .C(n1099), .Q(n1098) );
  INV3 U248 ( .A(n1100), .Q(n1965) );
  NAND31 U249 ( .A(n1067), .B(i_con_RegWr), .C(n1099), .Q(n1100) );
  INV3 U250 ( .A(n1101), .Q(n1964) );
  NAND31 U251 ( .A(n1069), .B(i_con_RegWr), .C(n1099), .Q(n1101) );
  INV3 U252 ( .A(n1102), .Q(n1963) );
  NAND31 U253 ( .A(n1071), .B(i_con_RegWr), .C(n1099), .Q(n1102) );
  INV3 U254 ( .A(n1103), .Q(n1962) );
  NAND31 U255 ( .A(n1073), .B(i_con_RegWr), .C(n1099), .Q(n1103) );
  INV3 U256 ( .A(n1104), .Q(n1961) );
  NAND31 U257 ( .A(n1075), .B(i_con_RegWr), .C(n1099), .Q(n1104) );
  INV3 U258 ( .A(n1105), .Q(n1960) );
  NAND31 U259 ( .A(n1077), .B(i_con_RegWr), .C(n1099), .Q(n1105) );
  INV3 U260 ( .A(n1106), .Q(n1959) );
  NAND31 U261 ( .A(n1079), .B(i_con_RegWr), .C(n1099), .Q(n1106) );
  INV3 U262 ( .A(n1066), .Q(n1982) );
  NAND31 U263 ( .A(i_con_RegWr), .B(n1065), .C(n1067), .Q(n1066) );
  INV3 U264 ( .A(n1068), .Q(n1981) );
  NAND31 U265 ( .A(i_con_RegWr), .B(n1065), .C(n1069), .Q(n1068) );
  INV3 U266 ( .A(n1070), .Q(n1980) );
  NAND31 U267 ( .A(i_con_RegWr), .B(n1065), .C(n1071), .Q(n1070) );
  INV3 U268 ( .A(n1072), .Q(n1979) );
  NAND31 U269 ( .A(i_con_RegWr), .B(n1065), .C(n1073), .Q(n1072) );
  INV3 U270 ( .A(n1074), .Q(n1978) );
  NAND31 U271 ( .A(i_con_RegWr), .B(n1065), .C(n1075), .Q(n1074) );
  INV3 U272 ( .A(n1076), .Q(n1977) );
  NAND31 U273 ( .A(i_con_RegWr), .B(n1065), .C(n1077), .Q(n1076) );
  INV3 U274 ( .A(n1078), .Q(n1976) );
  NAND31 U275 ( .A(i_con_RegWr), .B(n1065), .C(n1079), .Q(n1078) );
  BUF2 U276 ( .A(n1427), .Q(n1425) );
  BUF2 U277 ( .A(n1427), .Q(n1426) );
  BUF2 U278 ( .A(i_addr_Rs[0]), .Q(n1822) );
  BUF2 U279 ( .A(i_addr_Rt[0]), .Q(n1449) );
  BUF2 U280 ( .A(i_addr_Rt[0]), .Q(n1450) );
  BUF2 U281 ( .A(n1429), .Q(n1408) );
  BUF2 U282 ( .A(n1429), .Q(n1407) );
  BUF2 U283 ( .A(n1428), .Q(n1406) );
  BUF2 U284 ( .A(n1428), .Q(n1405) );
  BUF2 U285 ( .A(n1428), .Q(n1404) );
  MUX22 U286 ( .A(n1616), .B(n1611), .S(i_addr_Rs[4]), .Q(o_data_Rs[16]) );
  IMUX40 U287 ( .A(n1617), .B(n1618), .C(n1619), .D(n1620), .S0(n1775), .S1(
        n1778), .Q(n1616) );
  IMUX40 U288 ( .A(n1612), .B(n1613), .C(n1614), .D(n1615), .S0(n1775), .S1(
        n1778), .Q(n1611) );
  IMUX40 U289 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n1819), .S1(n1799), .Q(n1617) );
  IMUX40 U290 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n1818), .S1(n1789), .Q(n1460) );
  IMUX40 U291 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n1818), .S1(n1789), .Q(n1458) );
  IMUX40 U292 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n1818), .S1(n1789), .Q(n1457) );
  IMUX40 U293 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(n1822), .S1(n1788), .Q(n1455) );
  IMUX40 U294 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(n1822), .S1(n1788), .Q(n1453) );
  IMUX40 U295 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(n1822), .S1(n1788), .Q(n1452) );
  IMUX40 U296 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n1818), .S1(n1789), .Q(n1465) );
  IMUX40 U297 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n1), .S1(n1789), .Q(n1463) );
  IMUX40 U298 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n1817), .S1(n1789), .Q(n1462) );
  IMUX40 U299 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n1818), .S1(n1789), .Q(n1470) );
  IMUX40 U300 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n1819), .S1(n1790), .Q(n1468) );
  IMUX40 U301 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n1815), .S1(n1790), .Q(n1475) );
  IMUX40 U302 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n1815), .S1(n1790), .Q(n1473) );
  IMUX40 U303 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n1818), .S1(n1790), .Q(n1472) );
  IMUX40 U304 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n1818), .S1(n1790), .Q(n1480) );
  IMUX40 U305 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n1818), .S1(n1790), .Q(n1478) );
  IMUX40 U306 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n1815), .S1(n1791), .Q(n1485) );
  IMUX40 U307 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n1815), .S1(n1791), .Q(n1483) );
  IMUX40 U308 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n1818), .S1(n1791), .Q(n1482) );
  IMUX40 U309 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n1816), .S1(n1791), .Q(n1490) );
  IMUX40 U310 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n1816), .S1(n1791), .Q(n1488) );
  IMUX40 U311 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n1816), .S1(n1792), .Q(n1495) );
  IMUX40 U312 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n1816), .S1(n1792), .Q(n1493) );
  IMUX40 U313 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n1816), .S1(n1792), .Q(n1492) );
  IMUX40 U314 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n1816), .S1(n1792), .Q(n1500) );
  IMUX40 U315 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n1816), .S1(n1792), .Q(n1498) );
  IMUX40 U316 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n1822), .S1(n1793), .Q(n1505) );
  IMUX40 U317 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n1817), .S1(n1793), .Q(n1503) );
  IMUX40 U318 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n1822), .S1(n1793), .Q(n1502) );
  IMUX40 U319 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n1818), .S1(n1793), .Q(n1510) );
  IMUX40 U320 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n1817), .S1(n1793), .Q(n1508) );
  IMUX40 U321 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n1822), .S1(n1793), .Q(n1515) );
  IMUX40 U322 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n1822), .S1(n1785), .Q(n1513) );
  IMUX40 U323 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n1818), .S1(n1785), .Q(n1512) );
  IMUX40 U324 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n1817), .S1(n1785), .Q(n1520) );
  IMUX40 U325 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n1817), .S1(n1785), .Q(n1518) );
  IMUX40 U326 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n1817), .S1(n1785), .Q(n1525) );
  IMUX40 U327 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n1817), .S1(n1794), .Q(n1523) );
  IMUX40 U328 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n1817), .S1(n1788), .Q(n1522) );
  IMUX40 U329 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n1817), .S1(n1788), .Q(n1530) );
  IMUX40 U330 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n1817), .S1(n1811), .Q(n1528) );
  IMUX40 U331 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n1818), .S1(n1811), .Q(n1535) );
  IMUX40 U332 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n1818), .S1(n1811), .Q(n1533) );
  IMUX40 U333 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n1818), .S1(n1785), .Q(n1532) );
  IMUX40 U334 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n1818), .S1(n1787), .Q(n1540) );
  IMUX40 U335 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n1818), .S1(n1783), .Q(n1538) );
  IMUX40 U336 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n1818), .S1(n1806), .Q(n1545) );
  IMUX40 U337 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n1818), .S1(n1797), .Q(n1543) );
  IMUX40 U338 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n1818), .S1(n1801), .Q(n1542) );
  IMUX40 U339 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n1820), .S1(n1794), .Q(n1550) );
  IMUX40 U340 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n1820), .S1(n1794), .Q(n1548) );
  IMUX40 U341 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n1820), .S1(n1794), .Q(n1555) );
  IMUX40 U342 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n1820), .S1(n1794), .Q(n1553) );
  IMUX40 U343 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n1820), .S1(n1794), .Q(n1552) );
  IMUX40 U344 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n1820), .S1(n1794), .Q(n1560) );
  IMUX40 U345 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n1820), .S1(n1795), .Q(n1558) );
  IMUX40 U346 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n1818), .S1(n1795), .Q(n1565) );
  IMUX40 U347 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n1818), .S1(n1795), .Q(n1563) );
  IMUX40 U348 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n1817), .S1(n1795), .Q(n1562) );
  IMUX40 U349 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n1818), .S1(n1795), .Q(n1570) );
  IMUX40 U350 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n1818), .S1(n1795), .Q(n1568) );
  IMUX40 U351 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n1817), .S1(n1796), .Q(n1575) );
  IMUX40 U352 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n1818), .S1(n1796), .Q(n1573) );
  IMUX40 U353 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n1818), .S1(n1796), .Q(n1572) );
  IMUX40 U354 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n1), .S1(n1796), .Q(n1580) );
  IMUX40 U355 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n1818), .S1(n1796), .Q(n1578) );
  IMUX40 U356 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n1), .S1(n1792), .Q(n1585) );
  IMUX40 U357 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n1), .S1(n1784), .Q(n1583) );
  IMUX40 U358 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n1), .S1(n1783), .Q(n1582) );
  IMUX40 U359 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n1), .S1(n1787), .Q(n1590) );
  IMUX40 U360 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n1), .S1(n1791), .Q(n1588) );
  IMUX40 U361 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n1819), .S1(n1797), .Q(n1595) );
  IMUX40 U362 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n1), .S1(n1797), .Q(n1593) );
  IMUX40 U363 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n1818), .S1(n1797), .Q(n1592) );
  IMUX40 U364 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n1), .S1(n1797), .Q(n1600) );
  IMUX40 U365 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n1819), .S1(n1797), .Q(n1598) );
  IMUX40 U366 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n1817), .S1(n1797), .Q(n1605) );
  IMUX40 U367 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n1818), .S1(n1798), .Q(n1603) );
  IMUX40 U368 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n1816), .S1(n1798), .Q(n1602) );
  IMUX40 U369 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n1819), .S1(n1798), .Q(n1610) );
  IMUX40 U370 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n1817), .S1(n1798), .Q(n1608) );
  IMUX40 U371 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n1817), .S1(n1798), .Q(n1615) );
  IMUX40 U372 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n1819), .S1(n1798), .Q(n1613) );
  IMUX40 U373 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n1817), .S1(n1799), .Q(n1612) );
  IMUX40 U374 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n1819), .S1(n1799), .Q(n1620) );
  IMUX40 U375 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n1819), .S1(n1799), .Q(n1618) );
  IMUX40 U376 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n1820), .S1(n1799), .Q(n1625) );
  IMUX40 U377 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n1820), .S1(n1799), .Q(n1623) );
  IMUX40 U378 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n1820), .S1(n1800), .Q(n1622) );
  IMUX40 U379 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n1820), .S1(n1800), .Q(n1630) );
  IMUX40 U380 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n1820), .S1(n1800), .Q(n1628) );
  IMUX40 U381 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n1820), .S1(n1800), .Q(n1635) );
  IMUX40 U382 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n1820), .S1(n1800), .Q(n1633) );
  IMUX40 U383 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n1820), .S1(n1800), .Q(n1632) );
  IMUX40 U384 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n1819), .S1(n1801), .Q(n1640) );
  IMUX40 U385 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n1), .S1(n1801), .Q(n1638) );
  IMUX40 U386 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n1819), .S1(n1801), .Q(n1645) );
  IMUX40 U387 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n1), .S1(n1801), .Q(n1643) );
  IMUX40 U388 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n1818), .S1(n1801), .Q(n1642) );
  IMUX40 U389 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n1819), .S1(n1801), .Q(n1650) );
  IMUX40 U390 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n1819), .S1(n1802), .Q(n1648) );
  IMUX40 U391 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n1819), .S1(n1802), .Q(n1655) );
  IMUX40 U392 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n1819), .S1(n1802), .Q(n1653) );
  IMUX40 U393 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n1819), .S1(n1802), .Q(n1652) );
  IMUX40 U394 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n1819), .S1(n1802), .Q(n1660) );
  IMUX40 U395 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n1817), .S1(n1802), .Q(n1658) );
  IMUX40 U396 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n1818), .S1(n1803), .Q(n1665) );
  IMUX40 U397 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n1819), .S1(n1803), .Q(n1663) );
  IMUX40 U398 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n1818), .S1(n1803), .Q(n1662) );
  IMUX40 U399 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n1), .S1(n1803), .Q(n1670) );
  IMUX40 U400 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n1), .S1(n1803), .Q(n1668) );
  IMUX40 U401 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n1), .S1(n1804), .Q(n1675) );
  IMUX40 U402 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n1), .S1(n1804), .Q(n1673) );
  IMUX40 U403 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n1), .S1(n1804), .Q(n1672) );
  IMUX40 U404 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n1), .S1(n1804), .Q(n1680) );
  IMUX40 U405 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n1), .S1(n1804), .Q(n1678) );
  IMUX40 U406 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n1817), .S1(n1805), .Q(n1685) );
  IMUX40 U407 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n2), .S1(n1805), .Q(n1683) );
  IMUX40 U408 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n2), .S1(n1805), .Q(n1682) );
  IMUX40 U409 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n1818), .S1(n1805), .Q(n1690) );
  IMUX40 U410 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n1818), .S1(n1805), .Q(n1688) );
  IMUX40 U411 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n1820), .S1(n1805), .Q(n1695) );
  IMUX40 U412 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n1817), .S1(n1806), .Q(n1693) );
  IMUX40 U413 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n1819), .S1(n1806), .Q(n1692) );
  IMUX40 U414 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n1816), .S1(n1806), .Q(n1700) );
  IMUX40 U415 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n1820), .S1(n1806), .Q(n1698) );
  IMUX40 U416 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n1820), .S1(n1806), .Q(n1705) );
  IMUX40 U417 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n1820), .S1(n1806), .Q(n1703) );
  IMUX40 U418 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n1), .S1(n1807), .Q(n1702) );
  IMUX40 U419 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n1818), .S1(n1807), .Q(n1710) );
  IMUX40 U420 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n1817), .S1(n1807), .Q(n1708) );
  IMUX40 U421 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n1818), .S1(n1807), .Q(n1715) );
  IMUX40 U422 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n1818), .S1(n1807), .Q(n1713) );
  IMUX40 U423 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n1818), .S1(n1808), .Q(n1712) );
  IMUX40 U424 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n1818), .S1(n1808), .Q(n1720) );
  IMUX40 U425 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n1818), .S1(n1808), .Q(n1718) );
  IMUX40 U426 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n1818), .S1(n1808), .Q(n1725) );
  IMUX40 U427 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n1818), .S1(n1808), .Q(n1723) );
  IMUX40 U428 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n1818), .S1(n1808), .Q(n1722) );
  IMUX40 U429 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n2), .S1(n1809), .Q(n1730) );
  IMUX40 U430 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n2), .S1(n1809), .Q(n1728) );
  IMUX40 U431 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n2), .S1(n1809), .Q(n1735) );
  IMUX40 U432 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n2), .S1(n1809), .Q(n1733) );
  IMUX40 U433 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n2), .S1(n1809), .Q(n1732) );
  IMUX40 U434 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n2), .S1(n1809), .Q(n1740) );
  IMUX40 U435 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n2), .S1(n1810), .Q(n1738) );
  IMUX40 U436 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n1821), .S1(n1810), .Q(n1745) );
  IMUX40 U437 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n2), .S1(n1810), .Q(n1743) );
  IMUX40 U438 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n1821), .S1(n1810), .Q(n1742) );
  IMUX40 U439 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n2), .S1(n1810), .Q(n1750) );
  IMUX40 U440 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n1821), .S1(n1810), .Q(n1748) );
  IMUX40 U441 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n2), .S1(n1794), .Q(n1755) );
  IMUX40 U442 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n1821), .S1(n1795), .Q(n1753) );
  IMUX40 U443 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n2), .S1(n1811), .Q(n1752) );
  IMUX40 U444 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n1816), .S1(n1794), .Q(n1760) );
  IMUX40 U445 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n2), .S1(n1795), .Q(n1758) );
  IMUX40 U446 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n1821), .S1(n1785), .Q(n1765) );
  IMUX40 U447 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n2), .S1(n1794), .Q(n1763) );
  IMUX40 U448 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n2), .S1(n1794), .Q(n1762) );
  IMUX40 U449 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n2), .S1(n1785), .Q(n1770) );
  IMUX40 U450 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n2), .S1(n1797), .Q(n1768) );
  IMUX40 U451 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n1815), .S1(n1789), .Q(n1459) );
  IMUX40 U452 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(n1822), .S1(n1788), .Q(n1454) );
  IMUX40 U453 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n1819), .S1(n1789), .Q(n1464) );
  IMUX40 U454 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n1816), .S1(n1790), .Q(n1469) );
  IMUX40 U455 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n1815), .S1(n1790), .Q(n1474) );
  IMUX40 U456 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n1818), .S1(n1791), .Q(n1479) );
  IMUX40 U457 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n1815), .S1(n1791), .Q(n1484) );
  IMUX40 U458 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n1816), .S1(n1791), .Q(n1489) );
  IMUX40 U459 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n1816), .S1(n1792), .Q(n1494) );
  IMUX40 U460 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n1816), .S1(n1792), .Q(n1499) );
  IMUX40 U461 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n1822), .S1(n1793), .Q(n1504) );
  IMUX40 U462 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n1817), .S1(n1793), .Q(n1509) );
  IMUX40 U463 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n1822), .S1(n1785), .Q(n1514) );
  IMUX40 U464 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n1817), .S1(n1785), .Q(n1519) );
  IMUX40 U465 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n1817), .S1(n1788), .Q(n1524) );
  IMUX40 U466 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n1817), .S1(n1788), .Q(n1529) );
  IMUX40 U467 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n1818), .S1(n1811), .Q(n1534) );
  IMUX40 U468 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n1818), .S1(n1785), .Q(n1539) );
  IMUX40 U469 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n1818), .S1(n1805), .Q(n1544) );
  IMUX40 U470 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n1820), .S1(n1794), .Q(n1549) );
  IMUX40 U471 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n1820), .S1(n1794), .Q(n1554) );
  IMUX40 U472 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n1820), .S1(n1795), .Q(n1559) );
  IMUX40 U473 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n1817), .S1(n1795), .Q(n1564) );
  IMUX40 U474 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n1817), .S1(n1796), .Q(n1569) );
  IMUX40 U475 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n1818), .S1(n1796), .Q(n1574) );
  IMUX40 U476 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n1820), .S1(n1796), .Q(n1579) );
  IMUX40 U477 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n1818), .S1(n1795), .Q(n1584) );
  IMUX40 U478 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n1820), .S1(n1782), .Q(n1589) );
  IMUX40 U479 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n1817), .S1(n1797), .Q(n1594) );
  IMUX40 U480 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n1818), .S1(n1797), .Q(n1599) );
  IMUX40 U481 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n1819), .S1(n1798), .Q(n1604) );
  IMUX40 U482 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n1819), .S1(n1798), .Q(n1609) );
  IMUX40 U483 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n1817), .S1(n1799), .Q(n1614) );
  IMUX40 U484 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n1819), .S1(n1799), .Q(n1619) );
  IMUX40 U485 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n1820), .S1(n1799), .Q(n1624) );
  IMUX40 U486 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n1820), .S1(n1800), .Q(n1629) );
  IMUX40 U487 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n1820), .S1(n1800), .Q(n1634) );
  IMUX40 U488 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n1816), .S1(n1801), .Q(n1639) );
  IMUX40 U489 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n1815), .S1(n1801), .Q(n1644) );
  IMUX40 U490 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n1), .S1(n1802), .Q(n1649) );
  IMUX40 U491 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n1819), .S1(n1802), .Q(n1654) );
  IMUX40 U492 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n1), .S1(n1803), .Q(n1659) );
  IMUX40 U493 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n1819), .S1(n1803), .Q(n1664) );
  IMUX40 U494 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n1), .S1(n1803), .Q(n1669) );
  IMUX40 U495 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n1), .S1(n1804), .Q(n1674) );
  IMUX40 U496 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n1), .S1(n1804), .Q(n1679) );
  IMUX40 U497 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n1821), .S1(n1805), .Q(n1684) );
  IMUX40 U498 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n1), .S1(n1805), .Q(n1689) );
  IMUX40 U499 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n1), .S1(n1806), .Q(n1694) );
  IMUX40 U500 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n1820), .S1(n1806), .Q(n1699) );
  IMUX40 U501 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n1820), .S1(n1807), .Q(n1704) );
  IMUX40 U502 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n1820), .S1(n1807), .Q(n1709) );
  IMUX40 U503 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n1818), .S1(n1807), .Q(n1714) );
  IMUX40 U504 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n1818), .S1(n1808), .Q(n1719) );
  IMUX40 U505 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n1818), .S1(n1808), .Q(n1724) );
  IMUX40 U506 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n2), .S1(n1809), .Q(n1729) );
  IMUX40 U507 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n2), .S1(n1809), .Q(n1734) );
  IMUX40 U508 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n2), .S1(n1810), .Q(n1739) );
  IMUX40 U509 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n1821), .S1(n1810), .Q(n1744) );
  IMUX40 U510 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n2), .S1(n1811), .Q(n1749) );
  IMUX40 U511 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n1821), .S1(n1796), .Q(n1754) );
  IMUX40 U512 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n1817), .S1(n1785), .Q(n1759) );
  IMUX40 U513 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n1), .S1(n1795), .Q(n1764) );
  IMUX40 U514 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n1818), .S1(n1795), .Q(n1769) );
  MUX22 U515 ( .A(n1556), .B(n1551), .S(i_addr_Rs[4]), .Q(o_data_Rs[10]) );
  IMUX40 U516 ( .A(n1557), .B(n1558), .C(n1559), .D(n1560), .S0(n1774), .S1(
        n1777), .Q(n1556) );
  IMUX40 U517 ( .A(n1552), .B(n1553), .C(n1554), .D(n1555), .S0(n1774), .S1(
        n1777), .Q(n1551) );
  IMUX40 U518 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n1820), .S1(n1795), .Q(n1557) );
  MUX22 U519 ( .A(n1566), .B(n1561), .S(n1771), .Q(o_data_Rs[11]) );
  IMUX40 U520 ( .A(n1567), .B(n1568), .C(n1569), .D(n1570), .S0(n1774), .S1(
        n1777), .Q(n1566) );
  IMUX40 U521 ( .A(n1562), .B(n1563), .C(n1564), .D(n1565), .S0(n1774), .S1(
        n1777), .Q(n1561) );
  IMUX40 U522 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n1818), .S1(n1796), .Q(n1567) );
  MUX22 U523 ( .A(n1596), .B(n1591), .S(i_addr_Rs[4]), .Q(o_data_Rs[14]) );
  IMUX40 U524 ( .A(n1597), .B(n1598), .C(n1599), .D(n1600), .S0(n1775), .S1(
        n1778), .Q(n1596) );
  IMUX40 U525 ( .A(n1592), .B(n1593), .C(n1594), .D(n1595), .S0(n1775), .S1(
        n1778), .Q(n1591) );
  IMUX40 U526 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n1), .S1(n1797), .Q(n1597) );
  MUX22 U527 ( .A(n1606), .B(n1601), .S(i_addr_Rs[4]), .Q(o_data_Rs[15]) );
  IMUX40 U528 ( .A(n1607), .B(n1608), .C(n1609), .D(n1610), .S0(n1775), .S1(
        n1778), .Q(n1606) );
  IMUX40 U529 ( .A(n1602), .B(n1603), .C(n1604), .D(n1605), .S0(n1775), .S1(
        n1778), .Q(n1601) );
  IMUX40 U530 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n1817), .S1(n1798), .Q(n1607) );
  MUX22 U531 ( .A(n1626), .B(n1621), .S(i_addr_Rs[4]), .Q(o_data_Rs[17]) );
  IMUX40 U532 ( .A(n1627), .B(n1628), .C(n1629), .D(n1630), .S0(n1775), .S1(
        n1778), .Q(n1626) );
  IMUX40 U533 ( .A(n1622), .B(n1623), .C(n1624), .D(n1625), .S0(n1775), .S1(
        n1778), .Q(n1621) );
  IMUX40 U534 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n1820), .S1(n1800), .Q(n1627) );
  MUX22 U535 ( .A(n1636), .B(n1631), .S(i_addr_Rs[4]), .Q(o_data_Rs[18]) );
  IMUX40 U536 ( .A(n1637), .B(n1638), .C(n1639), .D(n1640), .S0(n1775), .S1(
        n1779), .Q(n1636) );
  IMUX40 U537 ( .A(n1632), .B(n1633), .C(n1634), .D(n1635), .S0(n1775), .S1(
        n1778), .Q(n1631) );
  IMUX40 U538 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n1818), .S1(n1801), .Q(n1637) );
  MUX22 U539 ( .A(n1646), .B(n1641), .S(n1772), .Q(o_data_Rs[19]) );
  IMUX40 U540 ( .A(n1647), .B(n1648), .C(n1649), .D(n1650), .S0(n1775), .S1(
        n1779), .Q(n1646) );
  IMUX40 U541 ( .A(n1642), .B(n1643), .C(n1644), .D(n1645), .S0(n1775), .S1(
        n1779), .Q(n1641) );
  IMUX40 U542 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n1), .S1(n1802), .Q(n1647) );
  MUX22 U543 ( .A(n1656), .B(n1651), .S(n1772), .Q(o_data_Rs[20]) );
  IMUX40 U544 ( .A(n1657), .B(n1658), .C(n1659), .D(n1660), .S0(n1776), .S1(
        n1779), .Q(n1656) );
  IMUX40 U545 ( .A(n1652), .B(n1653), .C(n1654), .D(n1655), .S0(n1776), .S1(
        n1779), .Q(n1651) );
  IMUX40 U546 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n1819), .S1(n1803), .Q(n1657) );
  MUX22 U547 ( .A(n1666), .B(n1661), .S(n1772), .Q(o_data_Rs[21]) );
  IMUX40 U548 ( .A(n1667), .B(n1668), .C(n1669), .D(n1670), .S0(n1776), .S1(
        n1779), .Q(n1666) );
  IMUX40 U549 ( .A(n1662), .B(n1663), .C(n1664), .D(n1665), .S0(n1776), .S1(
        n1779), .Q(n1661) );
  IMUX40 U550 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n1), .S1(n1804), .Q(n1667) );
  MUX22 U551 ( .A(n1676), .B(n1671), .S(n1772), .Q(o_data_Rs[22]) );
  IMUX40 U552 ( .A(n1677), .B(n1678), .C(n1679), .D(n1680), .S0(n1776), .S1(
        n1779), .Q(n1676) );
  IMUX40 U553 ( .A(n1672), .B(n1673), .C(n1674), .D(n1675), .S0(n1776), .S1(
        n1779), .Q(n1671) );
  IMUX40 U554 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n1), .S1(n1804), .Q(n1677) );
  MUX22 U555 ( .A(n1686), .B(n1681), .S(n1772), .Q(o_data_Rs[23]) );
  IMUX40 U556 ( .A(n1687), .B(n1688), .C(n1689), .D(n1690), .S0(n1776), .S1(
        i_addr_Rs[2]), .Q(n1686) );
  IMUX40 U557 ( .A(n1682), .B(n1683), .C(n1684), .D(n1685), .S0(n1776), .S1(
        i_addr_Rs[2]), .Q(n1681) );
  IMUX40 U558 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n1820), .S1(n1805), .Q(n1687) );
  MUX22 U559 ( .A(n1696), .B(n1691), .S(n1772), .Q(o_data_Rs[24]) );
  IMUX40 U560 ( .A(n1697), .B(n1698), .C(n1699), .D(n1700), .S0(n1776), .S1(
        i_addr_Rs[2]), .Q(n1696) );
  IMUX40 U561 ( .A(n1692), .B(n1693), .C(n1694), .D(n1695), .S0(n1776), .S1(
        i_addr_Rs[2]), .Q(n1691) );
  IMUX40 U562 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n1818), .S1(n1806), .Q(n1697) );
  MUX22 U563 ( .A(n1706), .B(n1701), .S(n1772), .Q(o_data_Rs[25]) );
  IMUX40 U564 ( .A(n1707), .B(n1708), .C(n1709), .D(n1710), .S0(n1776), .S1(
        i_addr_Rs[2]), .Q(n1706) );
  IMUX40 U565 ( .A(n1702), .B(n1703), .C(n1704), .D(n1705), .S0(n1776), .S1(
        i_addr_Rs[2]), .Q(n1701) );
  IMUX40 U566 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n1818), .S1(n1807), .Q(n1707) );
  MUX22 U567 ( .A(n1716), .B(n1711), .S(n1772), .Q(o_data_Rs[26]) );
  IMUX40 U568 ( .A(n1717), .B(n1718), .C(n1719), .D(n1720), .S0(n1774), .S1(
        i_addr_Rs[2]), .Q(n1716) );
  IMUX40 U569 ( .A(n1712), .B(n1713), .C(n1714), .D(n1715), .S0(n1774), .S1(
        n1779), .Q(n1711) );
  IMUX40 U570 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n1818), .S1(n1808), .Q(n1717) );
  MUX22 U571 ( .A(n1726), .B(n1721), .S(n1772), .Q(o_data_Rs[27]) );
  IMUX40 U572 ( .A(n1727), .B(n1728), .C(n1729), .D(n1730), .S0(n1773), .S1(
        n1780), .Q(n1726) );
  IMUX40 U573 ( .A(n1722), .B(n1723), .C(n1724), .D(n1725), .S0(n1774), .S1(
        i_addr_Rs[2]), .Q(n1721) );
  IMUX40 U574 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n2), .S1(n1809), .Q(n1727) );
  MUX22 U575 ( .A(n1736), .B(n1731), .S(n1772), .Q(o_data_Rs[28]) );
  IMUX40 U576 ( .A(n1737), .B(n1738), .C(n1739), .D(n1740), .S0(n1774), .S1(
        n1780), .Q(n1736) );
  IMUX40 U577 ( .A(n1732), .B(n1733), .C(n1734), .D(n1735), .S0(n1774), .S1(
        n1780), .Q(n1731) );
  IMUX40 U578 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n2), .S1(n1810), .Q(n1737) );
  MUX22 U579 ( .A(n1746), .B(n1741), .S(n1772), .Q(o_data_Rs[29]) );
  IMUX40 U580 ( .A(n1747), .B(n1748), .C(n1749), .D(n1750), .S0(n1774), .S1(
        n1780), .Q(n1746) );
  IMUX40 U581 ( .A(n1742), .B(n1743), .C(n1744), .D(n1745), .S0(n1773), .S1(
        n1780), .Q(n1741) );
  IMUX40 U582 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n1), .S1(n1785), .Q(n1747) );
  MUX22 U583 ( .A(n1756), .B(n1751), .S(n1772), .Q(o_data_Rs[30]) );
  IMUX40 U584 ( .A(n1757), .B(n1758), .C(n1759), .D(n1760), .S0(n1774), .S1(
        n1780), .Q(n1756) );
  IMUX40 U585 ( .A(n1752), .B(n1753), .C(n1754), .D(n1755), .S0(n1774), .S1(
        n1780), .Q(n1751) );
  IMUX40 U586 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n1816), .S1(n1795), .Q(n1757) );
  MUX22 U587 ( .A(n1766), .B(n1761), .S(n1772), .Q(o_data_Rs[31]) );
  IMUX40 U588 ( .A(n1767), .B(n1768), .C(n1769), .D(n1770), .S0(n1774), .S1(
        n1780), .Q(n1766) );
  IMUX40 U589 ( .A(n1762), .B(n1763), .C(n1764), .D(n1765), .S0(n1773), .S1(
        n1780), .Q(n1761) );
  IMUX40 U590 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n1819), .S1(n1785), .Q(n1767) );
  BUF2 U591 ( .A(i_addr_Rs[1]), .Q(n1814) );
  BUF2 U592 ( .A(i_addr_Rs[1]), .Q(n1813) );
  BUF2 U593 ( .A(i_addr_Rs[1]), .Q(n1812) );
  MUX22 U594 ( .A(n1456), .B(n1451), .S(n1771), .Q(o_data_Rs[0]) );
  IMUX40 U595 ( .A(n1452), .B(n1453), .C(n1454), .D(n1455), .S0(n1773), .S1(
        n1778), .Q(n1451) );
  IMUX40 U596 ( .A(n1457), .B(n1458), .C(n1459), .D(n1460), .S0(n1773), .S1(
        i_addr_Rs[2]), .Q(n1456) );
  MUX22 U597 ( .A(n1466), .B(n1461), .S(n1771), .Q(o_data_Rs[1]) );
  IMUX40 U598 ( .A(n1467), .B(n1468), .C(n1469), .D(n1470), .S0(n1773), .S1(
        n1780), .Q(n1466) );
  IMUX40 U599 ( .A(n1462), .B(n1463), .C(n1464), .D(n1465), .S0(n1773), .S1(
        n1778), .Q(n1461) );
  IMUX40 U600 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(n2), 
        .S1(n1790), .Q(n1467) );
  MUX22 U601 ( .A(n1476), .B(n1471), .S(n1771), .Q(o_data_Rs[2]) );
  IMUX40 U602 ( .A(n1477), .B(n1478), .C(n1479), .D(n1480), .S0(n1774), .S1(
        i_addr_Rs[2]), .Q(n1476) );
  IMUX40 U603 ( .A(n1472), .B(n1473), .C(n1474), .D(n1475), .S0(n1774), .S1(
        n1780), .Q(n1471) );
  IMUX40 U604 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n1818), .S1(n1791), .Q(n1477) );
  MUX22 U605 ( .A(n1486), .B(n1481), .S(n1771), .Q(o_data_Rs[3]) );
  IMUX40 U606 ( .A(n1487), .B(n1488), .C(n1489), .D(n1490), .S0(n1774), .S1(
        n1779), .Q(n1486) );
  IMUX40 U607 ( .A(n1482), .B(n1483), .C(n1484), .D(n1485), .S0(n1774), .S1(
        n1779), .Q(n1481) );
  IMUX40 U608 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n1816), .S1(n1792), .Q(n1487) );
  MUX22 U609 ( .A(n1496), .B(n1491), .S(n1771), .Q(o_data_Rs[4]) );
  IMUX40 U610 ( .A(n1497), .B(n1498), .C(n1499), .D(n1500), .S0(n1774), .S1(
        n1780), .Q(n1496) );
  IMUX40 U611 ( .A(n1492), .B(n1493), .C(n1494), .D(n1495), .S0(n1774), .S1(
        n1778), .Q(n1491) );
  IMUX40 U612 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n1816), .S1(n1792), .Q(n1497) );
  MUX22 U613 ( .A(n1506), .B(n1501), .S(n1771), .Q(o_data_Rs[5]) );
  IMUX40 U614 ( .A(n1507), .B(n1508), .C(n1509), .D(n1510), .S0(n1773), .S1(
        i_addr_Rs[2]), .Q(n1506) );
  IMUX40 U615 ( .A(n1502), .B(n1503), .C(n1504), .D(n1505), .S0(n1774), .S1(
        n1777), .Q(n1501) );
  IMUX40 U616 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n1815), .S1(n1793), .Q(n1507) );
  MUX22 U617 ( .A(n1516), .B(n1511), .S(n1771), .Q(o_data_Rs[6]) );
  IMUX40 U618 ( .A(n1517), .B(n1518), .C(n1519), .D(n1520), .S0(n1774), .S1(
        i_addr_Rs[2]), .Q(n1516) );
  IMUX40 U619 ( .A(n1512), .B(n1513), .C(n1514), .D(n1515), .S0(n1774), .S1(
        i_addr_Rs[2]), .Q(n1511) );
  IMUX40 U620 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n1817), .S1(n1785), .Q(n1517) );
  MUX22 U621 ( .A(n1526), .B(n1521), .S(i_addr_Rs[4]), .Q(o_data_Rs[7]) );
  IMUX40 U622 ( .A(n1527), .B(n1528), .C(n1529), .D(n1530), .S0(n1773), .S1(
        n1779), .Q(n1526) );
  IMUX40 U623 ( .A(n1522), .B(n1523), .C(n1524), .D(n1525), .S0(n1773), .S1(
        n1780), .Q(n1521) );
  IMUX40 U624 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n1817), .S1(n1783), .Q(n1527) );
  MUX22 U625 ( .A(n1536), .B(n1531), .S(n1771), .Q(o_data_Rs[8]) );
  IMUX40 U626 ( .A(n1537), .B(n1538), .C(n1539), .D(n1540), .S0(n1774), .S1(
        i_addr_Rs[2]), .Q(n1536) );
  IMUX40 U627 ( .A(n1532), .B(n1533), .C(n1534), .D(n1535), .S0(n1774), .S1(
        i_addr_Rs[2]), .Q(n1531) );
  IMUX40 U628 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n1818), .S1(n1781), .Q(n1537) );
  MUX22 U629 ( .A(n1546), .B(n1541), .S(i_addr_Rs[4]), .Q(o_data_Rs[9]) );
  IMUX40 U630 ( .A(n1547), .B(n1548), .C(n1549), .D(n1550), .S0(n1774), .S1(
        n1777), .Q(n1546) );
  IMUX40 U631 ( .A(n1542), .B(n1543), .C(n1544), .D(n1545), .S0(n1774), .S1(
        n1778), .Q(n1541) );
  IMUX40 U632 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n1820), .S1(n1794), .Q(n1547) );
  MUX22 U633 ( .A(n1576), .B(n1571), .S(n1771), .Q(o_data_Rs[12]) );
  IMUX40 U634 ( .A(n1572), .B(n1573), .C(n1574), .D(n1575), .S0(n1774), .S1(
        n1777), .Q(n1571) );
  IMUX40 U635 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n1818), .S1(n1784), .Q(n1577) );
  MUX22 U636 ( .A(n1586), .B(n1581), .S(n1771), .Q(o_data_Rs[13]) );
  IMUX40 U637 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n1818), .S1(n1794), .Q(n1587) );
  BUF2 U638 ( .A(i_addr_Rs[1]), .Q(n1811) );
  NOR21 U639 ( .A(n1984), .B(i_addr_Rd[4]), .Q(n1081) );
  NOR21 U640 ( .A(n1967), .B(i_addr_Rd[3]), .Q(n1090) );
  NOR21 U641 ( .A(i_addr_Rd[4]), .B(i_addr_Rd[3]), .Q(n1065) );
  IMUX40 U642 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n1430), .S1(n1427), .Q(n1036) );
  IMUX40 U643 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n1430), .S1(n1428), .Q(n1034) );
  IMUX40 U644 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n1430), .S1(n1427), .Q(n1033) );
  IMUX40 U645 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(i_addr_Rt[0]), .S1(n1428), .Q(n1031) );
  IMUX40 U646 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(i_addr_Rt[0]), .S1(n1408), .Q(n1029) );
  IMUX40 U647 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(i_addr_Rt[0]), .S1(n1412), .Q(n1028) );
  IMUX40 U648 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n1430), .S1(n1404), .Q(n1041) );
  IMUX40 U649 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n1430), .S1(n1427), .Q(n1039) );
  IMUX40 U650 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n1430), .S1(n1407), .Q(n1038) );
  IMUX40 U651 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n1430), .S1(n1426), .Q(n1046) );
  IMUX40 U652 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n1430), .S1(n1405), .Q(n1044) );
  IMUX40 U653 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n1431), .S1(n1406), .Q(n1051) );
  IMUX40 U654 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n1431), .S1(n1405), .Q(n1049) );
  IMUX40 U655 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n1431), .S1(n1411), .Q(n1048) );
  IMUX40 U656 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n1431), .S1(n1428), .Q(n1056) );
  IMUX40 U657 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n1431), .S1(n1410), .Q(n1054) );
  IMUX40 U658 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n1431), .S1(n1426), .Q(n1061) );
  IMUX40 U659 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n1431), .S1(n1411), .Q(n1059) );
  IMUX40 U660 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n1431), .S1(i_addr_Rt[1]), .Q(n1058) );
  IMUX40 U661 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n1432), .S1(n1429), .Q(n1110) );
  IMUX40 U662 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n1432), .S1(i_addr_Rt[1]), .Q(n1108) );
  IMUX40 U663 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n1432), .S1(n1409), .Q(n1115) );
  IMUX40 U664 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n1432), .S1(n1404), .Q(n1113) );
  IMUX40 U665 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n1432), .S1(n1411), .Q(n1112) );
  IMUX40 U666 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n1432), .S1(n1412), .Q(n1120) );
  IMUX40 U667 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n1432), .S1(n1410), .Q(n1118) );
  IMUX40 U668 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n1433), .S1(n1407), .Q(n1125) );
  IMUX40 U669 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n1433), .S1(n1426), .Q(n1123) );
  IMUX40 U670 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n1433), .S1(n1414), .Q(n1122) );
  IMUX40 U671 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n1433), .S1(n1427), .Q(n1130) );
  IMUX40 U672 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n1433), .S1(n1413), .Q(n1128) );
  IMUX40 U673 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n1433), .S1(n1425), .Q(n1135) );
  IMUX40 U674 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n1433), .S1(n1409), .Q(n1133) );
  IMUX40 U675 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n1433), .S1(n1409), .Q(n1132) );
  IMUX40 U676 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n1434), .S1(n1409), .Q(n1140) );
  IMUX40 U677 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n1434), .S1(n1409), .Q(n1138) );
  IMUX40 U678 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n1434), .S1(n1409), .Q(n1145) );
  IMUX40 U679 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n1434), .S1(n1409), .Q(n1143) );
  IMUX40 U680 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n1434), .S1(n1408), .Q(n1142) );
  IMUX40 U681 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n1434), .S1(n1408), .Q(n1150) );
  IMUX40 U682 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n1434), .S1(n1426), .Q(n1148) );
  IMUX40 U683 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n1435), .S1(n1410), .Q(n1155) );
  IMUX40 U684 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n1435), .S1(n1408), .Q(n1153) );
  IMUX40 U685 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n1435), .S1(n1409), .Q(n1152) );
  IMUX40 U686 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n1435), .S1(n1407), .Q(n1160) );
  IMUX40 U687 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n1435), .S1(n1425), .Q(n1158) );
  IMUX40 U688 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n1435), .S1(n1409), .Q(n1165) );
  IMUX40 U689 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n1435), .S1(n1409), .Q(n1163) );
  IMUX40 U690 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n1435), .S1(n1406), .Q(n1162) );
  IMUX40 U691 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n1436), .S1(n1410), .Q(n1170) );
  IMUX40 U692 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n1436), .S1(n1410), .Q(n1168) );
  IMUX40 U693 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n1436), .S1(n1410), .Q(n1175) );
  IMUX40 U694 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n1436), .S1(n1410), .Q(n1173) );
  IMUX40 U695 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n1436), .S1(n1410), .Q(n1172) );
  IMUX40 U696 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n1436), .S1(n1410), .Q(n1180) );
  IMUX40 U697 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n1436), .S1(n1411), .Q(n1178) );
  IMUX40 U698 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n1437), .S1(n1411), .Q(n1185) );
  IMUX40 U699 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n1437), .S1(n1411), .Q(n1183) );
  IMUX40 U700 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n1437), .S1(n1411), .Q(n1182) );
  IMUX40 U701 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n1437), .S1(n1411), .Q(n1190) );
  IMUX40 U702 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n1437), .S1(n1411), .Q(n1188) );
  IMUX40 U703 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n1437), .S1(n1425), .Q(n1195) );
  IMUX40 U704 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n1437), .S1(n1406), .Q(n1193) );
  IMUX40 U705 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n1437), .S1(n1429), .Q(n1192) );
  IMUX40 U706 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n1438), .S1(n1428), .Q(n1200) );
  IMUX40 U707 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n1438), .S1(n1407), .Q(n1198) );
  IMUX40 U708 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n1438), .S1(n1406), .Q(n1205) );
  IMUX40 U709 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n1438), .S1(n1405), .Q(n1203) );
  IMUX40 U710 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n1438), .S1(n1410), .Q(n1202) );
  IMUX40 U711 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n1438), .S1(n1428), .Q(n1210) );
  IMUX40 U712 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n1438), .S1(n1425), .Q(n1208) );
  IMUX40 U713 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n1439), .S1(n1412), .Q(n1215) );
  IMUX40 U714 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n1439), .S1(n1412), .Q(n1213) );
  IMUX40 U715 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n1439), .S1(n1412), .Q(n1212) );
  IMUX40 U716 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n1439), .S1(n1412), .Q(n1220) );
  IMUX40 U717 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n1439), .S1(n1412), .Q(n1218) );
  IMUX40 U718 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n1439), .S1(n1412), .Q(n1225) );
  IMUX40 U719 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n1439), .S1(n1413), .Q(n1223) );
  IMUX40 U720 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n1439), .S1(n1413), .Q(n1222) );
  IMUX40 U721 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n1440), .S1(n1413), .Q(n1230) );
  IMUX40 U722 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n1440), .S1(n1413), .Q(n1228) );
  IMUX40 U723 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n1440), .S1(n1413), .Q(n1235) );
  IMUX40 U724 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n1440), .S1(n1413), .Q(n1233) );
  IMUX40 U725 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n1440), .S1(n1414), .Q(n1232) );
  IMUX40 U726 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n1440), .S1(n1414), .Q(n1240) );
  IMUX40 U727 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n1440), .S1(n1414), .Q(n1238) );
  IMUX40 U728 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n1441), .S1(n1414), .Q(n1245) );
  IMUX40 U729 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n1441), .S1(n1414), .Q(n1243) );
  IMUX40 U730 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n1441), .S1(n1409), .Q(n1242) );
  IMUX40 U731 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n1441), .S1(n1427), .Q(n1250) );
  IMUX40 U732 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n1441), .S1(n1427), .Q(n1248) );
  IMUX40 U733 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n1441), .S1(n1427), .Q(n1255) );
  IMUX40 U734 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n1441), .S1(n1427), .Q(n1253) );
  IMUX40 U735 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n1441), .S1(n1413), .Q(n1252) );
  IMUX40 U736 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n1438), .S1(n1415), .Q(n1260) );
  IMUX40 U737 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n1435), .S1(n1415), .Q(n1258) );
  IMUX40 U738 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n1435), .S1(n1415), .Q(n1265) );
  IMUX40 U739 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n1431), .S1(n1415), .Q(n1263) );
  IMUX40 U740 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n1432), .S1(n1415), .Q(n1262) );
  IMUX40 U741 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n1433), .S1(n1415), .Q(n1270) );
  IMUX40 U742 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n1431), .S1(n1416), .Q(n1268) );
  IMUX40 U743 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n1437), .S1(n1416), .Q(n1275) );
  IMUX40 U744 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n1431), .S1(n1416), .Q(n1273) );
  IMUX40 U745 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n1430), .S1(n1416), .Q(n1272) );
  IMUX40 U746 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n1433), .S1(n1416), .Q(n1280) );
  IMUX40 U747 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n1438), .S1(n1416), .Q(n1278) );
  IMUX40 U748 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n1434), .S1(n1417), .Q(n1285) );
  IMUX40 U749 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n1432), .S1(n1417), .Q(n1283) );
  IMUX40 U750 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n1436), .S1(n1417), .Q(n1282) );
  IMUX40 U751 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n1442), .S1(n1417), .Q(n1290) );
  IMUX40 U752 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n1442), .S1(n1417), .Q(n1288) );
  IMUX40 U753 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n1442), .S1(n1418), .Q(n1295) );
  IMUX40 U754 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n1442), .S1(n1418), .Q(n1293) );
  IMUX40 U755 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n1442), .S1(n1418), .Q(n1292) );
  IMUX40 U756 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n1442), .S1(n1418), .Q(n1300) );
  IMUX40 U757 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n1442), .S1(n1418), .Q(n1298) );
  IMUX40 U758 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n1443), .S1(n1419), .Q(n1305) );
  IMUX40 U759 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n1443), .S1(n1419), .Q(n1303) );
  IMUX40 U760 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n1443), .S1(n1419), .Q(n1302) );
  IMUX40 U761 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n1443), .S1(n1419), .Q(n1310) );
  IMUX40 U762 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n1443), .S1(n1419), .Q(n1308) );
  IMUX40 U763 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n1443), .S1(n1419), .Q(n1315) );
  IMUX40 U764 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n1443), .S1(n1420), .Q(n1313) );
  IMUX40 U765 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n1443), .S1(n1420), .Q(n1312) );
  IMUX40 U766 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n1444), .S1(n1420), .Q(n1320) );
  IMUX40 U767 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n1444), .S1(n1420), .Q(n1318) );
  IMUX40 U768 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n1444), .S1(n1420), .Q(n1325) );
  IMUX40 U769 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n1444), .S1(n1420), .Q(n1323) );
  IMUX40 U770 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n1444), .S1(n1421), .Q(n1322) );
  IMUX40 U771 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n1444), .S1(n1421), .Q(n1330) );
  IMUX40 U772 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n1444), .S1(n1421), .Q(n1328) );
  IMUX40 U773 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n1445), .S1(n1421), .Q(n1335) );
  IMUX40 U774 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n1445), .S1(n1421), .Q(n1333) );
  IMUX40 U775 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n1445), .S1(n1422), .Q(n1332) );
  IMUX40 U776 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n1445), .S1(n1422), .Q(n1340) );
  IMUX40 U777 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n1445), .S1(n1422), .Q(n1338) );
  IMUX40 U778 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n1445), .S1(n1422), .Q(n1345) );
  IMUX40 U779 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n1445), .S1(n1422), .Q(n1343) );
  IMUX40 U780 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n1445), .S1(n1422), .Q(n1342) );
  IMUX40 U781 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n1446), .S1(n1423), .Q(n1350) );
  IMUX40 U782 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n1446), .S1(n1423), .Q(n1348) );
  IMUX40 U783 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n1446), .S1(n1423), .Q(n1355) );
  IMUX40 U784 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n1446), .S1(n1423), .Q(n1353) );
  IMUX40 U785 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n1446), .S1(n1423), .Q(n1352) );
  IMUX40 U786 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n1446), .S1(n1423), .Q(n1360) );
  IMUX40 U787 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n1446), .S1(n1424), .Q(n1358) );
  IMUX40 U788 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n1447), .S1(n1424), .Q(n1365) );
  IMUX40 U789 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n1447), .S1(n1424), .Q(n1363) );
  IMUX40 U790 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n1447), .S1(n1424), .Q(n1362) );
  IMUX40 U791 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n1447), .S1(n1424), .Q(n1370) );
  IMUX40 U792 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n1447), .S1(n1424), .Q(n1368) );
  IMUX40 U793 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n1447), .S1(n1425), .Q(n1375) );
  IMUX40 U794 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n1447), .S1(n1425), .Q(n1373) );
  IMUX40 U795 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n1447), .S1(n1425), .Q(n1372) );
  IMUX40 U796 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n1448), .S1(n1425), .Q(n1380) );
  IMUX40 U797 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n1448), .S1(n1425), .Q(n1378) );
  IMUX40 U798 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n1448), .S1(n1426), .Q(n1385) );
  IMUX40 U799 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n1448), .S1(n1426), .Q(n1383) );
  IMUX40 U800 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n1448), .S1(n1426), .Q(n1382) );
  IMUX40 U801 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n1448), .S1(n1426), .Q(n1390) );
  IMUX40 U802 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n1448), .S1(n1426), .Q(n1388) );
  IMUX40 U803 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n1430), .S1(n1428), .Q(n1035) );
  IMUX40 U804 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(i_addr_Rt[0]), .S1(n1409), .Q(n1030) );
  IMUX40 U805 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n1430), .S1(n1406), .Q(n1040) );
  IMUX40 U806 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n1430), .S1(n1415), .Q(n1045) );
  IMUX40 U807 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n1431), .S1(n1405), .Q(n1050) );
  IMUX40 U808 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n1431), .S1(n1411), .Q(n1055) );
  IMUX40 U809 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n1431), .S1(n1409), .Q(n1060) );
  IMUX40 U810 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n1432), .S1(n1407), .Q(n1109) );
  IMUX40 U811 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n1432), .S1(n1409), .Q(n1114) );
  IMUX40 U812 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n1432), .S1(n1408), .Q(n1119) );
  IMUX40 U813 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n1433), .S1(n1409), .Q(n1124) );
  IMUX40 U814 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n1433), .S1(n1427), .Q(n1129) );
  IMUX40 U815 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n1433), .S1(n1409), .Q(n1134) );
  IMUX40 U816 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n1434), .S1(n1409), .Q(n1139) );
  IMUX40 U817 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n1434), .S1(n1407), .Q(n1144) );
  IMUX40 U818 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n1434), .S1(n1407), .Q(n1149) );
  IMUX40 U819 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n1435), .S1(n1409), .Q(n1154) );
  IMUX40 U820 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n1435), .S1(n1409), .Q(n1159) );
  IMUX40 U821 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n1435), .S1(n1409), .Q(n1164) );
  IMUX40 U822 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n1436), .S1(n1410), .Q(n1169) );
  IMUX40 U823 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n1436), .S1(n1410), .Q(n1174) );
  IMUX40 U824 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n1436), .S1(n1411), .Q(n1179) );
  IMUX40 U825 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n1437), .S1(n1411), .Q(n1184) );
  IMUX40 U826 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n1437), .S1(n1405), .Q(n1189) );
  IMUX40 U827 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n1437), .S1(n1408), .Q(n1194) );
  IMUX40 U828 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n1438), .S1(n1404), .Q(n1199) );
  IMUX40 U829 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n1438), .S1(n1409), .Q(n1204) );
  IMUX40 U830 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n1438), .S1(n1404), .Q(n1209) );
  IMUX40 U831 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n1439), .S1(n1412), .Q(n1214) );
  IMUX40 U832 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n1439), .S1(n1412), .Q(n1219) );
  IMUX40 U833 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n1439), .S1(n1413), .Q(n1224) );
  IMUX40 U834 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n1440), .S1(n1413), .Q(n1229) );
  IMUX40 U835 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n1440), .S1(n1414), .Q(n1234) );
  IMUX40 U836 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n1440), .S1(n1414), .Q(n1239) );
  IMUX40 U837 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n1441), .S1(n1414), .Q(n1244) );
  IMUX40 U838 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n1441), .S1(n1427), .Q(n1249) );
  IMUX40 U839 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n1441), .S1(n1427), .Q(n1254) );
  IMUX40 U840 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n1432), .S1(n1415), .Q(n1259) );
  IMUX40 U841 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n1433), .S1(n1415), .Q(n1264) );
  IMUX40 U842 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n1434), .S1(n1416), .Q(n1269) );
  IMUX40 U843 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n1430), .S1(n1416), .Q(n1274) );
  IMUX40 U844 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n1435), .S1(n1417), .Q(n1279) );
  IMUX40 U845 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n1436), .S1(n1417), .Q(n1284) );
  IMUX40 U846 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n1442), .S1(n1417), .Q(n1289) );
  IMUX40 U847 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n1442), .S1(n1418), .Q(n1294) );
  IMUX40 U848 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n1442), .S1(n1418), .Q(n1299) );
  IMUX40 U849 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n1443), .S1(n1419), .Q(n1304) );
  IMUX40 U850 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n1443), .S1(n1419), .Q(n1309) );
  IMUX40 U851 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n1443), .S1(n1420), .Q(n1314) );
  IMUX40 U852 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n1444), .S1(n1420), .Q(n1319) );
  IMUX40 U853 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n1444), .S1(n1421), .Q(n1324) );
  IMUX40 U854 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n1444), .S1(n1421), .Q(n1329) );
  IMUX40 U855 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n1445), .S1(n1421), .Q(n1334) );
  IMUX40 U856 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n1445), .S1(n1422), .Q(n1339) );
  IMUX40 U857 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n1445), .S1(n1422), .Q(n1344) );
  IMUX40 U858 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n1446), .S1(n1423), .Q(n1349) );
  IMUX40 U859 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n1446), .S1(n1423), .Q(n1354) );
  IMUX40 U860 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n1446), .S1(n1424), .Q(n1359) );
  IMUX40 U861 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n1447), .S1(n1424), .Q(n1364) );
  IMUX40 U862 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n1447), .S1(n1425), .Q(n1369) );
  IMUX40 U863 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n1447), .S1(n1425), .Q(n1374) );
  IMUX40 U864 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n1448), .S1(n1425), .Q(n1379) );
  IMUX40 U865 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n1448), .S1(n1426), .Q(n1384) );
  IMUX40 U866 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n1448), .S1(n1426), .Q(n1389) );
  NOR31 U867 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n1985), .Q(n1073) );
  NOR31 U868 ( .A(n1987), .B(i_addr_Rd[1]), .C(n1985), .Q(n1075) );
  NOR31 U869 ( .A(n1986), .B(i_addr_Rd[0]), .C(n1985), .Q(n1077) );
  NOR31 U870 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(n1987), .Q(n1067) );
  NOR31 U871 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[2]), .C(n1986), .Q(n1069) );
  NOR31 U872 ( .A(n1987), .B(i_addr_Rd[2]), .C(n1986), .Q(n1071) );
  NOR31 U873 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(i_addr_Rd[0]), .Q(n1064)
         );
  BUF2 U874 ( .A(i_addr_Rt[3]), .Q(n1394) );
  BUF2 U875 ( .A(i_addr_Rt[3]), .Q(n1395) );
  BUF2 U876 ( .A(i_addr_Rt[3]), .Q(n1396) );
  BUF2 U877 ( .A(i_addr_Rt[3]), .Q(n1397) );
  BUF2 U878 ( .A(i_addr_Rs[3]), .Q(n1775) );
  BUF2 U879 ( .A(i_addr_Rs[3]), .Q(n1776) );
  INV3 U880 ( .A(i_addr_Rd[0]), .Q(n1987) );
  INV3 U881 ( .A(i_addr_Rd[1]), .Q(n1986) );
  INV3 U882 ( .A(i_addr_Rd[2]), .Q(n1985) );
  BUF2 U883 ( .A(i_addr_Rs[4]), .Q(n1771) );
  BUF2 U884 ( .A(i_addr_Rt[2]), .Q(n1398) );
  BUF2 U885 ( .A(i_addr_Rt[2]), .Q(n1399) );
  BUF2 U886 ( .A(i_addr_Rt[2]), .Q(n1400) );
  BUF2 U887 ( .A(i_addr_Rt[2]), .Q(n1401) );
  BUF2 U888 ( .A(i_addr_Rt[2]), .Q(n1402) );
  BUF2 U889 ( .A(i_addr_Rt[2]), .Q(n1403) );
  BUF2 U890 ( .A(i_addr_Rs[2]), .Q(n1777) );
  BUF2 U891 ( .A(i_addr_Rs[2]), .Q(n1778) );
  BUF2 U892 ( .A(i_addr_Rs[2]), .Q(n1779) );
  BUF2 U893 ( .A(i_addr_Rs[2]), .Q(n1780) );
  INV3 U894 ( .A(i_addr_Rd[4]), .Q(n1967) );
  INV3 U895 ( .A(i_addr_Rd[3]), .Q(n1984) );
  BUF2 U896 ( .A(i_addr_Rt[3]), .Q(n1393) );
  BUF2 U897 ( .A(i_addr_Rs[3]), .Q(n1773) );
  BUF2 U898 ( .A(i_addr_Rt[1]), .Q(n1429) );
  BUF2 U899 ( .A(i_addr_Rt[1]), .Q(n1428) );
  BUF2 U900 ( .A(i_addr_Rt[1]), .Q(n1427) );
  MUX22 U901 ( .A(n1032), .B(n1027), .S(n1391), .Q(o_data_Rt[0]) );
  IMUX40 U902 ( .A(n1028), .B(n1029), .C(n1030), .D(n1031), .S0(n1393), .S1(
        i_addr_Rt[2]), .Q(n1027) );
  IMUX40 U903 ( .A(n1033), .B(n1034), .C(n1035), .D(n1036), .S0(n1393), .S1(
        n1398), .Q(n1032) );
  MUX22 U904 ( .A(n1042), .B(n1037), .S(n1391), .Q(o_data_Rt[1]) );
  IMUX40 U905 ( .A(n1043), .B(n1044), .C(n1045), .D(n1046), .S0(n1393), .S1(
        n1398), .Q(n1042) );
  IMUX40 U906 ( .A(n1038), .B(n1039), .C(n1040), .D(n1041), .S0(n1393), .S1(
        n1398), .Q(n1037) );
  IMUX40 U907 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n1430), .S1(i_addr_Rt[1]), .Q(n1043) );
  MUX22 U908 ( .A(n1052), .B(n1047), .S(n1391), .Q(o_data_Rt[2]) );
  IMUX40 U909 ( .A(n1053), .B(n1054), .C(n1055), .D(n1056), .S0(n1394), .S1(
        n1398), .Q(n1052) );
  IMUX40 U910 ( .A(n1048), .B(n1049), .C(n1050), .D(n1051), .S0(n1394), .S1(
        n1398), .Q(n1047) );
  IMUX40 U911 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n1431), .S1(i_addr_Rt[1]), .Q(n1053) );
  MUX22 U912 ( .A(n1062), .B(n1057), .S(n1391), .Q(o_data_Rt[3]) );
  IMUX40 U913 ( .A(n1107), .B(n1108), .C(n1109), .D(n1110), .S0(n1394), .S1(
        n1398), .Q(n1062) );
  IMUX40 U914 ( .A(n1058), .B(n1059), .C(n1060), .D(n1061), .S0(n1394), .S1(
        n1398), .Q(n1057) );
  IMUX40 U915 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n1432), .S1(i_addr_Rt[1]), .Q(n1107) );
  MUX22 U916 ( .A(n1116), .B(n1111), .S(n1391), .Q(o_data_Rt[4]) );
  IMUX40 U917 ( .A(n1117), .B(n1118), .C(n1119), .D(n1120), .S0(n1394), .S1(
        n1398), .Q(n1116) );
  IMUX40 U918 ( .A(n1112), .B(n1113), .C(n1114), .D(n1115), .S0(n1394), .S1(
        n1398), .Q(n1111) );
  IMUX40 U919 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n1432), .S1(n1427), .Q(n1117) );
  MUX22 U920 ( .A(n1126), .B(n1121), .S(n1391), .Q(o_data_Rt[5]) );
  IMUX40 U921 ( .A(n1127), .B(n1128), .C(n1129), .D(n1130), .S0(n1394), .S1(
        n1399), .Q(n1126) );
  IMUX40 U922 ( .A(n1122), .B(n1123), .C(n1124), .D(n1125), .S0(n1394), .S1(
        n1399), .Q(n1121) );
  IMUX40 U923 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n1433), .S1(n1427), .Q(n1127) );
  MUX22 U924 ( .A(n1136), .B(n1131), .S(n1392), .Q(o_data_Rt[6]) );
  IMUX40 U925 ( .A(n1137), .B(n1138), .C(n1139), .D(n1140), .S0(n1394), .S1(
        n1399), .Q(n1136) );
  IMUX40 U926 ( .A(n1132), .B(n1133), .C(n1134), .D(n1135), .S0(n1394), .S1(
        n1399), .Q(n1131) );
  IMUX40 U927 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n1434), .S1(n1409), .Q(n1137) );
  MUX22 U928 ( .A(n1146), .B(n1141), .S(n1392), .Q(o_data_Rt[7]) );
  IMUX40 U929 ( .A(n1147), .B(n1148), .C(n1149), .D(n1150), .S0(n1394), .S1(
        n1399), .Q(n1146) );
  IMUX40 U930 ( .A(n1142), .B(n1143), .C(n1144), .D(n1145), .S0(n1394), .S1(
        n1399), .Q(n1141) );
  IMUX40 U931 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n1434), .S1(n1427), .Q(n1147) );
  MUX22 U932 ( .A(n1156), .B(n1151), .S(n1392), .Q(o_data_Rt[8]) );
  IMUX40 U933 ( .A(n1157), .B(n1158), .C(n1159), .D(n1160), .S0(n1395), .S1(
        n1399), .Q(n1156) );
  IMUX40 U934 ( .A(n1152), .B(n1153), .C(n1154), .D(n1155), .S0(n1395), .S1(
        n1399), .Q(n1151) );
  IMUX40 U935 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n1435), .S1(n1407), .Q(n1157) );
  MUX22 U936 ( .A(n1166), .B(n1161), .S(n1392), .Q(o_data_Rt[9]) );
  IMUX40 U937 ( .A(n1167), .B(n1168), .C(n1169), .D(n1170), .S0(n1395), .S1(
        n1400), .Q(n1166) );
  IMUX40 U938 ( .A(n1162), .B(n1163), .C(n1164), .D(n1165), .S0(n1395), .S1(
        n1399), .Q(n1161) );
  IMUX40 U939 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n1436), .S1(n1410), .Q(n1167) );
  MUX22 U940 ( .A(n1176), .B(n1171), .S(n1392), .Q(o_data_Rt[10]) );
  IMUX40 U941 ( .A(n1177), .B(n1178), .C(n1179), .D(n1180), .S0(n1395), .S1(
        n1400), .Q(n1176) );
  IMUX40 U942 ( .A(n1172), .B(n1173), .C(n1174), .D(n1175), .S0(n1395), .S1(
        n1400), .Q(n1171) );
  IMUX40 U943 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n1436), .S1(n1411), .Q(n1177) );
  MUX22 U944 ( .A(n1186), .B(n1181), .S(n1392), .Q(o_data_Rt[11]) );
  IMUX40 U945 ( .A(n1187), .B(n1188), .C(n1189), .D(n1190), .S0(n1395), .S1(
        n1400), .Q(n1186) );
  IMUX40 U946 ( .A(n1182), .B(n1183), .C(n1184), .D(n1185), .S0(n1395), .S1(
        n1400), .Q(n1181) );
  IMUX40 U947 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n1437), .S1(i_addr_Rt[1]), .Q(n1187) );
  MUX22 U948 ( .A(n1196), .B(n1191), .S(n1392), .Q(o_data_Rt[12]) );
  IMUX40 U949 ( .A(n1197), .B(n1198), .C(n1199), .D(n1200), .S0(n1395), .S1(
        n1400), .Q(n1196) );
  IMUX40 U950 ( .A(n1192), .B(n1193), .C(n1194), .D(n1195), .S0(n1395), .S1(
        n1400), .Q(n1191) );
  IMUX40 U951 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n1438), .S1(n1404), .Q(n1197) );
  MUX22 U952 ( .A(n1206), .B(n1201), .S(n1392), .Q(o_data_Rt[13]) );
  IMUX40 U953 ( .A(n1207), .B(n1208), .C(n1209), .D(n1210), .S0(n1395), .S1(
        n1400), .Q(n1206) );
  IMUX40 U954 ( .A(n1202), .B(n1203), .C(n1204), .D(n1205), .S0(n1395), .S1(
        n1400), .Q(n1201) );
  IMUX40 U955 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n1438), .S1(n1428), .Q(n1207) );
  MUX22 U956 ( .A(n1216), .B(n1211), .S(n1392), .Q(o_data_Rt[14]) );
  IMUX40 U957 ( .A(n1217), .B(n1218), .C(n1219), .D(n1220), .S0(n1396), .S1(
        n1401), .Q(n1216) );
  IMUX40 U958 ( .A(n1212), .B(n1213), .C(n1214), .D(n1215), .S0(n1396), .S1(
        n1401), .Q(n1211) );
  IMUX40 U959 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n1439), .S1(n1412), .Q(n1217) );
  MUX22 U960 ( .A(n1226), .B(n1221), .S(n1392), .Q(o_data_Rt[15]) );
  IMUX40 U961 ( .A(n1227), .B(n1228), .C(n1229), .D(n1230), .S0(n1396), .S1(
        n1401), .Q(n1226) );
  IMUX40 U962 ( .A(n1222), .B(n1223), .C(n1224), .D(n1225), .S0(n1396), .S1(
        n1401), .Q(n1221) );
  IMUX40 U963 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n1440), .S1(n1413), .Q(n1227) );
  MUX22 U964 ( .A(n1236), .B(n1231), .S(n1392), .Q(o_data_Rt[16]) );
  IMUX40 U965 ( .A(n1237), .B(n1238), .C(n1239), .D(n1240), .S0(n1396), .S1(
        n1401), .Q(n1236) );
  IMUX40 U966 ( .A(n1232), .B(n1233), .C(n1234), .D(n1235), .S0(n1396), .S1(
        n1401), .Q(n1231) );
  IMUX40 U967 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n1440), .S1(n1414), .Q(n1237) );
  MUX22 U968 ( .A(n1246), .B(n1241), .S(n1392), .Q(o_data_Rt[17]) );
  IMUX40 U969 ( .A(n1247), .B(n1248), .C(n1249), .D(n1250), .S0(n1396), .S1(
        n1401), .Q(n1246) );
  IMUX40 U970 ( .A(n1242), .B(n1243), .C(n1244), .D(n1245), .S0(n1396), .S1(
        n1401), .Q(n1241) );
  IMUX40 U971 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n1441), .S1(n1414), .Q(n1247) );
  MUX22 U972 ( .A(n1256), .B(n1251), .S(n1392), .Q(o_data_Rt[18]) );
  IMUX40 U973 ( .A(n1257), .B(n1258), .C(n1259), .D(n1260), .S0(n1396), .S1(
        n1402), .Q(n1256) );
  IMUX40 U974 ( .A(n1252), .B(n1253), .C(n1254), .D(n1255), .S0(n1396), .S1(
        n1401), .Q(n1251) );
  IMUX40 U975 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n1434), .S1(n1415), .Q(n1257) );
  MUX22 U976 ( .A(n1266), .B(n1261), .S(n1391), .Q(o_data_Rt[19]) );
  IMUX40 U977 ( .A(n1267), .B(n1268), .C(n1269), .D(n1270), .S0(n1396), .S1(
        n1402), .Q(n1266) );
  IMUX40 U978 ( .A(n1262), .B(n1263), .C(n1264), .D(n1265), .S0(n1396), .S1(
        n1402), .Q(n1261) );
  IMUX40 U979 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n1442), .S1(n1416), .Q(n1267) );
  MUX22 U980 ( .A(n1276), .B(n1271), .S(n1391), .Q(o_data_Rt[20]) );
  IMUX40 U981 ( .A(n1277), .B(n1278), .C(n1279), .D(n1280), .S0(n1397), .S1(
        n1402), .Q(n1276) );
  IMUX40 U982 ( .A(n1272), .B(n1273), .C(n1274), .D(n1275), .S0(n1397), .S1(
        n1402), .Q(n1271) );
  IMUX40 U983 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n1437), .S1(n1417), .Q(n1277) );
  MUX22 U984 ( .A(n1286), .B(n1281), .S(n1391), .Q(o_data_Rt[21]) );
  IMUX40 U985 ( .A(n1287), .B(n1288), .C(n1289), .D(n1290), .S0(n1397), .S1(
        n1402), .Q(n1286) );
  IMUX40 U986 ( .A(n1282), .B(n1283), .C(n1284), .D(n1285), .S0(n1397), .S1(
        n1402), .Q(n1281) );
  IMUX40 U987 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n1442), .S1(n1418), .Q(n1287) );
  MUX22 U988 ( .A(n1296), .B(n1291), .S(n1391), .Q(o_data_Rt[22]) );
  IMUX40 U989 ( .A(n1297), .B(n1298), .C(n1299), .D(n1300), .S0(n1397), .S1(
        n1402), .Q(n1296) );
  IMUX40 U990 ( .A(n1292), .B(n1293), .C(n1294), .D(n1295), .S0(n1397), .S1(
        n1402), .Q(n1291) );
  IMUX40 U991 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n1442), .S1(n1418), .Q(n1297) );
  MUX22 U992 ( .A(n1306), .B(n1301), .S(n1391), .Q(o_data_Rt[23]) );
  IMUX40 U993 ( .A(n1307), .B(n1308), .C(n1309), .D(n1310), .S0(n1397), .S1(
        n1403), .Q(n1306) );
  IMUX40 U994 ( .A(n1302), .B(n1303), .C(n1304), .D(n1305), .S0(n1397), .S1(
        n1403), .Q(n1301) );
  IMUX40 U995 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n1443), .S1(n1419), .Q(n1307) );
  MUX22 U996 ( .A(n1316), .B(n1311), .S(n1391), .Q(o_data_Rt[24]) );
  IMUX40 U997 ( .A(n1317), .B(n1318), .C(n1319), .D(n1320), .S0(n1397), .S1(
        n1403), .Q(n1316) );
  IMUX40 U998 ( .A(n1312), .B(n1313), .C(n1314), .D(n1315), .S0(n1397), .S1(
        n1403), .Q(n1311) );
  IMUX40 U999 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n1444), .S1(n1420), .Q(n1317) );
  MUX22 U1000 ( .A(n1326), .B(n1321), .S(n1391), .Q(o_data_Rt[25]) );
  IMUX40 U1001 ( .A(n1327), .B(n1328), .C(n1329), .D(n1330), .S0(n1397), .S1(
        n1403), .Q(n1326) );
  IMUX40 U1002 ( .A(n1322), .B(n1323), .C(n1324), .D(n1325), .S0(n1397), .S1(
        n1403), .Q(n1321) );
  IMUX40 U1003 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n1444), .S1(n1421), .Q(n1327) );
  MUX22 U1004 ( .A(n1336), .B(n1331), .S(i_addr_Rt[4]), .Q(o_data_Rt[26]) );
  IMUX40 U1005 ( .A(n1337), .B(n1338), .C(n1339), .D(n1340), .S0(n1393), .S1(
        n1403), .Q(n1336) );
  IMUX40 U1006 ( .A(n1332), .B(n1333), .C(n1334), .D(n1335), .S0(n1393), .S1(
        n1403), .Q(n1331) );
  IMUX40 U1007 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n1445), .S1(n1422), .Q(n1337) );
  MUX22 U1008 ( .A(n1346), .B(n1341), .S(i_addr_Rt[4]), .Q(o_data_Rt[27]) );
  IMUX40 U1009 ( .A(n1347), .B(n1348), .C(n1349), .D(n1350), .S0(n1393), .S1(
        i_addr_Rt[2]), .Q(n1346) );
  IMUX40 U1010 ( .A(n1342), .B(n1343), .C(n1344), .D(n1345), .S0(n1393), .S1(
        n1403), .Q(n1341) );
  IMUX40 U1011 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n1446), .S1(n1423), .Q(n1347) );
  MUX22 U1012 ( .A(n1356), .B(n1351), .S(i_addr_Rt[4]), .Q(o_data_Rt[28]) );
  IMUX40 U1013 ( .A(n1357), .B(n1358), .C(n1359), .D(n1360), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n1356) );
  IMUX40 U1014 ( .A(n1352), .B(n1353), .C(n1354), .D(n1355), .S0(n1393), .S1(
        i_addr_Rt[2]), .Q(n1351) );
  IMUX40 U1015 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n1446), .S1(n1424), .Q(n1357) );
  MUX22 U1016 ( .A(n1366), .B(n1361), .S(i_addr_Rt[4]), .Q(o_data_Rt[29]) );
  IMUX40 U1017 ( .A(n1367), .B(n1368), .C(n1369), .D(n1370), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n1366) );
  IMUX40 U1018 ( .A(n1362), .B(n1363), .C(n1364), .D(n1365), .S0(n1393), .S1(
        i_addr_Rt[2]), .Q(n1361) );
  IMUX40 U1019 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n1447), .S1(n1425), .Q(n1367) );
  MUX22 U1020 ( .A(n1376), .B(n1371), .S(i_addr_Rt[4]), .Q(o_data_Rt[30]) );
  IMUX40 U1021 ( .A(n1377), .B(n1378), .C(n1379), .D(n1380), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n1376) );
  IMUX40 U1022 ( .A(n1372), .B(n1373), .C(n1374), .D(n1375), .S0(n1393), .S1(
        i_addr_Rt[2]), .Q(n1371) );
  IMUX40 U1023 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n1448), .S1(n1426), .Q(n1377) );
  MUX22 U1024 ( .A(n1386), .B(n1381), .S(i_addr_Rt[4]), .Q(o_data_Rt[31]) );
  IMUX40 U1025 ( .A(n1387), .B(n1388), .C(n1389), .D(n1390), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n1386) );
  IMUX40 U1026 ( .A(n1382), .B(n1383), .C(n1384), .D(n1385), .S0(n1393), .S1(
        i_addr_Rt[2]), .Q(n1381) );
  IMUX40 U1027 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n1448), .S1(n1426), .Q(n1387) );
  BUF2 U1028 ( .A(i_addr_Rt[4]), .Q(n1391) );
endmodule


module D_shiftleft ( i_data_immE, o_data_immshiftl );
  input [15:0] i_data_immE;
  output [31:0] o_data_immshiftl;
  wire   n_Logic0_, i_data_immE_15_, i_data_immE_14_, i_data_immE_13_,
         i_data_immE_12_, i_data_immE_11_, i_data_immE_10_, i_data_immE_9_,
         i_data_immE_8_, i_data_immE_7_, i_data_immE_6_, i_data_immE_5_,
         i_data_immE_4_, i_data_immE_3_, i_data_immE_2_, i_data_immE_1_,
         i_data_immE_0_, n1, o_data_immshiftl_23_, o_data_immshiftl_17_;
  assign o_data_immshiftl[0] = n_Logic0_;
  assign o_data_immshiftl[1] = n_Logic0_;
  assign o_data_immshiftl[25] = i_data_immE_15_;
  assign o_data_immshiftl[22] = i_data_immE_15_;
  assign o_data_immshiftl[18] = i_data_immE_15_;
  assign o_data_immshiftl[31] = i_data_immE_15_;
  assign i_data_immE_15_ = i_data_immE[15];
  assign o_data_immshiftl[16] = i_data_immE_14_;
  assign i_data_immE_14_ = i_data_immE[14];
  assign o_data_immshiftl[15] = i_data_immE_13_;
  assign i_data_immE_13_ = i_data_immE[13];
  assign o_data_immshiftl[14] = i_data_immE_12_;
  assign i_data_immE_12_ = i_data_immE[12];
  assign o_data_immshiftl[13] = i_data_immE_11_;
  assign i_data_immE_11_ = i_data_immE[11];
  assign o_data_immshiftl[12] = i_data_immE_10_;
  assign i_data_immE_10_ = i_data_immE[10];
  assign o_data_immshiftl[11] = i_data_immE_9_;
  assign i_data_immE_9_ = i_data_immE[9];
  assign o_data_immshiftl[10] = i_data_immE_8_;
  assign i_data_immE_8_ = i_data_immE[8];
  assign o_data_immshiftl[9] = i_data_immE_7_;
  assign i_data_immE_7_ = i_data_immE[7];
  assign o_data_immshiftl[8] = i_data_immE_6_;
  assign i_data_immE_6_ = i_data_immE[6];
  assign o_data_immshiftl[7] = i_data_immE_5_;
  assign i_data_immE_5_ = i_data_immE[5];
  assign o_data_immshiftl[6] = i_data_immE_4_;
  assign i_data_immE_4_ = i_data_immE[4];
  assign o_data_immshiftl[5] = i_data_immE_3_;
  assign i_data_immE_3_ = i_data_immE[3];
  assign o_data_immshiftl[4] = i_data_immE_2_;
  assign i_data_immE_2_ = i_data_immE[2];
  assign o_data_immshiftl[3] = i_data_immE_1_;
  assign i_data_immE_1_ = i_data_immE[1];
  assign o_data_immshiftl[2] = i_data_immE_0_;
  assign i_data_immE_0_ = i_data_immE[0];
  assign o_data_immshiftl[19] = o_data_immshiftl_23_;
  assign o_data_immshiftl[30] = o_data_immshiftl_23_;
  assign o_data_immshiftl[24] = o_data_immshiftl_23_;
  assign o_data_immshiftl[20] = o_data_immshiftl_23_;
  assign o_data_immshiftl[23] = o_data_immshiftl_23_;
  assign o_data_immshiftl[27] = o_data_immshiftl_17_;
  assign o_data_immshiftl[28] = o_data_immshiftl_17_;
  assign o_data_immshiftl[29] = o_data_immshiftl_17_;
  assign o_data_immshiftl[26] = o_data_immshiftl_17_;
  assign o_data_immshiftl[21] = o_data_immshiftl_17_;
  assign o_data_immshiftl[17] = o_data_immshiftl_17_;

  CLKIN3 U2 ( .A(i_data_immE_15_), .Q(n1) );
  INV3 U3 ( .A(n1), .Q(o_data_immshiftl_17_) );
  INV3 U4 ( .A(n1), .Q(o_data_immshiftl_23_) );
  LOGIC0 U5 ( .Q(n_Logic0_) );
endmodule


module D_sign_extend ( i_data_immD, i_con_signext, o_data_immD );
  input [15:0] i_data_immD;
  output [31:0] o_data_immD;
  input i_con_signext;
  wire   n3, o_data_immD_31_;
  assign o_data_immD[15] = i_data_immD[15];
  assign o_data_immD[14] = i_data_immD[14];
  assign o_data_immD[13] = i_data_immD[13];
  assign o_data_immD[12] = i_data_immD[12];
  assign o_data_immD[11] = i_data_immD[11];
  assign o_data_immD[10] = i_data_immD[10];
  assign o_data_immD[9] = i_data_immD[9];
  assign o_data_immD[8] = i_data_immD[8];
  assign o_data_immD[7] = i_data_immD[7];
  assign o_data_immD[6] = i_data_immD[6];
  assign o_data_immD[5] = i_data_immD[5];
  assign o_data_immD[4] = i_data_immD[4];
  assign o_data_immD[3] = i_data_immD[3];
  assign o_data_immD[2] = i_data_immD[2];
  assign o_data_immD[1] = i_data_immD[1];
  assign o_data_immD[0] = i_data_immD[0];
  assign o_data_immD[16] = o_data_immD_31_;
  assign o_data_immD[17] = o_data_immD_31_;
  assign o_data_immD[18] = o_data_immD_31_;
  assign o_data_immD[19] = o_data_immD_31_;
  assign o_data_immD[20] = o_data_immD_31_;
  assign o_data_immD[21] = o_data_immD_31_;
  assign o_data_immD[22] = o_data_immD_31_;
  assign o_data_immD[23] = o_data_immD_31_;
  assign o_data_immD[24] = o_data_immD_31_;
  assign o_data_immD[25] = o_data_immD_31_;
  assign o_data_immD[26] = o_data_immD_31_;
  assign o_data_immD[27] = o_data_immD_31_;
  assign o_data_immD[28] = o_data_immD_31_;
  assign o_data_immD[29] = o_data_immD_31_;
  assign o_data_immD[30] = o_data_immD_31_;
  assign o_data_immD[31] = o_data_immD_31_;

  NAND20 U2 ( .A(i_con_signext), .B(i_data_immD[15]), .Q(n3) );
  INV3 U3 ( .A(n3), .Q(o_data_immD_31_) );
endmodule


module D_jump_ext ( i_addr_j, i_PC4_j, o_addr_j );
  input [25:0] i_addr_j;
  input [3:0] i_PC4_j;
  output [31:0] o_addr_j;
  wire   n_Logic0_, i_PC4_j_3_, i_PC4_j_2_, i_PC4_j_1_, i_PC4_j_0_,
         i_addr_j_25_, i_addr_j_24_, i_addr_j_23_, i_addr_j_22_, i_addr_j_21_,
         i_addr_j_20_, i_addr_j_19_, i_addr_j_18_, i_addr_j_17_, i_addr_j_16_,
         i_addr_j_15_, i_addr_j_14_, i_addr_j_13_, i_addr_j_12_, i_addr_j_11_,
         i_addr_j_10_, i_addr_j_9_, i_addr_j_8_, i_addr_j_7_, i_addr_j_6_,
         i_addr_j_5_, i_addr_j_4_, i_addr_j_3_, i_addr_j_2_, i_addr_j_1_,
         i_addr_j_0_;
  assign o_addr_j[0] = n_Logic0_;
  assign o_addr_j[1] = n_Logic0_;
  assign o_addr_j[31] = i_PC4_j_3_;
  assign i_PC4_j_3_ = i_PC4_j[3];
  assign o_addr_j[30] = i_PC4_j_2_;
  assign i_PC4_j_2_ = i_PC4_j[2];
  assign o_addr_j[29] = i_PC4_j_1_;
  assign i_PC4_j_1_ = i_PC4_j[1];
  assign o_addr_j[28] = i_PC4_j_0_;
  assign i_PC4_j_0_ = i_PC4_j[0];
  assign o_addr_j[27] = i_addr_j_25_;
  assign i_addr_j_25_ = i_addr_j[25];
  assign o_addr_j[26] = i_addr_j_24_;
  assign i_addr_j_24_ = i_addr_j[24];
  assign o_addr_j[25] = i_addr_j_23_;
  assign i_addr_j_23_ = i_addr_j[23];
  assign o_addr_j[24] = i_addr_j_22_;
  assign i_addr_j_22_ = i_addr_j[22];
  assign o_addr_j[23] = i_addr_j_21_;
  assign i_addr_j_21_ = i_addr_j[21];
  assign o_addr_j[22] = i_addr_j_20_;
  assign i_addr_j_20_ = i_addr_j[20];
  assign o_addr_j[21] = i_addr_j_19_;
  assign i_addr_j_19_ = i_addr_j[19];
  assign o_addr_j[20] = i_addr_j_18_;
  assign i_addr_j_18_ = i_addr_j[18];
  assign o_addr_j[19] = i_addr_j_17_;
  assign i_addr_j_17_ = i_addr_j[17];
  assign o_addr_j[18] = i_addr_j_16_;
  assign i_addr_j_16_ = i_addr_j[16];
  assign o_addr_j[17] = i_addr_j_15_;
  assign i_addr_j_15_ = i_addr_j[15];
  assign o_addr_j[16] = i_addr_j_14_;
  assign i_addr_j_14_ = i_addr_j[14];
  assign o_addr_j[15] = i_addr_j_13_;
  assign i_addr_j_13_ = i_addr_j[13];
  assign o_addr_j[14] = i_addr_j_12_;
  assign i_addr_j_12_ = i_addr_j[12];
  assign o_addr_j[13] = i_addr_j_11_;
  assign i_addr_j_11_ = i_addr_j[11];
  assign o_addr_j[12] = i_addr_j_10_;
  assign i_addr_j_10_ = i_addr_j[10];
  assign o_addr_j[11] = i_addr_j_9_;
  assign i_addr_j_9_ = i_addr_j[9];
  assign o_addr_j[10] = i_addr_j_8_;
  assign i_addr_j_8_ = i_addr_j[8];
  assign o_addr_j[9] = i_addr_j_7_;
  assign i_addr_j_7_ = i_addr_j[7];
  assign o_addr_j[8] = i_addr_j_6_;
  assign i_addr_j_6_ = i_addr_j[6];
  assign o_addr_j[7] = i_addr_j_5_;
  assign i_addr_j_5_ = i_addr_j[5];
  assign o_addr_j[6] = i_addr_j_4_;
  assign i_addr_j_4_ = i_addr_j[4];
  assign o_addr_j[5] = i_addr_j_3_;
  assign i_addr_j_3_ = i_addr_j[3];
  assign o_addr_j[4] = i_addr_j_2_;
  assign i_addr_j_2_ = i_addr_j[2];
  assign o_addr_j[3] = i_addr_j_1_;
  assign i_addr_j_1_ = i_addr_j[1];
  assign o_addr_j[2] = i_addr_j_0_;
  assign i_addr_j_0_ = i_addr_j[0];

  LOGIC0 U2 ( .Q(n_Logic0_) );
endmodule


module E_forward ( i_addr_rs, i_addr_rt, i_addr_rdM, i_addr_rdW, i_addr_rtM, 
        i_addr_rtW, i_con_regwriteM, i_con_regwriteW, i_con_memreadM, 
        i_con_memreadW, o_con_fa, o_con_fb, o_con_cmpalu, o_con_cmpmem );
  input [4:0] i_addr_rs;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rdM;
  input [4:0] i_addr_rdW;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  output [2:0] o_con_fa;
  output [2:0] o_con_fb;
  input i_con_regwriteM, i_con_regwriteW, i_con_memreadM, i_con_memreadW;
  output o_con_cmpalu, o_con_cmpmem;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87;

  INV3 U1 ( .A(n1), .Q(n19) );
  OAI212 U2 ( .A(o_con_cmpmem), .B(n50), .C(n51), .Q(o_con_fa[0]) );
  NOR31 U3 ( .A(i_addr_rs[0]), .B(i_addr_rs[1]), .C(n86), .Q(n72) );
  NOR31 U4 ( .A(i_addr_rs[2]), .B(i_addr_rs[4]), .C(i_addr_rs[3]), .Q(n87) );
  NAND41 U5 ( .A(n23), .B(n24), .C(n25), .D(n26), .Q(n1) );
  NOR31 U6 ( .A(i_addr_rt[2]), .B(i_addr_rt[4]), .C(i_addr_rt[3]), .Q(n47) );
  NOR31 U7 ( .A(i_addr_rt[0]), .B(i_addr_rt[1]), .C(n46), .Q(n13) );
  NAND22 U8 ( .A(n61), .B(n50), .Q(o_con_fa[2]) );
  NAND41 U9 ( .A(n68), .B(n69), .C(n70), .D(n71), .Q(n50) );
  NAND41 U10 ( .A(n75), .B(n76), .C(n77), .D(n78), .Q(n61) );
  INV2 U11 ( .A(n87), .Q(n86) );
  INV3 U12 ( .A(n47), .Q(n46) );
  NOR20 U13 ( .A(o_con_fb[2]), .B(n1), .Q(o_con_fb[1]) );
  NAND20 U14 ( .A(n2), .B(n3), .Q(o_con_fb[2]) );
  NOR20 U15 ( .A(n4), .B(n5), .Q(o_con_fb[0]) );
  AOI210 U16 ( .A(n6), .B(n7), .C(n8), .Q(n5) );
  CLKIN0 U17 ( .A(n3), .Q(n8) );
  NAND40 U18 ( .A(n9), .B(n10), .C(n11), .D(n12), .Q(n3) );
  NOR40 U19 ( .A(n13), .B(n14), .C(n15), .D(n16), .Q(n12) );
  XNR20 U20 ( .A(n17), .B(i_addr_rt[1]), .Q(n16) );
  XNR20 U21 ( .A(n18), .B(i_addr_rt[0]), .Q(n15) );
  XNR20 U22 ( .A(i_addr_rt[3]), .B(i_addr_rtW[3]), .Q(n11) );
  XNR20 U23 ( .A(i_addr_rt[4]), .B(i_addr_rtW[4]), .Q(n10) );
  XNR20 U24 ( .A(i_addr_rt[2]), .B(i_addr_rtW[2]), .Q(n9) );
  NOR40 U25 ( .A(n13), .B(n19), .C(n20), .D(n21), .Q(n7) );
  XNR20 U26 ( .A(n22), .B(i_addr_rt[0]), .Q(n21) );
  NOR40 U27 ( .A(n13), .B(n27), .C(n28), .D(n29), .Q(n26) );
  XOR20 U28 ( .A(i_addr_rdM[1]), .B(i_addr_rt[1]), .Q(n29) );
  XOR20 U29 ( .A(i_addr_rdM[0]), .B(i_addr_rt[0]), .Q(n28) );
  XNR20 U30 ( .A(i_addr_rt[3]), .B(i_addr_rdM[3]), .Q(n25) );
  XNR20 U31 ( .A(i_addr_rt[4]), .B(i_addr_rdM[4]), .Q(n24) );
  XNR20 U32 ( .A(i_addr_rt[2]), .B(i_addr_rdM[2]), .Q(n23) );
  NOR40 U33 ( .A(n30), .B(n31), .C(n32), .D(n33), .Q(n6) );
  XOR20 U34 ( .A(i_addr_rdW[4]), .B(i_addr_rt[4]), .Q(n33) );
  XNR20 U35 ( .A(n34), .B(i_addr_rt[3]), .Q(n32) );
  XNR20 U36 ( .A(n35), .B(i_addr_rt[2]), .Q(n31) );
  XNR20 U37 ( .A(n36), .B(i_addr_rt[1]), .Q(n30) );
  CLKIN0 U38 ( .A(n2), .Q(n4) );
  NAND40 U39 ( .A(n37), .B(n38), .C(n39), .D(n40), .Q(n2) );
  NOR40 U40 ( .A(n13), .B(n41), .C(n42), .D(n43), .Q(n40) );
  XNR20 U41 ( .A(n44), .B(i_addr_rt[1]), .Q(n43) );
  XNR20 U42 ( .A(n45), .B(i_addr_rt[0]), .Q(n42) );
  XNR20 U43 ( .A(i_addr_rt[3]), .B(i_addr_rtM[3]), .Q(n39) );
  XNR20 U44 ( .A(i_addr_rt[4]), .B(i_addr_rtM[4]), .Q(n38) );
  XNR20 U45 ( .A(i_addr_rt[2]), .B(i_addr_rtM[2]), .Q(n37) );
  NOR20 U46 ( .A(o_con_fa[2]), .B(n48), .Q(o_con_fa[1]) );
  CLKIN0 U47 ( .A(n49), .Q(n48) );
  NAND20 U48 ( .A(n52), .B(n53), .Q(n51) );
  NOR40 U49 ( .A(o_con_fa[2]), .B(n49), .C(n20), .D(n54), .Q(n53) );
  XNR20 U50 ( .A(n22), .B(i_addr_rs[0]), .Q(n54) );
  CLKIN0 U51 ( .A(i_addr_rdW[0]), .Q(n22) );
  CLKIN0 U52 ( .A(i_con_regwriteW), .Q(n20) );
  NOR40 U53 ( .A(n55), .B(n56), .C(n57), .D(n58), .Q(n49) );
  OAI310 U54 ( .A(i_addr_rdM[0]), .B(i_addr_rdM[1]), .C(n59), .D(
        i_con_regwriteM), .Q(n57) );
  CLKIN0 U55 ( .A(n60), .Q(n59) );
  NOR30 U56 ( .A(i_addr_rdM[2]), .B(i_addr_rdM[4]), .C(i_addr_rdM[3]), .Q(n60)
         );
  NOR40 U57 ( .A(n62), .B(n63), .C(n64), .D(n65), .Q(n52) );
  IMUX20 U58 ( .A(n66), .B(i_addr_rs[4]), .S(i_addr_rdW[4]), .Q(n65) );
  NOR20 U59 ( .A(n67), .B(i_addr_rs[4]), .Q(n66) );
  NOR40 U60 ( .A(i_addr_rdW[3]), .B(i_addr_rdW[2]), .C(i_addr_rdW[1]), .D(
        i_addr_rdW[0]), .Q(n67) );
  XNR20 U61 ( .A(n34), .B(i_addr_rs[3]), .Q(n64) );
  CLKIN0 U62 ( .A(i_addr_rdW[3]), .Q(n34) );
  XNR20 U63 ( .A(n35), .B(i_addr_rs[2]), .Q(n63) );
  CLKIN0 U64 ( .A(i_addr_rdW[2]), .Q(n35) );
  XNR20 U65 ( .A(n36), .B(i_addr_rs[1]), .Q(n62) );
  CLKIN0 U66 ( .A(i_addr_rdW[1]), .Q(n36) );
  NOR40 U67 ( .A(n72), .B(n14), .C(n73), .D(n74), .Q(n71) );
  XNR20 U68 ( .A(n17), .B(i_addr_rs[1]), .Q(n74) );
  CLKIN0 U69 ( .A(i_addr_rtW[1]), .Q(n17) );
  XNR20 U70 ( .A(n18), .B(i_addr_rs[0]), .Q(n73) );
  CLKIN0 U71 ( .A(i_addr_rtW[0]), .Q(n18) );
  CLKIN0 U72 ( .A(i_con_memreadW), .Q(n14) );
  XNR20 U73 ( .A(i_addr_rtW[3]), .B(i_addr_rs[3]), .Q(n70) );
  XNR20 U74 ( .A(i_addr_rtW[4]), .B(i_addr_rs[4]), .Q(n69) );
  XNR20 U75 ( .A(i_addr_rtW[2]), .B(i_addr_rs[2]), .Q(n68) );
  CLKIN0 U76 ( .A(n61), .Q(o_con_cmpmem) );
  NOR40 U77 ( .A(n72), .B(n41), .C(n79), .D(n80), .Q(n78) );
  XNR20 U78 ( .A(n44), .B(i_addr_rs[1]), .Q(n80) );
  CLKIN0 U79 ( .A(i_addr_rtM[1]), .Q(n44) );
  XNR20 U80 ( .A(n45), .B(i_addr_rs[0]), .Q(n79) );
  CLKIN0 U81 ( .A(i_addr_rtM[0]), .Q(n45) );
  CLKIN0 U82 ( .A(i_con_memreadM), .Q(n41) );
  XNR20 U83 ( .A(i_addr_rtM[3]), .B(i_addr_rs[3]), .Q(n77) );
  XNR20 U84 ( .A(i_addr_rtM[4]), .B(i_addr_rs[4]), .Q(n76) );
  XNR20 U85 ( .A(i_addr_rtM[2]), .B(i_addr_rs[2]), .Q(n75) );
  NOR40 U86 ( .A(n58), .B(n81), .C(n56), .D(n55), .Q(o_con_cmpalu) );
  XOR20 U87 ( .A(i_addr_rs[4]), .B(i_addr_rdM[4]), .Q(n55) );
  NAND30 U88 ( .A(n82), .B(n83), .C(n84), .Q(n56) );
  XNR20 U89 ( .A(i_addr_rs[1]), .B(i_addr_rdM[1]), .Q(n84) );
  XNR20 U90 ( .A(i_addr_rs[2]), .B(i_addr_rdM[2]), .Q(n83) );
  XNR20 U91 ( .A(i_addr_rs[0]), .B(i_addr_rdM[0]), .Q(n82) );
  CLKIN0 U92 ( .A(n85), .Q(n81) );
  NOR20 U93 ( .A(n27), .B(n72), .Q(n85) );
  CLKIN0 U94 ( .A(i_con_regwriteM), .Q(n27) );
  XOR20 U95 ( .A(i_addr_rs[3]), .B(i_addr_rdM[3]), .Q(n58) );
endmodule


module decode ( i_clk, i_nrst, i_addr_pc4, i_data_instr, i_con_Wregwrite, 
        i_data_Wregwrite, i_addr_Wregwrite, i_addr_Erd, i_addr_Mrd, 
        i_con_Eregwrite, i_con_Mregwrite, i_addr_rtM, i_addr_rtW, 
        i_con_memreadM, i_con_memreadW, i_data_aluresE, i_data_memoutM, 
        o_data_rs, o_data_rt, o_addr_rd, o_addr_rt, o_data_jr, o_con_jump, 
        o_addr_pc4, o_addr_branch, o_addr_jump, o_con_Ealuop, o_con_Ealusrc, 
        o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite, o_con_Wloadmux, 
        o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall, 
        o_con_Ebop, o_data_signext, o_con_Efamux, o_con_Efbmux, o_data_Fmemout
 );
  input [31:0] i_addr_pc4;
  input [31:0] i_data_instr;
  input [31:0] i_data_Wregwrite;
  input [4:0] i_addr_Wregwrite;
  input [4:0] i_addr_Erd;
  input [4:0] i_addr_Mrd;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  input [31:0] i_data_aluresE;
  input [31:0] i_data_memoutM;
  output [31:0] o_data_rs;
  output [31:0] o_data_rt;
  output [4:0] o_addr_rd;
  output [4:0] o_addr_rt;
  output [31:0] o_data_jr;
  output [1:0] o_con_jump;
  output [31:0] o_addr_pc4;
  output [31:0] o_addr_branch;
  output [31:0] o_addr_jump;
  output [5:0] o_con_Ealuop;
  output [1:0] o_con_Wloadmux;
  output [2:0] o_con_Ebop;
  output [31:0] o_data_signext;
  output [2:0] o_con_Efamux;
  output [2:0] o_con_Efbmux;
  output [31:0] o_data_Fmemout;
  input i_clk, i_nrst, i_con_Wregwrite, i_con_Eregwrite, i_con_Mregwrite,
         i_con_memreadM, i_con_memreadW;
  output o_con_Ealusrc, o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite,
         o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall;
  wire   control_o_con_alusrc, control_o_con_regdst, jbcon_o_con_aluPC4,
         control_o_con_regwrite, signext_i_con_signext, o_con_Wmemtoreg, n122,
         n123;
  wire   [31:0] regbank_o_data_Rt;
  wire   [5:0] control_o_con_aluop;
  wire   [31:0] signext_o_data_immD;
  wire   [2:0] for_o_con_fa;
  wire   [2:0] for_o_con_fb;
  wire   [31:0] pcadd_o_addr_pcbranchE;
  wire   [2:0] jbcon_o_con_bop;
  wire   [31:2] pcadd_i_data_immshiftl;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign o_addr_jump[1] = o_con_Wmemtoreg;
  assign o_addr_jump[0] = o_con_Wmemtoreg;
  assign o_con_Mmemread = o_con_Wmemtoreg;
  assign o_con_Mmemwrite = o_con_Wmemtoreg;
  assign o_con_Wloadmux[1] = o_con_Wmemtoreg;
  assign o_con_Wloadmux[0] = o_con_Wmemtoreg;

  DFC3 pipe_bop_reg_2_ ( .D(jbcon_o_con_bop[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[2]) );
  DFC3 pipe_bop_reg_1_ ( .D(jbcon_o_con_bop[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[1]) );
  DFC3 pipe_bop_reg_0_ ( .D(jbcon_o_con_bop[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[0]) );
  DFC3 pipe_addr_rd_reg_3_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[3]) );
  DFC3 pipe_addr_rd_reg_2_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[2]) );
  DFC3 pipe_addr_rd_reg_1_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[1]) );
  DFC3 pipe_addr_rd_reg_0_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[0]) );
  DFC3 pipe_addr_rt_reg_4_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(n122), .C(i_clk), .RN(i_nrst), .Q(o_addr_rt[0]) );
  DFC3 pipe_addr_pc4_reg_31_ ( .D(i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_addr_pc4_reg_30_ ( .D(i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_addr_pc4_reg_29_ ( .D(i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_addr_pc4_reg_28_ ( .D(i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_addr_pc4_reg_27_ ( .D(i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_addr_pc4_reg_26_ ( .D(i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_addr_pc4_reg_25_ ( .D(i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_addr_pc4_reg_24_ ( .D(i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_addr_pc4_reg_23_ ( .D(i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_addr_pc4_reg_22_ ( .D(i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_addr_pc4_reg_21_ ( .D(i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_addr_pc4_reg_20_ ( .D(i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_addr_pc4_reg_19_ ( .D(i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_addr_pc4_reg_18_ ( .D(i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_addr_pc4_reg_17_ ( .D(i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_addr_pc4_reg_16_ ( .D(i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_addr_pc4_reg_15_ ( .D(i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_addr_pc4_reg_14_ ( .D(i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_addr_pc4_reg_13_ ( .D(i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_addr_pc4_reg_11_ ( .D(i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_addr_pc4_reg_10_ ( .D(i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_addr_pc4_reg_9_ ( .D(i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_addr_pc4_reg_8_ ( .D(i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_addr_pc4_reg_7_ ( .D(i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_addr_pc4_reg_4_ ( .D(i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_addr_pc4_reg_2_ ( .D(i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_addr_pc4_reg_1_ ( .D(i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_addr_pc4_reg_0_ ( .D(i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  DFC3 pipe_con_Ealuop_reg_5_ ( .D(control_o_con_aluop[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[5]) );
  DFC3 pipe_con_Ealuop_reg_4_ ( .D(control_o_con_aluop[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[4]) );
  DFC3 pipe_con_Ealuop_reg_3_ ( .D(control_o_con_aluop[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[3]) );
  DFC3 pipe_con_Ealuop_reg_2_ ( .D(control_o_con_aluop[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[2]) );
  DFC3 pipe_con_Ealuop_reg_1_ ( .D(control_o_con_aluop[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[1]) );
  DFC3 pipe_con_Ealuop_reg_0_ ( .D(control_o_con_aluop[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[0]) );
  DFC3 pipe_con_Ealusrc_reg ( .D(control_o_con_alusrc), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Ealusrc) );
  DFC3 pipe_con_Eregdst_reg ( .D(control_o_con_regdst), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Eregdst) );
  DFC3 pipe_con_EaluPC4_reg ( .D(jbcon_o_con_aluPC4), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Walupc8) );
  DFC3 pipe_con_Wregwrite_reg ( .D(control_o_con_regwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wregwrite) );
  DFC3 pipe_signext_o_data_immD_reg_31_ ( .D(signext_o_data_immD[31]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[31]) );
  DFC3 pipe_signext_o_data_immD_reg_30_ ( .D(signext_o_data_immD[30]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[30]) );
  DFC3 pipe_signext_o_data_immD_reg_29_ ( .D(signext_o_data_immD[29]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[29]) );
  DFC3 pipe_signext_o_data_immD_reg_28_ ( .D(signext_o_data_immD[28]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[28]) );
  DFC3 pipe_signext_o_data_immD_reg_27_ ( .D(signext_o_data_immD[27]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[27]) );
  DFC3 pipe_signext_o_data_immD_reg_26_ ( .D(signext_o_data_immD[26]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[26]) );
  DFC3 pipe_signext_o_data_immD_reg_25_ ( .D(signext_o_data_immD[25]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[25]) );
  DFC3 pipe_signext_o_data_immD_reg_24_ ( .D(signext_o_data_immD[24]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[24]) );
  DFC3 pipe_signext_o_data_immD_reg_23_ ( .D(signext_o_data_immD[23]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[23]) );
  DFC3 pipe_signext_o_data_immD_reg_22_ ( .D(signext_o_data_immD[22]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[22]) );
  DFC3 pipe_signext_o_data_immD_reg_21_ ( .D(signext_o_data_immD[21]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[21]) );
  DFC3 pipe_signext_o_data_immD_reg_20_ ( .D(signext_o_data_immD[20]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[20]) );
  DFC3 pipe_signext_o_data_immD_reg_19_ ( .D(signext_o_data_immD[19]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[19]) );
  DFC3 pipe_signext_o_data_immD_reg_18_ ( .D(signext_o_data_immD[18]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[18]) );
  DFC3 pipe_signext_o_data_immD_reg_17_ ( .D(signext_o_data_immD[17]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[17]) );
  DFC3 pipe_signext_o_data_immD_reg_16_ ( .D(signext_o_data_immD[16]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[16]) );
  DFC3 pipe_signext_o_data_immD_reg_14_ ( .D(signext_o_data_immD[14]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[14]) );
  DFC3 pipe_signext_o_data_immD_reg_13_ ( .D(signext_o_data_immD[13]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[13]) );
  DFC3 pipe_signext_o_data_immD_reg_12_ ( .D(signext_o_data_immD[12]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[12]) );
  DFC3 pipe_signext_o_data_immD_reg_11_ ( .D(signext_o_data_immD[11]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[11]) );
  DFC3 pipe_signext_o_data_immD_reg_10_ ( .D(signext_o_data_immD[10]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[10]) );
  DFC3 pipe_signext_o_data_immD_reg_9_ ( .D(signext_o_data_immD[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[9]) );
  DFC3 pipe_signext_o_data_immD_reg_8_ ( .D(signext_o_data_immD[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[8]) );
  DFC3 pipe_signext_o_data_immD_reg_7_ ( .D(signext_o_data_immD[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[7]) );
  DFC3 pipe_signext_o_data_immD_reg_6_ ( .D(signext_o_data_immD[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[6]) );
  DFC3 pipe_signext_o_data_immD_reg_5_ ( .D(signext_o_data_immD[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[5]) );
  DFC3 pipe_signext_o_data_immD_reg_4_ ( .D(signext_o_data_immD[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[4]) );
  DFC3 pipe_signext_o_data_immD_reg_3_ ( .D(signext_o_data_immD[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[3]) );
  DFC3 pipe_signext_o_data_immD_reg_2_ ( .D(signext_o_data_immD[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[2]) );
  DFC3 pipe_signext_o_data_immD_reg_1_ ( .D(signext_o_data_immD[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[1]) );
  DFC3 pipe_signext_o_data_immD_reg_0_ ( .D(signext_o_data_immD[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[0]) );
  DFC3 pipe_con_Efamux_reg_2_ ( .D(for_o_con_fa[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[2]) );
  DFC3 pipe_con_Efamux_reg_1_ ( .D(for_o_con_fa[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[1]) );
  DFC3 pipe_con_Efbmux_reg_2_ ( .D(for_o_con_fb[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[2]) );
  DFC3 pipe_con_Efbmux_reg_1_ ( .D(for_o_con_fb[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[1]) );
  DFC3 pipe_addr_branch_reg_31_ ( .D(pcadd_o_addr_pcbranchE[31]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[31]) );
  DFC3 pipe_addr_branch_reg_27_ ( .D(pcadd_o_addr_pcbranchE[27]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[27]) );
  DFC3 pipe_addr_branch_reg_23_ ( .D(pcadd_o_addr_pcbranchE[23]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[23]) );
  DFC3 pipe_addr_branch_reg_19_ ( .D(pcadd_o_addr_pcbranchE[19]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[19]) );
  DFC3 pipe_addr_branch_reg_16_ ( .D(pcadd_o_addr_pcbranchE[16]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[16]) );
  DFC3 pipe_addr_branch_reg_13_ ( .D(pcadd_o_addr_pcbranchE[13]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[13]) );
  DFC3 pipe_addr_branch_reg_12_ ( .D(pcadd_o_addr_pcbranchE[12]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[12]) );
  DFC3 pipe_addr_branch_reg_9_ ( .D(pcadd_o_addr_pcbranchE[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[9]) );
  DFC3 pipe_addr_branch_reg_8_ ( .D(pcadd_o_addr_pcbranchE[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[8]) );
  DFC3 pipe_addr_branch_reg_5_ ( .D(pcadd_o_addr_pcbranchE[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[5]) );
  DFC3 pipe_addr_branch_reg_4_ ( .D(pcadd_o_addr_pcbranchE[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[4]) );
  DFC3 pipe_addr_branch_reg_3_ ( .D(pcadd_o_addr_pcbranchE[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[3]) );
  DFC3 pipe_addr_branch_reg_2_ ( .D(pcadd_o_addr_pcbranchE[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[2]) );
  DFC3 pipe_addr_branch_reg_1_ ( .D(pcadd_o_addr_pcbranchE[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[1]) );
  DFC3 pipe_addr_branch_reg_0_ ( .D(pcadd_o_addr_pcbranchE[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[0]) );
  D_control u_control ( .o_con_regdst(control_o_con_regdst), .o_con_alusrc(
        control_o_con_alusrc), .o_con_regwrite(control_o_con_regwrite), 
        .o_con_ifsign(signext_i_con_signext), .o_con_aluop(control_o_con_aluop), .i_con_instru(i_data_instr[31:26]) );
  D_jb_control u_jb_control ( .o_con_jump(o_con_jump), .o_con_bop(
        jbcon_o_con_bop), .o_con_aluPC4(jbcon_o_con_aluPC4), .o_con_ifstall(
        o_con_ifstall), .i_con_instru(i_data_instr[31:26]), .i_con_func(
        i_data_instr[5:0]), .i_con_rt(o_con_Wmemtoreg) );
  D_pcadd u_pcadd ( .i_addr_pcadd4E(i_addr_pc4), .i_data_immshiftl({
        pcadd_i_data_immshiftl, o_con_Wmemtoreg, o_con_Wmemtoreg}), 
        .o_addr_pcbranchE(pcadd_o_addr_pcbranchE) );
  D_register_bank u_regbank ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_addr_Rs({
        i_data_instr[25:22], n123}), .i_addr_Rt({i_data_instr[20:17], n122}), 
        .i_con_RegWr(i_con_Wregwrite), .i_addr_Rd(i_addr_Wregwrite), 
        .i_data_Rd(i_data_Wregwrite), .o_data_Rs(o_data_jr), .o_data_Rt(
        regbank_o_data_Rt) );
  D_shiftleft u_sl ( .i_data_immE(i_data_instr[15:0]), .o_data_immshiftl({
        pcadd_i_data_immshiftl, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}) );
  D_sign_extend u_signext ( .i_data_immD(i_data_instr[15:0]), .i_con_signext(
        signext_i_con_signext), .o_data_immD(signext_o_data_immD) );
  D_jump_ext u_jump_ext ( .i_addr_j({i_data_instr[25:22], n123, 
        i_data_instr[20:17], n122, i_data_instr[15:0]}), .i_PC4_j(
        i_addr_pc4[31:28]), .o_addr_j({o_addr_jump[31:2], 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3}) );
  E_forward u_forward ( .i_addr_rs({i_data_instr[25:22], n123}), .i_addr_rt({
        i_data_instr[20:17], n122}), .i_addr_rdM(i_addr_Erd), .i_addr_rdW(
        i_addr_Mrd), .i_addr_rtM(i_addr_rtM), .i_addr_rtW(i_addr_rtW), 
        .i_con_regwriteM(i_con_Eregwrite), .i_con_regwriteW(i_con_Mregwrite), 
        .i_con_memreadM(i_con_memreadM), .i_con_memreadW(i_con_memreadW), 
        .o_con_fa(for_o_con_fa), .o_con_fb(for_o_con_fb) );
  DFC1 pipe_data_rs_reg_31_ ( .D(o_data_jr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[31]) );
  DFC1 pipe_data_rs_reg_30_ ( .D(o_data_jr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[30]) );
  DFC1 pipe_data_rs_reg_29_ ( .D(o_data_jr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[29]) );
  DFC1 pipe_data_rs_reg_28_ ( .D(o_data_jr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[28]) );
  DFC1 pipe_data_rs_reg_27_ ( .D(o_data_jr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[27]) );
  DFC1 pipe_data_rs_reg_26_ ( .D(o_data_jr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[26]) );
  DFC1 pipe_data_rs_reg_25_ ( .D(o_data_jr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[25]) );
  DFC1 pipe_data_rs_reg_24_ ( .D(o_data_jr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[24]) );
  DFC1 pipe_data_rs_reg_23_ ( .D(o_data_jr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[23]) );
  DFC1 pipe_data_rs_reg_22_ ( .D(o_data_jr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[22]) );
  DFC1 pipe_data_rs_reg_21_ ( .D(o_data_jr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[21]) );
  DFC1 pipe_data_rs_reg_20_ ( .D(o_data_jr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[20]) );
  DFC1 pipe_data_rs_reg_19_ ( .D(o_data_jr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[19]) );
  DFC1 pipe_data_rs_reg_18_ ( .D(o_data_jr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[18]) );
  DFC1 pipe_data_rs_reg_17_ ( .D(o_data_jr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[17]) );
  DFC1 pipe_data_rs_reg_16_ ( .D(o_data_jr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[16]) );
  DFC1 pipe_data_rs_reg_15_ ( .D(o_data_jr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[15]) );
  DFC1 pipe_data_rs_reg_14_ ( .D(o_data_jr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[14]) );
  DFC1 pipe_data_rs_reg_13_ ( .D(o_data_jr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[13]) );
  DFC1 pipe_data_rs_reg_12_ ( .D(o_data_jr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[12]) );
  DFC1 pipe_data_rs_reg_11_ ( .D(o_data_jr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[11]) );
  DFC1 pipe_data_rs_reg_10_ ( .D(o_data_jr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[10]) );
  DFC1 pipe_data_rs_reg_9_ ( .D(o_data_jr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[9]) );
  DFC1 pipe_data_rs_reg_8_ ( .D(o_data_jr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[8]) );
  DFC1 pipe_data_rs_reg_7_ ( .D(o_data_jr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[7]) );
  DFC1 pipe_data_rs_reg_6_ ( .D(o_data_jr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[6]) );
  DFC1 pipe_data_rs_reg_5_ ( .D(o_data_jr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[5]) );
  DFC1 pipe_data_rs_reg_4_ ( .D(o_data_jr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[4]) );
  DFC1 pipe_data_rs_reg_3_ ( .D(o_data_jr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[3]) );
  DFC1 pipe_data_rs_reg_2_ ( .D(o_data_jr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[2]) );
  DFC1 pipe_data_rs_reg_1_ ( .D(o_data_jr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[1]) );
  DFC1 pipe_data_rs_reg_0_ ( .D(o_data_jr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[0]) );
  DFC1 pipe_data_rt_reg_31_ ( .D(regbank_o_data_Rt[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[31]) );
  DFC1 pipe_data_rt_reg_30_ ( .D(regbank_o_data_Rt[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC1 pipe_data_rt_reg_29_ ( .D(regbank_o_data_Rt[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[29]) );
  DFC1 pipe_data_rt_reg_28_ ( .D(regbank_o_data_Rt[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28]) );
  DFC1 pipe_data_rt_reg_27_ ( .D(regbank_o_data_Rt[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27]) );
  DFC1 pipe_data_rt_reg_26_ ( .D(regbank_o_data_Rt[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26]) );
  DFC1 pipe_data_rt_reg_25_ ( .D(regbank_o_data_Rt[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25]) );
  DFC1 pipe_data_rt_reg_24_ ( .D(regbank_o_data_Rt[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24]) );
  DFC1 pipe_data_rt_reg_23_ ( .D(regbank_o_data_Rt[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23]) );
  DFC1 pipe_data_rt_reg_22_ ( .D(regbank_o_data_Rt[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC1 pipe_data_rt_reg_21_ ( .D(regbank_o_data_Rt[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21]) );
  DFC1 pipe_data_rt_reg_20_ ( .D(regbank_o_data_Rt[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20]) );
  DFC1 pipe_data_rt_reg_19_ ( .D(regbank_o_data_Rt[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19]) );
  DFC1 pipe_data_rt_reg_18_ ( .D(regbank_o_data_Rt[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18]) );
  DFC1 pipe_data_rt_reg_17_ ( .D(regbank_o_data_Rt[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17]) );
  DFC1 pipe_data_rt_reg_16_ ( .D(regbank_o_data_Rt[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC1 pipe_data_rt_reg_15_ ( .D(regbank_o_data_Rt[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15]) );
  DFC1 pipe_data_rt_reg_14_ ( .D(regbank_o_data_Rt[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14]) );
  DFC1 pipe_data_rt_reg_13_ ( .D(regbank_o_data_Rt[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC1 pipe_data_rt_reg_12_ ( .D(regbank_o_data_Rt[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12]) );
  DFC1 pipe_data_rt_reg_11_ ( .D(regbank_o_data_Rt[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11]) );
  DFC1 pipe_data_rt_reg_10_ ( .D(regbank_o_data_Rt[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC1 pipe_data_rt_reg_9_ ( .D(regbank_o_data_Rt[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[9]) );
  DFC1 pipe_data_rt_reg_8_ ( .D(regbank_o_data_Rt[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[8]) );
  DFC1 pipe_data_rt_reg_7_ ( .D(regbank_o_data_Rt[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[7]) );
  DFC1 pipe_data_rt_reg_6_ ( .D(regbank_o_data_Rt[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[6]) );
  DFC1 pipe_data_rt_reg_5_ ( .D(regbank_o_data_Rt[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[5]) );
  DFC1 pipe_data_rt_reg_4_ ( .D(regbank_o_data_Rt[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[4]) );
  DFC1 pipe_data_rt_reg_3_ ( .D(regbank_o_data_Rt[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[3]) );
  DFC1 pipe_data_rt_reg_2_ ( .D(regbank_o_data_Rt[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[2]) );
  DFC1 pipe_data_rt_reg_1_ ( .D(regbank_o_data_Rt[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[1]) );
  DFC1 pipe_data_rt_reg_0_ ( .D(regbank_o_data_Rt[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[0]) );
  DFC1 pipe_memout_reg_31_ ( .D(i_data_Wregwrite[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[31]) );
  DFC1 pipe_memout_reg_30_ ( .D(i_data_Wregwrite[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[30]) );
  DFC1 pipe_memout_reg_29_ ( .D(i_data_Wregwrite[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[29]) );
  DFC1 pipe_memout_reg_28_ ( .D(i_data_Wregwrite[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[28]) );
  DFC1 pipe_memout_reg_27_ ( .D(i_data_Wregwrite[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[27]) );
  DFC1 pipe_memout_reg_26_ ( .D(i_data_Wregwrite[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[26]) );
  DFC1 pipe_memout_reg_25_ ( .D(i_data_Wregwrite[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[25]) );
  DFC1 pipe_memout_reg_24_ ( .D(i_data_Wregwrite[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[24]) );
  DFC1 pipe_memout_reg_23_ ( .D(i_data_Wregwrite[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[23]) );
  DFC1 pipe_memout_reg_22_ ( .D(i_data_Wregwrite[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[22]) );
  DFC1 pipe_memout_reg_21_ ( .D(i_data_Wregwrite[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[21]) );
  DFC1 pipe_memout_reg_20_ ( .D(i_data_Wregwrite[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[20]) );
  DFC1 pipe_memout_reg_19_ ( .D(i_data_Wregwrite[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[19]) );
  DFC1 pipe_memout_reg_18_ ( .D(i_data_Wregwrite[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[18]) );
  DFC1 pipe_memout_reg_17_ ( .D(i_data_Wregwrite[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[17]) );
  DFC1 pipe_memout_reg_16_ ( .D(i_data_Wregwrite[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[16]) );
  DFC1 pipe_memout_reg_15_ ( .D(i_data_Wregwrite[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[15]) );
  DFC1 pipe_memout_reg_14_ ( .D(i_data_Wregwrite[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[14]) );
  DFC1 pipe_memout_reg_13_ ( .D(i_data_Wregwrite[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[13]) );
  DFC1 pipe_memout_reg_12_ ( .D(i_data_Wregwrite[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[12]) );
  DFC1 pipe_memout_reg_11_ ( .D(i_data_Wregwrite[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[11]) );
  DFC1 pipe_memout_reg_10_ ( .D(i_data_Wregwrite[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[10]) );
  DFC1 pipe_memout_reg_9_ ( .D(i_data_Wregwrite[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[9]) );
  DFC1 pipe_memout_reg_8_ ( .D(i_data_Wregwrite[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[8]) );
  DFC1 pipe_memout_reg_7_ ( .D(i_data_Wregwrite[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[7]) );
  DFC1 pipe_memout_reg_6_ ( .D(i_data_Wregwrite[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[6]) );
  DFC1 pipe_memout_reg_5_ ( .D(i_data_Wregwrite[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[5]) );
  DFC1 pipe_memout_reg_4_ ( .D(i_data_Wregwrite[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[4]) );
  DFC1 pipe_memout_reg_3_ ( .D(i_data_Wregwrite[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[3]) );
  DFC1 pipe_memout_reg_2_ ( .D(i_data_Wregwrite[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[2]) );
  DFC1 pipe_memout_reg_1_ ( .D(i_data_Wregwrite[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[1]) );
  DFC1 pipe_memout_reg_0_ ( .D(i_data_Wregwrite[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[0]) );
  DFC1 pipe_con_Efamux_reg_0_ ( .D(for_o_con_fa[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[0]) );
  DFC1 pipe_con_Efbmux_reg_0_ ( .D(for_o_con_fb[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[0]) );
  DFC1 pipe_addr_branch_reg_30_ ( .D(pcadd_o_addr_pcbranchE[30]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[30]) );
  DFC1 pipe_addr_branch_reg_29_ ( .D(pcadd_o_addr_pcbranchE[29]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[29]) );
  DFC1 pipe_addr_branch_reg_28_ ( .D(pcadd_o_addr_pcbranchE[28]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[28]) );
  DFC1 pipe_addr_branch_reg_26_ ( .D(pcadd_o_addr_pcbranchE[26]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[26]) );
  DFC1 pipe_addr_branch_reg_25_ ( .D(pcadd_o_addr_pcbranchE[25]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[25]) );
  DFC1 pipe_addr_branch_reg_22_ ( .D(pcadd_o_addr_pcbranchE[22]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[22]) );
  DFC1 pipe_addr_branch_reg_7_ ( .D(pcadd_o_addr_pcbranchE[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[7]) );
  DFC1 pipe_addr_branch_reg_6_ ( .D(pcadd_o_addr_pcbranchE[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[6]) );
  DFC1 pipe_addr_branch_reg_24_ ( .D(pcadd_o_addr_pcbranchE[24]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[24]) );
  DFC1 pipe_addr_branch_reg_21_ ( .D(pcadd_o_addr_pcbranchE[21]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[21]) );
  DFC1 pipe_addr_branch_reg_20_ ( .D(pcadd_o_addr_pcbranchE[20]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[20]) );
  DFC1 pipe_addr_branch_reg_18_ ( .D(pcadd_o_addr_pcbranchE[18]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[18]) );
  DFC1 pipe_addr_branch_reg_17_ ( .D(pcadd_o_addr_pcbranchE[17]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[17]) );
  DFC1 pipe_addr_branch_reg_15_ ( .D(pcadd_o_addr_pcbranchE[15]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[15]) );
  DFC1 pipe_addr_branch_reg_14_ ( .D(pcadd_o_addr_pcbranchE[14]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[14]) );
  DFC1 pipe_addr_branch_reg_11_ ( .D(pcadd_o_addr_pcbranchE[11]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[11]) );
  DFC1 pipe_addr_branch_reg_10_ ( .D(pcadd_o_addr_pcbranchE[10]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[10]) );
  DFC1 pipe_addr_pc4_reg_12_ ( .D(i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC1 pipe_addr_pc4_reg_6_ ( .D(i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC1 pipe_addr_pc4_reg_5_ ( .D(i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC1 pipe_addr_pc4_reg_3_ ( .D(i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC1 pipe_addr_rd_reg_4_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[4]) );
  DFC3 pipe_signext_o_data_immD_reg_15_ ( .D(signext_o_data_immD[15]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[15]) );
  BUF15 U3 ( .A(i_data_instr[21]), .Q(n123) );
  BUF6 U4 ( .A(i_data_instr[16]), .Q(n122) );
  LOGIC0 U5 ( .Q(o_con_Wmemtoreg) );
endmodule


module E_alu_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   ML_int_1__31_, ML_int_1__30_, ML_int_1__29_, ML_int_1__28_,
         ML_int_1__27_, ML_int_1__26_, ML_int_1__25_, ML_int_1__24_,
         ML_int_1__23_, ML_int_1__22_, ML_int_1__21_, ML_int_1__20_,
         ML_int_1__19_, ML_int_1__18_, ML_int_1__17_, ML_int_1__16_,
         ML_int_1__15_, ML_int_1__14_, ML_int_1__13_, ML_int_1__12_,
         ML_int_1__11_, ML_int_1__10_, ML_int_1__9_, ML_int_1__8_,
         ML_int_1__7_, ML_int_1__6_, ML_int_1__5_, ML_int_1__4_, ML_int_1__3_,
         ML_int_1__2_, ML_int_1__1_, ML_int_1__0_, ML_int_2__31_,
         ML_int_2__30_, ML_int_2__29_, ML_int_2__28_, ML_int_2__27_,
         ML_int_2__26_, ML_int_2__25_, ML_int_2__24_, ML_int_2__23_,
         ML_int_2__22_, ML_int_2__21_, ML_int_2__20_, ML_int_2__19_,
         ML_int_2__18_, ML_int_2__17_, ML_int_2__16_, ML_int_2__15_,
         ML_int_2__14_, ML_int_2__13_, ML_int_2__12_, ML_int_2__11_,
         ML_int_2__10_, ML_int_2__9_, ML_int_2__8_, ML_int_2__7_, ML_int_2__6_,
         ML_int_2__5_, ML_int_2__4_, ML_int_2__3_, ML_int_2__2_, ML_int_3__31_,
         ML_int_3__30_, ML_int_3__29_, ML_int_3__28_, ML_int_3__27_,
         ML_int_3__26_, ML_int_3__25_, ML_int_3__24_, ML_int_3__23_,
         ML_int_3__22_, ML_int_3__21_, ML_int_3__20_, ML_int_3__19_,
         ML_int_3__18_, ML_int_3__17_, ML_int_3__16_, ML_int_3__15_,
         ML_int_3__14_, ML_int_3__13_, ML_int_3__12_, ML_int_3__11_,
         ML_int_3__10_, ML_int_3__9_, ML_int_3__8_, ML_int_3__7_, ML_int_3__6_,
         ML_int_3__5_, ML_int_3__4_, ML_int_3__1_, ML_int_3__0_, ML_int_4__31_,
         ML_int_4__30_, ML_int_4__29_, ML_int_4__28_, ML_int_4__27_,
         ML_int_4__26_, ML_int_4__25_, ML_int_4__24_, ML_int_4__21_,
         ML_int_4__15_, ML_int_4__14_, ML_int_4__13_, ML_int_4__12_,
         ML_int_4__11_, ML_int_4__10_, ML_int_4__9_, ML_int_4__8_, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51;

  MUX21 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n1), .Q(ML_int_1__4_) );
  MUX21 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n16), .Q(ML_int_1__3_) );
  MUX22 M1_2_6 ( .A(ML_int_2__6_), .B(ML_int_2__2_), .S(n21), .Q(ML_int_3__6_)
         );
  MUX21 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n1), .Q(ML_int_1__6_) );
  MUX21 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n16), .Q(ML_int_1__20_) );
  MUX21 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n16), .Q(ML_int_1__19_) );
  MUX21 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n1), .Q(ML_int_1__11_) );
  MUX21 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n1), .Q(ML_int_1__10_) );
  MUX22 M1_1_7 ( .A(ML_int_1__7_), .B(ML_int_1__5_), .S(n17), .Q(ML_int_2__7_)
         );
  MUX22 M1_1_6 ( .A(ML_int_1__6_), .B(ML_int_1__4_), .S(n17), .Q(ML_int_2__6_)
         );
  MUX22 M1_1_4 ( .A(ML_int_1__4_), .B(ML_int_1__2_), .S(n17), .Q(ML_int_2__4_)
         );
  MUX21 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n1), .Q(ML_int_1__17_) );
  MUX21 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n1), .Q(ML_int_1__16_) );
  MUX22 M1_2_4 ( .A(ML_int_2__4_), .B(n38), .S(n20), .Q(ML_int_3__4_) );
  MUX22 M1_2_31 ( .A(ML_int_2__31_), .B(ML_int_2__27_), .S(n20), .Q(
        ML_int_3__31_) );
  MUX22 M1_3_31 ( .A(ML_int_3__31_), .B(ML_int_3__23_), .S(SH[3]), .Q(
        ML_int_4__31_) );
  MUX22 M1_4_31 ( .A(ML_int_4__31_), .B(ML_int_4__15_), .S(n25), .Q(B[31]) );
  MUX22 M1_2_30 ( .A(ML_int_2__30_), .B(ML_int_2__26_), .S(n20), .Q(
        ML_int_3__30_) );
  MUX22 M1_3_30 ( .A(ML_int_3__30_), .B(ML_int_3__22_), .S(SH[3]), .Q(
        ML_int_4__30_) );
  MUX22 M1_4_30 ( .A(ML_int_4__30_), .B(ML_int_4__14_), .S(n25), .Q(B[30]) );
  MUX22 M1_2_27 ( .A(ML_int_2__27_), .B(ML_int_2__23_), .S(n20), .Q(
        ML_int_3__27_) );
  MUX22 M1_3_27 ( .A(ML_int_3__27_), .B(ML_int_3__19_), .S(n23), .Q(
        ML_int_4__27_) );
  MUX22 M1_4_27 ( .A(ML_int_4__27_), .B(ML_int_4__11_), .S(n25), .Q(B[27]) );
  MUX22 M1_3_25 ( .A(ML_int_3__25_), .B(ML_int_3__17_), .S(SH[3]), .Q(
        ML_int_4__25_) );
  MUX22 M1_4_25 ( .A(ML_int_4__25_), .B(ML_int_4__9_), .S(n25), .Q(B[25]) );
  MUX22 M1_2_26 ( .A(ML_int_2__26_), .B(ML_int_2__22_), .S(n20), .Q(
        ML_int_3__26_) );
  MUX22 M1_3_26 ( .A(ML_int_3__26_), .B(ML_int_3__18_), .S(SH[3]), .Q(
        ML_int_4__26_) );
  MUX22 M1_4_26 ( .A(ML_int_4__26_), .B(ML_int_4__10_), .S(n25), .Q(B[26]) );
  MUX22 M1_2_29 ( .A(ML_int_2__29_), .B(ML_int_2__25_), .S(n20), .Q(
        ML_int_3__29_) );
  MUX22 M1_4_24 ( .A(ML_int_4__24_), .B(ML_int_4__8_), .S(n25), .Q(B[24]) );
  MUX22 M1_4_28 ( .A(ML_int_4__28_), .B(ML_int_4__12_), .S(n25), .Q(B[28]) );
  MUX22 M1_4_21 ( .A(ML_int_4__21_), .B(n34), .S(n25), .Q(B[21]) );
  MUX22 M1_1_28 ( .A(ML_int_1__28_), .B(ML_int_1__26_), .S(n18), .Q(
        ML_int_2__28_) );
  MUX22 M1_2_28 ( .A(ML_int_2__28_), .B(ML_int_2__24_), .S(n20), .Q(
        ML_int_3__28_) );
  MUX22 M1_3_28 ( .A(ML_int_3__28_), .B(ML_int_3__20_), .S(SH[3]), .Q(
        ML_int_4__28_) );
  MUX22 M1_1_3 ( .A(ML_int_1__3_), .B(ML_int_1__1_), .S(n17), .Q(ML_int_2__3_)
         );
  MUX22 M1_3_13 ( .A(ML_int_3__13_), .B(ML_int_3__5_), .S(n23), .Q(
        ML_int_4__13_) );
  MUX22 M1_3_10 ( .A(ML_int_3__10_), .B(n36), .S(n23), .Q(ML_int_4__10_) );
  MUX22 M1_3_12 ( .A(ML_int_3__12_), .B(ML_int_3__4_), .S(n23), .Q(
        ML_int_4__12_) );
  MUX22 M1_3_8 ( .A(ML_int_3__8_), .B(ML_int_3__0_), .S(n23), .Q(ML_int_4__8_)
         );
  MUX22 M1_3_9 ( .A(ML_int_3__9_), .B(ML_int_3__1_), .S(n23), .Q(ML_int_4__9_)
         );
  MUX22 M1_3_14 ( .A(ML_int_3__14_), .B(ML_int_3__6_), .S(n23), .Q(
        ML_int_4__14_) );
  MUX22 M1_2_15 ( .A(ML_int_2__15_), .B(ML_int_2__11_), .S(n21), .Q(
        ML_int_3__15_) );
  MUX22 M1_2_23 ( .A(ML_int_2__23_), .B(ML_int_2__19_), .S(n20), .Q(
        ML_int_3__23_) );
  MUX22 M1_1_26 ( .A(ML_int_1__26_), .B(ML_int_1__24_), .S(n18), .Q(
        ML_int_2__26_) );
  MUX22 M1_1_15 ( .A(ML_int_1__15_), .B(ML_int_1__13_), .S(n18), .Q(
        ML_int_2__15_) );
  MUX22 M1_1_25 ( .A(ML_int_1__25_), .B(ML_int_1__23_), .S(n18), .Q(
        ML_int_2__25_) );
  MUX22 M1_1_23 ( .A(ML_int_1__23_), .B(ML_int_1__21_), .S(n18), .Q(
        ML_int_2__23_) );
  MUX22 M1_1_27 ( .A(ML_int_1__27_), .B(ML_int_1__25_), .S(n18), .Q(
        ML_int_2__27_) );
  MUX22 M1_1_24 ( .A(ML_int_1__24_), .B(ML_int_1__22_), .S(n18), .Q(
        ML_int_2__24_) );
  MUX22 M1_2_13 ( .A(ML_int_2__13_), .B(ML_int_2__9_), .S(n21), .Q(
        ML_int_3__13_) );
  MUX22 M1_2_22 ( .A(ML_int_2__22_), .B(ML_int_2__18_), .S(n20), .Q(
        ML_int_3__22_) );
  MUX22 M1_2_14 ( .A(ML_int_2__14_), .B(ML_int_2__10_), .S(n21), .Q(
        ML_int_3__14_) );
  MUX22 M1_2_20 ( .A(ML_int_2__20_), .B(ML_int_2__16_), .S(n20), .Q(
        ML_int_3__20_) );
  MUX22 M1_2_12 ( .A(ML_int_2__12_), .B(ML_int_2__8_), .S(n21), .Q(
        ML_int_3__12_) );
  MUX22 M1_2_11 ( .A(ML_int_2__11_), .B(ML_int_2__7_), .S(n21), .Q(
        ML_int_3__11_) );
  MUX22 M1_2_9 ( .A(ML_int_2__9_), .B(ML_int_2__5_), .S(n21), .Q(ML_int_3__9_)
         );
  MUX22 M1_1_8 ( .A(ML_int_1__8_), .B(ML_int_1__6_), .S(n17), .Q(ML_int_2__8_)
         );
  MUX22 M1_2_7 ( .A(ML_int_2__7_), .B(ML_int_2__3_), .S(n21), .Q(ML_int_3__7_)
         );
  MUX22 M1_1_13 ( .A(ML_int_1__13_), .B(ML_int_1__11_), .S(n17), .Q(
        ML_int_2__13_) );
  MUX22 M1_1_22 ( .A(ML_int_1__22_), .B(ML_int_1__20_), .S(n18), .Q(
        ML_int_2__22_) );
  MUX22 M1_1_18 ( .A(ML_int_1__18_), .B(ML_int_1__16_), .S(n18), .Q(
        ML_int_2__18_) );
  MUX22 M1_1_14 ( .A(ML_int_1__14_), .B(ML_int_1__12_), .S(n17), .Q(
        ML_int_2__14_) );
  MUX22 M1_1_17 ( .A(ML_int_1__17_), .B(ML_int_1__15_), .S(n18), .Q(
        ML_int_2__17_) );
  MUX22 M1_1_16 ( .A(ML_int_1__16_), .B(ML_int_1__14_), .S(n18), .Q(
        ML_int_2__16_) );
  MUX22 M1_1_11 ( .A(ML_int_1__11_), .B(ML_int_1__9_), .S(n17), .Q(
        ML_int_2__11_) );
  MUX22 M1_1_10 ( .A(ML_int_1__10_), .B(ML_int_1__8_), .S(n17), .Q(
        ML_int_2__10_) );
  MUX22 M1_1_20 ( .A(ML_int_1__20_), .B(ML_int_1__18_), .S(n18), .Q(
        ML_int_2__20_) );
  MUX22 M1_1_12 ( .A(ML_int_1__12_), .B(ML_int_1__10_), .S(n17), .Q(
        ML_int_2__12_) );
  MUX22 M1_1_19 ( .A(ML_int_1__19_), .B(ML_int_1__17_), .S(n18), .Q(
        ML_int_2__19_) );
  MUX22 M1_2_5 ( .A(ML_int_2__5_), .B(n37), .S(n21), .Q(ML_int_3__5_) );
  MUX21 M1_2_25 ( .A(ML_int_2__25_), .B(ML_int_2__21_), .S(n20), .Q(
        ML_int_3__25_) );
  MUX21 M1_2_24 ( .A(ML_int_2__24_), .B(ML_int_2__20_), .S(n20), .Q(
        ML_int_3__24_) );
  MUX21 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n16), .Q(ML_int_1__30_) );
  MUX21 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n16), .Q(ML_int_1__31_) );
  MUX21 M1_3_29 ( .A(ML_int_3__29_), .B(ML_int_3__21_), .S(SH[3]), .Q(
        ML_int_4__29_) );
  MUX21 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n16), .Q(ML_int_1__24_) );
  MUX21 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n1), .Q(ML_int_1__18_) );
  MUX21 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n1), .Q(ML_int_1__14_) );
  MUX21 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n16), .Q(ML_int_1__23_) );
  MUX21 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n1), .Q(ML_int_1__15_) );
  MUX21 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n16), .Q(ML_int_1__22_) );
  MUX21 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n16), .Q(ML_int_1__26_) );
  MUX21 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n16), .Q(ML_int_1__28_) );
  MUX21 M1_3_21 ( .A(ML_int_3__21_), .B(ML_int_3__13_), .S(SH[3]), .Q(
        ML_int_4__21_) );
  MUX21 M1_2_16 ( .A(ML_int_2__16_), .B(ML_int_2__12_), .S(n21), .Q(
        ML_int_3__16_) );
  MUX21 M1_2_17 ( .A(ML_int_2__17_), .B(ML_int_2__13_), .S(n21), .Q(
        ML_int_3__17_) );
  MUX21 M1_2_8 ( .A(ML_int_2__8_), .B(ML_int_2__4_), .S(n21), .Q(ML_int_3__8_)
         );
  MUX21 M1_2_18 ( .A(ML_int_2__18_), .B(ML_int_2__14_), .S(n21), .Q(
        ML_int_3__18_) );
  MUX22 M1_1_30 ( .A(ML_int_1__30_), .B(ML_int_1__28_), .S(n18), .Q(
        ML_int_2__30_) );
  MUX22 M1_2_10 ( .A(ML_int_2__10_), .B(ML_int_2__6_), .S(n21), .Q(
        ML_int_3__10_) );
  MUX22 M1_2_19 ( .A(ML_int_2__19_), .B(ML_int_2__15_), .S(n20), .Q(
        ML_int_3__19_) );
  MUX22 M1_3_24 ( .A(ML_int_3__24_), .B(ML_int_3__16_), .S(SH[3]), .Q(
        ML_int_4__24_) );
  MUX22 M1_1_29 ( .A(ML_int_1__29_), .B(ML_int_1__27_), .S(n18), .Q(
        ML_int_2__29_) );
  MUX21 M1_1_31 ( .A(ML_int_1__31_), .B(ML_int_1__29_), .S(n18), .Q(
        ML_int_2__31_) );
  MUX22 M1_1_2 ( .A(ML_int_1__2_), .B(ML_int_1__0_), .S(n17), .Q(ML_int_2__2_)
         );
  MUX22 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n16), .Q(ML_int_1__29_) );
  MUX22 M1_1_21 ( .A(ML_int_1__21_), .B(ML_int_1__19_), .S(n18), .Q(
        ML_int_2__21_) );
  MUX22 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n1), .Q(ML_int_1__7_) );
  MUX24 M1_3_11 ( .A(ML_int_3__11_), .B(n35), .S(n23), .Q(ML_int_4__11_) );
  MUX21 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n16), .Q(ML_int_1__2_) );
  MUX22 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n1), .Q(ML_int_1__8_) );
  MUX21 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n1), .Q(ML_int_1__12_) );
  MUX22 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n16), .Q(ML_int_1__1_) );
  MUX22 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n16), .Q(ML_int_1__21_) );
  MUX22 M1_4_29 ( .A(ML_int_4__29_), .B(ML_int_4__13_), .S(n25), .Q(B[29]) );
  MUX22 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n16), .Q(ML_int_1__27_) );
  MUX22 M1_1_9 ( .A(ML_int_1__9_), .B(ML_int_1__7_), .S(n17), .Q(ML_int_2__9_)
         );
  MUX22 M1_1_5 ( .A(ML_int_1__5_), .B(ML_int_1__3_), .S(n17), .Q(ML_int_2__5_)
         );
  MUX22 M1_3_15 ( .A(ML_int_3__15_), .B(ML_int_3__7_), .S(n23), .Q(
        ML_int_4__15_) );
  MUX21 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n1), .Q(ML_int_1__9_) );
  MUX21 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n1), .Q(ML_int_1__13_) );
  MUX22 M1_2_21 ( .A(ML_int_2__21_), .B(ML_int_2__17_), .S(n20), .Q(
        ML_int_3__21_) );
  BUF6 U3 ( .A(SH[0]), .Q(n1) );
  INV3 U4 ( .A(n26), .Q(n8) );
  NOR21 U5 ( .A(n26), .B(n27), .Q(B[14]) );
  INV3 U6 ( .A(n7), .Q(B[15]) );
  NAND22 U7 ( .A(n8), .B(ML_int_4__15_), .Q(n7) );
  BUF6 U8 ( .A(SH[0]), .Q(n16) );
  INV3 U9 ( .A(SH[1]), .Q(n19) );
  CLKIN3 U10 ( .A(ML_int_4__14_), .Q(n27) );
  NAND22 U11 ( .A(ML_int_1__0_), .B(n19), .Q(n51) );
  NOR21 U12 ( .A(n39), .B(SH[0]), .Q(ML_int_1__0_) );
  NOR21 U13 ( .A(n26), .B(n33), .Q(B[8]) );
  NAND21 U14 ( .A(A[25]), .B(n2), .Q(n3) );
  NAND20 U15 ( .A(A[24]), .B(n16), .Q(n4) );
  NAND22 U16 ( .A(n3), .B(n4), .Q(ML_int_1__25_) );
  INV0 U17 ( .A(n16), .Q(n2) );
  NAND20 U18 ( .A(A[5]), .B(n2), .Q(n5) );
  NAND21 U19 ( .A(A[4]), .B(SH[0]), .Q(n6) );
  NAND22 U20 ( .A(n5), .B(n6), .Q(ML_int_1__5_) );
  CLKIN1 U21 ( .A(SH[2]), .Q(n22) );
  NAND22 U22 ( .A(ML_int_3__0_), .B(n24), .Q(n47) );
  NOR20 U23 ( .A(n51), .B(SH[2]), .Q(ML_int_3__0_) );
  NAND21 U24 ( .A(ML_int_2__2_), .B(n22), .Q(n49) );
  INV3 U25 ( .A(n19), .Q(n18) );
  INV1 U26 ( .A(n42), .Q(n34) );
  INV2 U27 ( .A(A[0]), .Q(n39) );
  CLKIN3 U28 ( .A(ML_int_4__10_), .Q(n31) );
  CLKIN3 U29 ( .A(ML_int_4__8_), .Q(n33) );
  NOR20 U30 ( .A(n50), .B(n21), .Q(ML_int_3__1_) );
  INV3 U31 ( .A(ML_int_4__9_), .Q(n32) );
  IMUX21 U32 ( .A(n15), .B(n45), .S(n26), .Q(B[18]) );
  IMUX21 U33 ( .A(ML_int_3__16_), .B(ML_int_3__8_), .S(n23), .Q(n13) );
  NAND20 U34 ( .A(ML_int_3__1_), .B(n24), .Q(n46) );
  IMUX20 U35 ( .A(ML_int_3__22_), .B(ML_int_3__14_), .S(SH[3]), .Q(n11) );
  IMUX20 U36 ( .A(ML_int_3__23_), .B(ML_int_3__15_), .S(SH[3]), .Q(n12) );
  IMUX20 U37 ( .A(ML_int_3__19_), .B(ML_int_3__11_), .S(n23), .Q(n14) );
  IMUX20 U38 ( .A(ML_int_3__18_), .B(ML_int_3__10_), .S(n23), .Q(n15) );
  IMUX20 U39 ( .A(ML_int_3__17_), .B(ML_int_3__9_), .S(n23), .Q(n9) );
  IMUX20 U40 ( .A(ML_int_3__20_), .B(ML_int_3__12_), .S(n23), .Q(n10) );
  NAND21 U41 ( .A(ML_int_3__6_), .B(n24), .Q(n41) );
  CLKIN3 U42 ( .A(ML_int_4__11_), .Q(n30) );
  NOR21 U43 ( .A(n26), .B(n30), .Q(B[11]) );
  CLKIN3 U44 ( .A(ML_int_4__12_), .Q(n29) );
  NOR21 U45 ( .A(n26), .B(n29), .Q(B[12]) );
  BUF2 U46 ( .A(SH[4]), .Q(n25) );
  INV3 U47 ( .A(n51), .Q(n38) );
  INV3 U48 ( .A(ML_int_4__13_), .Q(n28) );
  INV3 U49 ( .A(n22), .Q(n20) );
  INV3 U50 ( .A(n22), .Q(n21) );
  INV3 U51 ( .A(n19), .Q(n17) );
  NOR21 U52 ( .A(n26), .B(n47), .Q(B[0]) );
  NAND22 U53 ( .A(ML_int_3__5_), .B(n24), .Q(n42) );
  INV3 U54 ( .A(n48), .Q(n35) );
  IMUX21 U55 ( .A(n9), .B(n46), .S(n26), .Q(B[17]) );
  IMUX21 U56 ( .A(n10), .B(n43), .S(n25), .Q(B[20]) );
  IMUX21 U57 ( .A(n11), .B(n41), .S(n25), .Q(B[22]) );
  IMUX21 U58 ( .A(n12), .B(n40), .S(n25), .Q(B[23]) );
  IMUX21 U59 ( .A(n13), .B(n47), .S(n26), .Q(B[16]) );
  IMUX21 U60 ( .A(n14), .B(n44), .S(n25), .Q(B[19]) );
  INV3 U61 ( .A(n24), .Q(n23) );
  INV3 U62 ( .A(SH[3]), .Q(n24) );
  BUF2 U63 ( .A(SH[4]), .Q(n26) );
  NAND22 U64 ( .A(ML_int_3__4_), .B(n24), .Q(n43) );
  NAND22 U65 ( .A(ML_int_1__1_), .B(n19), .Q(n50) );
  NAND22 U66 ( .A(ML_int_3__7_), .B(n24), .Q(n40) );
  NAND21 U67 ( .A(ML_int_2__3_), .B(n22), .Q(n48) );
  NAND21 U68 ( .A(n35), .B(n24), .Q(n44) );
  INV3 U69 ( .A(n50), .Q(n37) );
  NAND22 U70 ( .A(n36), .B(n24), .Q(n45) );
  CLKIN3 U71 ( .A(n49), .Q(n36) );
  NOR20 U72 ( .A(n26), .B(n32), .Q(B[9]) );
  NOR20 U73 ( .A(n26), .B(n40), .Q(B[7]) );
  NOR20 U74 ( .A(n26), .B(n41), .Q(B[6]) );
  NOR20 U75 ( .A(n26), .B(n42), .Q(B[5]) );
  NOR20 U76 ( .A(n26), .B(n43), .Q(B[4]) );
  NOR20 U77 ( .A(n26), .B(n44), .Q(B[3]) );
  NOR20 U78 ( .A(n26), .B(n45), .Q(B[2]) );
  NOR20 U79 ( .A(n26), .B(n46), .Q(B[1]) );
  NOR20 U80 ( .A(n26), .B(n28), .Q(B[13]) );
  NOR20 U81 ( .A(n26), .B(n31), .Q(B[10]) );
endmodule


module E_alu_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263;

  NAND30 U1 ( .A(n92), .B(n55), .C(B[7]), .Q(n168) );
  INV3 U2 ( .A(n55), .Q(n73) );
  INV3 U3 ( .A(n175), .Q(n92) );
  NAND24 U4 ( .A(A[23]), .B(n13), .Q(n55) );
  NOR21 U5 ( .A(n255), .B(n148), .Q(n247) );
  INV0 U6 ( .A(B[19]), .Q(n11) );
  AOI221 U7 ( .A(n49), .B(n50), .C(n51), .D(n50), .Q(n48) );
  NOR22 U8 ( .A(n234), .B(n235), .Q(n233) );
  NAND43 U9 ( .A(n45), .B(n46), .C(n47), .D(n48), .Q(n44) );
  CLKIN1 U10 ( .A(B[8]), .Q(n7) );
  INV0 U11 ( .A(B[20]), .Q(n12) );
  CLKIN3 U12 ( .A(B[27]), .Q(n16) );
  NOR21 U13 ( .A(n173), .B(n174), .Q(n172) );
  NAND22 U14 ( .A(n224), .B(n2), .Q(n192) );
  INV3 U15 ( .A(n1), .Q(n2) );
  NAND31 U16 ( .A(n223), .B(n222), .C(n191), .Q(n1) );
  NOR21 U17 ( .A(B[27]), .B(n23), .Q(n148) );
  NOR22 U18 ( .A(n256), .B(n257), .Q(n246) );
  NAND26 U19 ( .A(A[22]), .B(n262), .Q(n81) );
  NOR22 U20 ( .A(n68), .B(n69), .Q(n67) );
  AOI2111 U21 ( .A(n118), .B(n50), .C(n119), .D(n120), .Q(n25) );
  NOR22 U22 ( .A(n143), .B(n144), .Q(n142) );
  NOR21 U23 ( .A(n73), .B(n10), .Q(n65) );
  NOR22 U24 ( .A(n156), .B(n157), .Q(n24) );
  NAND21 U25 ( .A(A[11]), .B(n198), .Q(n96) );
  AOI310 U26 ( .A(n98), .B(n99), .C(n50), .D(n100), .Q(n87) );
  NOR21 U27 ( .A(n83), .B(n101), .Q(n100) );
  INV3 U28 ( .A(n146), .Q(n83) );
  AOI221 U29 ( .A(n136), .B(n76), .C(n137), .D(n138), .Q(n127) );
  INV3 U30 ( .A(n81), .Q(n60) );
  NOR33 U31 ( .A(n3), .B(n4), .C(n5), .Q(n6) );
  CLKIN3 U32 ( .A(n50), .Q(n5) );
  NAND21 U33 ( .A(A[9]), .B(n114), .Q(n176) );
  NOR24 U34 ( .A(n43), .B(n44), .Q(n26) );
  NOR23 U35 ( .A(n6), .B(n67), .Q(n47) );
  CLKIN3 U36 ( .A(B[17]), .Q(n261) );
  NOR23 U37 ( .A(n14), .B(n22), .Q(n143) );
  NOR20 U38 ( .A(n83), .B(n141), .Q(n137) );
  INV12 U39 ( .A(n123), .Q(n50) );
  INV2 U40 ( .A(B[30]), .Q(n36) );
  INV2 U41 ( .A(B[22]), .Q(n262) );
  NAND20 U42 ( .A(B[18]), .B(n55), .Q(n242) );
  NOR20 U43 ( .A(B[18]), .B(n244), .Q(n250) );
  NOR20 U44 ( .A(B[2]), .B(n209), .Q(n215) );
  NAND22 U45 ( .A(n172), .B(n50), .Q(n159) );
  NAND43 U46 ( .A(n246), .B(n247), .C(n248), .D(n249), .Q(n123) );
  OAI311 U47 ( .A(n192), .B(n193), .C(n194), .D(n195), .Q(n158) );
  NAND21 U48 ( .A(B[6]), .B(n202), .Q(n191) );
  CLKIN3 U49 ( .A(B[23]), .Q(n13) );
  INV3 U50 ( .A(n225), .Q(n224) );
  INV2 U51 ( .A(n66), .Q(n4) );
  INV2 U52 ( .A(n65), .Q(n3) );
  NOR21 U53 ( .A(B[0]), .B(n218), .Q(n220) );
  NAND31 U54 ( .A(n89), .B(n50), .C(n90), .Q(n88) );
  NOR21 U55 ( .A(B[25]), .B(n145), .Q(n144) );
  INV6 U56 ( .A(n15), .Q(n14) );
  NAND41 U57 ( .A(n107), .B(n108), .C(n109), .D(n50), .Q(n86) );
  NAND30 U58 ( .A(n95), .B(n96), .C(n72), .Q(n197) );
  NAND30 U59 ( .A(n92), .B(n55), .C(B[8]), .Q(n91) );
  INV1 U60 ( .A(n41), .Q(n39) );
  INV3 U61 ( .A(n82), .Q(n253) );
  INV1 U62 ( .A(B[2]), .Q(n228) );
  INV2 U63 ( .A(B[9]), .Q(n114) );
  NOR21 U64 ( .A(n250), .B(n251), .Q(n249) );
  NOR22 U65 ( .A(n252), .B(n253), .Q(n248) );
  INV1 U66 ( .A(n37), .Q(n34) );
  INV2 U67 ( .A(n191), .Q(n184) );
  NOR21 U68 ( .A(n91), .B(n54), .Q(n90) );
  AOI311 U69 ( .A(n161), .B(n50), .C(n162), .D(n41), .Q(n160) );
  CLKIN1 U70 ( .A(B[14]), .Q(n239) );
  NAND20 U71 ( .A(n134), .B(n20), .Q(n132) );
  NAND24 U72 ( .A(A[16]), .B(n10), .Q(n95) );
  NOR30 U73 ( .A(n114), .B(n60), .C(n73), .Q(n108) );
  NAND20 U74 ( .A(n142), .B(B[21]), .Q(n141) );
  NOR20 U75 ( .A(n83), .B(n84), .Q(n77) );
  NAND20 U76 ( .A(n142), .B(B[20]), .Q(n84) );
  NOR20 U77 ( .A(n73), .B(n83), .Q(n130) );
  NOR20 U78 ( .A(n135), .B(n11), .Q(n129) );
  NOR20 U79 ( .A(B[26]), .B(n149), .Q(n147) );
  NOR22 U80 ( .A(n147), .B(n148), .Q(n146) );
  NAND30 U81 ( .A(n72), .B(n95), .C(n81), .Q(n170) );
  NOR20 U82 ( .A(n60), .B(n71), .Q(n66) );
  NAND20 U83 ( .A(n55), .B(n81), .Q(n80) );
  NAND20 U84 ( .A(n182), .B(n181), .Q(n238) );
  NOR20 U85 ( .A(n104), .B(n54), .Q(n99) );
  NAND20 U86 ( .A(n72), .B(n95), .Q(n110) );
  NAND20 U87 ( .A(B[31]), .B(n165), .Q(n37) );
  XNR20 U88 ( .A(B[31]), .B(A[31]), .Q(n33) );
  OAI2110 U89 ( .A(n184), .B(n185), .C(n55), .D(n81), .Q(n173) );
  NAND30 U90 ( .A(n72), .B(n95), .C(n81), .Q(n94) );
  NAND20 U91 ( .A(B[15]), .B(n55), .Q(n258) );
  NAND20 U92 ( .A(n233), .B(n50), .Q(n232) );
  NAND30 U93 ( .A(B[13]), .B(n81), .C(n55), .Q(n235) );
  NAND20 U94 ( .A(n81), .B(n72), .Q(n105) );
  NAND20 U95 ( .A(n126), .B(n76), .Q(n121) );
  NAND40 U96 ( .A(n81), .B(n125), .C(B[17]), .D(n55), .Q(n124) );
  NAND20 U97 ( .A(B[22]), .B(n142), .Q(n122) );
  NAND20 U98 ( .A(n241), .B(n50), .Q(n231) );
  NAND20 U99 ( .A(n81), .B(n244), .Q(n243) );
  NAND20 U100 ( .A(n81), .B(n82), .Q(n133) );
  NAND20 U101 ( .A(n72), .B(n19), .Q(n71) );
  NAND20 U102 ( .A(B[29]), .B(n166), .Q(n164) );
  INV2 U103 ( .A(n167), .Q(n163) );
  INV0 U104 ( .A(B[28]), .Q(n117) );
  INV1 U105 ( .A(B[12]), .Q(n9) );
  NOR20 U106 ( .A(B[13]), .B(n181), .Q(n180) );
  INV0 U107 ( .A(B[25]), .Q(n150) );
  INV2 U108 ( .A(n227), .Q(n226) );
  NOR20 U109 ( .A(B[5]), .B(n189), .Q(n187) );
  NAND20 U110 ( .A(B[12]), .B(n55), .Q(n53) );
  NAND20 U111 ( .A(n81), .B(n140), .Q(n139) );
  NAND30 U112 ( .A(B[14]), .B(n81), .C(n55), .Q(n152) );
  NAND20 U113 ( .A(A[30]), .B(n36), .Q(n35) );
  NAND20 U114 ( .A(B[23]), .B(n70), .Q(n69) );
  NOR20 U115 ( .A(B[29]), .B(n166), .Q(n38) );
  NOR20 U116 ( .A(B[28]), .B(n42), .Q(n40) );
  INV2 U117 ( .A(n102), .Q(n101) );
  INV0 U118 ( .A(B[26]), .Q(n103) );
  NAND22 U119 ( .A(n142), .B(n76), .Q(n68) );
  INV3 U120 ( .A(n95), .Q(n58) );
  NAND22 U121 ( .A(A[20]), .B(n12), .Q(n134) );
  NOR21 U122 ( .A(n59), .B(n60), .Q(n63) );
  NOR21 U123 ( .A(n59), .B(n60), .Q(n56) );
  NOR21 U124 ( .A(A[27]), .B(n16), .Q(n115) );
  NOR21 U125 ( .A(A[24]), .B(n15), .Q(n74) );
  NAND31 U126 ( .A(n230), .B(n231), .C(n232), .Q(n156) );
  NOR21 U127 ( .A(n211), .B(n212), .Q(n193) );
  NAND22 U128 ( .A(n219), .B(B[0]), .Q(n211) );
  NAND22 U129 ( .A(n213), .B(n214), .Q(n212) );
  NOR21 U130 ( .A(B[19]), .B(n20), .Q(n251) );
  INV3 U131 ( .A(A[8]), .Q(n17) );
  INV3 U132 ( .A(A[24]), .Q(n22) );
  INV3 U133 ( .A(A[19]), .Q(n20) );
  INV3 U134 ( .A(A[27]), .Q(n23) );
  INV3 U135 ( .A(n207), .Q(n206) );
  NAND22 U136 ( .A(n77), .B(n78), .Q(n45) );
  NAND22 U137 ( .A(n74), .B(n75), .Q(n46) );
  NAND31 U138 ( .A(n28), .B(n29), .C(n30), .Q(n27) );
  NAND42 U139 ( .A(n85), .B(n86), .C(n87), .D(n88), .Q(n43) );
  NOR21 U140 ( .A(n115), .B(n116), .Q(n85) );
  NAND22 U141 ( .A(A[10]), .B(n8), .Q(n97) );
  NAND31 U142 ( .A(n96), .B(n171), .C(n97), .Q(n169) );
  NOR21 U143 ( .A(n169), .B(n170), .Q(n161) );
  INV3 U144 ( .A(A[31]), .Q(n165) );
  NOR31 U145 ( .A(n110), .B(n111), .C(n112), .Q(n109) );
  NAND22 U146 ( .A(n96), .B(n113), .Q(n112) );
  INV3 U147 ( .A(A[16]), .Q(n19) );
  NOR21 U148 ( .A(B[26]), .B(n149), .Q(n255) );
  NAND22 U149 ( .A(n182), .B(n183), .Q(n179) );
  NAND22 U150 ( .A(n236), .B(n237), .Q(n234) );
  NOR21 U151 ( .A(n155), .B(n238), .Q(n237) );
  NOR21 U152 ( .A(n93), .B(n94), .Q(n89) );
  NAND31 U153 ( .A(n96), .B(n17), .C(n97), .Q(n93) );
  NAND22 U154 ( .A(n96), .B(n18), .Q(n106) );
  INV3 U155 ( .A(A[10]), .Q(n18) );
  NAND22 U156 ( .A(n107), .B(n92), .Q(n174) );
  NOR21 U157 ( .A(B[25]), .B(n145), .Q(n257) );
  NOR22 U158 ( .A(n14), .B(n22), .Q(n256) );
  NOR21 U159 ( .A(n79), .B(n80), .Q(n78) );
  NAND22 U160 ( .A(n82), .B(n21), .Q(n79) );
  INV3 U161 ( .A(A[20]), .Q(n21) );
  INV3 U162 ( .A(B[5]), .Q(n188) );
  NOR21 U163 ( .A(n242), .B(n243), .Q(n241) );
  NAND22 U164 ( .A(n127), .B(n128), .Q(n119) );
  NAND31 U165 ( .A(n129), .B(n130), .C(n131), .Q(n128) );
  NOR21 U166 ( .A(n132), .B(n133), .Q(n131) );
  NOR21 U167 ( .A(n31), .B(n32), .Q(n30) );
  NOR21 U168 ( .A(n33), .B(n34), .Q(n32) );
  NOR21 U169 ( .A(n34), .B(n35), .Q(n31) );
  NAND22 U170 ( .A(n245), .B(n50), .Q(n230) );
  NOR31 U171 ( .A(n258), .B(n259), .C(n260), .Q(n245) );
  NAND22 U172 ( .A(n81), .B(n72), .Q(n260) );
  NAND22 U173 ( .A(n95), .B(n263), .Q(n259) );
  INV3 U174 ( .A(B[24]), .Q(n15) );
  INV3 U175 ( .A(n142), .Q(n135) );
  NOR21 U176 ( .A(n196), .B(n197), .Q(n195) );
  NAND22 U177 ( .A(n97), .B(n199), .Q(n196) );
  INV3 U178 ( .A(n229), .Q(n222) );
  INV3 U179 ( .A(n215), .Q(n214) );
  NAND22 U180 ( .A(A[15]), .B(n240), .Q(n183) );
  INV3 U181 ( .A(B[15]), .Q(n240) );
  NOR21 U182 ( .A(A[2]), .B(n228), .Q(n227) );
  NOR21 U183 ( .A(A[30]), .B(n36), .Q(n167) );
  NAND22 U184 ( .A(A[21]), .B(n254), .Q(n82) );
  INV3 U185 ( .A(B[21]), .Q(n254) );
  INV3 U186 ( .A(A[5]), .Q(n189) );
  NAND22 U187 ( .A(n63), .B(n64), .Q(n61) );
  NOR21 U188 ( .A(A[11]), .B(n58), .Q(n64) );
  NOR21 U189 ( .A(A[5]), .B(n188), .Q(n229) );
  NOR21 U190 ( .A(A[22]), .B(n73), .Q(n126) );
  NAND22 U191 ( .A(A[14]), .B(n239), .Q(n182) );
  NAND31 U192 ( .A(n163), .B(n164), .C(n37), .Q(n41) );
  INV3 U193 ( .A(A[29]), .Q(n166) );
  NAND22 U194 ( .A(n176), .B(n177), .Q(n175) );
  NAND22 U195 ( .A(A[8]), .B(n7), .Q(n177) );
  INV3 U196 ( .A(A[23]), .Q(n70) );
  NOR21 U197 ( .A(n73), .B(n139), .Q(n138) );
  INV3 U198 ( .A(A[21]), .Q(n140) );
  NOR31 U199 ( .A(n52), .B(n53), .C(n54), .Q(n51) );
  NAND22 U200 ( .A(n56), .B(n57), .Q(n52) );
  NAND22 U201 ( .A(n38), .B(n39), .Q(n29) );
  NAND22 U202 ( .A(n40), .B(n39), .Q(n28) );
  INV3 U203 ( .A(A[28]), .Q(n42) );
  NOR21 U204 ( .A(n151), .B(n152), .Q(n118) );
  NAND22 U205 ( .A(n153), .B(n154), .Q(n151) );
  NOR21 U206 ( .A(A[14]), .B(n155), .Q(n154) );
  NOR21 U207 ( .A(A[28]), .B(n117), .Q(n116) );
  NOR21 U208 ( .A(A[26]), .B(n103), .Q(n102) );
  NOR21 U209 ( .A(A[25]), .B(n150), .Q(n136) );
  INV3 U210 ( .A(A[25]), .Q(n145) );
  INV3 U211 ( .A(A[26]), .Q(n149) );
  INV3 U212 ( .A(A[15]), .Q(n263) );
  INV3 U213 ( .A(A[18]), .Q(n244) );
  INV3 U214 ( .A(A[9]), .Q(n113) );
  INV3 U215 ( .A(A[13]), .Q(n181) );
  INV3 U216 ( .A(A[17]), .Q(n125) );
  INV3 U217 ( .A(A[0]), .Q(n218) );
  INV3 U218 ( .A(A[7]), .Q(n171) );
  INV3 U219 ( .A(A[4]), .Q(n190) );
  INV3 U220 ( .A(A[3]), .Q(n217) );
  INV3 U221 ( .A(A[2]), .Q(n209) );
  INV3 U222 ( .A(A[6]), .Q(n202) );
  INV3 U223 ( .A(A[1]), .Q(n210) );
  NAND20 U224 ( .A(B[10]), .B(n55), .Q(n104) );
  INV0 U225 ( .A(B[10]), .Q(n8) );
  INV3 U226 ( .A(B[16]), .Q(n10) );
  NOR21 U227 ( .A(A[12]), .B(n58), .Q(n57) );
  NOR31 U228 ( .A(n105), .B(n58), .C(n106), .Q(n98) );
  NOR21 U229 ( .A(n58), .B(n59), .Q(n153) );
  NOR21 U230 ( .A(n58), .B(n59), .Q(n236) );
  NAND20 U231 ( .A(B[4]), .B(n190), .Q(n223) );
  NOR20 U232 ( .A(B[7]), .B(n171), .Q(n200) );
  NOR20 U233 ( .A(A[3]), .B(n208), .Q(n207) );
  NOR21 U234 ( .A(A[0]), .B(n216), .Q(n213) );
  OAI311 U235 ( .A(n203), .B(n204), .C(n205), .D(n206), .Q(n194) );
  NOR21 U236 ( .A(n204), .B(n226), .Q(n225) );
  NOR21 U237 ( .A(n220), .B(n221), .Q(n219) );
  NOR21 U238 ( .A(n200), .B(n201), .Q(n199) );
  NOR20 U239 ( .A(n168), .B(n54), .Q(n162) );
  CLKIN0 U240 ( .A(B[1]), .Q(n205) );
  NOR20 U241 ( .A(B[1]), .B(n210), .Q(n221) );
  CLKIN0 U242 ( .A(B[11]), .Q(n198) );
  NAND20 U243 ( .A(B[11]), .B(n55), .Q(n62) );
  NOR31 U244 ( .A(n61), .B(n62), .C(n54), .Q(n49) );
  INV0 U245 ( .A(B[3]), .Q(n208) );
  NOR20 U246 ( .A(B[3]), .B(n217), .Q(n216) );
  NOR20 U247 ( .A(B[3]), .B(n217), .Q(n204) );
  NOR20 U248 ( .A(B[4]), .B(n190), .Q(n186) );
  NOR20 U249 ( .A(B[6]), .B(n202), .Q(n201) );
  OAI210 U250 ( .A(B[2]), .B(n209), .C(n210), .Q(n203) );
  AOI312 U251 ( .A(n24), .B(n25), .C(n26), .D(n27), .Q(LT_LE) );
  CLKIN3 U252 ( .A(n68), .Q(n75) );
  CLKIN3 U253 ( .A(n97), .Q(n111) );
  OAI222 U254 ( .A(n121), .B(n122), .C(n5), .D(n124), .Q(n120) );
  CLKIN3 U255 ( .A(n83), .Q(n76) );
  OAI212 U256 ( .A(n158), .B(n159), .C(n160), .Q(n157) );
  CLKIN3 U257 ( .A(n54), .Q(n107) );
  CLKIN6 U258 ( .A(n178), .Q(n54) );
  AOI2112 U259 ( .A(A[12]), .B(n9), .C(n179), .D(n180), .Q(n178) );
  OAI222 U260 ( .A(n186), .B(n187), .C(A[5]), .D(n188), .Q(n185) );
  CLKIN3 U261 ( .A(n183), .Q(n155) );
  CLKIN3 U262 ( .A(n72), .Q(n59) );
  CLKIN3 U263 ( .A(n134), .Q(n252) );
  NAND24 U264 ( .A(A[17]), .B(n261), .Q(n72) );
endmodule


module E_alu_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222;

  NAND21 U3 ( .A(n55), .B(n44), .Q(n53) );
  INV1 U4 ( .A(n44), .Q(n129) );
  NAND22 U5 ( .A(n89), .B(n90), .Q(n88) );
  NOR24 U6 ( .A(A[11]), .B(n171), .Q(n170) );
  NOR23 U7 ( .A(A[15]), .B(n103), .Q(n102) );
  INV8 U8 ( .A(B[15]), .Q(n103) );
  NOR23 U9 ( .A(n113), .B(n102), .Q(n112) );
  NOR24 U10 ( .A(n218), .B(n219), .Q(n217) );
  NOR24 U11 ( .A(A[4]), .B(n65), .Q(n218) );
  NOR24 U12 ( .A(A[7]), .B(n193), .Q(n219) );
  NAND24 U13 ( .A(n89), .B(n2), .Q(n85) );
  NAND33 U14 ( .A(n35), .B(n37), .C(n217), .Q(n128) );
  INV6 U15 ( .A(n128), .Q(n13) );
  NOR22 U16 ( .A(A[3]), .B(n204), .Q(n203) );
  INV6 U17 ( .A(B[9]), .Q(n167) );
  NOR23 U18 ( .A(n104), .B(n105), .Q(n86) );
  NAND22 U19 ( .A(n107), .B(n44), .Q(n104) );
  NAND23 U20 ( .A(A[5]), .B(n196), .Q(n56) );
  NAND24 U21 ( .A(n160), .B(n161), .Q(n90) );
  NAND22 U22 ( .A(n182), .B(n183), .Q(n25) );
  NAND22 U23 ( .A(B[9]), .B(n216), .Q(n21) );
  INV6 U24 ( .A(B[3]), .Q(n204) );
  NAND21 U25 ( .A(n21), .B(n22), .Q(n10) );
  OAI2110 U26 ( .A(n180), .B(n19), .C(n172), .D(n22), .Q(n177) );
  OAI2110 U27 ( .A(n17), .B(n190), .C(n191), .D(n22), .Q(n189) );
  NAND34 U28 ( .A(n82), .B(n69), .C(n211), .Q(n106) );
  NAND34 U29 ( .A(n208), .B(n69), .C(n209), .Q(n45) );
  INV6 U30 ( .A(n147), .Q(n99) );
  NOR21 U31 ( .A(n141), .B(n142), .Q(n139) );
  NAND22 U32 ( .A(A[4]), .B(n65), .Q(n38) );
  INV3 U33 ( .A(B[8]), .Q(n5) );
  INV3 U34 ( .A(n17), .Q(n124) );
  NAND23 U35 ( .A(A[12]), .B(n7), .Q(n147) );
  NAND33 U36 ( .A(n201), .B(n69), .C(n202), .Q(n44) );
  NOR22 U37 ( .A(A[12]), .B(n7), .Q(n113) );
  NAND33 U38 ( .A(n162), .B(n163), .C(n164), .Q(n161) );
  NOR23 U39 ( .A(n174), .B(n175), .Q(n108) );
  NAND22 U40 ( .A(A[7]), .B(n193), .Q(n109) );
  NAND22 U41 ( .A(n69), .B(n75), .Q(n71) );
  AOI211 U42 ( .A(n38), .B(n51), .C(n52), .Q(n50) );
  AOI211 U43 ( .A(n29), .B(n30), .C(n31), .Q(n28) );
  AOI221 U44 ( .A(n177), .B(n178), .C(n25), .D(n179), .Q(n176) );
  NAND22 U45 ( .A(A[10]), .B(n6), .Q(n172) );
  CLKIN6 U46 ( .A(B[12]), .Q(n7) );
  INV3 U47 ( .A(n82), .Q(n72) );
  INV3 U48 ( .A(n35), .Q(n36) );
  AOI310 U49 ( .A(n12), .B(n13), .C(n14), .D(n15), .Q(n11) );
  NOR22 U50 ( .A(A[9]), .B(n167), .Q(n166) );
  NAND20 U51 ( .A(n109), .B(n17), .Q(n140) );
  NAND23 U52 ( .A(n194), .B(n195), .Q(n17) );
  CLKIN3 U53 ( .A(n106), .Q(n40) );
  OAI211 U54 ( .A(n40), .B(n41), .C(n42), .Q(n39) );
  NOR22 U55 ( .A(n203), .B(n210), .Q(n209) );
  NOR22 U56 ( .A(B[0]), .B(n72), .Q(n208) );
  OAI212 U57 ( .A(B[8]), .B(n8), .C(n22), .Q(n163) );
  CLKIN3 U58 ( .A(B[10]), .Q(n6) );
  NAND24 U59 ( .A(A[9]), .B(n167), .Q(n22) );
  AOI312 U60 ( .A(n56), .B(n33), .C(n38), .D(n36), .Q(n195) );
  NOR21 U61 ( .A(n124), .B(n20), .Q(n182) );
  NAND24 U62 ( .A(n108), .B(n13), .Q(n1) );
  CLKIN6 U63 ( .A(n131), .Q(n47) );
  OAI312 U64 ( .A(n53), .B(n54), .C(n40), .D(n42), .Q(n51) );
  CLKIN3 U65 ( .A(B[11]), .Q(n171) );
  CLKIN6 U66 ( .A(n170), .Q(n164) );
  XNR22 U67 ( .A(n114), .B(n4), .Q(DIFF[15]) );
  AOI312 U68 ( .A(n91), .B(n92), .C(n93), .D(n94), .Q(n87) );
  NOR22 U69 ( .A(n165), .B(n166), .Q(n162) );
  NAND21 U70 ( .A(n146), .B(n147), .Q(n145) );
  CLKIN1 U71 ( .A(n108), .Q(n141) );
  OAI2112 U72 ( .A(n124), .B(n125), .C(n126), .D(n115), .Q(n123) );
  INV3 U73 ( .A(n127), .Q(n126) );
  INV2 U74 ( .A(n45), .Q(n54) );
  NAND30 U75 ( .A(n43), .B(n44), .C(n45), .Q(n41) );
  INV2 U76 ( .A(n14), .Q(n63) );
  AOI211 U77 ( .A(n42), .B(n14), .C(n59), .Q(n58) );
  AOI2111 U78 ( .A(n152), .B(n14), .C(n153), .D(n116), .Q(n151) );
  AOI311 U79 ( .A(n13), .B(n188), .C(n14), .D(n189), .Q(n187) );
  NAND43 U80 ( .A(n106), .B(n45), .C(n200), .D(n44), .Q(n14) );
  NAND24 U81 ( .A(n106), .B(n45), .Q(n105) );
  NAND32 U82 ( .A(n13), .B(n139), .C(n14), .Q(n138) );
  CLKIN4 U83 ( .A(n203), .Q(n202) );
  NAND22 U84 ( .A(n146), .B(n147), .Q(n116) );
  NAND31 U85 ( .A(n185), .B(n44), .C(n45), .Q(n184) );
  INV3 U86 ( .A(B[7]), .Q(n193) );
  NAND22 U87 ( .A(n131), .B(n109), .Q(n130) );
  INV3 U88 ( .A(n109), .Q(n20) );
  OAI211 U89 ( .A(n16), .B(n109), .C(n19), .Q(n192) );
  AOI211 U90 ( .A(n108), .B(n25), .C(n90), .Q(n159) );
  AOI312 U91 ( .A(n120), .B(n121), .C(n122), .D(n123), .Q(n117) );
  NOR22 U92 ( .A(n54), .B(n40), .Q(n121) );
  OAI222 U93 ( .A(A[9]), .B(n167), .C(A[10]), .D(n6), .Q(n175) );
  INV0 U94 ( .A(n38), .Q(n59) );
  NAND22 U95 ( .A(n108), .B(n89), .Q(n110) );
  INV3 U96 ( .A(B[0]), .Q(n80) );
  NOR21 U97 ( .A(B[0]), .B(n210), .Q(n81) );
  NAND20 U98 ( .A(n210), .B(B[0]), .Q(n222) );
  NAND20 U99 ( .A(n20), .B(n12), .Q(n18) );
  OAI2112 U100 ( .A(n85), .B(n86), .C(n87), .D(n88), .Q(n84) );
  AOI211 U101 ( .A(n68), .B(n69), .C(n70), .Q(n67) );
  NAND22 U102 ( .A(n192), .B(n21), .Q(n191) );
  NAND20 U103 ( .A(n21), .B(n12), .Q(n190) );
  NAND22 U104 ( .A(B[13]), .B(n156), .Q(n100) );
  CLKIN1 U105 ( .A(B[14]), .Q(n148) );
  INV3 U106 ( .A(n21), .Q(n180) );
  NAND21 U107 ( .A(n100), .B(n143), .Q(n142) );
  INV3 U108 ( .A(n1), .Q(n2) );
  INV6 U109 ( .A(n111), .Q(n89) );
  NAND20 U110 ( .A(n178), .B(n172), .Q(n186) );
  NAND21 U111 ( .A(n139), .B(n140), .Q(n137) );
  NOR21 U112 ( .A(A[3]), .B(n204), .Q(n213) );
  NAND22 U113 ( .A(B[14]), .B(n149), .Q(n92) );
  CLKIN2 U114 ( .A(n81), .Q(n78) );
  INV0 U115 ( .A(n19), .Q(n27) );
  NOR20 U116 ( .A(n180), .B(n16), .Q(n188) );
  NOR30 U117 ( .A(n16), .B(n180), .C(n181), .Q(n179) );
  INV6 U118 ( .A(B[4]), .Q(n65) );
  IMUX20 U119 ( .A(n23), .B(n24), .S(n25), .Q(DIFF[8]) );
  XOR20 U120 ( .A(B[8]), .B(A[8]), .Q(n23) );
  NOR20 U121 ( .A(A[8]), .B(n5), .Q(n26) );
  AOI210 U122 ( .A(n109), .B(n17), .C(n127), .Q(n153) );
  NAND20 U123 ( .A(n100), .B(n101), .Q(n150) );
  NAND20 U124 ( .A(n37), .B(n56), .Q(n57) );
  OAI2110 U125 ( .A(n16), .B(n17), .C(n18), .D(n19), .Q(n15) );
  NAND20 U126 ( .A(n35), .B(n33), .Q(n48) );
  NAND20 U127 ( .A(n34), .B(n35), .Q(n32) );
  INV0 U128 ( .A(n37), .Q(n52) );
  XNR20 U129 ( .A(B[11]), .B(A[11]), .Q(n3) );
  XOR20 U130 ( .A(B[12]), .B(A[12]), .Q(n158) );
  AOI210 U131 ( .A(B[12]), .B(n154), .C(n99), .Q(n157) );
  NAND20 U132 ( .A(n32), .B(n33), .Q(n31) );
  XNR20 U133 ( .A(B[15]), .B(A[15]), .Q(n4) );
  NOR20 U134 ( .A(A[0]), .B(n80), .Q(n79) );
  NOR23 U135 ( .A(n212), .B(n213), .Q(n211) );
  NAND22 U136 ( .A(A[8]), .B(n5), .Q(n19) );
  INV3 U137 ( .A(n172), .Q(n169) );
  NAND22 U138 ( .A(B[8]), .B(n8), .Q(n12) );
  XOR21 U139 ( .A(n186), .B(n187), .Q(DIFF[10]) );
  NOR21 U140 ( .A(n26), .B(n27), .Q(n24) );
  NAND22 U141 ( .A(n90), .B(n143), .Q(n146) );
  INV3 U142 ( .A(A[8]), .Q(n8) );
  INV3 U143 ( .A(A[10]), .Q(n9) );
  NAND22 U144 ( .A(B[12]), .B(n154), .Q(n143) );
  NAND22 U145 ( .A(n222), .B(n78), .Q(DIFF[0]) );
  NOR21 U146 ( .A(n129), .B(n130), .Q(n120) );
  NOR21 U147 ( .A(n46), .B(n124), .Q(n122) );
  NOR21 U148 ( .A(B[15]), .B(n95), .Q(n94) );
  INV3 U149 ( .A(n102), .Q(n91) );
  NAND22 U150 ( .A(n96), .B(n97), .Q(n93) );
  XOR21 U151 ( .A(n150), .B(n151), .Q(DIFF[13]) );
  XOR21 U152 ( .A(n57), .B(n58), .Q(DIFF[5]) );
  NAND22 U153 ( .A(n108), .B(n143), .Q(n127) );
  XOR21 U154 ( .A(n133), .B(n134), .Q(DIFF[14]) );
  NAND22 U155 ( .A(n92), .B(n96), .Q(n133) );
  NOR21 U156 ( .A(n135), .B(n136), .Q(n134) );
  NAND22 U157 ( .A(n144), .B(n101), .Q(n135) );
  NAND22 U158 ( .A(n137), .B(n138), .Q(n136) );
  XNR21 U159 ( .A(n71), .B(n68), .Q(DIFF[2]) );
  INV3 U160 ( .A(B[5]), .Q(n196) );
  NAND22 U161 ( .A(n145), .B(n100), .Q(n144) );
  XOR21 U162 ( .A(n48), .B(n49), .Q(DIFF[6]) );
  NOR21 U163 ( .A(n34), .B(n50), .Q(n49) );
  NAND22 U164 ( .A(n38), .B(n39), .Q(n29) );
  NAND22 U165 ( .A(n92), .B(n100), .Q(n132) );
  NOR22 U166 ( .A(n46), .B(n47), .Q(n107) );
  XOR21 U167 ( .A(n76), .B(n73), .Q(DIFF[1]) );
  INV3 U168 ( .A(A[4]), .Q(n60) );
  INV3 U169 ( .A(A[2]), .Q(n214) );
  INV3 U170 ( .A(A[13]), .Q(n156) );
  NAND22 U171 ( .A(B[6]), .B(n221), .Q(n35) );
  INV3 U172 ( .A(A[6]), .Q(n221) );
  NOR23 U173 ( .A(A[0]), .B(n80), .Q(n212) );
  INV3 U174 ( .A(A[14]), .Q(n149) );
  NAND22 U175 ( .A(A[14]), .B(n148), .Q(n96) );
  NAND22 U176 ( .A(A[6]), .B(n199), .Q(n33) );
  INV3 U177 ( .A(B[6]), .Q(n199) );
  NAND22 U178 ( .A(B[5]), .B(n220), .Q(n37) );
  INV3 U179 ( .A(A[5]), .Q(n220) );
  INV3 U180 ( .A(A[9]), .Q(n216) );
  XNR21 U181 ( .A(n176), .B(n3), .Q(DIFF[11]) );
  NOR21 U182 ( .A(A[5]), .B(n196), .Q(n198) );
  NAND22 U183 ( .A(A[2]), .B(n206), .Q(n75) );
  INV3 U184 ( .A(A[7]), .Q(n197) );
  IMUX21 U185 ( .A(n157), .B(n158), .S(n159), .Q(DIFF[12]) );
  IMUX21 U186 ( .A(n61), .B(n62), .S(n63), .Q(DIFF[4]) );
  NOR21 U187 ( .A(n64), .B(n59), .Q(n61) );
  NAND22 U188 ( .A(A[1]), .B(n205), .Q(n74) );
  NAND22 U189 ( .A(n78), .B(n79), .Q(n77) );
  NOR21 U190 ( .A(n52), .B(n36), .Q(n30) );
  NAND22 U191 ( .A(B[1]), .B(n215), .Q(n82) );
  INV3 U192 ( .A(A[1]), .Q(n215) );
  XNR21 U193 ( .A(n66), .B(n67), .Q(DIFF[3]) );
  NOR21 U194 ( .A(A[10]), .B(n6), .Q(n165) );
  NAND22 U195 ( .A(A[13]), .B(n155), .Q(n101) );
  CLKIN3 U196 ( .A(B[13]), .Q(n155) );
  INV3 U197 ( .A(A[12]), .Q(n154) );
  INV3 U198 ( .A(A[15]), .Q(n95) );
  INV3 U199 ( .A(A[0]), .Q(n210) );
  INV3 U200 ( .A(A[11]), .Q(n173) );
  CLKIN6 U201 ( .A(n207), .Q(n46) );
  NAND21 U202 ( .A(A[3]), .B(n204), .Q(n207) );
  NAND20 U203 ( .A(B[10]), .B(n9), .Q(n178) );
  INV2 U204 ( .A(B[2]), .Q(n206) );
  NOR24 U205 ( .A(n83), .B(n84), .Q(DIFF[16]) );
  OAI222 U206 ( .A(n109), .B(n110), .C(n17), .D(n110), .Q(n83) );
  NAND20 U207 ( .A(B[4]), .B(n60), .Q(n42) );
  NAND20 U208 ( .A(n82), .B(n74), .Q(n76) );
  AOI221 U209 ( .A(B[7]), .B(n197), .C(n198), .D(n33), .Q(n194) );
  INV1 U210 ( .A(B[1]), .Q(n205) );
  NAND22 U211 ( .A(B[2]), .B(n214), .Q(n69) );
  NOR20 U212 ( .A(B[11]), .B(n173), .Q(n168) );
  NOR20 U213 ( .A(A[4]), .B(n65), .Q(n64) );
  XOR21 U214 ( .A(n10), .B(n11), .Q(DIFF[9]) );
  NOR21 U215 ( .A(n46), .B(n47), .Q(n55) );
  NOR21 U216 ( .A(n46), .B(n47), .Q(n43) );
  NOR21 U217 ( .A(n46), .B(n47), .Q(n185) );
  NOR22 U218 ( .A(n46), .B(n47), .Q(n200) );
  OAI212 U219 ( .A(n40), .B(n184), .C(n13), .Q(n183) );
  NOR20 U220 ( .A(n127), .B(n128), .Q(n152) );
  NAND20 U221 ( .A(n109), .B(n128), .Q(n125) );
  XNR20 U222 ( .A(B[3]), .B(A[3]), .Q(n66) );
  XOR20 U223 ( .A(B[4]), .B(A[4]), .Q(n62) );
  XOR31 U224 ( .A(B[7]), .B(A[7]), .C(n28), .Q(DIFF[7]) );
  CLKIN3 U225 ( .A(n56), .Q(n34) );
  OAI212 U226 ( .A(n72), .B(n73), .C(n74), .Q(n68) );
  CLKIN3 U227 ( .A(n77), .Q(n73) );
  OAI212 U228 ( .A(n98), .B(n99), .C(n100), .Q(n97) );
  CLKIN3 U229 ( .A(n101), .Q(n98) );
  NAND33 U230 ( .A(n92), .B(n100), .C(n112), .Q(n111) );
  AOI2112 U231 ( .A(n115), .B(n116), .C(n117), .D(n118), .Q(n114) );
  OAI212 U232 ( .A(n119), .B(n101), .C(n96), .Q(n118) );
  CLKIN3 U233 ( .A(n92), .Q(n119) );
  CLKIN3 U234 ( .A(n132), .Q(n115) );
  OAI212 U235 ( .A(n168), .B(n169), .C(n164), .Q(n160) );
  OAI222 U236 ( .A(A[8]), .B(n5), .C(A[11]), .D(n171), .Q(n174) );
  CLKIN3 U237 ( .A(n178), .Q(n181) );
  CLKIN3 U238 ( .A(n74), .Q(n201) );
  OAI212 U239 ( .A(A[3]), .B(n204), .C(n70), .Q(n131) );
  CLKIN3 U240 ( .A(n75), .Q(n70) );
  CLKIN3 U241 ( .A(n12), .Q(n16) );
endmodule


module E_alu_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173;

  INV8 U3 ( .A(B[3]), .Q(n16) );
  NOR23 U4 ( .A(n7), .B(n32), .Q(n8) );
  INV8 U5 ( .A(B[4]), .Q(n17) );
  XOR21 U6 ( .A(n22), .B(n23), .Q(DIFF[9]) );
  INV6 U7 ( .A(n4), .Q(n60) );
  NAND22 U8 ( .A(n158), .B(n3), .Q(n4) );
  INV3 U9 ( .A(n143), .Q(n95) );
  NAND31 U10 ( .A(n37), .B(n44), .C(n144), .Q(n143) );
  NAND22 U11 ( .A(n41), .B(n42), .Q(n36) );
  XNR21 U12 ( .A(n115), .B(n11), .Q(DIFF[12]) );
  INV2 U13 ( .A(B[0]), .Q(n15) );
  INV3 U14 ( .A(n88), .Q(n160) );
  NOR24 U15 ( .A(A[3]), .B(n16), .Q(n155) );
  XNR21 U16 ( .A(n40), .B(n36), .Q(DIFF[6]) );
  NAND21 U17 ( .A(A[3]), .B(n16), .Q(n159) );
  NAND33 U18 ( .A(n153), .B(n65), .C(n154), .Q(n58) );
  INV2 U19 ( .A(n155), .Q(n154) );
  NOR21 U20 ( .A(n150), .B(n21), .Q(n149) );
  NAND23 U21 ( .A(n122), .B(n123), .Q(n109) );
  AOI211 U22 ( .A(A[11]), .B(n20), .C(n129), .Q(n122) );
  NAND22 U23 ( .A(n37), .B(n39), .Q(n40) );
  INV3 U24 ( .A(B[5]), .Q(n167) );
  NOR21 U25 ( .A(n43), .B(n47), .Q(n164) );
  NOR21 U26 ( .A(A[4]), .B(n17), .Q(n145) );
  NAND22 U27 ( .A(A[4]), .B(n17), .Q(n53) );
  NAND22 U28 ( .A(B[5]), .B(n147), .Q(n44) );
  INV6 U29 ( .A(n53), .Q(n43) );
  NAND24 U30 ( .A(n56), .B(n2), .Q(n46) );
  NAND23 U31 ( .A(n57), .B(n58), .Q(n1) );
  INV3 U32 ( .A(n15), .Q(n14) );
  AOI211 U33 ( .A(n64), .B(n65), .C(n66), .Q(n63) );
  NAND22 U34 ( .A(B[6]), .B(n168), .Q(n37) );
  NOR22 U35 ( .A(n8), .B(n106), .Q(n105) );
  INV3 U36 ( .A(n139), .Q(n26) );
  INV3 U37 ( .A(B[7]), .Q(n18) );
  INV3 U38 ( .A(n48), .Q(n47) );
  NAND22 U39 ( .A(n83), .B(n84), .Q(n82) );
  INV3 U40 ( .A(n56), .Q(n94) );
  XOR20 U41 ( .A(B[4]), .B(A[4]), .Q(n54) );
  INV1 U42 ( .A(B[10]), .Q(n172) );
  NAND21 U43 ( .A(n80), .B(n104), .Q(n106) );
  OAI211 U44 ( .A(n93), .B(n94), .C(n95), .Q(n89) );
  NAND24 U45 ( .A(n108), .B(n109), .Q(n80) );
  NOR23 U46 ( .A(n120), .B(n121), .Q(n119) );
  NAND32 U47 ( .A(n118), .B(n28), .C(n119), .Q(n117) );
  INV4 U48 ( .A(n117), .Q(n113) );
  INV6 U49 ( .A(n112), .Q(n91) );
  CLKIN2 U50 ( .A(n91), .Q(n7) );
  NOR24 U51 ( .A(n156), .B(n155), .Q(n3) );
  NOR24 U52 ( .A(A[11]), .B(n20), .Q(n120) );
  INV2 U53 ( .A(B[11]), .Q(n20) );
  AOI312 U54 ( .A(n87), .B(n88), .C(n89), .D(n90), .Q(n77) );
  XNR21 U55 ( .A(n68), .B(n64), .Q(DIFF[2]) );
  AOI212 U56 ( .A(n132), .B(n25), .C(n135), .Q(n137) );
  NAND28 U57 ( .A(n6), .B(n95), .Q(n141) );
  AOI222 U58 ( .A(n109), .B(n116), .C(n113), .D(n25), .Q(n115) );
  AOI312 U59 ( .A(n118), .B(n132), .C(n25), .D(n133), .Q(n131) );
  NAND22 U60 ( .A(n45), .B(n46), .Q(n52) );
  INV2 U61 ( .A(n25), .Q(n32) );
  XNR22 U62 ( .A(n131), .B(n9), .Q(DIFF[11]) );
  NAND22 U63 ( .A(n84), .B(n91), .Q(n90) );
  AOI311 U64 ( .A(n44), .B(n45), .C(n46), .D(n47), .Q(n41) );
  NAND21 U65 ( .A(n52), .B(n53), .Q(n51) );
  INV6 U66 ( .A(n1), .Q(n2) );
  NOR22 U67 ( .A(n59), .B(n60), .Q(n57) );
  NAND33 U68 ( .A(n148), .B(n65), .C(n149), .Q(n56) );
  INV2 U69 ( .A(B[2]), .Q(n158) );
  NAND23 U70 ( .A(n5), .B(n56), .Q(n6) );
  CLKIN3 U71 ( .A(n142), .Q(n5) );
  NAND28 U72 ( .A(n140), .B(n141), .Q(n25) );
  NAND21 U73 ( .A(n65), .B(n67), .Q(n68) );
  NAND22 U74 ( .A(B[2]), .B(n156), .Q(n65) );
  XNR22 U75 ( .A(n105), .B(n10), .Q(DIFF[13]) );
  NOR21 U76 ( .A(n59), .B(n60), .Q(n152) );
  INV3 U77 ( .A(n111), .Q(n114) );
  NAND22 U78 ( .A(B[10]), .B(n173), .Q(n118) );
  INV0 U79 ( .A(n97), .Q(n87) );
  INV2 U80 ( .A(n104), .Q(n86) );
  NOR21 U81 ( .A(n145), .B(n146), .Q(n144) );
  INV2 U82 ( .A(B[14]), .Q(n85) );
  NAND21 U83 ( .A(n96), .B(n58), .Q(n93) );
  NOR21 U84 ( .A(n110), .B(n111), .Q(n108) );
  NAND22 U85 ( .A(B[9]), .B(n171), .Q(n28) );
  NAND20 U86 ( .A(A[12]), .B(n107), .Q(n104) );
  INV2 U87 ( .A(n169), .Q(n162) );
  INV2 U88 ( .A(n73), .Q(n72) );
  NOR20 U89 ( .A(A[4]), .B(n17), .Q(n49) );
  NOR20 U90 ( .A(A[8]), .B(n19), .Q(n27) );
  NOR20 U91 ( .A(A[11]), .B(n20), .Q(n110) );
  NAND20 U92 ( .A(A[8]), .B(n19), .Q(n139) );
  NOR20 U93 ( .A(A[4]), .B(n17), .Q(n61) );
  NOR20 U94 ( .A(n59), .B(n60), .Q(n96) );
  IMUX20 U95 ( .A(n54), .B(n55), .S(n46), .Q(DIFF[4]) );
  NOR20 U96 ( .A(A[8]), .B(n19), .Q(n33) );
  NOR23 U97 ( .A(n160), .B(n97), .Q(n140) );
  NOR20 U98 ( .A(B[13]), .B(n103), .Q(n83) );
  XNR20 U99 ( .A(B[11]), .B(A[11]), .Q(n9) );
  NAND22 U100 ( .A(B[13]), .B(n103), .Q(n92) );
  XOR20 U101 ( .A(n71), .B(n72), .Q(DIFF[1]) );
  NAND20 U102 ( .A(n74), .B(n70), .Q(n71) );
  NAND20 U103 ( .A(n118), .B(n130), .Q(n136) );
  NAND20 U104 ( .A(n43), .B(n44), .Q(n42) );
  NAND20 U105 ( .A(n44), .B(n48), .Q(n50) );
  INV0 U106 ( .A(n67), .Q(n66) );
  INV2 U107 ( .A(B[6]), .Q(n166) );
  XNR20 U108 ( .A(B[14]), .B(A[14]), .Q(n13) );
  XNR20 U109 ( .A(B[13]), .B(A[13]), .Q(n10) );
  XNR20 U110 ( .A(B[12]), .B(A[12]), .Q(n11) );
  NOR20 U111 ( .A(A[7]), .B(n18), .Q(n169) );
  NOR21 U112 ( .A(n14), .B(n21), .Q(n73) );
  MUX22 U113 ( .A(B[0]), .B(n15), .S(n21), .Q(DIFF[0]) );
  INV3 U114 ( .A(n61), .Q(n45) );
  NOR21 U115 ( .A(n49), .B(n43), .Q(n55) );
  NOR21 U116 ( .A(A[8]), .B(n19), .Q(n121) );
  INV3 U117 ( .A(B[12]), .Q(n107) );
  INV3 U118 ( .A(B[9]), .Q(n128) );
  NAND22 U119 ( .A(n86), .B(n92), .Q(n101) );
  INV3 U120 ( .A(n83), .Q(n102) );
  INV3 U121 ( .A(A[0]), .Q(n21) );
  XNR21 U122 ( .A(n75), .B(n76), .Q(DIFF[15]) );
  XNR21 U123 ( .A(B[15]), .B(A[15]), .Q(n75) );
  NAND22 U124 ( .A(n152), .B(n58), .Q(n142) );
  NOR21 U125 ( .A(n14), .B(n69), .Q(n148) );
  NOR21 U126 ( .A(A[3]), .B(n16), .Q(n150) );
  XNR21 U127 ( .A(n62), .B(n63), .Q(DIFF[3]) );
  NAND22 U128 ( .A(n113), .B(n114), .Q(n112) );
  NAND22 U129 ( .A(n138), .B(n29), .Q(n135) );
  NAND22 U130 ( .A(n26), .B(n28), .Q(n138) );
  XOR21 U131 ( .A(n136), .B(n137), .Q(DIFF[10]) );
  XNR21 U132 ( .A(n50), .B(n51), .Q(DIFF[5]) );
  NAND22 U133 ( .A(n134), .B(n130), .Q(n133) );
  NAND22 U134 ( .A(n28), .B(n29), .Q(n22) );
  AOI211 U135 ( .A(n24), .B(n25), .C(n26), .Q(n23) );
  INV3 U136 ( .A(n27), .Q(n24) );
  IMUX21 U137 ( .A(n30), .B(n31), .S(n32), .Q(DIFF[8]) );
  XOR21 U138 ( .A(B[8]), .B(A[8]), .Q(n31) );
  NOR21 U139 ( .A(n33), .B(n26), .Q(n30) );
  NOR21 U140 ( .A(n27), .B(n170), .Q(n132) );
  NOR22 U141 ( .A(n77), .B(n78), .Q(n76) );
  OAI2111 U142 ( .A(n79), .B(n80), .C(n81), .D(n82), .Q(n78) );
  INV3 U143 ( .A(B[8]), .Q(n19) );
  NAND22 U144 ( .A(n135), .B(n118), .Q(n134) );
  NOR21 U145 ( .A(A[7]), .B(n18), .Q(n146) );
  AOI221 U146 ( .A(A[14]), .B(n85), .C(n86), .D(n84), .Q(n81) );
  NOR21 U147 ( .A(A[12]), .B(n107), .Q(n111) );
  NAND22 U148 ( .A(A[9]), .B(n128), .Q(n29) );
  NAND22 U149 ( .A(A[10]), .B(n172), .Q(n130) );
  NAND22 U150 ( .A(A[5]), .B(n167), .Q(n48) );
  NAND22 U151 ( .A(A[2]), .B(n158), .Q(n67) );
  NAND22 U152 ( .A(A[1]), .B(n157), .Q(n70) );
  INV3 U153 ( .A(B[1]), .Q(n157) );
  INV3 U154 ( .A(A[10]), .Q(n173) );
  NAND22 U155 ( .A(A[6]), .B(n166), .Q(n39) );
  INV3 U156 ( .A(A[5]), .Q(n147) );
  XNR21 U157 ( .A(n98), .B(n13), .Q(DIFF[14]) );
  INV3 U158 ( .A(A[9]), .Q(n171) );
  INV3 U159 ( .A(A[2]), .Q(n156) );
  INV3 U160 ( .A(A[6]), .Q(n168) );
  NOR21 U161 ( .A(B[7]), .B(n161), .Q(n97) );
  INV3 U162 ( .A(A[7]), .Q(n161) );
  XNR21 U163 ( .A(n34), .B(n35), .Q(DIFF[7]) );
  XNR21 U164 ( .A(B[7]), .B(A[7]), .Q(n34) );
  AOI211 U165 ( .A(n36), .B(n37), .C(n38), .Q(n35) );
  NAND22 U166 ( .A(B[1]), .B(n151), .Q(n74) );
  INV3 U167 ( .A(A[1]), .Q(n151) );
  NAND22 U168 ( .A(n162), .B(n163), .Q(n88) );
  INV3 U169 ( .A(n110), .Q(n116) );
  NOR21 U170 ( .A(n126), .B(n127), .Q(n125) );
  NOR21 U171 ( .A(A[9]), .B(n128), .Q(n126) );
  INV3 U172 ( .A(A[13]), .Q(n103) );
  XNR20 U173 ( .A(B[3]), .B(A[3]), .Q(n62) );
  CLKIN3 U174 ( .A(n39), .Q(n38) );
  OAI212 U175 ( .A(n69), .B(n72), .C(n70), .Q(n64) );
  CLKIN3 U176 ( .A(n79), .Q(n84) );
  OAI212 U177 ( .A(A[14]), .B(n85), .C(n92), .Q(n79) );
  AOI312 U178 ( .A(n92), .B(n91), .C(n25), .D(n99), .Q(n98) );
  OAI2112 U179 ( .A(n100), .B(n80), .C(n101), .D(n102), .Q(n99) );
  CLKIN3 U180 ( .A(n92), .Q(n100) );
  OAI212 U181 ( .A(n124), .B(n26), .C(n125), .Q(n123) );
  CLKIN3 U182 ( .A(n118), .Q(n127) );
  CLKIN3 U183 ( .A(n29), .Q(n124) );
  CLKIN3 U184 ( .A(n130), .Q(n129) );
  CLKIN3 U185 ( .A(n74), .Q(n69) );
  CLKIN3 U186 ( .A(n70), .Q(n153) );
  CLKIN3 U187 ( .A(n159), .Q(n59) );
  OAI212 U188 ( .A(n164), .B(n165), .C(n39), .Q(n163) );
  OAI212 U189 ( .A(A[5]), .B(n167), .C(n37), .Q(n165) );
  CLKIN3 U190 ( .A(n28), .Q(n170) );
endmodule


module E_alu_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178;

  CLKIN6 U3 ( .A(n143), .Q(n94) );
  NAND23 U4 ( .A(n164), .B(n165), .Q(n86) );
  CLKIN0 U5 ( .A(n21), .Q(n28) );
  NAND23 U6 ( .A(A[4]), .B(n13), .Q(n47) );
  NAND24 U7 ( .A(n37), .B(n38), .Q(n32) );
  NAND24 U8 ( .A(n154), .B(n53), .Q(n142) );
  INV8 U9 ( .A(B[3]), .Q(n12) );
  NOR22 U10 ( .A(n39), .B(n171), .Q(n166) );
  NOR22 U11 ( .A(A[11]), .B(n16), .Q(n120) );
  CLKIN3 U12 ( .A(n131), .Q(n2) );
  NAND22 U13 ( .A(B[2]), .B(n158), .Q(n60) );
  NOR22 U14 ( .A(n75), .B(n76), .Q(n74) );
  CLKIN6 U15 ( .A(n47), .Q(n39) );
  NOR24 U16 ( .A(A[3]), .B(n12), .Q(n157) );
  CLKIN4 U17 ( .A(B[4]), .Q(n13) );
  NOR22 U18 ( .A(A[8]), .B(n15), .Q(n121) );
  INV2 U19 ( .A(B[5]), .Q(n169) );
  NOR22 U20 ( .A(n148), .B(n149), .Q(n147) );
  NAND22 U21 ( .A(A[10]), .B(n175), .Q(n130) );
  NAND23 U22 ( .A(B[10]), .B(n176), .Q(n118) );
  INV3 U23 ( .A(n8), .Q(n3) );
  NOR22 U24 ( .A(n43), .B(n145), .Q(n144) );
  INV3 U25 ( .A(n110), .Q(n116) );
  NAND22 U26 ( .A(n33), .B(n35), .Q(n36) );
  INV3 U27 ( .A(n118), .Q(n127) );
  NOR21 U28 ( .A(A[4]), .B(n13), .Q(n43) );
  NOR21 U29 ( .A(A[12]), .B(n107), .Q(n111) );
  NAND22 U30 ( .A(A[2]), .B(n160), .Q(n62) );
  NAND23 U31 ( .A(B[6]), .B(n170), .Q(n33) );
  NAND22 U32 ( .A(B[9]), .B(n174), .Q(n24) );
  NAND22 U33 ( .A(n4), .B(n5), .Q(DIFF[11]) );
  NAND22 U34 ( .A(n1), .B(n8), .Q(n4) );
  NAND22 U35 ( .A(n2), .B(n3), .Q(n5) );
  NAND22 U36 ( .A(n138), .B(n25), .Q(n135) );
  INV3 U37 ( .A(n72), .Q(n64) );
  AOI211 U38 ( .A(n59), .B(n60), .C(n61), .Q(n58) );
  NAND28 U39 ( .A(n140), .B(n141), .Q(n21) );
  AOI312 U40 ( .A(n118), .B(n132), .C(n21), .D(n133), .Q(n1) );
  AOI212 U41 ( .A(n20), .B(n21), .C(n22), .Q(n19) );
  CLKIN6 U42 ( .A(n66), .Q(n155) );
  NAND21 U43 ( .A(n46), .B(n47), .Q(n45) );
  CLKIN4 U44 ( .A(B[2]), .Q(n160) );
  NAND21 U45 ( .A(n95), .B(n53), .Q(n91) );
  NOR22 U46 ( .A(A[0]), .B(n11), .Q(n148) );
  INV6 U47 ( .A(B[0]), .Q(n11) );
  NAND32 U48 ( .A(n72), .B(n60), .C(n147), .Q(n51) );
  NAND33 U49 ( .A(n33), .B(n40), .C(n144), .Q(n143) );
  INV6 U50 ( .A(n51), .Q(n93) );
  XNR21 U51 ( .A(n36), .B(n32), .Q(DIFF[6]) );
  NOR24 U52 ( .A(n162), .B(n96), .Q(n140) );
  CLKIN6 U53 ( .A(n86), .Q(n162) );
  NOR22 U54 ( .A(n54), .B(n55), .Q(n154) );
  INV6 U55 ( .A(n52), .Q(n92) );
  NAND24 U56 ( .A(n52), .B(n95), .Q(n6) );
  NAND22 U57 ( .A(B[1]), .B(n153), .Q(n72) );
  INV6 U58 ( .A(B[8]), .Q(n15) );
  NAND22 U59 ( .A(A[8]), .B(n15), .Q(n139) );
  NOR23 U60 ( .A(A[7]), .B(n14), .Q(n145) );
  NAND22 U61 ( .A(A[3]), .B(n12), .Q(n161) );
  NAND33 U62 ( .A(n150), .B(n60), .C(n151), .Q(n52) );
  NOR22 U63 ( .A(n152), .B(n17), .Q(n151) );
  NAND21 U64 ( .A(n135), .B(n118), .Q(n134) );
  NAND33 U65 ( .A(n118), .B(n24), .C(n119), .Q(n117) );
  INV1 U66 ( .A(B[10]), .Q(n175) );
  INV3 U67 ( .A(B[14]), .Q(n83) );
  INV2 U68 ( .A(B[6]), .Q(n168) );
  INV2 U69 ( .A(B[11]), .Q(n16) );
  INV2 U70 ( .A(B[12]), .Q(n107) );
  NAND33 U71 ( .A(n53), .B(n51), .C(n7), .Q(n41) );
  INV6 U72 ( .A(n6), .Q(n7) );
  NAND34 U73 ( .A(n155), .B(n60), .C(n156), .Q(n53) );
  IMUX21 U74 ( .A(n49), .B(n50), .S(n41), .Q(DIFF[4]) );
  NAND21 U75 ( .A(n48), .B(n41), .Q(n46) );
  NOR23 U76 ( .A(n54), .B(n55), .Q(n95) );
  INV0 U77 ( .A(n62), .Q(n61) );
  NAND20 U78 ( .A(n60), .B(n62), .Q(n63) );
  NOR24 U79 ( .A(n157), .B(n62), .Q(n55) );
  NAND22 U80 ( .A(B[5]), .B(n146), .Q(n40) );
  NAND22 U81 ( .A(n84), .B(n90), .Q(n100) );
  INV1 U82 ( .A(n96), .Q(n85) );
  INV1 U83 ( .A(B[1]), .Q(n159) );
  NAND21 U84 ( .A(A[12]), .B(n107), .Q(n103) );
  NAND22 U85 ( .A(A[5]), .B(n169), .Q(n42) );
  NAND21 U86 ( .A(n81), .B(n82), .Q(n80) );
  OAI2111 U87 ( .A(n77), .B(n78), .C(n79), .D(n80), .Q(n76) );
  INV1 U88 ( .A(n43), .Q(n48) );
  OAI310 U89 ( .A(n91), .B(n92), .C(n93), .D(n94), .Q(n87) );
  XOR20 U90 ( .A(B[4]), .B(A[4]), .Q(n49) );
  NOR20 U91 ( .A(A[4]), .B(n13), .Q(n56) );
  INV2 U92 ( .A(n11), .Q(n178) );
  INV2 U93 ( .A(n71), .Q(n69) );
  NOR20 U94 ( .A(A[0]), .B(n11), .Q(n70) );
  NOR20 U95 ( .A(A[8]), .B(n15), .Q(n29) );
  NOR20 U96 ( .A(B[13]), .B(n102), .Q(n81) );
  XOR20 U97 ( .A(n67), .B(n65), .Q(DIFF[1]) );
  NAND20 U98 ( .A(n72), .B(n66), .Q(n67) );
  NAND20 U99 ( .A(n118), .B(n130), .Q(n136) );
  XNR20 U100 ( .A(B[11]), .B(A[11]), .Q(n8) );
  CLKIN3 U101 ( .A(n23), .Q(n20) );
  XNR20 U102 ( .A(n63), .B(n59), .Q(DIFF[2]) );
  CLKIN2 U103 ( .A(B[7]), .Q(n14) );
  AOI212 U104 ( .A(A[11]), .B(n16), .C(n129), .Q(n122) );
  XOR20 U105 ( .A(B[13]), .B(A[13]), .Q(n105) );
  XNR20 U106 ( .A(B[14]), .B(A[14]), .Q(n9) );
  XNR20 U107 ( .A(B[12]), .B(A[12]), .Q(n10) );
  NOR21 U108 ( .A(n178), .B(n17), .Q(n71) );
  NAND22 U109 ( .A(n177), .B(n69), .Q(DIFF[0]) );
  NAND22 U110 ( .A(n17), .B(n178), .Q(n177) );
  XNR21 U111 ( .A(n57), .B(n58), .Q(DIFF[3]) );
  NOR21 U112 ( .A(A[8]), .B(n15), .Q(n23) );
  NAND22 U113 ( .A(n69), .B(n70), .Q(n68) );
  NOR21 U114 ( .A(A[11]), .B(n16), .Q(n110) );
  NOR21 U115 ( .A(n56), .B(n39), .Q(n50) );
  INV3 U116 ( .A(B[9]), .Q(n128) );
  NAND22 U117 ( .A(n82), .B(n89), .Q(n88) );
  INV3 U118 ( .A(n81), .Q(n101) );
  INV3 U119 ( .A(A[0]), .Q(n17) );
  INV3 U120 ( .A(n157), .Q(n156) );
  NOR21 U121 ( .A(A[3]), .B(n12), .Q(n149) );
  NAND22 U122 ( .A(B[13]), .B(n102), .Q(n90) );
  NOR22 U123 ( .A(n178), .B(n64), .Q(n150) );
  NOR21 U124 ( .A(A[3]), .B(n12), .Q(n152) );
  AOI211 U125 ( .A(n89), .B(n21), .C(n106), .Q(n104) );
  NAND22 U126 ( .A(n78), .B(n103), .Q(n106) );
  NAND22 U127 ( .A(n113), .B(n114), .Q(n112) );
  INV3 U128 ( .A(n111), .Q(n114) );
  NAND22 U129 ( .A(n108), .B(n109), .Q(n78) );
  NOR21 U130 ( .A(n110), .B(n111), .Q(n108) );
  NAND22 U131 ( .A(n22), .B(n24), .Q(n138) );
  NAND22 U132 ( .A(n122), .B(n123), .Q(n109) );
  NOR22 U133 ( .A(n120), .B(n121), .Q(n119) );
  XOR21 U134 ( .A(n136), .B(n137), .Q(DIFF[10]) );
  NAND22 U135 ( .A(n134), .B(n130), .Q(n133) );
  XOR21 U136 ( .A(n18), .B(n19), .Q(DIFF[9]) );
  NAND22 U137 ( .A(n24), .B(n25), .Q(n18) );
  IMUX21 U138 ( .A(n26), .B(n27), .S(n28), .Q(DIFF[8]) );
  XOR21 U139 ( .A(B[8]), .B(A[8]), .Q(n27) );
  NOR21 U140 ( .A(n29), .B(n22), .Q(n26) );
  XNR21 U141 ( .A(n73), .B(n74), .Q(DIFF[15]) );
  XNR21 U142 ( .A(B[15]), .B(A[15]), .Q(n73) );
  AOI311 U143 ( .A(n85), .B(n86), .C(n87), .D(n88), .Q(n75) );
  AOI311 U144 ( .A(n40), .B(n48), .C(n41), .D(n171), .Q(n37) );
  XNR21 U145 ( .A(n44), .B(n45), .Q(DIFF[5]) );
  NAND22 U146 ( .A(n40), .B(n42), .Q(n44) );
  NOR21 U147 ( .A(n23), .B(n173), .Q(n132) );
  INV3 U148 ( .A(n42), .Q(n171) );
  NAND22 U149 ( .A(A[9]), .B(n128), .Q(n25) );
  AOI221 U150 ( .A(A[14]), .B(n83), .C(n84), .D(n82), .Q(n79) );
  NAND22 U151 ( .A(A[1]), .B(n159), .Q(n66) );
  INV3 U152 ( .A(A[10]), .Q(n176) );
  INV3 U153 ( .A(A[2]), .Q(n158) );
  NAND22 U154 ( .A(A[6]), .B(n168), .Q(n35) );
  INV3 U155 ( .A(A[9]), .Q(n174) );
  INV3 U156 ( .A(A[5]), .Q(n146) );
  INV3 U157 ( .A(A[6]), .Q(n170) );
  NOR21 U158 ( .A(B[7]), .B(n163), .Q(n96) );
  INV3 U159 ( .A(A[7]), .Q(n163) );
  INV3 U160 ( .A(A[1]), .Q(n153) );
  INV3 U161 ( .A(n172), .Q(n164) );
  NOR21 U162 ( .A(A[7]), .B(n14), .Q(n172) );
  XNR21 U163 ( .A(n97), .B(n9), .Q(DIFF[14]) );
  XOR21 U164 ( .A(n104), .B(n105), .Q(DIFF[13]) );
  XNR21 U165 ( .A(n115), .B(n10), .Q(DIFF[12]) );
  NOR21 U166 ( .A(n126), .B(n127), .Q(n125) );
  NOR21 U167 ( .A(A[9]), .B(n128), .Q(n126) );
  XNR21 U168 ( .A(n30), .B(n31), .Q(DIFF[7]) );
  XNR21 U169 ( .A(B[7]), .B(A[7]), .Q(n30) );
  AOI211 U170 ( .A(n32), .B(n33), .C(n34), .Q(n31) );
  INV3 U171 ( .A(A[13]), .Q(n102) );
  NAND22 U172 ( .A(n39), .B(n40), .Q(n38) );
  XNR20 U173 ( .A(B[3]), .B(A[3]), .Q(n57) );
  CLKIN3 U174 ( .A(n35), .Q(n34) );
  OAI212 U175 ( .A(n64), .B(n65), .C(n66), .Q(n59) );
  CLKIN3 U176 ( .A(n68), .Q(n65) );
  CLKIN3 U177 ( .A(n77), .Q(n82) );
  OAI212 U178 ( .A(A[14]), .B(n83), .C(n90), .Q(n77) );
  AOI312 U179 ( .A(n90), .B(n89), .C(n21), .D(n98), .Q(n97) );
  OAI2112 U180 ( .A(n99), .B(n78), .C(n100), .D(n101), .Q(n98) );
  CLKIN3 U181 ( .A(n103), .Q(n84) );
  CLKIN3 U182 ( .A(n90), .Q(n99) );
  CLKIN3 U183 ( .A(n112), .Q(n89) );
  AOI222 U184 ( .A(n109), .B(n116), .C(n113), .D(n21), .Q(n115) );
  CLKIN3 U185 ( .A(n117), .Q(n113) );
  OAI212 U186 ( .A(n124), .B(n22), .C(n125), .Q(n123) );
  CLKIN3 U187 ( .A(n25), .Q(n124) );
  CLKIN3 U188 ( .A(n130), .Q(n129) );
  AOI312 U189 ( .A(n118), .B(n132), .C(n21), .D(n133), .Q(n131) );
  AOI212 U190 ( .A(n132), .B(n21), .C(n135), .Q(n137) );
  CLKIN3 U191 ( .A(n139), .Q(n22) );
  OAI312 U192 ( .A(n142), .B(n92), .C(n93), .D(n94), .Q(n141) );
  CLKIN3 U193 ( .A(n161), .Q(n54) );
  OAI212 U194 ( .A(n166), .B(n167), .C(n35), .Q(n165) );
  OAI212 U195 ( .A(A[5]), .B(n169), .C(n33), .Q(n167) );
  CLKIN3 U196 ( .A(n24), .Q(n173) );
endmodule


module E_alu_DW01_add_8 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  INV6 U2 ( .A(n20), .Q(n13) );
  NAND33 U3 ( .A(n26), .B(n27), .C(n28), .Q(n12) );
  NOR24 U4 ( .A(n7), .B(n8), .Q(n67) );
  BUF15 U5 ( .A(B[2]), .Q(n7) );
  NAND28 U6 ( .A(n11), .B(n10), .Q(SUM[8]) );
  NAND33 U7 ( .A(n21), .B(n22), .C(n59), .Q(n20) );
  NOR32 U8 ( .A(n65), .B(n66), .C(n67), .Q(n64) );
  NAND24 U9 ( .A(n54), .B(n55), .Q(n39) );
  NOR23 U10 ( .A(n23), .B(n66), .Q(n59) );
  NOR24 U11 ( .A(A[1]), .B(B[1]), .Q(n23) );
  NOR24 U12 ( .A(A[3]), .B(B[3]), .Q(n66) );
  NOR23 U13 ( .A(n16), .B(n17), .Q(n15) );
  OAI2112 U14 ( .A(n18), .B(n36), .C(n37), .D(n38), .Q(n30) );
  INV3 U15 ( .A(n70), .Q(n1) );
  OAI2111 U16 ( .A(n48), .B(n49), .C(n50), .D(n39), .Q(n47) );
  NAND22 U17 ( .A(n3), .B(n4), .Q(SUM[3]) );
  NAND22 U18 ( .A(n1), .B(n71), .Q(n4) );
  NOR21 U19 ( .A(n18), .B(n19), .Q(n14) );
  INV6 U20 ( .A(B[0]), .Q(n82) );
  NAND22 U21 ( .A(n72), .B(n73), .Q(n70) );
  NAND22 U22 ( .A(n58), .B(n6), .Q(n49) );
  AOI211 U23 ( .A(n59), .B(n60), .C(n61), .Q(n58) );
  NOR21 U24 ( .A(B[4]), .B(A[4]), .Q(n19) );
  INV6 U25 ( .A(n64), .Q(n28) );
  NAND23 U26 ( .A(A[1]), .B(B[1]), .Q(n65) );
  NAND21 U27 ( .A(B[0]), .B(A[0]), .Q(n63) );
  NAND21 U28 ( .A(n70), .B(n2), .Q(n3) );
  INV0 U29 ( .A(n71), .Q(n2) );
  NAND21 U30 ( .A(A[4]), .B(B[4]), .Q(n36) );
  NAND22 U31 ( .A(n28), .B(n26), .Q(n5) );
  OAI2111 U32 ( .A(A[3]), .B(B[3]), .C(n9), .D(n7), .Q(n26) );
  INV2 U33 ( .A(n5), .Q(n6) );
  INV4 U34 ( .A(B[5]), .Q(n54) );
  IMUX20 U35 ( .A(n56), .B(n57), .S(n49), .Q(SUM[4]) );
  AOI210 U36 ( .A(n50), .B(n49), .C(n48), .Q(n52) );
  CLKIN1 U37 ( .A(n63), .Q(n78) );
  NAND22 U38 ( .A(n47), .B(n38), .Q(n42) );
  NOR20 U39 ( .A(n43), .B(n16), .Q(n44) );
  OAI2112 U40 ( .A(n12), .B(n13), .C(n14), .D(n15), .Q(n11) );
  NOR20 U41 ( .A(n7), .B(n8), .Q(n62) );
  NAND20 U42 ( .A(n39), .B(n38), .Q(n51) );
  NAND20 U43 ( .A(n7), .B(n9), .Q(n72) );
  INV0 U44 ( .A(n37), .Q(n43) );
  CLKIN3 U45 ( .A(n35), .Q(n31) );
  XNR21 U46 ( .A(n74), .B(n75), .Q(SUM[2]) );
  XOR21 U47 ( .A(n42), .B(n44), .Q(SUM[6]) );
  NAND22 U48 ( .A(n76), .B(n77), .Q(n74) );
  NAND22 U49 ( .A(n78), .B(n79), .Q(n77) );
  XOR21 U50 ( .A(n51), .B(n52), .Q(SUM[5]) );
  NOR21 U51 ( .A(n7), .B(n8), .Q(n24) );
  INV3 U52 ( .A(n39), .Q(n18) );
  NAND22 U53 ( .A(n22), .B(n74), .Q(n73) );
  XOR21 U54 ( .A(n78), .B(n80), .Q(SUM[1]) );
  INV3 U55 ( .A(n24), .Q(n22) );
  NAND22 U56 ( .A(B[5]), .B(A[5]), .Q(n38) );
  NAND22 U57 ( .A(n45), .B(n46), .Q(n29) );
  INV3 U58 ( .A(A[6]), .Q(n46) );
  INV3 U59 ( .A(B[6]), .Q(n45) );
  AOI211 U60 ( .A(n42), .B(n29), .C(n43), .Q(n41) );
  NOR21 U61 ( .A(n68), .B(n48), .Q(n57) );
  INV3 U62 ( .A(n53), .Q(n50) );
  INV3 U63 ( .A(A[5]), .Q(n55) );
  INV3 U64 ( .A(n84), .Q(n83) );
  INV3 U65 ( .A(A[0]), .Q(n25) );
  INV3 U66 ( .A(A[7]), .Q(n33) );
  BUF2 U67 ( .A(A[2]), .Q(n8) );
  BUF2 U68 ( .A(A[2]), .Q(n9) );
  NAND20 U69 ( .A(B[4]), .B(A[4]), .Q(n69) );
  XNR20 U70 ( .A(B[7]), .B(A[7]), .Q(n40) );
  CLKIN1 U71 ( .A(B[7]), .Q(n34) );
  NOR20 U72 ( .A(n81), .B(n23), .Q(n80) );
  CLKIN0 U73 ( .A(n23), .Q(n79) );
  NOR21 U74 ( .A(A[7]), .B(B[7]), .Q(n35) );
  NOR21 U75 ( .A(B[7]), .B(A[7]), .Q(n17) );
  NOR21 U76 ( .A(n25), .B(n82), .Q(n21) );
  NOR21 U77 ( .A(n62), .B(n63), .Q(n60) );
  XOR21 U78 ( .A(n40), .B(n41), .Q(SUM[7]) );
  NOR21 U79 ( .A(n33), .B(n34), .Q(n32) );
  NAND20 U80 ( .A(B[1]), .B(A[1]), .Q(n76) );
  NAND21 U81 ( .A(B[3]), .B(A[3]), .Q(n27) );
  NOR20 U82 ( .A(B[4]), .B(A[4]), .Q(n68) );
  NOR20 U83 ( .A(A[4]), .B(B[4]), .Q(n53) );
  NAND22 U84 ( .A(B[6]), .B(A[6]), .Q(n37) );
  XOR20 U85 ( .A(B[3]), .B(A[3]), .Q(n71) );
  NOR20 U86 ( .A(B[0]), .B(n25), .Q(n84) );
  XNR20 U87 ( .A(B[4]), .B(A[4]), .Q(n56) );
  AOI312 U88 ( .A(n29), .B(n30), .C(n31), .D(n32), .Q(n10) );
  CLKIN3 U89 ( .A(n29), .Q(n16) );
  CLKIN3 U90 ( .A(n27), .Q(n61) );
  CLKIN3 U91 ( .A(n69), .Q(n48) );
  OAI212 U92 ( .A(n7), .B(n9), .C(n72), .Q(n75) );
  CLKIN3 U93 ( .A(n76), .Q(n81) );
  OAI212 U94 ( .A(A[0]), .B(n82), .C(n83), .Q(SUM[0]) );
endmodule


module E_alu_DW01_add_7 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97;

  CLKIN3 U2 ( .A(n36), .Q(n80) );
  INV6 U3 ( .A(n21), .Q(n1) );
  NOR21 U4 ( .A(n36), .B(n37), .Q(n35) );
  NAND42 U5 ( .A(A[1]), .B(B[1]), .C(n79), .D(n80), .Q(n39) );
  INV8 U6 ( .A(n9), .Q(n8) );
  NAND23 U7 ( .A(n32), .B(n33), .Q(n31) );
  INV3 U8 ( .A(n39), .Q(n77) );
  AOI212 U9 ( .A(n70), .B(n71), .C(n40), .Q(n69) );
  NOR20 U10 ( .A(n36), .B(n73), .Q(n71) );
  AOI212 U11 ( .A(n10), .B(n9), .C(n34), .Q(n70) );
  INV2 U12 ( .A(n34), .Q(n75) );
  NOR20 U13 ( .A(A[0]), .B(B[0]), .Q(n95) );
  NOR21 U14 ( .A(B[0]), .B(A[0]), .Q(n43) );
  NAND22 U15 ( .A(B[0]), .B(A[0]), .Q(n37) );
  NAND21 U16 ( .A(B[0]), .B(A[0]), .Q(n73) );
  NAND33 U17 ( .A(n67), .B(n68), .C(n69), .Q(n60) );
  INV8 U18 ( .A(B[2]), .Q(n9) );
  INV3 U19 ( .A(n35), .Q(n30) );
  INV3 U20 ( .A(n60), .Q(n54) );
  INV3 U21 ( .A(n51), .Q(n17) );
  NAND23 U22 ( .A(n54), .B(n55), .Q(n49) );
  NAND23 U23 ( .A(A[2]), .B(n8), .Q(n78) );
  NOR22 U24 ( .A(n8), .B(A[2]), .Q(n44) );
  NAND23 U25 ( .A(n56), .B(n57), .Q(n18) );
  NAND22 U26 ( .A(n63), .B(n64), .Q(n21) );
  INV3 U27 ( .A(n62), .Q(n48) );
  CLKIN6 U28 ( .A(n34), .Q(n33) );
  NAND24 U29 ( .A(n38), .B(n39), .Q(n28) );
  NOR21 U30 ( .A(n77), .B(n41), .Q(n67) );
  NOR23 U31 ( .A(n36), .B(n78), .Q(n41) );
  AOI311 U32 ( .A(n47), .B(n48), .C(n49), .D(n50), .Q(n46) );
  NOR21 U33 ( .A(B[3]), .B(A[3]), .Q(n42) );
  NOR22 U34 ( .A(n42), .B(n43), .Q(n74) );
  OAI210 U35 ( .A(n25), .B(n51), .C(n20), .Q(n50) );
  NAND20 U36 ( .A(B[1]), .B(A[1]), .Q(n89) );
  NAND21 U37 ( .A(n91), .B(n75), .Q(n90) );
  NOR22 U38 ( .A(n40), .B(n41), .Q(n38) );
  NOR22 U39 ( .A(n34), .B(n44), .Q(n27) );
  AOI211 U40 ( .A(n48), .B(n60), .C(n61), .Q(n59) );
  NAND22 U41 ( .A(B[4]), .B(A[4]), .Q(n55) );
  NAND21 U42 ( .A(B[0]), .B(A[0]), .Q(n94) );
  NOR24 U43 ( .A(A[3]), .B(B[3]), .Q(n36) );
  NAND22 U44 ( .A(B[3]), .B(A[3]), .Q(n72) );
  AOI2112 U45 ( .A(n27), .B(n74), .C(n28), .D(n29), .Q(n11) );
  NOR24 U46 ( .A(n30), .B(n31), .Q(n29) );
  OAI2112 U47 ( .A(n12), .B(n11), .C(n13), .D(n14), .Q(SUM[8]) );
  NOR32 U48 ( .A(n62), .B(n1), .C(n2), .Q(n3) );
  NOR22 U49 ( .A(n3), .B(n17), .Q(n53) );
  CLKIN2 U50 ( .A(n49), .Q(n2) );
  XOR22 U51 ( .A(n52), .B(n53), .Q(SUM[6]) );
  NOR20 U52 ( .A(n93), .B(n34), .Q(n92) );
  NOR24 U53 ( .A(A[1]), .B(B[1]), .Q(n34) );
  OAI312 U54 ( .A(n25), .B(n55), .C(n1), .D(n16), .Q(n15) );
  CLKIN3 U55 ( .A(B[6]), .Q(n56) );
  NAND22 U56 ( .A(B[5]), .B(A[5]), .Q(n51) );
  INV2 U57 ( .A(n55), .Q(n61) );
  NAND20 U58 ( .A(n8), .B(A[2]), .Q(n84) );
  NOR20 U59 ( .A(n1), .B(n25), .Q(n47) );
  INV0 U60 ( .A(B[0]), .Q(n97) );
  NAND20 U61 ( .A(n18), .B(n20), .Q(n52) );
  NAND20 U62 ( .A(n21), .B(n51), .Q(n58) );
  NOR20 U63 ( .A(B[7]), .B(A[7]), .Q(n26) );
  XNR20 U64 ( .A(B[7]), .B(A[7]), .Q(n45) );
  IMUX20 U65 ( .A(n65), .B(n66), .S(n54), .Q(SUM[4]) );
  XNR20 U66 ( .A(B[4]), .B(A[4]), .Q(n66) );
  NOR20 U67 ( .A(B[4]), .B(A[4]), .Q(n81) );
  NAND20 U68 ( .A(B[7]), .B(A[7]), .Q(n14) );
  NOR20 U69 ( .A(A[4]), .B(B[4]), .Q(n62) );
  NAND22 U70 ( .A(n96), .B(n94), .Q(SUM[0]) );
  INV3 U71 ( .A(n88), .Q(n87) );
  INV3 U72 ( .A(n44), .Q(n76) );
  XOR21 U73 ( .A(n91), .B(n92), .Q(SUM[1]) );
  XOR21 U74 ( .A(n86), .B(n87), .Q(SUM[2]) );
  NAND22 U75 ( .A(n94), .B(n95), .Q(n91) );
  NAND22 U76 ( .A(n4), .B(n97), .Q(n96) );
  INV3 U77 ( .A(A[0]), .Q(n4) );
  INV3 U78 ( .A(A[2]), .Q(n10) );
  NAND31 U79 ( .A(n74), .B(n75), .C(n76), .Q(n68) );
  NAND22 U80 ( .A(n89), .B(n90), .Q(n86) );
  XOR21 U81 ( .A(n58), .B(n59), .Q(SUM[5]) );
  AOI211 U82 ( .A(n17), .B(n18), .C(n19), .Q(n16) );
  INV3 U83 ( .A(n20), .Q(n19) );
  NAND22 U84 ( .A(n10), .B(n9), .Q(n32) );
  NAND22 U85 ( .A(n10), .B(n9), .Q(n79) );
  NAND22 U86 ( .A(B[6]), .B(A[6]), .Q(n20) );
  INV3 U87 ( .A(A[6]), .Q(n57) );
  INV3 U88 ( .A(A[5]), .Q(n64) );
  INV3 U89 ( .A(B[5]), .Q(n63) );
  XOR21 U90 ( .A(n45), .B(n46), .Q(SUM[7]) );
  NOR21 U91 ( .A(n81), .B(n61), .Q(n65) );
  NAND22 U92 ( .A(n22), .B(n23), .Q(n12) );
  NOR21 U93 ( .A(n1), .B(n24), .Q(n23) );
  NOR21 U94 ( .A(n25), .B(n26), .Q(n22) );
  NOR21 U95 ( .A(B[4]), .B(A[4]), .Q(n24) );
  NAND22 U96 ( .A(n84), .B(n85), .Q(n82) );
  NAND22 U97 ( .A(n76), .B(n86), .Q(n85) );
  NAND22 U98 ( .A(n5), .B(n6), .Q(n7) );
  NAND22 U99 ( .A(n7), .B(n15), .Q(n13) );
  INV3 U100 ( .A(A[7]), .Q(n5) );
  INV0 U101 ( .A(B[7]), .Q(n6) );
  XOR20 U102 ( .A(B[3]), .B(A[3]), .Q(n83) );
  XOR21 U103 ( .A(n82), .B(n83), .Q(SUM[3]) );
  CLKIN3 U104 ( .A(n18), .Q(n25) );
  CLKIN3 U105 ( .A(n72), .Q(n40) );
  OAI212 U106 ( .A(n8), .B(A[2]), .C(n84), .Q(n88) );
  CLKIN3 U107 ( .A(n89), .Q(n93) );
endmodule


module E_alu_DW01_add_9 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  INV3 U2 ( .A(n37), .Q(n74) );
  INV3 U3 ( .A(n36), .Q(n31) );
  OAI311 U4 ( .A(n16), .B(n17), .C(n18), .D(n19), .Q(n15) );
  XOR21 U5 ( .A(n50), .B(n51), .Q(SUM[6]) );
  INV6 U6 ( .A(n35), .Q(n34) );
  CLKIN3 U7 ( .A(n24), .Q(n18) );
  NAND33 U8 ( .A(B[1]), .B(n73), .C(A[1]), .Q(n3) );
  NAND20 U9 ( .A(B[0]), .B(A[0]), .Q(n70) );
  NAND22 U10 ( .A(n39), .B(n40), .Q(n29) );
  NOR22 U11 ( .A(n37), .B(n38), .Q(n36) );
  NOR21 U12 ( .A(n18), .B(n27), .Q(n26) );
  NAND22 U13 ( .A(n74), .B(n4), .Q(n40) );
  INV3 U14 ( .A(n3), .Q(n4) );
  NAND22 U15 ( .A(n10), .B(n9), .Q(n73) );
  NOR21 U16 ( .A(n2), .B(n70), .Q(n68) );
  INV3 U17 ( .A(n69), .Q(n41) );
  CLKIN10 U18 ( .A(B[2]), .Q(n9) );
  NAND23 U19 ( .A(B[5]), .B(A[5]), .Q(n49) );
  NAND23 U20 ( .A(n54), .B(n55), .Q(n21) );
  NAND22 U21 ( .A(B[0]), .B(A[0]), .Q(n38) );
  AOI211 U22 ( .A(n20), .B(n21), .C(n22), .Q(n19) );
  NOR23 U23 ( .A(n29), .B(n30), .Q(n11) );
  NAND22 U24 ( .A(n65), .B(n66), .Q(n58) );
  INV3 U25 ( .A(n21), .Q(n16) );
  INV3 U26 ( .A(n9), .Q(n8) );
  NAND23 U27 ( .A(n52), .B(n53), .Q(n47) );
  AOI211 U28 ( .A(n10), .B(n9), .C(n35), .Q(n67) );
  NOR22 U29 ( .A(A[1]), .B(B[1]), .Q(n35) );
  NAND22 U30 ( .A(n61), .B(n62), .Q(n24) );
  MUX22 U31 ( .A(B[0]), .B(n90), .S(A[0]), .Q(SUM[0]) );
  NOR24 U32 ( .A(n41), .B(n42), .Q(n39) );
  INV2 U33 ( .A(B[5]), .Q(n61) );
  NOR20 U34 ( .A(n18), .B(n16), .Q(n45) );
  NAND20 U35 ( .A(B[1]), .B(A[1]), .Q(n84) );
  NAND22 U36 ( .A(B[3]), .B(A[3]), .Q(n69) );
  NAND24 U37 ( .A(n33), .B(n34), .Q(n32) );
  NOR24 U38 ( .A(n37), .B(n72), .Q(n42) );
  INV2 U39 ( .A(n74), .Q(n2) );
  NAND23 U40 ( .A(A[2]), .B(n8), .Q(n72) );
  NAND22 U41 ( .A(n25), .B(n26), .Q(n12) );
  NOR22 U42 ( .A(n16), .B(n28), .Q(n25) );
  NOR21 U43 ( .A(B[7]), .B(A[7]), .Q(n28) );
  NOR21 U44 ( .A(n71), .B(n42), .Q(n65) );
  INV1 U45 ( .A(n40), .Q(n71) );
  AOI312 U46 ( .A(n45), .B(n46), .C(n47), .D(n48), .Q(n44) );
  NOR24 U47 ( .A(n31), .B(n32), .Q(n30) );
  AOI311 U48 ( .A(n46), .B(n24), .C(n47), .D(n20), .Q(n51) );
  XOR20 U49 ( .A(n86), .B(n87), .Q(SUM[1]) );
  INV2 U50 ( .A(n53), .Q(n59) );
  NAND20 U51 ( .A(B[7]), .B(A[7]), .Q(n14) );
  NAND22 U52 ( .A(B[4]), .B(A[4]), .Q(n17) );
  NAND20 U53 ( .A(n8), .B(A[2]), .Q(n78) );
  INV0 U54 ( .A(B[0]), .Q(n90) );
  XNR20 U55 ( .A(n81), .B(n83), .Q(SUM[2]) );
  NOR20 U56 ( .A(n8), .B(A[2]), .Q(n82) );
  NAND20 U57 ( .A(B[0]), .B(A[0]), .Q(n89) );
  NOR20 U58 ( .A(n88), .B(n35), .Q(n87) );
  NAND20 U59 ( .A(n24), .B(n49), .Q(n56) );
  NAND20 U60 ( .A(n21), .B(n23), .Q(n50) );
  NOR24 U61 ( .A(A[3]), .B(B[3]), .Q(n37) );
  NAND20 U62 ( .A(B[4]), .B(A[4]), .Q(n53) );
  XNR20 U63 ( .A(B[7]), .B(A[7]), .Q(n43) );
  IMUX20 U64 ( .A(n63), .B(n64), .S(n52), .Q(SUM[4]) );
  XNR20 U65 ( .A(B[4]), .B(A[4]), .Q(n64) );
  NOR20 U66 ( .A(B[4]), .B(A[4]), .Q(n75) );
  INV2 U67 ( .A(B[6]), .Q(n54) );
  NOR20 U68 ( .A(A[4]), .B(B[4]), .Q(n60) );
  NAND22 U69 ( .A(n10), .B(n9), .Q(n33) );
  INV3 U70 ( .A(n89), .Q(n86) );
  NAND22 U71 ( .A(n78), .B(n79), .Q(n76) );
  NAND22 U72 ( .A(n80), .B(n81), .Q(n79) );
  INV3 U73 ( .A(n82), .Q(n80) );
  INV3 U74 ( .A(A[2]), .Q(n10) );
  XOR21 U75 ( .A(n56), .B(n57), .Q(SUM[5]) );
  AOI211 U76 ( .A(n46), .B(n58), .C(n59), .Q(n57) );
  NAND22 U77 ( .A(n84), .B(n85), .Q(n81) );
  NAND22 U78 ( .A(n86), .B(n34), .Q(n85) );
  INV3 U79 ( .A(n23), .Q(n22) );
  AOI211 U80 ( .A(n67), .B(n68), .C(n41), .Q(n66) );
  NAND22 U81 ( .A(B[6]), .B(A[6]), .Q(n23) );
  INV3 U82 ( .A(A[6]), .Q(n55) );
  INV3 U83 ( .A(A[5]), .Q(n62) );
  INV3 U84 ( .A(n60), .Q(n46) );
  XOR21 U85 ( .A(n43), .B(n44), .Q(SUM[7]) );
  NOR21 U86 ( .A(n75), .B(n59), .Q(n63) );
  NOR21 U87 ( .A(B[4]), .B(A[4]), .Q(n27) );
  NAND22 U88 ( .A(n5), .B(n6), .Q(n7) );
  NAND22 U89 ( .A(n15), .B(n7), .Q(n13) );
  INV3 U90 ( .A(A[7]), .Q(n5) );
  INV0 U91 ( .A(B[7]), .Q(n6) );
  XOR20 U92 ( .A(B[3]), .B(A[3]), .Q(n77) );
  XOR21 U93 ( .A(n76), .B(n77), .Q(SUM[3]) );
  OAI2112 U94 ( .A(n11), .B(n12), .C(n13), .D(n14), .Q(SUM[8]) );
  OAI212 U95 ( .A(n16), .B(n49), .C(n23), .Q(n48) );
  CLKIN3 U96 ( .A(n49), .Q(n20) );
  CLKIN3 U97 ( .A(n58), .Q(n52) );
  OAI212 U98 ( .A(n8), .B(A[2]), .C(n78), .Q(n83) );
  CLKIN3 U99 ( .A(n84), .Q(n88) );
endmodule


module E_alu_DW01_add_10 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  NOR23 U2 ( .A(A[2]), .B(B[2]), .Q(n55) );
  NAND22 U3 ( .A(n12), .B(n13), .Q(SUM[8]) );
  NAND22 U4 ( .A(n21), .B(n32), .Q(n33) );
  NOR21 U5 ( .A(n61), .B(n62), .Q(n50) );
  INV3 U6 ( .A(n16), .Q(n34) );
  INV3 U7 ( .A(n22), .Q(n40) );
  XNR20 U8 ( .A(B[4]), .B(A[4]), .Q(n49) );
  NAND21 U9 ( .A(A[4]), .B(B[4]), .Q(n24) );
  NAND21 U10 ( .A(B[4]), .B(A[4]), .Q(n67) );
  NOR20 U11 ( .A(A[4]), .B(B[4]), .Q(n39) );
  NOR20 U12 ( .A(B[4]), .B(A[4]), .Q(n20) );
  INV6 U13 ( .A(B[3]), .Q(n6) );
  NOR22 U14 ( .A(n10), .B(n5), .Q(n63) );
  INV6 U15 ( .A(n6), .Q(n5) );
  NAND33 U16 ( .A(n50), .B(n51), .C(n52), .Q(n16) );
  NAND21 U17 ( .A(B[5]), .B(A[5]), .Q(n28) );
  INV1 U18 ( .A(B[5]), .Q(n46) );
  NOR21 U19 ( .A(n55), .B(n60), .Q(n59) );
  INV6 U20 ( .A(n4), .Q(n3) );
  NOR20 U21 ( .A(B[4]), .B(A[4]), .Q(n66) );
  CLKIN1 U22 ( .A(B[7]), .Q(n8) );
  NAND22 U23 ( .A(n21), .B(n22), .Q(n19) );
  INV2 U24 ( .A(n75), .Q(n80) );
  NAND20 U25 ( .A(n7), .B(A[7]), .Q(n13) );
  XNR20 U26 ( .A(n7), .B(A[7]), .Q(n2) );
  IMUX20 U27 ( .A(n48), .B(n49), .S(n34), .Q(SUM[4]) );
  NAND20 U28 ( .A(n37), .B(n22), .Q(n36) );
  INV2 U29 ( .A(n38), .Q(n35) );
  AOI210 U30 ( .A(n6), .B(n11), .C(n57), .Q(n58) );
  NAND20 U31 ( .A(n22), .B(n28), .Q(n43) );
  AOI210 U32 ( .A(n45), .B(n16), .C(n37), .Q(n44) );
  INV0 U33 ( .A(n39), .Q(n45) );
  NOR20 U34 ( .A(n74), .B(n55), .Q(n73) );
  XOR20 U35 ( .A(n71), .B(n73), .Q(SUM[2]) );
  NOR20 U36 ( .A(n80), .B(n57), .Q(n79) );
  XOR20 U37 ( .A(n77), .B(n79), .Q(SUM[1]) );
  CLKIN0 U38 ( .A(n57), .Q(n78) );
  INV3 U39 ( .A(n32), .Q(n27) );
  INV0 U40 ( .A(n55), .Q(n72) );
  INV2 U41 ( .A(n21), .Q(n23) );
  XNR21 U42 ( .A(n68), .B(n1), .Q(SUM[3]) );
  XNR20 U43 ( .A(n5), .B(n10), .Q(n1) );
  NAND20 U44 ( .A(B[1]), .B(A[1]), .Q(n65) );
  NAND20 U45 ( .A(B[1]), .B(A[1]), .Q(n75) );
  NAND20 U46 ( .A(B[2]), .B(A[2]), .Q(n69) );
  NAND20 U47 ( .A(A[2]), .B(B[2]), .Q(n64) );
  XOR21 U48 ( .A(n2), .B(n30), .Q(SUM[7]) );
  NAND22 U49 ( .A(n83), .B(n81), .Q(SUM[0]) );
  NAND22 U50 ( .A(n9), .B(n84), .Q(n83) );
  NAND22 U51 ( .A(n81), .B(n82), .Q(n77) );
  NOR21 U52 ( .A(A[0]), .B(n3), .Q(n82) );
  NAND22 U53 ( .A(n3), .B(A[0]), .Q(n81) );
  INV3 U54 ( .A(n3), .Q(n84) );
  INV3 U55 ( .A(n11), .Q(n10) );
  NOR21 U56 ( .A(n66), .B(n37), .Q(n48) );
  INV3 U57 ( .A(n8), .Q(n7) );
  INV3 U58 ( .A(A[3]), .Q(n11) );
  INV3 U59 ( .A(A[0]), .Q(n9) );
  OAI2111 U60 ( .A(n34), .B(n35), .C(n36), .D(n28), .Q(n31) );
  NOR21 U61 ( .A(n39), .B(n40), .Q(n38) );
  AOI221 U62 ( .A(n5), .B(n10), .C(n53), .D(n54), .Q(n52) );
  NAND22 U63 ( .A(n58), .B(n59), .Q(n51) );
  AOI221 U64 ( .A(n14), .B(n15), .C(n16), .D(n17), .Q(n12) );
  INV3 U65 ( .A(n29), .Q(n14) );
  AOI2111 U66 ( .A(n18), .B(n8), .C(n19), .D(n20), .Q(n17) );
  OAI311 U67 ( .A(n23), .B(n24), .C(n40), .D(n25), .Q(n15) );
  AOI211 U68 ( .A(n9), .B(n4), .C(n57), .Q(n53) );
  NAND22 U69 ( .A(n3), .B(A[0]), .Q(n60) );
  XOR21 U70 ( .A(n43), .B(n44), .Q(SUM[5]) );
  NAND22 U71 ( .A(n75), .B(n76), .Q(n71) );
  NAND22 U72 ( .A(n77), .B(n78), .Q(n76) );
  NOR21 U73 ( .A(n55), .B(n56), .Q(n54) );
  NOR21 U74 ( .A(n5), .B(n10), .Q(n56) );
  AOI211 U75 ( .A(n26), .B(n21), .C(n27), .Q(n25) );
  INV3 U76 ( .A(n28), .Q(n26) );
  XNR21 U77 ( .A(n33), .B(n31), .Q(SUM[6]) );
  NAND22 U78 ( .A(n71), .B(n72), .Q(n70) );
  NAND22 U79 ( .A(n69), .B(n70), .Q(n68) );
  NOR21 U80 ( .A(A[7]), .B(n7), .Q(n29) );
  NOR22 U81 ( .A(A[1]), .B(B[1]), .Q(n57) );
  NAND22 U82 ( .A(n46), .B(n47), .Q(n22) );
  INV3 U83 ( .A(A[5]), .Q(n47) );
  NAND22 U84 ( .A(B[6]), .B(A[6]), .Q(n32) );
  NOR31 U85 ( .A(n65), .B(n55), .C(n63), .Q(n61) );
  NOR21 U86 ( .A(n63), .B(n64), .Q(n62) );
  NAND22 U87 ( .A(n41), .B(n42), .Q(n21) );
  INV3 U88 ( .A(A[6]), .Q(n42) );
  INV3 U89 ( .A(B[6]), .Q(n41) );
  INV3 U90 ( .A(A[7]), .Q(n18) );
  INV2 U91 ( .A(B[0]), .Q(n4) );
  AOI212 U92 ( .A(n31), .B(n21), .C(n27), .Q(n30) );
  CLKIN3 U93 ( .A(n67), .Q(n37) );
  CLKIN3 U94 ( .A(n69), .Q(n74) );
endmodule


module E_alu_DW01_add_11 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78;

  NOR23 U2 ( .A(A[3]), .B(n7), .Q(n59) );
  NOR22 U3 ( .A(A[2]), .B(B[2]), .Q(n52) );
  AOI221 U4 ( .A(n13), .B(n14), .C(n15), .D(n16), .Q(n11) );
  CLKIN6 U5 ( .A(n8), .Q(n7) );
  NOR21 U6 ( .A(n52), .B(n56), .Q(n55) );
  INV3 U7 ( .A(B[3]), .Q(n8) );
  AOI211 U8 ( .A(n44), .B(n15), .C(n36), .Q(n43) );
  NAND22 U9 ( .A(n20), .B(n31), .Q(n32) );
  INV3 U10 ( .A(n31), .Q(n26) );
  NAND22 U11 ( .A(n40), .B(n41), .Q(n20) );
  INV3 U12 ( .A(n20), .Q(n22) );
  INV3 U13 ( .A(n6), .Q(n78) );
  XNR21 U14 ( .A(n32), .B(n30), .Q(SUM[6]) );
  CLKIN3 U15 ( .A(n38), .Q(n44) );
  CLKIN3 U16 ( .A(n37), .Q(n34) );
  INV6 U17 ( .A(n15), .Q(n33) );
  NAND34 U18 ( .A(n49), .B(n50), .C(n51), .Q(n15) );
  INV3 U19 ( .A(n30), .Q(n1) );
  NOR22 U20 ( .A(n57), .B(n58), .Q(n49) );
  NOR24 U21 ( .A(n1), .B(n22), .Q(n2) );
  NOR24 U22 ( .A(n2), .B(n26), .Q(n29) );
  XNR22 U23 ( .A(n5), .B(n29), .Q(SUM[7]) );
  OAI2112 U24 ( .A(n33), .B(n34), .C(n35), .D(n27), .Q(n30) );
  NOR31 U25 ( .A(n61), .B(n52), .C(n59), .Q(n57) );
  INV1 U26 ( .A(B[5]), .Q(n45) );
  NAND20 U27 ( .A(n20), .B(n21), .Q(n18) );
  IMUX20 U28 ( .A(n6), .B(n78), .S(A[0]), .Q(SUM[0]) );
  NAND20 U29 ( .A(B[7]), .B(A[7]), .Q(n12) );
  NOR20 U30 ( .A(A[4]), .B(B[4]), .Q(n38) );
  NOR20 U31 ( .A(B[4]), .B(A[4]), .Q(n19) );
  NOR20 U32 ( .A(n62), .B(n36), .Q(n47) );
  XNR20 U33 ( .A(B[4]), .B(A[4]), .Q(n48) );
  NOR20 U34 ( .A(B[4]), .B(A[4]), .Q(n62) );
  NAND20 U35 ( .A(A[4]), .B(B[4]), .Q(n23) );
  NAND20 U36 ( .A(B[4]), .B(A[4]), .Q(n63) );
  NAND20 U37 ( .A(n36), .B(n21), .Q(n35) );
  AOI210 U38 ( .A(n8), .B(n10), .C(n53), .Q(n54) );
  XNR21 U39 ( .A(n64), .B(n4), .Q(SUM[3]) );
  XNR20 U40 ( .A(n7), .B(A[3]), .Q(n4) );
  NOR20 U41 ( .A(n76), .B(n53), .Q(n75) );
  INV0 U42 ( .A(n53), .Q(n74) );
  INV1 U43 ( .A(B[7]), .Q(n9) );
  INV0 U44 ( .A(n52), .Q(n68) );
  INV0 U45 ( .A(n21), .Q(n39) );
  NAND20 U46 ( .A(n21), .B(n27), .Q(n42) );
  NAND21 U47 ( .A(B[5]), .B(A[5]), .Q(n27) );
  NAND20 U48 ( .A(B[1]), .B(A[1]), .Q(n61) );
  NAND20 U49 ( .A(B[1]), .B(A[1]), .Q(n71) );
  NAND20 U50 ( .A(B[2]), .B(A[2]), .Q(n65) );
  XOR20 U51 ( .A(B[7]), .B(A[7]), .Q(n5) );
  NAND20 U52 ( .A(A[2]), .B(B[2]), .Q(n60) );
  IMUX21 U53 ( .A(n47), .B(n48), .S(n33), .Q(SUM[4]) );
  INV3 U54 ( .A(n77), .Q(n73) );
  NAND22 U55 ( .A(n78), .B(A[0]), .Q(n77) );
  INV3 U56 ( .A(A[3]), .Q(n10) );
  NOR21 U57 ( .A(n38), .B(n39), .Q(n37) );
  NAND22 U58 ( .A(n7), .B(A[3]), .Q(n51) );
  NAND22 U59 ( .A(n54), .B(n55), .Q(n50) );
  INV3 U60 ( .A(n28), .Q(n13) );
  AOI2111 U61 ( .A(n17), .B(n9), .C(n18), .D(n19), .Q(n16) );
  OAI311 U62 ( .A(n22), .B(n23), .C(n39), .D(n24), .Q(n14) );
  NAND22 U63 ( .A(n78), .B(A[0]), .Q(n56) );
  XOR21 U64 ( .A(n67), .B(n69), .Q(SUM[2]) );
  NOR21 U65 ( .A(n70), .B(n52), .Q(n69) );
  NAND22 U66 ( .A(n71), .B(n72), .Q(n67) );
  NAND22 U67 ( .A(n73), .B(n74), .Q(n72) );
  AOI211 U68 ( .A(n25), .B(n20), .C(n26), .Q(n24) );
  INV3 U69 ( .A(n27), .Q(n25) );
  NAND22 U70 ( .A(n65), .B(n66), .Q(n64) );
  NAND22 U71 ( .A(n67), .B(n68), .Q(n66) );
  XOR21 U72 ( .A(n42), .B(n43), .Q(SUM[5]) );
  XOR21 U73 ( .A(n73), .B(n75), .Q(SUM[1]) );
  NOR21 U74 ( .A(A[7]), .B(B[7]), .Q(n28) );
  NOR21 U75 ( .A(A[1]), .B(B[1]), .Q(n53) );
  NAND22 U76 ( .A(n45), .B(n46), .Q(n21) );
  INV3 U77 ( .A(A[5]), .Q(n46) );
  NAND22 U78 ( .A(B[6]), .B(A[6]), .Q(n31) );
  NAND22 U79 ( .A(n11), .B(n12), .Q(SUM[8]) );
  NOR21 U80 ( .A(n59), .B(n60), .Q(n58) );
  INV3 U81 ( .A(A[6]), .Q(n41) );
  INV3 U82 ( .A(B[6]), .Q(n40) );
  INV3 U83 ( .A(A[7]), .Q(n17) );
  INV3 U84 ( .A(B[0]), .Q(n6) );
  CLKIN3 U85 ( .A(n63), .Q(n36) );
  CLKIN3 U86 ( .A(n65), .Q(n70) );
  CLKIN3 U87 ( .A(n71), .Q(n76) );
endmodule


module E_alu_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277;

  AOI211 U3 ( .A(n21), .B(n113), .C(n179), .Q(n178) );
  NAND24 U4 ( .A(n192), .B(n193), .Q(n125) );
  NAND22 U5 ( .A(n139), .B(n140), .Q(n81) );
  AOI221 U6 ( .A(A[29]), .B(n11), .C(A[30]), .D(n184), .Q(n193) );
  NOR21 U7 ( .A(n21), .B(n122), .Q(B[25]) );
  AOI221 U8 ( .A(A[27]), .B(n10), .C(A[28]), .D(n184), .Q(n218) );
  NAND21 U9 ( .A(n99), .B(n125), .Q(n124) );
  NOR21 U10 ( .A(n167), .B(n216), .Q(n215) );
  NOR21 U11 ( .A(SH[3]), .B(SH[2]), .Q(n15) );
  NAND22 U12 ( .A(n229), .B(n230), .Q(n121) );
  NAND22 U13 ( .A(n237), .B(n238), .Q(n105) );
  NAND23 U14 ( .A(n256), .B(n257), .Q(n129) );
  INV3 U15 ( .A(n118), .Q(B[27]) );
  AOI221 U16 ( .A(A[26]), .B(n185), .C(A[27]), .D(n186), .Q(n258) );
  AOI221 U17 ( .A(A[20]), .B(n10), .C(A[21]), .D(n184), .Q(n261) );
  INV3 U18 ( .A(n13), .Q(n14) );
  INV2 U19 ( .A(n183), .Q(n13) );
  INV3 U20 ( .A(SH[4]), .Q(n22) );
  NAND22 U21 ( .A(n99), .B(n22), .Q(n245) );
  NAND22 U22 ( .A(n232), .B(n233), .Q(n107) );
  AOI221 U23 ( .A(A[28]), .B(n185), .C(A[29]), .D(n186), .Q(n232) );
  NAND22 U24 ( .A(n197), .B(n198), .Q(n33) );
  AOI221 U25 ( .A(A[28]), .B(n12), .C(A[29]), .D(n184), .Q(n257) );
  NAND22 U26 ( .A(n97), .B(n22), .Q(n239) );
  NAND21 U27 ( .A(n21), .B(n53), .Q(n52) );
  NAND21 U28 ( .A(n21), .B(n67), .Q(n66) );
  NAND21 U29 ( .A(n227), .B(n228), .Q(B[10]) );
  NAND21 U30 ( .A(n21), .B(n119), .Q(n209) );
  NAND21 U31 ( .A(n21), .B(n116), .Q(n205) );
  NAND21 U32 ( .A(n21), .B(n25), .Q(n24) );
  NAND21 U33 ( .A(n21), .B(n81), .Q(n80) );
  INV6 U34 ( .A(n277), .Q(n185) );
  NAND21 U35 ( .A(SH[1]), .B(n17), .Q(n277) );
  NAND20 U36 ( .A(A[31]), .B(n185), .Q(n192) );
  INV6 U37 ( .A(n276), .Q(n184) );
  INV1 U38 ( .A(n6), .Q(n7) );
  INV2 U39 ( .A(n5), .Q(n6) );
  AOI221 U40 ( .A(A[26]), .B(n14), .C(A[27]), .D(n184), .Q(n233) );
  NAND22 U41 ( .A(SH[2]), .B(n20), .Q(n216) );
  CLKIN2 U42 ( .A(n13), .Q(n11) );
  NAND20 U43 ( .A(n39), .B(n31), .Q(n180) );
  CLKIN2 U44 ( .A(n180), .Q(n179) );
  NAND21 U45 ( .A(n16), .B(n117), .Q(n127) );
  NAND21 U46 ( .A(n30), .B(n46), .Q(n90) );
  CLKIN1 U47 ( .A(n6), .Q(n10) );
  NAND22 U48 ( .A(n99), .B(n129), .Q(n128) );
  CLKIN1 U49 ( .A(n6), .Q(n8) );
  AOI221 U50 ( .A(n96), .B(n117), .C(n97), .D(n129), .Q(n255) );
  NAND21 U51 ( .A(A[31]), .B(n11), .Q(n167) );
  NAND22 U52 ( .A(n39), .B(n45), .Q(n91) );
  NAND22 U53 ( .A(n34), .B(n63), .Q(n62) );
  NAND20 U54 ( .A(n96), .B(n22), .Q(n242) );
  INV3 U55 ( .A(SH[0]), .Q(n17) );
  NAND20 U56 ( .A(n98), .B(n125), .Q(n191) );
  NOR21 U57 ( .A(SH[3]), .B(SH[2]), .Q(n16) );
  AOI220 U58 ( .A(n34), .B(n46), .C(n39), .D(n47), .Q(n203) );
  AOI221 U59 ( .A(n16), .B(n47), .C(n99), .D(n48), .Q(n254) );
  NAND22 U60 ( .A(n96), .B(n125), .Q(n140) );
  AOI220 U61 ( .A(n98), .B(n103), .C(n99), .D(n101), .Q(n131) );
  AOI2110 U62 ( .A(n34), .B(n49), .C(n87), .D(n88), .Q(n86) );
  INV3 U63 ( .A(n22), .Q(n21) );
  AOI220 U64 ( .A(A[21]), .B(n14), .C(A[22]), .D(n184), .Q(n198) );
  AOI220 U65 ( .A(A[23]), .B(n185), .C(A[24]), .D(n186), .Q(n197) );
  NOR21 U66 ( .A(n21), .B(n126), .Q(B[24]) );
  CLKIN1 U67 ( .A(n6), .Q(n9) );
  NAND20 U68 ( .A(n98), .B(n133), .Q(n166) );
  NOR21 U69 ( .A(n21), .B(n85), .Q(B[20]) );
  NAND20 U70 ( .A(SH[3]), .B(SH[2]), .Q(n268) );
  AOI221 U71 ( .A(n16), .B(n105), .C(n99), .D(n107), .Q(n135) );
  NAND21 U72 ( .A(n96), .B(n137), .Q(n136) );
  NAND20 U73 ( .A(n96), .B(n133), .Q(n132) );
  AOI220 U74 ( .A(n99), .B(n37), .C(n98), .D(n38), .Q(n146) );
  CLKIN2 U75 ( .A(n175), .Q(n171) );
  AOI220 U76 ( .A(n15), .B(n68), .C(n99), .D(n77), .Q(n110) );
  NAND20 U77 ( .A(n32), .B(n60), .Q(n57) );
  NAND20 U78 ( .A(n30), .B(n59), .Q(n58) );
  NAND20 U79 ( .A(n34), .B(n59), .Q(n165) );
  CLKIN3 U80 ( .A(n248), .Q(n34) );
  NAND21 U81 ( .A(n15), .B(n22), .Q(n248) );
  CLKIN3 U82 ( .A(n239), .Q(n32) );
  CLKIN3 U83 ( .A(n242), .Q(n30) );
  NAND22 U84 ( .A(n113), .B(n22), .Q(n112) );
  CLKIN1 U85 ( .A(SH[2]), .Q(n19) );
  NAND20 U86 ( .A(n21), .B(n121), .Q(n228) );
  CLKIN3 U87 ( .A(n206), .Q(n116) );
  CLKIN3 U88 ( .A(n191), .Q(n113) );
  INV3 U89 ( .A(n67), .Q(n134) );
  INV0 U90 ( .A(n44), .Q(n126) );
  AOI220 U91 ( .A(A[30]), .B(n185), .C(A[31]), .D(n186), .Q(n256) );
  AOI220 U92 ( .A(A[14]), .B(n185), .C(A[15]), .D(n186), .Q(n266) );
  AOI220 U93 ( .A(A[12]), .B(n9), .C(A[13]), .D(n184), .Q(n267) );
  AOI220 U94 ( .A(A[13]), .B(n185), .C(A[14]), .D(n186), .Q(n225) );
  AOI220 U95 ( .A(n97), .B(n40), .C(n96), .D(n35), .Q(n147) );
  CLKIN3 U96 ( .A(n231), .Q(n137) );
  AOI220 U97 ( .A(A[30]), .B(n11), .C(A[31]), .D(n184), .Q(n231) );
  NOR20 U98 ( .A(SH[1]), .B(SH[0]), .Q(n5) );
  NOR20 U99 ( .A(SH[1]), .B(SH[0]), .Q(n183) );
  CLKIN3 U100 ( .A(n214), .Q(n119) );
  AOI220 U101 ( .A(n30), .B(n48), .C(n32), .D(n117), .Q(n204) );
  AOI220 U102 ( .A(n32), .B(n114), .C(n30), .D(n33), .Q(n177) );
  NAND20 U103 ( .A(n98), .B(n114), .Q(n123) );
  AOI220 U104 ( .A(n96), .B(n107), .C(n97), .D(n137), .Q(n153) );
  AOI220 U105 ( .A(n96), .B(n101), .C(n97), .D(n133), .Q(n150) );
  AOI220 U106 ( .A(n16), .B(n60), .C(n99), .D(n103), .Q(n149) );
  AOI220 U107 ( .A(n98), .B(n31), .C(n99), .D(n33), .Q(n155) );
  AOI220 U108 ( .A(n96), .B(n114), .C(n97), .D(n125), .Q(n156) );
  NAND21 U109 ( .A(n39), .B(n40), .Q(n36) );
  NAND21 U110 ( .A(n30), .B(n73), .Q(n72) );
  NAND20 U111 ( .A(n34), .B(n73), .Q(n175) );
  MUX22 U112 ( .A(n92), .B(n93), .S(n21), .Q(B[3]) );
  NAND20 U113 ( .A(n30), .B(n103), .Q(n164) );
  NAND20 U114 ( .A(n34), .B(n40), .Q(n176) );
  AOI220 U115 ( .A(n98), .B(n48), .C(n99), .D(n117), .Q(n142) );
  NAND20 U116 ( .A(n96), .B(n129), .Q(n143) );
  AOI220 U117 ( .A(n39), .B(n74), .C(n21), .D(n106), .Q(n169) );
  NAND20 U118 ( .A(n32), .B(n47), .Q(n89) );
  NAND20 U119 ( .A(n32), .B(n101), .Q(n163) );
  NAND20 U120 ( .A(n39), .B(n64), .Q(n61) );
  NAND21 U121 ( .A(n30), .B(n31), .Q(n29) );
  AOI220 U122 ( .A(n32), .B(n33), .C(n34), .D(n35), .Q(n28) );
  NAND20 U123 ( .A(n30), .B(n105), .Q(n174) );
  NAND20 U124 ( .A(n32), .B(n107), .Q(n173) );
  AOI220 U125 ( .A(n39), .B(n60), .C(n21), .D(n102), .Q(n159) );
  INV3 U126 ( .A(n81), .Q(n138) );
  MUX21 U127 ( .A(n108), .B(n109), .S(n21), .Q(B[2]) );
  MUX21 U128 ( .A(n144), .B(n145), .S(n21), .Q(B[1]) );
  INV3 U129 ( .A(n53), .Q(n130) );
  MUX22 U130 ( .A(n253), .B(n158), .S(n21), .Q(B[0]) );
  AOI220 U131 ( .A(A[20]), .B(n185), .C(A[21]), .D(n186), .Q(n240) );
  AOI220 U132 ( .A(A[13]), .B(n14), .C(A[14]), .D(n184), .Q(n202) );
  AOI220 U133 ( .A(n185), .B(A[17]), .C(A[18]), .D(n186), .Q(n223) );
  AOI220 U134 ( .A(A[29]), .B(n185), .C(A[30]), .D(n186), .Q(n217) );
  AOI220 U135 ( .A(A[17]), .B(n12), .C(A[18]), .D(n184), .Q(n188) );
  AOI220 U136 ( .A(A[14]), .B(n14), .C(A[15]), .D(n184), .Q(n244) );
  AOI220 U137 ( .A(A[21]), .B(n185), .C(A[22]), .D(n186), .Q(n221) );
  AOI220 U138 ( .A(A[27]), .B(n185), .C(A[28]), .D(n186), .Q(n199) );
  AOI220 U139 ( .A(A[24]), .B(n11), .C(A[25]), .D(n184), .Q(n259) );
  AOI220 U140 ( .A(A[23]), .B(n8), .C(A[24]), .D(n184), .Q(n220) );
  AOI220 U141 ( .A(A[25]), .B(n185), .C(A[26]), .D(n186), .Q(n219) );
  AOI220 U142 ( .A(A[24]), .B(n185), .C(A[25]), .D(n186), .Q(n237) );
  AOI220 U143 ( .A(A[22]), .B(n12), .C(A[23]), .D(n184), .Q(n238) );
  AOI220 U144 ( .A(A[22]), .B(n185), .C(A[23]), .D(n186), .Q(n260) );
  AOI220 U145 ( .A(A[12]), .B(n185), .C(A[13]), .D(n186), .Q(n246) );
  AOI220 U146 ( .A(A[8]), .B(n8), .C(A[9]), .D(n184), .Q(n270) );
  CLKIN3 U147 ( .A(n104), .Q(B[30]) );
  AOI220 U148 ( .A(A[8]), .B(n185), .C(A[9]), .D(n186), .Q(n249) );
  CLKIN3 U149 ( .A(n115), .Q(B[28]) );
  INV3 U150 ( .A(n167), .Q(n133) );
  INV3 U151 ( .A(n234), .Q(n227) );
  NAND22 U152 ( .A(n235), .B(n236), .Q(n234) );
  NAND22 U153 ( .A(n23), .B(n24), .Q(B[9]) );
  NOR21 U154 ( .A(n26), .B(n27), .Q(n23) );
  INV3 U155 ( .A(n36), .Q(n26) );
  NAND22 U156 ( .A(n51), .B(n52), .Q(B[7]) );
  NOR21 U157 ( .A(n55), .B(n56), .Q(n51) );
  NAND22 U158 ( .A(n61), .B(n62), .Q(n55) );
  NAND22 U159 ( .A(n16), .B(n129), .Q(n206) );
  NAND22 U160 ( .A(n79), .B(n80), .Q(B[5]) );
  INV3 U161 ( .A(n82), .Q(n79) );
  NAND22 U162 ( .A(n83), .B(n84), .Q(n82) );
  INV3 U163 ( .A(n6), .Q(n12) );
  INV3 U164 ( .A(n166), .Q(n102) );
  INV3 U165 ( .A(n170), .Q(n106) );
  NAND22 U166 ( .A(n16), .B(n137), .Q(n170) );
  INV3 U167 ( .A(n194), .Q(n186) );
  NAND22 U168 ( .A(SH[1]), .B(SH[0]), .Q(n194) );
  NAND22 U169 ( .A(n152), .B(n153), .Q(n109) );
  AOI221 U170 ( .A(n34), .B(n37), .C(n39), .D(n35), .Q(n84) );
  AOI221 U171 ( .A(n96), .B(n78), .C(n97), .D(n73), .Q(n111) );
  NAND22 U172 ( .A(n266), .B(n267), .Q(n46) );
  NAND31 U173 ( .A(n42), .B(n43), .C(n41), .Q(B[8]) );
  AOI221 U174 ( .A(n34), .B(n45), .C(n39), .D(n46), .Q(n42) );
  NAND22 U175 ( .A(n21), .B(n44), .Q(n43) );
  AOI221 U176 ( .A(n30), .B(n47), .C(n32), .D(n48), .Q(n41) );
  INV3 U177 ( .A(n216), .Q(n99) );
  AOI221 U178 ( .A(n32), .B(n31), .C(n30), .D(n40), .Q(n83) );
  AOI221 U179 ( .A(n34), .B(n78), .C(n39), .D(n73), .Q(n235) );
  AOI221 U180 ( .A(n30), .B(n60), .C(n32), .D(n103), .Q(n208) );
  NAND22 U181 ( .A(n142), .B(n143), .Q(n141) );
  INV3 U182 ( .A(n91), .Q(n87) );
  NAND22 U183 ( .A(n89), .B(n90), .Q(n88) );
  AOI221 U184 ( .A(n15), .B(n33), .C(n99), .D(n114), .Q(n139) );
  NAND22 U185 ( .A(n127), .B(n128), .Q(n44) );
  NAND22 U186 ( .A(n123), .B(n124), .Q(n25) );
  NAND22 U187 ( .A(n99), .B(n137), .Q(n230) );
  NAND22 U188 ( .A(n15), .B(n107), .Q(n229) );
  NAND22 U189 ( .A(n135), .B(n136), .Q(n67) );
  NAND22 U190 ( .A(n131), .B(n132), .Q(n53) );
  NAND22 U191 ( .A(n254), .B(n255), .Q(n158) );
  NAND22 U192 ( .A(n149), .B(n150), .Q(n93) );
  NAND22 U193 ( .A(n155), .B(n156), .Q(n145) );
  NAND22 U194 ( .A(n94), .B(n95), .Q(n92) );
  INV3 U195 ( .A(n268), .Q(n97) );
  NAND31 U196 ( .A(n177), .B(n178), .C(n176), .Q(B[13]) );
  NAND22 U197 ( .A(n34), .B(n77), .Q(n76) );
  NAND22 U198 ( .A(n28), .B(n29), .Q(n27) );
  NAND22 U199 ( .A(n57), .B(n58), .Q(n56) );
  NAND22 U200 ( .A(n173), .B(n174), .Q(n172) );
  NOR21 U201 ( .A(n21), .B(n134), .Q(B[22]) );
  NOR21 U202 ( .A(n21), .B(n120), .Q(B[26]) );
  NOR21 U203 ( .A(n21), .B(n157), .Q(B[16]) );
  NOR21 U204 ( .A(n21), .B(n154), .Q(B[17]) );
  NOR21 U205 ( .A(n21), .B(n151), .Q(B[18]) );
  NOR21 U206 ( .A(n21), .B(n148), .Q(B[19]) );
  NAND22 U207 ( .A(n168), .B(n169), .Q(B[14]) );
  NOR21 U208 ( .A(n171), .B(n172), .Q(n168) );
  NOR21 U209 ( .A(n21), .B(n130), .Q(B[23]) );
  NOR21 U210 ( .A(n69), .B(n70), .Q(n65) );
  NAND22 U211 ( .A(n75), .B(n76), .Q(n69) );
  NAND22 U212 ( .A(n71), .B(n72), .Q(n70) );
  NAND22 U213 ( .A(n39), .B(n78), .Q(n75) );
  NAND22 U214 ( .A(n159), .B(n160), .Q(B[15]) );
  NOR21 U215 ( .A(n161), .B(n162), .Q(n160) );
  NAND22 U216 ( .A(n163), .B(n164), .Q(n162) );
  NOR21 U217 ( .A(n21), .B(n138), .Q(B[21]) );
  INV3 U218 ( .A(n165), .Q(n161) );
  NAND22 U219 ( .A(n264), .B(n265), .Q(n253) );
  AOI221 U220 ( .A(n96), .B(n45), .C(n97), .D(n46), .Q(n265) );
  NAND22 U221 ( .A(n110), .B(n111), .Q(n108) );
  NAND22 U222 ( .A(n146), .B(n147), .Q(n144) );
  NOR21 U223 ( .A(SH[3]), .B(SH[2]), .Q(n98) );
  NAND22 U224 ( .A(n223), .B(n224), .Q(n59) );
  NAND22 U225 ( .A(n249), .B(n250), .Q(n77) );
  NAND22 U226 ( .A(n246), .B(n247), .Q(n78) );
  NAND22 U227 ( .A(n187), .B(n188), .Q(n31) );
  NAND22 U228 ( .A(n119), .B(n22), .Q(n118) );
  NAND22 U229 ( .A(SH[0]), .B(n18), .Q(n276) );
  NAND22 U230 ( .A(n243), .B(n244), .Q(n73) );
  NAND22 U231 ( .A(n262), .B(n263), .Q(n47) );
  NAND22 U232 ( .A(n201), .B(n202), .Q(n40) );
  NAND22 U233 ( .A(n221), .B(n222), .Q(n60) );
  NAND22 U234 ( .A(n258), .B(n259), .Q(n117) );
  NAND22 U235 ( .A(n219), .B(n220), .Q(n103) );
  NAND22 U236 ( .A(n199), .B(n200), .Q(n114) );
  AOI221 U237 ( .A(A[25]), .B(n9), .C(A[26]), .D(n184), .Q(n200) );
  NAND22 U238 ( .A(n217), .B(n218), .Q(n101) );
  NAND22 U239 ( .A(n189), .B(n190), .Q(n37) );
  NAND22 U240 ( .A(n240), .B(n241), .Q(n74) );
  NAND22 U241 ( .A(n269), .B(n270), .Q(n45) );
  NAND22 U242 ( .A(n260), .B(n261), .Q(n48) );
  AOI221 U243 ( .A(n16), .B(n54), .C(n99), .D(n63), .Q(n94) );
  AOI221 U244 ( .A(n15), .B(n50), .C(n99), .D(n49), .Q(n264) );
  NAND22 U245 ( .A(n272), .B(n273), .Q(n49) );
  NAND22 U246 ( .A(n106), .B(n22), .Q(n104) );
  INV3 U247 ( .A(n245), .Q(n39) );
  INV3 U248 ( .A(n100), .Q(B[31]) );
  NAND22 U249 ( .A(n102), .B(n22), .Q(n100) );
  INV3 U250 ( .A(n271), .Q(n96) );
  NAND22 U251 ( .A(SH[3]), .B(n19), .Q(n271) );
  NAND22 U252 ( .A(n251), .B(n252), .Q(n68) );
  NAND31 U253 ( .A(n204), .B(n205), .C(n203), .Q(B[12]) );
  NAND31 U254 ( .A(n208), .B(n209), .C(n207), .Q(B[11]) );
  NAND22 U255 ( .A(n116), .B(n22), .Q(n115) );
  INV3 U256 ( .A(n112), .Q(B[29]) );
  NAND22 U257 ( .A(n65), .B(n66), .Q(B[6]) );
  INV3 U258 ( .A(SH[1]), .Q(n18) );
  INV3 U259 ( .A(SH[3]), .Q(n20) );
  OAI222 U260 ( .A(n15), .B(n215), .C(n101), .D(n215), .Q(n214) );
  AOI221 U261 ( .A(n34), .B(n64), .C(n39), .D(n59), .Q(n207) );
  AOI221 U262 ( .A(n96), .B(n64), .C(n97), .D(n59), .Q(n95) );
  AOI220 U263 ( .A(A[15]), .B(n185), .C(A[16]), .D(n186), .Q(n201) );
  AOI220 U264 ( .A(A[16]), .B(n12), .C(n184), .D(A[17]), .Q(n263) );
  AOI220 U265 ( .A(A[15]), .B(n14), .C(A[16]), .D(n184), .Q(n224) );
  AOI220 U266 ( .A(A[16]), .B(n185), .C(A[17]), .D(n186), .Q(n243) );
  AOI220 U267 ( .A(A[6]), .B(n8), .C(A[7]), .D(n184), .Q(n250) );
  AOI221 U268 ( .A(n15), .B(n74), .C(n99), .D(n105), .Q(n152) );
  AOI220 U269 ( .A(n30), .B(n74), .C(n32), .D(n105), .Q(n236) );
  NAND20 U270 ( .A(n32), .B(n74), .Q(n71) );
  AOI220 U271 ( .A(A[7]), .B(n12), .C(A[8]), .D(n184), .Q(n213) );
  AOI220 U272 ( .A(A[7]), .B(n185), .C(A[8]), .D(n186), .Q(n189) );
  AOI220 U273 ( .A(A[6]), .B(n185), .C(A[7]), .D(n186), .Q(n272) );
  NAND22 U274 ( .A(n210), .B(n211), .Q(n54) );
  NAND22 U275 ( .A(n195), .B(n196), .Q(n38) );
  NAND22 U276 ( .A(n274), .B(n275), .Q(n50) );
  NAND22 U277 ( .A(n212), .B(n213), .Q(n63) );
  AOI220 U278 ( .A(A[11]), .B(n11), .C(A[12]), .D(n184), .Q(n226) );
  AOI220 U279 ( .A(A[11]), .B(n185), .C(A[12]), .D(n186), .Q(n181) );
  NAND22 U280 ( .A(n225), .B(n226), .Q(n64) );
  NAND22 U281 ( .A(n181), .B(n182), .Q(n35) );
  AOI220 U282 ( .A(A[9]), .B(n185), .C(A[10]), .D(n186), .Q(n212) );
  AOI220 U283 ( .A(A[9]), .B(n14), .C(A[10]), .D(n184), .Q(n182) );
  AOI220 U284 ( .A(A[10]), .B(n185), .C(A[11]), .D(n186), .Q(n269) );
  AOI220 U285 ( .A(A[10]), .B(n9), .C(A[11]), .D(n184), .Q(n247) );
  AOI220 U286 ( .A(n185), .B(A[18]), .C(A[19]), .D(n186), .Q(n262) );
  AOI220 U287 ( .A(A[19]), .B(n185), .C(A[20]), .D(n186), .Q(n187) );
  AOI220 U288 ( .A(A[19]), .B(n7), .C(A[20]), .D(n184), .Q(n222) );
  AOI220 U289 ( .A(A[18]), .B(n14), .C(A[19]), .D(n184), .Q(n241) );
  AOI220 U290 ( .A(A[5]), .B(n185), .C(A[6]), .D(n186), .Q(n210) );
  AOI220 U291 ( .A(A[5]), .B(n12), .C(A[6]), .D(n184), .Q(n190) );
  AOI220 U292 ( .A(A[2]), .B(n185), .C(A[3]), .D(n186), .Q(n274) );
  AOI220 U293 ( .A(A[2]), .B(n7), .C(A[3]), .D(n184), .Q(n252) );
  AOI220 U294 ( .A(A[1]), .B(n10), .C(A[2]), .D(n184), .Q(n196) );
  AOI220 U295 ( .A(A[3]), .B(n7), .C(A[4]), .D(n184), .Q(n211) );
  AOI220 U296 ( .A(A[3]), .B(n185), .C(A[4]), .D(n186), .Q(n195) );
  AOI220 U297 ( .A(A[4]), .B(n185), .C(A[5]), .D(n186), .Q(n251) );
  AOI220 U298 ( .A(A[4]), .B(n7), .C(A[5]), .D(n184), .Q(n273) );
  AOI220 U299 ( .A(n12), .B(A[0]), .C(A[1]), .D(n184), .Q(n275) );
  OAI212 U300 ( .A(n85), .B(n22), .C(n86), .Q(B[4]) );
  CLKIN3 U301 ( .A(n121), .Q(n120) );
  CLKIN3 U302 ( .A(n25), .Q(n122) );
  CLKIN3 U303 ( .A(n141), .Q(n85) );
  CLKIN3 U304 ( .A(n93), .Q(n148) );
  CLKIN3 U305 ( .A(n109), .Q(n151) );
  CLKIN3 U306 ( .A(n145), .Q(n154) );
  CLKIN3 U307 ( .A(n158), .Q(n157) );
endmodule


module E_alu_DW01_add_13 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62;

  NOR23 U2 ( .A(A[2]), .B(B[2]), .Q(n36) );
  NAND21 U3 ( .A(n62), .B(n41), .Q(SUM[0]) );
  NAND33 U4 ( .A(n31), .B(n32), .C(n33), .Q(n23) );
  INV1 U5 ( .A(n23), .Q(n30) );
  NAND23 U6 ( .A(n17), .B(n18), .Q(n12) );
  NOR21 U7 ( .A(n36), .B(n41), .Q(n40) );
  NOR22 U8 ( .A(n42), .B(n43), .Q(n31) );
  NOR22 U9 ( .A(A[1]), .B(B[1]), .Q(n38) );
  NOR22 U10 ( .A(n5), .B(A[3]), .Q(n37) );
  CLKIN6 U11 ( .A(n6), .Q(n5) );
  CLKIN3 U12 ( .A(B[0]), .Q(n4) );
  AOI222 U13 ( .A(n5), .B(A[3]), .C(n34), .D(n35), .Q(n33) );
  AOI211 U14 ( .A(n27), .B(n23), .C(n28), .Q(n26) );
  NOR31 U15 ( .A(n46), .B(n36), .C(n44), .Q(n42) );
  NOR21 U16 ( .A(n44), .B(n45), .Q(n43) );
  NOR22 U17 ( .A(A[3]), .B(n5), .Q(n44) );
  NOR22 U18 ( .A(n36), .B(n37), .Q(n35) );
  XOR22 U19 ( .A(n25), .B(n26), .Q(SUM[5]) );
  XOR22 U20 ( .A(n9), .B(n10), .Q(SUM[7]) );
  AOI212 U21 ( .A(n11), .B(n12), .C(n13), .Q(n10) );
  INV1 U22 ( .A(n36), .Q(n51) );
  NOR20 U23 ( .A(n53), .B(n36), .Q(n52) );
  AOI222 U24 ( .A(B[5]), .B(A[5]), .C(n22), .D(n23), .Q(n17) );
  AOI210 U25 ( .A(n6), .B(n8), .C(n38), .Q(n39) );
  INV0 U26 ( .A(n21), .Q(n28) );
  XOR20 U27 ( .A(n56), .B(n58), .Q(SUM[1]) );
  CLKIN2 U28 ( .A(B[3]), .Q(n6) );
  NOR20 U29 ( .A(A[0]), .B(n3), .Q(n61) );
  NAND20 U30 ( .A(n3), .B(A[0]), .Q(n60) );
  INV0 U31 ( .A(B[6]), .Q(n15) );
  NOR20 U32 ( .A(n59), .B(n38), .Q(n58) );
  XNR21 U33 ( .A(n47), .B(n1), .Q(SUM[3]) );
  XNR20 U34 ( .A(n5), .B(A[3]), .Q(n1) );
  XOR20 U35 ( .A(n50), .B(n52), .Q(SUM[2]) );
  CLKIN0 U36 ( .A(n38), .Q(n57) );
  NOR20 U37 ( .A(A[4]), .B(B[4]), .Q(n24) );
  NAND20 U38 ( .A(B[1]), .B(A[1]), .Q(n46) );
  NAND20 U39 ( .A(B[4]), .B(A[4]), .Q(n21) );
  NAND20 U40 ( .A(B[1]), .B(A[1]), .Q(n54) );
  NAND20 U41 ( .A(B[2]), .B(A[2]), .Q(n48) );
  XNR20 U42 ( .A(n2), .B(n12), .Q(SUM[6]) );
  XNR20 U43 ( .A(B[6]), .B(A[6]), .Q(n2) );
  XNR20 U44 ( .A(B[5]), .B(A[5]), .Q(n25) );
  INV0 U45 ( .A(n24), .Q(n27) );
  NAND20 U46 ( .A(A[2]), .B(B[2]), .Q(n45) );
  XNR20 U47 ( .A(B[4]), .B(A[4]), .Q(n29) );
  NOR20 U48 ( .A(A[6]), .B(B[6]), .Q(n16) );
  NAND22 U49 ( .A(n60), .B(n61), .Q(n56) );
  NAND22 U50 ( .A(n7), .B(n4), .Q(n62) );
  INV3 U51 ( .A(n4), .Q(n3) );
  INV3 U52 ( .A(A[0]), .Q(n7) );
  INV3 U53 ( .A(A[3]), .Q(n8) );
  NAND22 U54 ( .A(n39), .B(n40), .Q(n32) );
  AOI211 U55 ( .A(n7), .B(n4), .C(n38), .Q(n34) );
  NAND22 U56 ( .A(n3), .B(A[0]), .Q(n41) );
  NAND22 U57 ( .A(n54), .B(n55), .Q(n50) );
  NAND22 U58 ( .A(n56), .B(n57), .Q(n55) );
  XNR21 U59 ( .A(B[7]), .B(A[7]), .Q(n9) );
  NOR21 U60 ( .A(n14), .B(n15), .Q(n13) );
  NOR21 U61 ( .A(n20), .B(n24), .Q(n22) );
  NAND22 U62 ( .A(n48), .B(n49), .Q(n47) );
  NAND22 U63 ( .A(n50), .B(n51), .Q(n49) );
  NOR21 U64 ( .A(A[5]), .B(B[5]), .Q(n20) );
  INV3 U65 ( .A(n19), .Q(n18) );
  NOR21 U66 ( .A(n20), .B(n21), .Q(n19) );
  XOR21 U67 ( .A(n29), .B(n30), .Q(SUM[4]) );
  INV3 U68 ( .A(n16), .Q(n11) );
  INV3 U69 ( .A(A[6]), .Q(n14) );
  CLKIN3 U70 ( .A(n48), .Q(n53) );
  CLKIN3 U71 ( .A(n54), .Q(n59) );
endmodule


module E_alu_DW01_add_12 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55;

  NAND22 U2 ( .A(B[1]), .B(A[1]), .Q(n48) );
  NOR21 U3 ( .A(A[3]), .B(B[3]), .Q(n39) );
  NOR21 U4 ( .A(n37), .B(n38), .Q(n29) );
  AOI211 U5 ( .A(n7), .B(n8), .C(n33), .Q(n34) );
  NOR22 U6 ( .A(n32), .B(n36), .Q(n35) );
  NAND23 U7 ( .A(n17), .B(n18), .Q(n12) );
  NOR22 U8 ( .A(A[1]), .B(B[1]), .Q(n33) );
  NOR20 U9 ( .A(n53), .B(n33), .Q(n52) );
  CLKIN3 U10 ( .A(n33), .Q(n51) );
  AOI222 U11 ( .A(B[5]), .B(A[5]), .C(n22), .D(n23), .Q(n17) );
  NOR31 U12 ( .A(n48), .B(n32), .C(n39), .Q(n37) );
  NOR20 U13 ( .A(n47), .B(n32), .Q(n46) );
  INV0 U14 ( .A(n32), .Q(n45) );
  AOI211 U15 ( .A(n27), .B(n23), .C(n28), .Q(n26) );
  NAND24 U16 ( .A(n29), .B(n2), .Q(n23) );
  NOR21 U17 ( .A(n20), .B(n21), .Q(n19) );
  NAND20 U18 ( .A(B[3]), .B(A[3]), .Q(n31) );
  NAND22 U19 ( .A(n30), .B(n31), .Q(n1) );
  CLKIN3 U20 ( .A(n1), .Q(n2) );
  NAND22 U21 ( .A(n34), .B(n35), .Q(n30) );
  CLKIN2 U22 ( .A(B[3]), .Q(n7) );
  INV0 U23 ( .A(n21), .Q(n28) );
  MUX21 U24 ( .A(B[0]), .B(n55), .S(A[0]), .Q(SUM[0]) );
  INV0 U25 ( .A(B[6]), .Q(n15) );
  NAND20 U26 ( .A(B[0]), .B(A[0]), .Q(n54) );
  INV0 U27 ( .A(B[0]), .Q(n55) );
  XNR21 U28 ( .A(n41), .B(n4), .Q(SUM[3]) );
  XNR20 U29 ( .A(B[3]), .B(A[3]), .Q(n4) );
  NOR22 U30 ( .A(A[2]), .B(B[2]), .Q(n32) );
  NOR20 U31 ( .A(A[4]), .B(B[4]), .Q(n24) );
  NOR20 U32 ( .A(A[5]), .B(B[5]), .Q(n20) );
  NAND20 U33 ( .A(B[4]), .B(A[4]), .Q(n21) );
  NAND20 U34 ( .A(B[2]), .B(A[2]), .Q(n42) );
  XNR20 U35 ( .A(n5), .B(n12), .Q(SUM[6]) );
  XNR20 U36 ( .A(B[6]), .B(A[6]), .Q(n5) );
  XNR20 U37 ( .A(B[5]), .B(A[5]), .Q(n25) );
  INV0 U38 ( .A(n24), .Q(n27) );
  XNR20 U39 ( .A(n6), .B(n23), .Q(SUM[4]) );
  XNR20 U40 ( .A(B[4]), .B(A[4]), .Q(n6) );
  NAND20 U41 ( .A(A[2]), .B(B[2]), .Q(n40) );
  NOR20 U42 ( .A(A[6]), .B(B[6]), .Q(n16) );
  INV3 U43 ( .A(n54), .Q(n50) );
  XOR21 U44 ( .A(n44), .B(n46), .Q(SUM[2]) );
  INV3 U45 ( .A(A[3]), .Q(n8) );
  NAND22 U46 ( .A(B[0]), .B(A[0]), .Q(n36) );
  XOR21 U47 ( .A(n9), .B(n10), .Q(SUM[7]) );
  XNR21 U48 ( .A(B[7]), .B(A[7]), .Q(n9) );
  AOI211 U49 ( .A(n11), .B(n12), .C(n13), .Q(n10) );
  NOR21 U50 ( .A(n14), .B(n15), .Q(n13) );
  NAND22 U51 ( .A(n42), .B(n43), .Q(n41) );
  NAND22 U52 ( .A(n44), .B(n45), .Q(n43) );
  NAND22 U53 ( .A(n48), .B(n49), .Q(n44) );
  NAND22 U54 ( .A(n50), .B(n51), .Q(n49) );
  NOR21 U55 ( .A(n20), .B(n24), .Q(n22) );
  XOR21 U56 ( .A(n50), .B(n52), .Q(SUM[1]) );
  XOR21 U57 ( .A(n25), .B(n26), .Q(SUM[5]) );
  NOR21 U58 ( .A(n39), .B(n40), .Q(n38) );
  INV3 U59 ( .A(n19), .Q(n18) );
  INV3 U60 ( .A(n16), .Q(n11) );
  INV3 U61 ( .A(A[6]), .Q(n14) );
  CLKIN3 U62 ( .A(n42), .Q(n47) );
  CLKIN3 U63 ( .A(n48), .Q(n53) );
endmodule


module E_alu ( o_data_AluRes, i_data_A, i_data_B, i_con_AluCtrl, i_data_shamt
 );
  output [31:0] o_data_AluRes;
  input [31:0] i_data_A;
  input [31:0] i_data_B;
  input [3:0] i_con_AluCtrl;
  input [4:0] i_data_shamt;
  wire   N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N321, n42, n43,
         n140, n220, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558;
  wire   [8:0] sum_1;
  wire   [8:0] pre_sum_2a;
  wire   [8:0] pre_sum_2b;
  wire   [8:0] pre_sum_3a;
  wire   [8:0] pre_sum_3b;
  wire   [7:0] pre_sum_4a;
  wire   [7:0] pre_sum_4b;
  wire   [16:0] half_sub;
  wire   [15:0] pre_suba;
  wire   [15:0] pre_subb;

  E_alu_DW01_ash_0 sll_55 ( .A({n70, n68, n67, n66, n82, n30, n65, n81, n80, 
        n63, n62, n79, n78, n61, n60, n77, n59, n57, n56, n76, n54, n75, n53, 
        n74, n38, i_data_B[6:5], n37, i_data_B[3], n41, i_data_B[1], n5}), 
        .DATA_TC(n43), .SH(i_data_shamt), .SH_TC(n43), .B({N239, N238, N237, 
        N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, 
        N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, 
        N212, N211, N210, N209, N208}) );
  E_alu_DW01_cmp2_1 r131 ( .A(i_data_A), .B({n69, n68, n67, n66, n82, n30, n64, 
        n81, n80, n63, n62, n79, n78, n61, n60, n77, n59, n57, n56, n76, n55, 
        n75, n53, n74, n38, i_data_B[6:5], n37, i_data_B[3], n41, i_data_B[1], 
        n5}), .LEQ(n43), .TC(n43), .LT_LE(N321) );
  E_alu_DW01_sub_3 sub_33 ( .A({n43, i_data_A[15:0]}), .B({n43, n58, n57, n56, 
        n76, n54, n75, n53, n74, i_data_B[7:5], n37, i_data_B[3:1], n5}), .CI(
        n43), .DIFF(half_sub) );
  E_alu_DW01_sub_5 sub_1_root_sub_35_2 ( .A(i_data_A[31:16]), .B({n70, n68, 
        n67, n66, n82, n31, n65, n81, n80, n63, n62, n79, n78, n61, n60, n77}), 
        .CI(n42), .DIFF(pre_subb) );
  E_alu_DW01_sub_4 sub_34 ( .A(i_data_A[31:16]), .B({n70, n68, n67, n66, n82, 
        n30, n65, n81, n80, n63, n62, n79, n78, n61, n60, n77}), .CI(n43), 
        .DIFF(pre_suba) );
  E_alu_DW01_add_8 add_25 ( .A({n43, i_data_A[7:0]}), .B({n43, i_data_B[7:5], 
        n37, i_data_B[3:1], n5}), .CI(n43), .SUM(sum_1) );
  E_alu_DW01_add_7 add_1_root_add_27_2 ( .A({n43, i_data_A[15:8]}), .B({n43, 
        n58, n57, n56, n76, n55, n75, n53, n74}), .CI(n42), .SUM(pre_sum_2b)
         );
  E_alu_DW01_add_9 add_26 ( .A({n43, i_data_A[15:8]}), .B({n43, n58, n57, n56, 
        n76, n54, n75, n53, n74}), .CI(n43), .SUM(pre_sum_2a) );
  E_alu_DW01_add_10 add_1_root_add_29_2 ( .A({n43, i_data_A[23:16]}), .B({n43, 
        n80, n63, n62, n79, n78, n61, n60, n77}), .CI(n42), .SUM(pre_sum_3b)
         );
  E_alu_DW01_add_11 add_28 ( .A({n43, i_data_A[23:16]}), .B({n43, n80, n63, 
        n62, n79, n78, n61, n60, n77}), .CI(n43), .SUM(pre_sum_3a) );
  E_alu_DW_rash_1 r130 ( .A({n69, n68, n67, n66, n82, n31, n65, n81, n80, n63, 
        n62, n79, n78, n61, n60, n77, n59, n57, n56, n76, n55, n75, n53, n74, 
        n38, i_data_B[6:5], n37, i_data_B[3], n41, i_data_B[1], n5}), 
        .DATA_TC(n43), .SH(i_data_shamt), .SH_TC(n43), .B({N271, N270, N269, 
        N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, 
        N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, 
        N244, N243, N242, N241, N240}) );
  E_alu_DW01_add_13 add_1_root_add_31_2 ( .A(i_data_A[31:24]), .B({n70, n68, 
        n67, n66, n82, n30, n64, n81}), .CI(n42), .SUM(pre_sum_4b) );
  E_alu_DW01_add_12 add_30 ( .A(i_data_A[31:24]), .B({n70, n68, n67, n66, n82, 
        n30, n64, n81}), .CI(n43), .SUM(pre_sum_4a) );
  AOI211 U3 ( .A(n521), .B(n73), .C(n71), .Q(n522) );
  NAND34 U4 ( .A(n39), .B(i_con_AluCtrl[1]), .C(n112), .Q(n548) );
  INV2 U5 ( .A(n111), .Q(n112) );
  IMUX20 U6 ( .A(n172), .B(n171), .S(i_data_B[5]), .Q(n181) );
  INV2 U7 ( .A(i_data_B[5]), .Q(n382) );
  OAI211 U8 ( .A(n356), .B(n71), .C(i_data_A[19]), .Q(n358) );
  CLKIN12 U9 ( .A(i_con_AluCtrl[3]), .Q(n103) );
  IMUX22 U10 ( .A(n475), .B(n474), .S(n82), .Q(n481) );
  NOR23 U11 ( .A(n530), .B(n529), .Q(n534) );
  NOR20 U12 ( .A(n135), .B(n98), .Q(n99) );
  OAI222 U13 ( .A(n210), .B(n83), .C(n271), .D(n209), .Q(n211) );
  IMUX22 U14 ( .A(n48), .B(n535), .S(n82), .Q(n476) );
  CLKBU4 U15 ( .A(n558), .Q(n48) );
  NAND22 U16 ( .A(n40), .B(n100), .Q(n135) );
  IMUX22 U17 ( .A(n72), .B(n489), .S(n61), .Q(n339) );
  AOI212 U18 ( .A(n3), .B(n383), .C(n390), .Q(n384) );
  INV6 U19 ( .A(n271), .Q(n233) );
  OAI2112 U20 ( .A(n548), .B(n452), .C(n451), .D(n450), .Q(n453) );
  AOI212 U21 ( .A(n52), .B(n108), .C(n107), .Q(n109) );
  NOR22 U22 ( .A(n454), .B(n453), .Q(n458) );
  NAND23 U23 ( .A(sum_1[8]), .B(n437), .Q(n243) );
  INV15 U24 ( .A(n440), .Q(n437) );
  NOR23 U25 ( .A(n381), .B(n341), .Q(n342) );
  NOR32 U26 ( .A(i_con_AluCtrl[3]), .B(i_con_AluCtrl[1]), .C(i_con_AluCtrl[2]), 
        .Q(n272) );
  NAND31 U27 ( .A(i_data_A[28]), .B(n489), .C(n66), .Q(n495) );
  NAND31 U28 ( .A(i_data_A[26]), .B(n489), .C(n31), .Q(n463) );
  IMUX21 U29 ( .A(n73), .B(n489), .S(n5), .Q(n108) );
  IMUX21 U30 ( .A(n73), .B(n489), .S(n79), .Q(n368) );
  INV8 U31 ( .A(n535), .Q(n489) );
  NAND26 U32 ( .A(half_sub[16]), .B(n486), .Q(n381) );
  NAND24 U33 ( .A(n310), .B(n100), .Q(n440) );
  CLKIN3 U34 ( .A(n90), .Q(n96) );
  IMUX21 U35 ( .A(n106), .B(n105), .S(n5), .Q(n110) );
  INV8 U36 ( .A(i_con_AluCtrl[1]), .Q(n97) );
  BUF8 U37 ( .A(i_data_B[29]), .Q(n67) );
  BUF8 U38 ( .A(i_data_B[2]), .Q(n41) );
  BUF6 U39 ( .A(i_data_B[15]), .Q(n58) );
  IMUX21 U40 ( .A(n319), .B(n318), .S(n77), .Q(n320) );
  INV8 U41 ( .A(n272), .Q(n535) );
  INV3 U42 ( .A(n243), .Q(n297) );
  AOI211 U43 ( .A(N226), .B(n499), .C(n348), .Q(n349) );
  INV12 U44 ( .A(n387), .Q(n538) );
  BUF12 U45 ( .A(i_data_B[4]), .Q(n37) );
  NOR23 U46 ( .A(n116), .B(n115), .Q(n117) );
  NOR21 U47 ( .A(n250), .B(n249), .Q(n251) );
  NOR21 U48 ( .A(n264), .B(n263), .Q(n265) );
  AOI211 U49 ( .A(half_sub[12]), .B(n486), .C(n255), .Q(n267) );
  INV3 U50 ( .A(n28), .Q(n29) );
  CLKBU4 U51 ( .A(i_data_B[26]), .Q(n31) );
  INV6 U52 ( .A(n8), .Q(n9) );
  INV6 U53 ( .A(sum_1[8]), .Q(n12) );
  OAI221 U54 ( .A(n542), .B(n46), .C(n541), .D(n540), .Q(n543) );
  NAND22 U55 ( .A(i_data_B[1]), .B(n524), .Q(n330) );
  BUF12 U56 ( .A(i_data_B[11]), .Q(n55) );
  NAND33 U57 ( .A(n429), .B(n428), .C(n427), .Q(o_data_AluRes[23]) );
  INV15 U58 ( .A(n308), .Q(n551) );
  NOR21 U59 ( .A(n208), .B(n71), .Q(n210) );
  AOI212 U60 ( .A(n107), .B(n72), .C(n71), .Q(n105) );
  NOR22 U61 ( .A(n110), .B(n109), .Q(n114) );
  CLKIN12 U62 ( .A(i_con_AluCtrl[2]), .Q(n310) );
  AOI220 U63 ( .A(pre_sum_3b[2]), .B(n418), .C(pre_suba[2]), .D(n551), .Q(n352) );
  AOI221 U64 ( .A(pre_sum_3b[7]), .B(n418), .C(pre_suba[7]), .D(n551), .Q(n428) );
  AOI220 U65 ( .A(pre_sum_3b[4]), .B(n418), .C(pre_suba[4]), .D(n551), .Q(n380) );
  CLKIN6 U66 ( .A(n541), .Q(n524) );
  CLKIN12 U67 ( .A(n438), .Q(n552) );
  OAI212 U68 ( .A(n476), .B(n71), .C(i_data_A[27]), .Q(n477) );
  NAND24 U69 ( .A(n12), .B(pre_sum_2a[8]), .Q(n13) );
  NAND21 U70 ( .A(n87), .B(n520), .Q(n375) );
  NAND23 U71 ( .A(n501), .B(n500), .Q(n502) );
  NAND32 U72 ( .A(n503), .B(n504), .C(n36), .Q(o_data_AluRes[28]) );
  CLKBU12 U73 ( .A(i_data_B[8]), .Q(n74) );
  OAI222 U74 ( .A(n177), .B(n176), .C(n387), .D(n175), .Q(n178) );
  NOR21 U75 ( .A(n174), .B(n71), .Q(n177) );
  CLKBU15 U76 ( .A(i_data_B[18]), .Q(n61) );
  INV10 U77 ( .A(n46), .Q(n72) );
  NAND21 U78 ( .A(n507), .B(n520), .Q(n509) );
  NAND21 U79 ( .A(n466), .B(n520), .Q(n468) );
  NAND24 U80 ( .A(n103), .B(n96), .Q(n387) );
  NAND21 U81 ( .A(n89), .B(n520), .Q(n475) );
  NAND21 U82 ( .A(n345), .B(n520), .Q(n347) );
  INV15 U83 ( .A(n49), .Q(n520) );
  BUF15 U84 ( .A(i_data_B[20]), .Q(n79) );
  NAND23 U85 ( .A(n311), .B(n15), .Q(n541) );
  NAND33 U86 ( .A(n397), .B(n396), .C(n398), .Q(n10) );
  BUF6 U87 ( .A(i_data_B[25]), .Q(n65) );
  INV3 U88 ( .A(n147), .Q(n150) );
  INV3 U89 ( .A(N238), .Q(n528) );
  BUF6 U90 ( .A(i_data_B[25]), .Q(n64) );
  BUF6 U91 ( .A(i_data_B[15]), .Q(n59) );
  BUF12 U92 ( .A(i_data_B[23]), .Q(n80) );
  NOR21 U93 ( .A(n50), .B(i_data_A[23]), .Q(n420) );
  BUF6 U94 ( .A(n140), .Q(n49) );
  BUF12 U95 ( .A(i_con_AluCtrl[0]), .Q(n39) );
  BUF6 U96 ( .A(i_data_B[7]), .Q(n38) );
  CLKBU12 U97 ( .A(i_data_B[11]), .Q(n54) );
  BUF12 U98 ( .A(i_data_B[14]), .Q(n57) );
  AOI221 U99 ( .A(pre_sum_3b[0]), .B(n418), .C(pre_suba[0]), .D(n551), .Q(n324) );
  NOR21 U100 ( .A(n164), .B(n163), .Q(n170) );
  NOR21 U101 ( .A(n157), .B(n156), .Q(n158) );
  NAND31 U102 ( .A(n267), .B(n266), .C(n265), .Q(o_data_AluRes[12]) );
  NAND22 U103 ( .A(n304), .B(n7), .Q(o_data_AluRes[15]) );
  AOI221 U104 ( .A(N255), .B(n538), .C(pre_sum_2b[7]), .D(n297), .Q(n304) );
  NAND22 U105 ( .A(n395), .B(n11), .Q(o_data_AluRes[21]) );
  AOI2111 U106 ( .A(N229), .B(n499), .C(n394), .D(n393), .Q(n395) );
  INV3 U107 ( .A(n10), .Q(n11) );
  NAND31 U108 ( .A(n412), .B(n411), .C(n410), .Q(o_data_AluRes[22]) );
  AOI211 U109 ( .A(pre_subb[8]), .B(n550), .C(n436), .Q(n443) );
  NAND22 U110 ( .A(pre_suba[15]), .B(n551), .Q(n556) );
  AOI221 U111 ( .A(sum_1[6]), .B(n437), .C(half_sub[6]), .D(n486), .Q(n193) );
  NOR22 U112 ( .A(n381), .B(n370), .Q(n371) );
  CLKBU12 U113 ( .A(i_data_B[30]), .Q(n68) );
  INV12 U114 ( .A(n4), .Q(n5) );
  INV6 U115 ( .A(n104), .Q(n51) );
  CLKBU12 U116 ( .A(i_data_B[12]), .Q(n76) );
  CLKBU12 U117 ( .A(i_data_B[17]), .Q(n60) );
  INV3 U118 ( .A(i_data_B[0]), .Q(n4) );
  IMUX22 U119 ( .A(n488), .B(n487), .S(n66), .Q(n498) );
  IMUX21 U120 ( .A(n46), .B(n535), .S(n65), .Q(n449) );
  OAI2112 U121 ( .A(n548), .B(n513), .C(n511), .D(n512), .Q(n514) );
  NOR22 U122 ( .A(n515), .B(n514), .Q(n519) );
  NOR23 U123 ( .A(n481), .B(n480), .Q(n485) );
  NAND24 U124 ( .A(pre_sum_4a[5]), .B(n552), .Q(n517) );
  AOI221 U125 ( .A(N258), .B(n538), .C(pre_sum_3a[2]), .D(n426), .Q(n350) );
  BUF8 U126 ( .A(n51), .Q(n3) );
  INV0 U127 ( .A(n103), .Q(n1) );
  OAI211 U128 ( .A(n510), .B(n71), .C(i_data_A[29]), .Q(n511) );
  AOI211 U129 ( .A(n87), .B(n73), .C(n71), .Q(n374) );
  CLKBU4 U130 ( .A(n553), .Q(n2) );
  IMUX21 U131 ( .A(n73), .B(n489), .S(n59), .Q(n295) );
  AOI212 U132 ( .A(pre_subb[15]), .B(n550), .C(n549), .Q(n557) );
  AOI211 U133 ( .A(n507), .B(n73), .C(n71), .Q(n508) );
  AOI210 U134 ( .A(n122), .B(n73), .C(n71), .Q(n123) );
  NAND26 U135 ( .A(n307), .B(n486), .Q(n308) );
  NAND22 U136 ( .A(n310), .B(n312), .Q(n14) );
  CLKIN3 U137 ( .A(n310), .Q(n40) );
  NAND24 U138 ( .A(n518), .B(n27), .Q(o_data_AluRes[29]) );
  OAI222 U139 ( .A(n243), .B(n217), .C(n387), .D(n216), .Q(n222) );
  OAI210 U140 ( .A(n46), .B(i_data_A[23]), .C(n51), .Q(n419) );
  IMUX20 U141 ( .A(n46), .B(n535), .S(i_data_B[5]), .Q(n174) );
  NAND31 U142 ( .A(n253), .B(n252), .C(n251), .Q(o_data_AluRes[11]) );
  NAND24 U143 ( .A(n517), .B(n516), .Q(n18) );
  AOI212 U144 ( .A(pre_sum_2a[6]), .B(n233), .C(n285), .Q(n293) );
  NAND21 U145 ( .A(n317), .B(n437), .Q(n361) );
  AOI211 U146 ( .A(n76), .B(n524), .C(n492), .Q(n493) );
  AOI212 U147 ( .A(N234), .B(n499), .C(n465), .Q(n473) );
  NAND26 U148 ( .A(n553), .B(pre_sum_4b[5]), .Q(n516) );
  OAI2112 U149 ( .A(n548), .B(n528), .C(n527), .D(n526), .Q(n529) );
  OAI211 U150 ( .A(n525), .B(n71), .C(i_data_A[30]), .Q(n526) );
  NAND32 U151 ( .A(n238), .B(n237), .C(n236), .Q(o_data_AluRes[10]) );
  AOI221 U152 ( .A(N218), .B(n499), .C(half_sub[10]), .D(n486), .Q(n236) );
  IMUX21 U153 ( .A(n73), .B(n489), .S(n62), .Q(n383) );
  OAI210 U154 ( .A(n47), .B(i_data_A[14]), .C(n52), .Q(n288) );
  OAI210 U155 ( .A(n47), .B(i_data_A[6]), .C(n3), .Q(n183) );
  OAI210 U156 ( .A(n47), .B(i_data_A[5]), .C(n52), .Q(n171) );
  OAI210 U157 ( .A(n47), .B(i_data_A[10]), .C(n52), .Q(n234) );
  OAI210 U158 ( .A(n47), .B(i_data_A[13]), .C(n52), .Q(n278) );
  OAI210 U159 ( .A(n47), .B(i_data_A[9]), .C(n3), .Q(n223) );
  OAI210 U160 ( .A(n47), .B(i_data_A[12]), .C(n3), .Q(n256) );
  AOI210 U161 ( .A(n3), .B(n219), .C(n218), .Q(n221) );
  AOI212 U162 ( .A(pre_sum_2a[7]), .B(n233), .C(n296), .Q(n305) );
  INV6 U163 ( .A(n26), .Q(n27) );
  IMUX22 U164 ( .A(n433), .B(n432), .S(n81), .Q(n434) );
  AOI211 U165 ( .A(half_sub[11]), .B(n486), .C(n240), .Q(n253) );
  INV3 U166 ( .A(n239), .Q(n240) );
  AOI221 U167 ( .A(N256), .B(n538), .C(pre_sum_3a[0]), .D(n426), .Q(n322) );
  IMUX20 U168 ( .A(n46), .B(n535), .S(n74), .Q(n208) );
  BUF6 U169 ( .A(n140), .Q(n50) );
  NAND33 U170 ( .A(n40), .B(n311), .C(n312), .Q(n140) );
  AOI221 U171 ( .A(n56), .B(n524), .C(N269), .D(n538), .Q(n512) );
  NAND21 U172 ( .A(pre_sum_4a[6]), .B(n552), .Q(n532) );
  AOI211 U173 ( .A(pre_sum_4a[4]), .B(n552), .C(n502), .Q(n503) );
  NAND21 U174 ( .A(pre_sum_4a[7]), .B(n552), .Q(n555) );
  NAND23 U175 ( .A(n441), .B(n437), .Q(n438) );
  OAI211 U176 ( .A(n329), .B(n71), .C(i_data_A[17]), .Q(n331) );
  INV4 U177 ( .A(n44), .Q(n45) );
  NAND24 U178 ( .A(n114), .B(n113), .Q(n115) );
  AOI221 U179 ( .A(half_sub[8]), .B(n486), .C(N216), .D(n499), .Q(n215) );
  CLKIN4 U180 ( .A(half_sub[16]), .Q(n307) );
  INV12 U181 ( .A(n39), .Q(n312) );
  NAND26 U182 ( .A(n310), .B(n103), .Q(n111) );
  AOI2111 U183 ( .A(pre_subb[6]), .B(n550), .C(n402), .D(n401), .Q(n412) );
  AOI222 U184 ( .A(N254), .B(n538), .C(pre_sum_2b[6]), .D(n297), .Q(n292) );
  NAND21 U185 ( .A(pre_sum_4b[6]), .B(n2), .Q(n531) );
  AOI220 U186 ( .A(pre_sum_4a[0]), .B(n552), .C(pre_sum_4b[0]), .D(n553), .Q(
        n442) );
  NAND21 U187 ( .A(n553), .B(pre_sum_4b[7]), .Q(n554) );
  AOI2111 U188 ( .A(N230), .B(n499), .C(n409), .D(n408), .Q(n410) );
  NOR23 U189 ( .A(n498), .B(n497), .Q(n501) );
  OAI210 U190 ( .A(n260), .B(n71), .C(i_data_A[12]), .Q(n262) );
  AOI210 U191 ( .A(n151), .B(n72), .C(n71), .Q(n152) );
  AOI210 U192 ( .A(n446), .B(n73), .C(n71), .Q(n447) );
  NAND21 U193 ( .A(n553), .B(pre_sum_4b[1]), .Q(n455) );
  NAND22 U194 ( .A(n52), .B(n339), .Q(n344) );
  AOI212 U195 ( .A(half_sub[15]), .B(n486), .C(n299), .Q(n303) );
  AOI212 U196 ( .A(half_sub[14]), .B(n486), .C(n287), .Q(n291) );
  NOR20 U197 ( .A(n381), .B(n313), .Q(n314) );
  CLKIN12 U198 ( .A(n381), .Q(n550) );
  AOI221 U199 ( .A(sum_1[7]), .B(n437), .C(half_sub[7]), .D(n486), .Q(n203) );
  AOI221 U200 ( .A(n54), .B(n524), .C(N267), .D(n538), .Q(n478) );
  IMUX22 U201 ( .A(N321), .B(i_data_A[31]), .S(n93), .Q(n120) );
  NAND21 U202 ( .A(n85), .B(n520), .Q(n319) );
  CLKIN3 U203 ( .A(N237), .Q(n513) );
  INV12 U204 ( .A(n317), .Q(n439) );
  NOR24 U205 ( .A(n440), .B(n441), .Q(n553) );
  AOI210 U206 ( .A(n3), .B(n148), .C(n151), .Q(n149) );
  NAND22 U207 ( .A(sum_1[3]), .B(n437), .Q(n154) );
  CLKBU15 U208 ( .A(i_data_B[27]), .Q(n82) );
  NAND21 U209 ( .A(n107), .B(n520), .Q(n106) );
  NAND21 U210 ( .A(n491), .B(n520), .Q(n488) );
  IMUX21 U211 ( .A(n347), .B(n346), .S(n61), .Q(n348) );
  NAND22 U212 ( .A(n505), .B(n506), .Q(n35) );
  AOI211 U213 ( .A(n85), .B(n73), .C(n71), .Q(n318) );
  CLKIN3 U214 ( .A(n104), .Q(n52) );
  NAND21 U215 ( .A(pre_sum_4a[3]), .B(n552), .Q(n483) );
  AOI2111 U216 ( .A(pre_suba[3]), .B(n551), .C(n363), .D(n362), .Q(n364) );
  AOI2112 U217 ( .A(pre_sum_3a[7]), .B(n426), .C(n425), .D(n424), .Q(n427) );
  OAI2112 U218 ( .A(n381), .B(n332), .C(n331), .D(n330), .Q(n335) );
  IMUX24 U219 ( .A(pre_sum_3b[8]), .B(pre_sum_3a[8]), .S(n439), .Q(n441) );
  NAND42 U220 ( .A(n464), .B(n463), .C(n462), .D(n461), .Q(n465) );
  AOI210 U221 ( .A(n75), .B(n524), .C(n460), .Q(n461) );
  NAND42 U222 ( .A(n496), .B(n495), .C(n494), .D(n493), .Q(n497) );
  NAND33 U223 ( .A(n350), .B(n349), .C(n351), .Q(n8) );
  BUF12 U224 ( .A(i_data_B[22]), .Q(n63) );
  NAND31 U225 ( .A(pre_subb[12]), .B(half_sub[16]), .C(n486), .Q(n505) );
  BUF8 U226 ( .A(i_data_B[26]), .Q(n30) );
  NAND26 U227 ( .A(n96), .B(n91), .Q(n558) );
  CLKBU4 U228 ( .A(n558), .Q(n47) );
  INV15 U229 ( .A(n46), .Q(n73) );
  BUF15 U230 ( .A(i_data_B[9]), .Q(n53) );
  AOI212 U231 ( .A(N224), .B(n499), .C(n320), .Q(n321) );
  BUF12 U232 ( .A(i_data_B[21]), .Q(n62) );
  NAND21 U233 ( .A(n535), .B(n60), .Q(n24) );
  AOI222 U234 ( .A(pre_suba[11]), .B(n551), .C(pre_subb[11]), .D(n550), .Q(
        n484) );
  NOR21 U235 ( .A(n50), .B(i_data_A[24]), .Q(n433) );
  NOR21 U236 ( .A(n50), .B(i_data_A[15]), .Q(n301) );
  OAI220 U237 ( .A(n47), .B(n137), .C(i_data_A[2]), .D(n50), .Q(n220) );
  AOI2112 U238 ( .A(i_data_A[18]), .B(n344), .C(n343), .D(n342), .Q(n351) );
  IMUX21 U239 ( .A(n46), .B(n535), .S(n67), .Q(n510) );
  NAND26 U240 ( .A(pre_sum_2b[8]), .B(sum_1[8]), .Q(n306) );
  BUF12 U241 ( .A(i_data_B[28]), .Q(n66) );
  CLKBU15 U242 ( .A(i_data_B[13]), .Q(n56) );
  NAND33 U243 ( .A(n303), .B(n305), .C(n302), .Q(n6) );
  CLKIN6 U244 ( .A(n6), .Q(n7) );
  NAND22 U245 ( .A(n352), .B(n9), .Q(o_data_AluRes[18]) );
  INV6 U246 ( .A(n34), .Q(n418) );
  NAND22 U247 ( .A(pre_sum_3b[5]), .B(n418), .Q(n397) );
  AOI2112 U248 ( .A(pre_subb[5]), .B(n550), .C(n385), .D(n384), .Q(n396) );
  OAI2112 U249 ( .A(n548), .B(n479), .C(n478), .D(n477), .Q(n480) );
  NAND28 U250 ( .A(n13), .B(n306), .Q(n317) );
  NAND22 U251 ( .A(i_con_AluCtrl[3]), .B(n97), .Q(n92) );
  CLKIN15 U252 ( .A(n51), .Q(n71) );
  INV3 U253 ( .A(n14), .Q(n15) );
  NOR24 U254 ( .A(i_con_AluCtrl[1]), .B(n111), .Q(n16) );
  NOR24 U255 ( .A(n17), .B(n312), .Q(n104) );
  INV6 U256 ( .A(n16), .Q(n17) );
  NAND24 U257 ( .A(n519), .B(n19), .Q(n26) );
  INV6 U258 ( .A(n18), .Q(n19) );
  AOI222 U259 ( .A(pre_suba[13]), .B(n551), .C(pre_subb[13]), .D(n550), .Q(
        n518) );
  NAND22 U260 ( .A(n95), .B(n94), .Q(n20) );
  NAND22 U261 ( .A(N321), .B(n21), .Q(n118) );
  INV3 U262 ( .A(n20), .Q(n21) );
  OAI2112 U263 ( .A(n120), .B(n119), .C(n118), .D(n117), .Q(o_data_AluRes[0])
         );
  NOR21 U264 ( .A(n34), .B(n333), .Q(n334) );
  NAND33 U265 ( .A(n483), .B(n485), .C(n484), .Q(n28) );
  NAND20 U266 ( .A(n558), .B(n22), .Q(n23) );
  NAND22 U267 ( .A(n23), .B(n24), .Q(n25) );
  INV0 U268 ( .A(n60), .Q(n22) );
  INV3 U269 ( .A(n25), .Q(n329) );
  CLKBU15 U270 ( .A(n558), .Q(n46) );
  AOI221 U271 ( .A(pre_suba[14]), .B(n551), .C(pre_subb[14]), .D(n550), .Q(
        n533) );
  NAND22 U272 ( .A(n482), .B(n29), .Q(o_data_AluRes[27]) );
  NAND20 U273 ( .A(pre_sum_4b[3]), .B(n553), .Q(n482) );
  NAND22 U274 ( .A(n323), .B(n33), .Q(o_data_AluRes[16]) );
  NAND33 U275 ( .A(n324), .B(n321), .C(n322), .Q(n32) );
  NAND22 U276 ( .A(n12), .B(n437), .Q(n271) );
  NAND42 U277 ( .A(n534), .B(n533), .C(n532), .D(n531), .Q(o_data_AluRes[30])
         );
  AOI2111 U278 ( .A(pre_subb[7]), .B(n550), .C(n417), .D(n416), .Q(n429) );
  AOI2111 U279 ( .A(i_data_A[16]), .B(n316), .C(n315), .D(n314), .Q(n323) );
  NAND20 U280 ( .A(n3), .B(n309), .Q(n316) );
  IMUX21 U281 ( .A(n448), .B(n447), .S(n65), .Q(n454) );
  IMUX20 U282 ( .A(n224), .B(n223), .S(n53), .Q(n226) );
  INV3 U283 ( .A(n32), .Q(n33) );
  NAND42 U284 ( .A(n367), .B(n366), .C(n365), .D(n364), .Q(o_data_AluRes[19])
         );
  NAND22 U285 ( .A(N253), .B(n538), .Q(n268) );
  NAND22 U286 ( .A(pre_suba[12]), .B(n551), .Q(n506) );
  AOI2111 U287 ( .A(pre_suba[1]), .B(n551), .C(n335), .D(n334), .Q(n336) );
  AOI221 U288 ( .A(N217), .B(n499), .C(half_sub[9]), .D(n486), .Q(n225) );
  CLKBU15 U289 ( .A(i_data_B[16]), .Q(n77) );
  NAND20 U290 ( .A(pre_sum_3a[3]), .B(n426), .Q(n367) );
  BUF6 U291 ( .A(n361), .Q(n34) );
  INV6 U292 ( .A(n389), .Q(n426) );
  INV12 U293 ( .A(n135), .Q(n486) );
  AOI211 U294 ( .A(N228), .B(n499), .C(n376), .Q(n377) );
  NAND20 U295 ( .A(pre_sum_4a[1]), .B(n552), .Q(n456) );
  CLKIN0 U296 ( .A(n31), .Q(n459) );
  CLKIN0 U297 ( .A(n41), .Q(n340) );
  AOI2111 U298 ( .A(N211), .B(n499), .C(n150), .D(n149), .Q(n159) );
  NAND22 U299 ( .A(pre_sum_2b[5]), .B(n297), .Q(n269) );
  INV6 U300 ( .A(n92), .Q(n311) );
  NOR31 U301 ( .A(n277), .B(n276), .C(n275), .Q(n282) );
  AOI221 U302 ( .A(N221), .B(n499), .C(half_sub[13]), .D(n486), .Q(n280) );
  NOR20 U303 ( .A(n70), .B(i_data_A[31]), .Q(n539) );
  NAND22 U304 ( .A(N242), .B(n538), .Q(n133) );
  NAND22 U305 ( .A(N252), .B(n538), .Q(n258) );
  NAND22 U306 ( .A(N251), .B(n538), .Q(n244) );
  NAND20 U307 ( .A(i_data_A[31]), .B(n70), .Q(n536) );
  NAND21 U308 ( .A(half_sub[3]), .B(n486), .Q(n155) );
  INV3 U309 ( .A(N233), .Q(n452) );
  IMUX21 U310 ( .A(n46), .B(n535), .S(n68), .Q(n525) );
  AOI211 U311 ( .A(n3), .B(n284), .C(n283), .Q(n285) );
  CLKBU15 U312 ( .A(i_data_B[24]), .Q(n81) );
  INV15 U313 ( .A(n548), .Q(n499) );
  NAND41 U314 ( .A(n380), .B(n379), .C(n378), .D(n377), .Q(o_data_AluRes[20])
         );
  AOI220 U315 ( .A(N260), .B(n538), .C(pre_sum_3a[4]), .D(n426), .Q(n378) );
  IMUX20 U316 ( .A(n205), .B(n204), .S(n74), .Q(n214) );
  IMUX20 U317 ( .A(n72), .B(n489), .S(n57), .Q(n284) );
  NOR20 U318 ( .A(n49), .B(i_data_A[8]), .Q(n205) );
  NOR20 U319 ( .A(n49), .B(i_data_A[10]), .Q(n235) );
  NOR20 U320 ( .A(n541), .B(n369), .Q(n372) );
  INV0 U321 ( .A(n66), .Q(n490) );
  AOI220 U322 ( .A(n553), .B(pre_sum_4b[2]), .C(pre_sum_4a[2]), .D(n552), .Q(
        n470) );
  INV2 U323 ( .A(pre_subb[4]), .Q(n370) );
  AOI220 U324 ( .A(n53), .B(n524), .C(N265), .D(n538), .Q(n451) );
  AOI220 U325 ( .A(N257), .B(n538), .C(pre_sum_3a[1]), .D(n426), .Q(n338) );
  NAND20 U326 ( .A(n405), .B(n520), .Q(n407) );
  NAND20 U327 ( .A(half_sub[2]), .B(n486), .Q(n145) );
  NAND20 U328 ( .A(n521), .B(n520), .Q(n523) );
  AOI210 U329 ( .A(n52), .B(n162), .C(n161), .Q(n163) );
  AOI220 U330 ( .A(n57), .B(n524), .C(N270), .D(n538), .Q(n527) );
  IMUX20 U331 ( .A(n279), .B(n278), .S(n56), .Q(n281) );
  AOI220 U332 ( .A(sum_1[4]), .B(n437), .C(half_sub[4]), .D(n486), .Q(n168) );
  NAND41 U333 ( .A(n170), .B(n169), .C(n168), .D(n167), .Q(o_data_AluRes[4])
         );
  AOI220 U334 ( .A(sum_1[5]), .B(n437), .C(half_sub[5]), .D(n486), .Q(n182) );
  IMUX20 U335 ( .A(n257), .B(n256), .S(n76), .Q(n266) );
  IMUX20 U336 ( .A(n73), .B(n489), .S(n63), .Q(n400) );
  AOI210 U337 ( .A(N271), .B(n538), .C(n537), .Q(n546) );
  NOR20 U338 ( .A(n536), .B(n535), .Q(n537) );
  IMUX20 U339 ( .A(n72), .B(n489), .S(n81), .Q(n430) );
  NAND20 U340 ( .A(n86), .B(n520), .Q(n354) );
  AOI210 U341 ( .A(n86), .B(n72), .C(n71), .Q(n353) );
  INV2 U342 ( .A(pre_sum_2a[5]), .Q(n270) );
  NOR20 U343 ( .A(n541), .B(n399), .Q(n402) );
  NOR20 U344 ( .A(n541), .B(n382), .Q(n385) );
  NAND20 U345 ( .A(n390), .B(n520), .Q(n392) );
  NAND20 U346 ( .A(n122), .B(n520), .Q(n124) );
  AOI220 U347 ( .A(n74), .B(n524), .C(N264), .D(n538), .Q(n435) );
  NAND20 U348 ( .A(n446), .B(n520), .Q(n448) );
  INV2 U349 ( .A(pre_subb[3]), .Q(n359) );
  NOR20 U350 ( .A(n50), .B(i_data_A[12]), .Q(n257) );
  IMUX20 U351 ( .A(n73), .B(n489), .S(i_data_A[2]), .Q(n141) );
  OAI210 U352 ( .A(n121), .B(n71), .C(i_data_A[1]), .Q(n132) );
  NOR20 U353 ( .A(n49), .B(i_data_A[9]), .Q(n224) );
  IMUX20 U354 ( .A(n72), .B(n489), .S(n80), .Q(n415) );
  IMUX20 U355 ( .A(n46), .B(n535), .S(n76), .Q(n260) );
  NOR20 U356 ( .A(n50), .B(i_data_A[11]), .Q(n242) );
  NOR20 U357 ( .A(n50), .B(i_data_A[13]), .Q(n279) );
  NOR20 U358 ( .A(n50), .B(i_data_A[14]), .Q(n289) );
  NOR20 U359 ( .A(n49), .B(i_data_A[5]), .Q(n172) );
  AOI210 U360 ( .A(n325), .B(n73), .C(n71), .Q(n326) );
  NAND20 U361 ( .A(n325), .B(n520), .Q(n327) );
  NOR20 U362 ( .A(n49), .B(i_data_A[4]), .Q(n166) );
  NOR20 U363 ( .A(n49), .B(i_data_A[6]), .Q(n184) );
  NOR20 U364 ( .A(n49), .B(i_data_A[7]), .Q(n195) );
  BUF15 U365 ( .A(i_data_B[19]), .Q(n78) );
  NOR20 U366 ( .A(n541), .B(n340), .Q(n343) );
  NAND20 U367 ( .A(sum_1[0]), .B(n437), .Q(n101) );
  OAI210 U368 ( .A(n186), .B(n71), .C(i_data_A[6]), .Q(n188) );
  INV3 U369 ( .A(n35), .Q(n36) );
  NAND20 U370 ( .A(pre_sum_4b[4]), .B(n553), .Q(n504) );
  NAND22 U371 ( .A(n439), .B(n437), .Q(n389) );
  INV3 U372 ( .A(N248), .Q(n206) );
  INV3 U373 ( .A(pre_sum_2b[1]), .Q(n217) );
  INV3 U374 ( .A(N249), .Q(n216) );
  NAND22 U375 ( .A(pre_suba[8]), .B(n551), .Q(n444) );
  AOI211 U376 ( .A(N232), .B(n499), .C(n431), .Q(n445) );
  NAND41 U377 ( .A(n458), .B(n457), .C(n456), .D(n455), .Q(o_data_AluRes[25])
         );
  INV3 U378 ( .A(pre_sum_2b[2]), .Q(n229) );
  INV3 U379 ( .A(N250), .Q(n228) );
  NAND41 U380 ( .A(n557), .B(n556), .C(n555), .D(n554), .Q(o_data_AluRes[31])
         );
  NAND22 U381 ( .A(pre_suba[5]), .B(n551), .Q(n398) );
  AOI211 U382 ( .A(N227), .B(n499), .C(n355), .Q(n365) );
  NOR21 U383 ( .A(n544), .B(n543), .Q(n545) );
  IMUX21 U384 ( .A(n51), .B(n50), .S(n539), .Q(n544) );
  INV3 U385 ( .A(n59), .Q(n540) );
  AOI2111 U386 ( .A(i_data_A[20]), .B(n373), .C(n372), .D(n371), .Q(n379) );
  NAND22 U387 ( .A(n52), .B(n368), .Q(n373) );
  NOR21 U388 ( .A(n34), .B(n360), .Q(n362) );
  OAI2111 U389 ( .A(n381), .B(n359), .C(n358), .D(n357), .Q(n363) );
  NAND31 U390 ( .A(n215), .B(n214), .C(n213), .Q(o_data_AluRes[8]) );
  NOR21 U391 ( .A(n212), .B(n211), .Q(n213) );
  NAND22 U392 ( .A(n159), .B(n158), .Q(o_data_AluRes[3]) );
  NAND22 U393 ( .A(n269), .B(n268), .Q(n277) );
  NAND22 U394 ( .A(n404), .B(n403), .Q(n409) );
  NAND22 U395 ( .A(pre_sum_3a[6]), .B(n426), .Q(n404) );
  NAND22 U396 ( .A(n470), .B(n45), .Q(o_data_AluRes[26]) );
  BUF2 U397 ( .A(i_data_B[31]), .Q(n70) );
  IMUX21 U398 ( .A(n301), .B(n300), .S(n59), .Q(n302) );
  AOI2111 U399 ( .A(N247), .B(n538), .C(n200), .D(n199), .Q(n201) );
  AOI211 U400 ( .A(N225), .B(n499), .C(n328), .Q(n337) );
  NAND41 U401 ( .A(n146), .B(n145), .C(n144), .D(n143), .Q(o_data_AluRes[2])
         );
  NOR21 U402 ( .A(n139), .B(n138), .Q(n144) );
  NAND42 U403 ( .A(n293), .B(n292), .C(n291), .D(n290), .Q(o_data_AluRes[14])
         );
  IMUX21 U404 ( .A(n289), .B(n288), .S(n57), .Q(n290) );
  AOI211 U405 ( .A(N210), .B(n499), .C(n134), .Q(n146) );
  XNR21 U406 ( .A(i_data_A[31]), .B(n70), .Q(n542) );
  AOI211 U407 ( .A(n3), .B(n230), .C(n84), .Q(n231) );
  AOI2111 U408 ( .A(pre_sum_2a[2]), .B(n233), .C(n232), .D(n231), .Q(n238) );
  NAND31 U409 ( .A(n227), .B(n226), .C(n225), .Q(o_data_AluRes[9]) );
  AOI2111 U410 ( .A(pre_sum_2a[1]), .B(n233), .C(n222), .D(n221), .Q(n227) );
  NAND31 U411 ( .A(n282), .B(n281), .C(n280), .Q(o_data_AluRes[13]) );
  NAND31 U412 ( .A(n182), .B(n181), .C(n180), .Q(o_data_AluRes[5]) );
  NOR21 U413 ( .A(n179), .B(n178), .Q(n180) );
  NAND31 U414 ( .A(n193), .B(n192), .C(n191), .Q(o_data_AluRes[6]) );
  NOR21 U415 ( .A(n190), .B(n189), .Q(n191) );
  IMUX21 U416 ( .A(n468), .B(n467), .S(n30), .Q(n469) );
  AOI211 U417 ( .A(n3), .B(n430), .C(n88), .Q(n431) );
  AOI211 U418 ( .A(n3), .B(n400), .C(n405), .Q(n401) );
  IMUX21 U419 ( .A(n523), .B(n522), .S(n68), .Q(n530) );
  NAND22 U420 ( .A(n259), .B(n258), .Q(n264) );
  NAND22 U421 ( .A(pre_sum_2b[4]), .B(n297), .Q(n259) );
  NAND22 U422 ( .A(n245), .B(n244), .Q(n250) );
  NAND22 U423 ( .A(pre_sum_2b[3]), .B(n297), .Q(n245) );
  NAND22 U424 ( .A(n155), .B(n154), .Q(n156) );
  NAND22 U425 ( .A(n435), .B(n434), .Q(n436) );
  NAND22 U426 ( .A(N236), .B(n499), .Q(n500) );
  BUF2 U427 ( .A(i_data_B[31]), .Q(n69) );
  INV3 U428 ( .A(N235), .Q(n479) );
  INV3 U429 ( .A(N239), .Q(n547) );
  AOI211 U430 ( .A(n52), .B(n198), .C(n197), .Q(n199) );
  INV3 U431 ( .A(i_data_A[7]), .Q(n197) );
  INV3 U432 ( .A(i_data_A[2]), .Q(n137) );
  NAND31 U433 ( .A(i_data_A[28]), .B(n73), .C(n490), .Q(n494) );
  NAND22 U434 ( .A(N268), .B(n538), .Q(n496) );
  INV3 U435 ( .A(i_data_A[5]), .Q(n176) );
  NAND31 U436 ( .A(i_data_A[26]), .B(n72), .C(n459), .Q(n462) );
  NAND22 U437 ( .A(N266), .B(n538), .Q(n464) );
  NAND42 U438 ( .A(n132), .B(n131), .C(n130), .D(n129), .Q(o_data_AluRes[1])
         );
  INV3 U439 ( .A(i_data_A[14]), .Q(n283) );
  IMUX21 U440 ( .A(n509), .B(n508), .S(n67), .Q(n515) );
  INV3 U441 ( .A(i_data_A[29]), .Q(n507) );
  AOI211 U442 ( .A(n274), .B(n3), .C(n273), .Q(n275) );
  INV3 U443 ( .A(i_data_A[13]), .Q(n273) );
  INV3 U444 ( .A(i_data_A[9]), .Q(n218) );
  AOI211 U445 ( .A(N240), .B(n538), .C(n99), .Q(n102) );
  NAND22 U446 ( .A(pre_sum_2a[3]), .B(n233), .Q(n247) );
  AOI211 U447 ( .A(n52), .B(n295), .C(n294), .Q(n296) );
  INV3 U448 ( .A(i_data_A[15]), .Q(n294) );
  AOI211 U449 ( .A(n3), .B(n415), .C(n414), .Q(n416) );
  INV3 U450 ( .A(i_data_A[23]), .Q(n414) );
  IMUX21 U451 ( .A(n327), .B(n326), .S(n60), .Q(n328) );
  INV3 U452 ( .A(i_data_A[17]), .Q(n325) );
  AOI211 U453 ( .A(n345), .B(n72), .C(n71), .Q(n346) );
  INV3 U454 ( .A(i_data_A[18]), .Q(n345) );
  NAND22 U455 ( .A(n262), .B(n261), .Q(n263) );
  NAND22 U456 ( .A(pre_sum_2a[4]), .B(n233), .Q(n261) );
  NAND22 U457 ( .A(n422), .B(n421), .Q(n425) );
  IMUX21 U458 ( .A(n420), .B(n419), .S(n80), .Q(n421) );
  NAND22 U459 ( .A(N231), .B(n499), .Q(n422) );
  NAND22 U460 ( .A(n52), .B(n141), .Q(n142) );
  INV3 U461 ( .A(i_data_A[28]), .Q(n491) );
  INV3 U462 ( .A(i_data_A[25]), .Q(n446) );
  INV3 U463 ( .A(i_data_A[26]), .Q(n466) );
  INV3 U464 ( .A(i_data_A[30]), .Q(n521) );
  INV3 U465 ( .A(i_data_A[21]), .Q(n390) );
  INV3 U466 ( .A(i_data_A[22]), .Q(n405) );
  INV3 U467 ( .A(i_data_A[0]), .Q(n107) );
  INV3 U468 ( .A(i_data_A[3]), .Q(n151) );
  INV3 U469 ( .A(i_data_A[4]), .Q(n161) );
  INV3 U470 ( .A(i_data_A[1]), .Q(n122) );
  INV3 U471 ( .A(i_data_A[16]), .Q(n85) );
  INV3 U472 ( .A(i_data_A[19]), .Q(n86) );
  INV3 U473 ( .A(i_data_A[27]), .Q(n89) );
  INV3 U474 ( .A(i_data_A[20]), .Q(n87) );
  INV3 U475 ( .A(i_data_A[10]), .Q(n84) );
  INV3 U476 ( .A(i_data_A[24]), .Q(n88) );
  INV3 U477 ( .A(i_data_A[8]), .Q(n83) );
  LOGIC0 U478 ( .Q(n43) );
  LOGIC1 U479 ( .Q(n42) );
  IMUX20 U480 ( .A(n73), .B(n272), .S(n56), .Q(n274) );
  NOR21 U481 ( .A(n271), .B(n270), .Q(n276) );
  IMUX20 U482 ( .A(n73), .B(n272), .S(n53), .Q(n219) );
  AOI211 U483 ( .A(n89), .B(n73), .C(n71), .Q(n474) );
  NAND31 U484 ( .A(n338), .B(n337), .C(n336), .Q(o_data_AluRes[17]) );
  NAND30 U485 ( .A(n39), .B(n311), .C(n310), .Q(n119) );
  OAI221 U486 ( .A(n389), .B(n388), .C(n387), .D(n386), .Q(n394) );
  IMUX20 U487 ( .A(n235), .B(n234), .S(n75), .Q(n237) );
  OAI212 U488 ( .A(n449), .B(n71), .C(i_data_A[25]), .Q(n450) );
  NOR20 U489 ( .A(n440), .B(n136), .Q(n139) );
  OAI220 U490 ( .A(n135), .B(n126), .C(n440), .D(n125), .Q(n127) );
  IMUX21 U491 ( .A(n375), .B(n374), .S(n79), .Q(n376) );
  NOR20 U492 ( .A(n97), .B(n1), .Q(n94) );
  IMUX21 U493 ( .A(n392), .B(n391), .S(n62), .Q(n393) );
  IMUX21 U494 ( .A(n72), .B(n489), .S(n77), .Q(n309) );
  IMUX20 U495 ( .A(n46), .B(n535), .S(i_data_B[6]), .Q(n186) );
  IMUX20 U496 ( .A(n46), .B(n535), .S(n55), .Q(n246) );
  OAI210 U497 ( .A(n246), .B(n71), .C(i_data_A[11]), .Q(n248) );
  CLKIN0 U498 ( .A(n37), .Q(n369) );
  CLKIN0 U499 ( .A(n38), .Q(n413) );
  IMUX20 U500 ( .A(n195), .B(n194), .S(n38), .Q(n202) );
  IMUX20 U501 ( .A(n124), .B(n123), .S(i_data_B[1]), .Q(n128) );
  NOR21 U502 ( .A(n128), .B(n127), .Q(n129) );
  NAND21 U503 ( .A(n151), .B(n520), .Q(n153) );
  AOI211 U504 ( .A(n491), .B(n73), .C(n71), .Q(n487) );
  IMUX20 U505 ( .A(n73), .B(n489), .S(n38), .Q(n198) );
  NOR20 U506 ( .A(n541), .B(n4), .Q(n315) );
  NOR20 U507 ( .A(n541), .B(n413), .Q(n417) );
  NAND31 U508 ( .A(n203), .B(n202), .C(n201), .Q(o_data_AluRes[7]) );
  IMUX20 U509 ( .A(n46), .B(n535), .S(i_data_B[1]), .Q(n121) );
  IMUX20 U510 ( .A(n242), .B(n241), .S(n54), .Q(n252) );
  IMUX20 U511 ( .A(n73), .B(n489), .S(n75), .Q(n230) );
  CLKBU15 U512 ( .A(i_data_B[10]), .Q(n75) );
  IMUX21 U513 ( .A(n153), .B(n152), .S(i_data_B[3]), .Q(n157) );
  NAND20 U514 ( .A(i_data_B[3]), .B(n524), .Q(n357) );
  IMUX20 U515 ( .A(n73), .B(n489), .S(i_data_B[3]), .Q(n148) );
  IMUX20 U516 ( .A(n166), .B(n165), .S(n37), .Q(n167) );
  IMUX20 U517 ( .A(n73), .B(n489), .S(n37), .Q(n162) );
  NOR21 U518 ( .A(n52), .B(n137), .Q(n138) );
  NOR21 U519 ( .A(n51), .B(n491), .Q(n492) );
  NOR21 U520 ( .A(n51), .B(n466), .Q(n460) );
  NOR20 U521 ( .A(n312), .B(n310), .Q(n95) );
  AOI211 U522 ( .A(n466), .B(n72), .C(n71), .Q(n467) );
  IMUX21 U523 ( .A(n354), .B(n353), .S(n78), .Q(n355) );
  IMUX21 U524 ( .A(n46), .B(n535), .S(n78), .Q(n356) );
  CLKIN0 U525 ( .A(i_data_B[6]), .Q(n399) );
  IMUX21 U526 ( .A(n184), .B(n183), .S(i_data_B[6]), .Q(n192) );
  NAND22 U527 ( .A(i_con_AluCtrl[2]), .B(n97), .Q(n90) );
  AOI221 U528 ( .A(pre_sum_3b[6]), .B(n418), .C(pre_suba[6]), .D(n551), .Q(
        n411) );
  AOI221 U529 ( .A(pre_suba[9]), .B(n551), .C(pre_subb[9]), .D(n550), .Q(n457)
         );
  IMUX21 U530 ( .A(n220), .B(n142), .S(n41), .Q(n143) );
  NOR32 U531 ( .A(n39), .B(n97), .C(i_con_AluCtrl[3]), .Q(n100) );
  NAND33 U532 ( .A(n471), .B(n473), .C(n472), .Q(n44) );
  NAND22 U533 ( .A(pre_suba[10]), .B(n551), .Q(n472) );
  IMUX21 U534 ( .A(n407), .B(n406), .S(n63), .Q(n408) );
  NAND42 U535 ( .A(n445), .B(n444), .C(n443), .D(n442), .Q(o_data_AluRes[24])
         );
  AOI210 U536 ( .A(n390), .B(n72), .C(n71), .Q(n391) );
  AOI210 U537 ( .A(n405), .B(n72), .C(n71), .Q(n406) );
  NOR24 U538 ( .A(n103), .B(n312), .Q(n91) );
  CLKIN3 U539 ( .A(n542), .Q(n93) );
  CLKIN3 U540 ( .A(half_sub[0]), .Q(n98) );
  NAND22 U541 ( .A(n102), .B(n101), .Q(n116) );
  NAND22 U542 ( .A(N208), .B(n499), .Q(n113) );
  NAND22 U543 ( .A(N241), .B(n538), .Q(n131) );
  NAND22 U544 ( .A(N209), .B(n499), .Q(n130) );
  CLKIN3 U545 ( .A(half_sub[1]), .Q(n126) );
  CLKIN3 U546 ( .A(sum_1[1]), .Q(n125) );
  CLKIN3 U547 ( .A(n133), .Q(n134) );
  CLKIN3 U548 ( .A(sum_1[2]), .Q(n136) );
  NAND22 U549 ( .A(N243), .B(n538), .Q(n147) );
  NAND22 U550 ( .A(N244), .B(n538), .Q(n160) );
  CLKIN3 U551 ( .A(n160), .Q(n164) );
  NAND22 U552 ( .A(N212), .B(n499), .Q(n169) );
  OAI212 U553 ( .A(n47), .B(i_data_A[4]), .C(n52), .Q(n165) );
  NAND22 U554 ( .A(N213), .B(n499), .Q(n173) );
  CLKIN3 U555 ( .A(n173), .Q(n179) );
  CLKIN3 U556 ( .A(N245), .Q(n175) );
  NAND22 U557 ( .A(N214), .B(n499), .Q(n185) );
  CLKIN3 U558 ( .A(n185), .Q(n190) );
  NAND22 U559 ( .A(N246), .B(n538), .Q(n187) );
  NAND22 U560 ( .A(n188), .B(n187), .Q(n189) );
  OAI212 U561 ( .A(n47), .B(i_data_A[7]), .C(n52), .Q(n194) );
  NAND22 U562 ( .A(N215), .B(n499), .Q(n196) );
  CLKIN3 U563 ( .A(n196), .Q(n200) );
  OAI212 U564 ( .A(n47), .B(i_data_A[8]), .C(n52), .Q(n204) );
  CLKIN3 U565 ( .A(pre_sum_2b[0]), .Q(n207) );
  OAI222 U566 ( .A(n243), .B(n207), .C(n387), .D(n206), .Q(n212) );
  CLKIN3 U567 ( .A(pre_sum_2a[0]), .Q(n209) );
  OAI222 U568 ( .A(n243), .B(n229), .C(n387), .D(n228), .Q(n232) );
  NAND22 U569 ( .A(N219), .B(n499), .Q(n239) );
  OAI212 U570 ( .A(n47), .B(i_data_A[11]), .C(n3), .Q(n241) );
  NAND22 U571 ( .A(n248), .B(n247), .Q(n249) );
  NAND22 U572 ( .A(N220), .B(n499), .Q(n254) );
  CLKIN3 U573 ( .A(n254), .Q(n255) );
  NAND22 U574 ( .A(N222), .B(n499), .Q(n286) );
  CLKIN3 U575 ( .A(n286), .Q(n287) );
  NAND22 U576 ( .A(N223), .B(n499), .Q(n298) );
  CLKIN3 U577 ( .A(n298), .Q(n299) );
  OAI212 U578 ( .A(n47), .B(i_data_A[15]), .C(n52), .Q(n300) );
  CLKIN3 U579 ( .A(pre_subb[0]), .Q(n313) );
  CLKIN3 U580 ( .A(pre_subb[1]), .Q(n332) );
  CLKIN3 U581 ( .A(pre_sum_3b[1]), .Q(n333) );
  CLKIN3 U582 ( .A(pre_subb[2]), .Q(n341) );
  NAND22 U583 ( .A(N259), .B(n538), .Q(n366) );
  CLKIN3 U584 ( .A(pre_sum_3b[3]), .Q(n360) );
  CLKIN3 U585 ( .A(pre_sum_3a[5]), .Q(n388) );
  CLKIN3 U586 ( .A(N261), .Q(n386) );
  NAND22 U587 ( .A(N262), .B(n538), .Q(n403) );
  NAND22 U588 ( .A(N263), .B(n538), .Q(n423) );
  CLKIN3 U589 ( .A(n423), .Q(n424) );
  OAI212 U590 ( .A(n46), .B(i_data_A[24]), .C(n3), .Q(n432) );
  AOI212 U591 ( .A(pre_subb[10]), .B(n550), .C(n469), .Q(n471) );
  OAI2112 U592 ( .A(n548), .B(n547), .C(n546), .D(n545), .Q(n549) );
endmodule


module E_alu_control ( o_con_AluCtrl, i_con_AluOp, i_con_FuncCode );
  output [3:0] o_con_AluCtrl;
  input [5:0] i_con_AluOp;
  input [5:0] i_con_FuncCode;
  wire   n20, n37, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68;

  NAND24 U3 ( .A(n56), .B(n45), .Q(n47) );
  OAI2112 U4 ( .A(n11), .B(n55), .C(n10), .D(n41), .Q(n18) );
  CLKIN8 U5 ( .A(i_con_FuncCode[2]), .Q(n25) );
  NAND28 U6 ( .A(n49), .B(n48), .Q(o_con_AluCtrl[1]) );
  IMUX24 U7 ( .A(n47), .B(n46), .S(i_con_AluOp[0]), .Q(n48) );
  CLKIN6 U8 ( .A(n55), .Q(n22) );
  NAND26 U9 ( .A(n29), .B(n28), .Q(n56) );
  NAND22 U10 ( .A(n54), .B(n24), .Q(n41) );
  CLKIN6 U11 ( .A(n19), .Q(n63) );
  CLKIN6 U12 ( .A(n14), .Q(n15) );
  INV3 U13 ( .A(i_con_AluOp[2]), .Q(n68) );
  NOR23 U14 ( .A(i_con_AluOp[3]), .B(n7), .Q(n8) );
  INV3 U15 ( .A(i_con_AluOp[0]), .Q(n30) );
  NAND24 U16 ( .A(i_con_FuncCode[1]), .B(n25), .Q(n14) );
  NAND31 U17 ( .A(n19), .B(n37), .C(n53), .Q(n17) );
  NAND23 U18 ( .A(n50), .B(n42), .Q(n27) );
  CLKIN3 U19 ( .A(i_con_FuncCode[3]), .Q(n13) );
  NOR22 U20 ( .A(n4), .B(n62), .Q(n65) );
  INV3 U21 ( .A(n31), .Q(n64) );
  INV2 U22 ( .A(n60), .Q(n1) );
  CLKIN12 U23 ( .A(n56), .Q(n60) );
  NOR32 U24 ( .A(n44), .B(n43), .C(n51), .Q(n45) );
  AOI312 U25 ( .A(n67), .B(n35), .C(n1), .D(n34), .Q(o_con_AluCtrl[0]) );
  OAI210 U26 ( .A(n52), .B(n51), .C(n64), .Q(n58) );
  CLKIN2 U27 ( .A(i_con_FuncCode[0]), .Q(n16) );
  NAND22 U28 ( .A(n53), .B(n42), .Q(n43) );
  CLKIN6 U29 ( .A(i_con_FuncCode[5]), .Q(n24) );
  NAND22 U30 ( .A(i_con_FuncCode[1]), .B(n25), .Q(n2) );
  NAND34 U31 ( .A(n67), .B(n66), .C(n65), .Q(o_con_AluCtrl[3]) );
  NAND24 U32 ( .A(i_con_FuncCode[5]), .B(i_con_FuncCode[0]), .Q(n12) );
  NOR22 U33 ( .A(n31), .B(n3), .Q(n4) );
  INV1 U34 ( .A(n63), .Q(n3) );
  NOR31 U35 ( .A(n17), .B(n51), .C(n18), .Q(n35) );
  INV2 U36 ( .A(n37), .Q(n32) );
  NAND22 U37 ( .A(i_con_AluOp[1]), .B(n30), .Q(n31) );
  OAI311 U38 ( .A(i_con_AluOp[5]), .B(n8), .C(n38), .D(i_con_AluOp[0]), .Q(n36) );
  NAND30 U39 ( .A(i_con_AluOp[0]), .B(i_con_AluOp[3]), .C(i_con_AluOp[2]), .Q(
        n20) );
  CLKIN3 U40 ( .A(i_con_FuncCode[4]), .Q(n53) );
  NOR24 U41 ( .A(n27), .B(n51), .Q(n28) );
  NOR24 U42 ( .A(n6), .B(n2), .Q(n51) );
  NOR20 U43 ( .A(i_con_AluOp[2]), .B(i_con_AluOp[3]), .Q(n46) );
  NAND40 U44 ( .A(i_con_AluOp[3]), .B(i_con_AluOp[2]), .C(i_con_AluOp[0]), .D(
        n7), .Q(n9) );
  CLKIN3 U45 ( .A(i_con_AluOp[1]), .Q(n38) );
  CLKIN3 U46 ( .A(i_con_AluOp[4]), .Q(n7) );
  NOR23 U47 ( .A(n12), .B(n13), .Q(n5) );
  CLKIN6 U48 ( .A(n5), .Q(n6) );
  INV3 U49 ( .A(n20), .Q(n62) );
  NOR31 U50 ( .A(n64), .B(n33), .C(n32), .Q(n34) );
  NAND31 U51 ( .A(i_con_AluOp[0]), .B(i_con_AluOp[4]), .C(n68), .Q(n59) );
  NOR31 U52 ( .A(n40), .B(n39), .C(n38), .Q(n49) );
  NAND22 U53 ( .A(n9), .B(n36), .Q(n33) );
  NAND31 U54 ( .A(i_con_AluOp[3]), .B(n68), .C(i_con_AluOp[0]), .Q(n37) );
  OAI211 U55 ( .A(n55), .B(n54), .C(n53), .Q(n61) );
  NAND20 U56 ( .A(n24), .B(i_con_FuncCode[0]), .Q(n10) );
  NAND22 U57 ( .A(n23), .B(i_con_FuncCode[1]), .Q(n50) );
  CLKIN2 U58 ( .A(i_con_FuncCode[1]), .Q(n54) );
  NAND23 U59 ( .A(n26), .B(n25), .Q(n42) );
  INV2 U60 ( .A(n50), .Q(n52) );
  NOR22 U61 ( .A(i_con_FuncCode[3]), .B(n24), .Q(n26) );
  NOR33 U62 ( .A(n63), .B(n22), .C(n21), .Q(n29) );
  NOR31 U63 ( .A(i_con_FuncCode[0]), .B(i_con_FuncCode[3]), .C(
        i_con_FuncCode[2]), .Q(n21) );
  XNR21 U64 ( .A(i_con_FuncCode[1]), .B(i_con_FuncCode[0]), .Q(n11) );
  NOR21 U65 ( .A(i_con_FuncCode[2]), .B(i_con_FuncCode[3]), .Q(n23) );
  NAND32 U66 ( .A(i_con_FuncCode[5]), .B(n13), .C(i_con_FuncCode[2]), .Q(n55)
         );
  CLKIN3 U67 ( .A(n33), .Q(n67) );
  NAND43 U68 ( .A(i_con_FuncCode[5]), .B(n16), .C(i_con_FuncCode[3]), .D(n15), 
        .Q(n19) );
  CLKIN3 U69 ( .A(n59), .Q(n40) );
  CLKIN3 U70 ( .A(n36), .Q(n39) );
  CLKIN3 U71 ( .A(n41), .Q(n44) );
  OAI212 U72 ( .A(n61), .B(n60), .C(n64), .Q(n57) );
  NAND43 U73 ( .A(n67), .B(n59), .C(n58), .D(n57), .Q(o_con_AluCtrl[2]) );
  AOI222 U74 ( .A(n64), .B(n61), .C(n64), .D(n60), .Q(n66) );
endmodule


module E_famux5 ( i_data_rs, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fa, o_data_alusra );
  input [31:0] i_data_rs;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fa;
  output [31:0] o_data_alusra;
  wire   N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N54, n2, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13;

  DLPQ3 o_data_alusra_reg_31_ ( .SN(n2), .D(N54), .GN(n46), .Q(
        o_data_alusra[31]) );
  DLPQ3 o_data_alusra_reg_30_ ( .SN(n2), .D(N52), .GN(n46), .Q(
        o_data_alusra[30]) );
  DLPQ3 o_data_alusra_reg_29_ ( .SN(n2), .D(N51), .GN(n46), .Q(
        o_data_alusra[29]) );
  DLPQ3 o_data_alusra_reg_28_ ( .SN(n2), .D(N50), .GN(n46), .Q(
        o_data_alusra[28]) );
  DLPQ3 o_data_alusra_reg_27_ ( .SN(n2), .D(N49), .GN(n46), .Q(
        o_data_alusra[27]) );
  DLPQ3 o_data_alusra_reg_26_ ( .SN(n2), .D(N48), .GN(n46), .Q(
        o_data_alusra[26]) );
  DLPQ3 o_data_alusra_reg_25_ ( .SN(n2), .D(N47), .GN(n8), .Q(
        o_data_alusra[25]) );
  DLPQ3 o_data_alusra_reg_24_ ( .SN(n2), .D(N46), .GN(n8), .Q(
        o_data_alusra[24]) );
  DLPQ3 o_data_alusra_reg_23_ ( .SN(n2), .D(N45), .GN(n8), .Q(
        o_data_alusra[23]) );
  DLPQ3 o_data_alusra_reg_22_ ( .SN(n2), .D(N44), .GN(n8), .Q(
        o_data_alusra[22]) );
  DLPQ3 o_data_alusra_reg_21_ ( .SN(n2), .D(N43), .GN(n8), .Q(
        o_data_alusra[21]) );
  DLPQ3 o_data_alusra_reg_20_ ( .SN(n2), .D(N42), .GN(n8), .Q(
        o_data_alusra[20]) );
  DLPQ3 o_data_alusra_reg_19_ ( .SN(n2), .D(N41), .GN(n8), .Q(
        o_data_alusra[19]) );
  DLPQ3 o_data_alusra_reg_18_ ( .SN(n2), .D(N40), .GN(n8), .Q(
        o_data_alusra[18]) );
  DLPQ3 o_data_alusra_reg_17_ ( .SN(n2), .D(N39), .GN(n8), .Q(
        o_data_alusra[17]) );
  DLPQ3 o_data_alusra_reg_16_ ( .SN(n2), .D(N38), .GN(n46), .Q(
        o_data_alusra[16]) );
  DLPQ3 o_data_alusra_reg_15_ ( .SN(n2), .D(N37), .GN(n8), .Q(
        o_data_alusra[15]) );
  DLPQ3 o_data_alusra_reg_14_ ( .SN(n2), .D(N36), .GN(n8), .Q(
        o_data_alusra[14]) );
  DLPQ3 o_data_alusra_reg_13_ ( .SN(n2), .D(N35), .GN(n46), .Q(
        o_data_alusra[13]) );
  DLPQ3 o_data_alusra_reg_12_ ( .SN(n2), .D(N34), .GN(n8), .Q(
        o_data_alusra[12]) );
  DLPQ3 o_data_alusra_reg_11_ ( .SN(n2), .D(N33), .GN(n8), .Q(
        o_data_alusra[11]) );
  DLPQ3 o_data_alusra_reg_10_ ( .SN(n2), .D(N32), .GN(n8), .Q(
        o_data_alusra[10]) );
  DLPQ3 o_data_alusra_reg_9_ ( .SN(n2), .D(N31), .GN(n8), .Q(o_data_alusra[9])
         );
  DLPQ3 o_data_alusra_reg_8_ ( .SN(n2), .D(N30), .GN(n8), .Q(o_data_alusra[8])
         );
  DLPQ3 o_data_alusra_reg_7_ ( .SN(n2), .D(N29), .GN(n8), .Q(o_data_alusra[7])
         );
  DLPQ3 o_data_alusra_reg_6_ ( .SN(n2), .D(N28), .GN(n8), .Q(o_data_alusra[6])
         );
  DLPQ3 o_data_alusra_reg_5_ ( .SN(n2), .D(N27), .GN(n8), .Q(o_data_alusra[5])
         );
  DLPQ3 o_data_alusra_reg_4_ ( .SN(n2), .D(N26), .GN(n8), .Q(o_data_alusra[4])
         );
  DLPQ3 o_data_alusra_reg_3_ ( .SN(n2), .D(N25), .GN(n8), .Q(o_data_alusra[3])
         );
  DLPQ3 o_data_alusra_reg_2_ ( .SN(n2), .D(N24), .GN(n8), .Q(o_data_alusra[2])
         );
  DLPQ3 o_data_alusra_reg_1_ ( .SN(n2), .D(N23), .GN(n8), .Q(o_data_alusra[1])
         );
  DLPQ3 o_data_alusra_reg_0_ ( .SN(n2), .D(N22), .GN(n8), .Q(o_data_alusra[0])
         );
  AOI220 U2 ( .A(i_data_writeres[0]), .B(n41), .C(i_data_rs[0]), .D(n42), .Q(
        n140) );
  AOI220 U3 ( .A(i_data_writeres[1]), .B(n41), .C(i_data_rs[1]), .D(n7), .Q(
        n137) );
  AOI220 U4 ( .A(i_data_writeres[3]), .B(n5), .C(i_data_rs[3]), .D(n42), .Q(
        n131) );
  AOI220 U5 ( .A(i_data_writeres[4]), .B(n41), .C(i_data_rs[4]), .D(n7), .Q(
        n128) );
  AOI220 U6 ( .A(i_data_writeres[6]), .B(n41), .C(i_data_rs[6]), .D(n42), .Q(
        n122) );
  AOI220 U7 ( .A(i_data_lwW[7]), .B(n44), .C(i_data_lwM[7]), .D(n3), .Q(n117)
         );
  AOI220 U8 ( .A(i_data_writeres[7]), .B(n41), .C(i_data_rs[7]), .D(n7), .Q(
        n119) );
  AOI220 U9 ( .A(i_data_writeres[9]), .B(n5), .C(i_data_rs[9]), .D(n42), .Q(
        n113) );
  AOI220 U10 ( .A(i_data_writeres[10]), .B(n41), .C(i_data_rs[10]), .D(n7), 
        .Q(n110) );
  AOI220 U11 ( .A(i_data_writeres[12]), .B(n41), .C(i_data_rs[12]), .D(n42), 
        .Q(n104) );
  AOI220 U12 ( .A(i_data_writeres[13]), .B(n41), .C(i_data_rs[13]), .D(n7), 
        .Q(n101) );
  AOI220 U13 ( .A(i_data_writeres[15]), .B(n5), .C(i_data_rs[15]), .D(n42), 
        .Q(n95) );
  AOI220 U14 ( .A(i_data_writeres[16]), .B(n41), .C(i_data_rs[16]), .D(n7), 
        .Q(n92) );
  AOI220 U15 ( .A(i_data_writeres[18]), .B(n41), .C(i_data_rs[18]), .D(n42), 
        .Q(n86) );
  AOI220 U16 ( .A(i_data_writeres[19]), .B(n41), .C(i_data_rs[19]), .D(n7), 
        .Q(n83) );
  AOI220 U17 ( .A(i_data_writeres[21]), .B(n5), .C(i_data_rs[21]), .D(n42), 
        .Q(n77) );
  AOI220 U18 ( .A(i_data_writeres[22]), .B(n41), .C(i_data_rs[22]), .D(n7), 
        .Q(n74) );
  AOI220 U19 ( .A(i_data_writeres[24]), .B(n41), .C(i_data_rs[24]), .D(n42), 
        .Q(n68) );
  AOI220 U20 ( .A(i_data_writeres[25]), .B(n41), .C(i_data_rs[25]), .D(n7), 
        .Q(n65) );
  AOI220 U21 ( .A(i_data_writeres[27]), .B(n5), .C(i_data_rs[27]), .D(n42), 
        .Q(n59) );
  AOI220 U22 ( .A(i_data_writeres[28]), .B(n41), .C(i_data_rs[28]), .D(n7), 
        .Q(n56) );
  AOI220 U23 ( .A(i_data_writeres[30]), .B(n41), .C(i_data_rs[30]), .D(n7), 
        .Q(n50) );
  AOI220 U24 ( .A(i_data_writeres[31]), .B(n5), .C(i_data_rs[31]), .D(n7), .Q(
        n40) );
  AOI220 U25 ( .A(i_data_writeres[2]), .B(n5), .C(i_data_rs[2]), .D(n7), .Q(
        n134) );
  AOI220 U26 ( .A(i_data_writeres[5]), .B(n5), .C(i_data_rs[5]), .D(n42), .Q(
        n125) );
  AOI220 U27 ( .A(i_data_writeres[8]), .B(n5), .C(i_data_rs[8]), .D(n7), .Q(
        n116) );
  AOI220 U28 ( .A(i_data_writeres[11]), .B(n5), .C(i_data_rs[11]), .D(n42), 
        .Q(n107) );
  AOI220 U29 ( .A(i_data_writeres[14]), .B(n5), .C(i_data_rs[14]), .D(n7), .Q(
        n98) );
  AOI220 U30 ( .A(i_data_writeres[17]), .B(n5), .C(i_data_rs[17]), .D(n42), 
        .Q(n89) );
  AOI220 U31 ( .A(i_data_writeres[20]), .B(n5), .C(i_data_rs[20]), .D(n7), .Q(
        n80) );
  AOI220 U32 ( .A(i_data_writeres[23]), .B(n5), .C(i_data_rs[23]), .D(n42), 
        .Q(n71) );
  AOI220 U33 ( .A(i_data_writeres[26]), .B(n5), .C(i_data_rs[26]), .D(n7), .Q(
        n62) );
  AOI220 U34 ( .A(i_data_writeres[29]), .B(n5), .C(i_data_rs[29]), .D(n42), 
        .Q(n53) );
  BUF2 U35 ( .A(n46), .Q(n8) );
  NOR40 U36 ( .A(n44), .B(n3), .C(n11), .D(n9), .Q(n46) );
  INV3 U37 ( .A(n47), .Q(n11) );
  NOR21 U38 ( .A(n42), .B(n5), .Q(n47) );
  BUF2 U39 ( .A(n44), .Q(n1) );
  BUF2 U40 ( .A(n45), .Q(n3) );
  INV3 U41 ( .A(n4), .Q(n5) );
  INV3 U42 ( .A(n6), .Q(n7) );
  BUF2 U43 ( .A(n43), .Q(n9) );
  NOR31 U44 ( .A(i_con_fa[0]), .B(i_con_fa[2]), .C(n12), .Q(n43) );
  INV3 U45 ( .A(i_con_fa[1]), .Q(n12) );
  NOR31 U46 ( .A(i_con_fa[0]), .B(i_con_fa[1]), .C(n10), .Q(n45) );
  NOR31 U47 ( .A(n13), .B(i_con_fa[1]), .C(n10), .Q(n44) );
  NAND31 U48 ( .A(n132), .B(n133), .C(n134), .Q(N24) );
  NAND22 U49 ( .A(i_data_alures[2]), .B(n9), .Q(n133) );
  AOI221 U50 ( .A(i_data_lwW[2]), .B(n44), .C(i_data_lwM[2]), .D(n3), .Q(n132)
         );
  NAND31 U51 ( .A(n123), .B(n124), .C(n125), .Q(N27) );
  NAND22 U52 ( .A(i_data_alures[5]), .B(n9), .Q(n124) );
  AOI221 U53 ( .A(i_data_lwW[5]), .B(n44), .C(i_data_lwM[5]), .D(n3), .Q(n123)
         );
  NAND31 U54 ( .A(n114), .B(n115), .C(n116), .Q(N30) );
  NAND22 U55 ( .A(i_data_alures[8]), .B(n43), .Q(n115) );
  AOI221 U56 ( .A(i_data_lwW[8]), .B(n44), .C(i_data_lwM[8]), .D(n3), .Q(n114)
         );
  NAND31 U57 ( .A(n105), .B(n106), .C(n107), .Q(N33) );
  NAND22 U58 ( .A(i_data_alures[11]), .B(n43), .Q(n106) );
  AOI221 U59 ( .A(i_data_lwW[11]), .B(n44), .C(i_data_lwM[11]), .D(n3), .Q(
        n105) );
  NAND31 U60 ( .A(n96), .B(n97), .C(n98), .Q(N36) );
  NAND22 U61 ( .A(i_data_alures[14]), .B(n43), .Q(n97) );
  AOI221 U62 ( .A(i_data_lwW[14]), .B(n44), .C(i_data_lwM[14]), .D(n3), .Q(n96) );
  NAND31 U63 ( .A(n87), .B(n88), .C(n89), .Q(N39) );
  NAND22 U64 ( .A(i_data_alures[17]), .B(n43), .Q(n88) );
  AOI221 U65 ( .A(i_data_lwW[17]), .B(n1), .C(i_data_lwM[17]), .D(n45), .Q(n87) );
  NAND31 U66 ( .A(n78), .B(n79), .C(n80), .Q(N42) );
  NAND22 U67 ( .A(i_data_alures[20]), .B(n43), .Q(n79) );
  AOI221 U68 ( .A(i_data_lwW[20]), .B(n1), .C(i_data_lwM[20]), .D(n45), .Q(n78) );
  NAND31 U69 ( .A(n69), .B(n70), .C(n71), .Q(N45) );
  NAND22 U70 ( .A(i_data_alures[23]), .B(n43), .Q(n70) );
  AOI221 U71 ( .A(i_data_lwW[23]), .B(n1), .C(i_data_lwM[23]), .D(n45), .Q(n69) );
  NAND31 U72 ( .A(n60), .B(n61), .C(n62), .Q(N48) );
  NAND22 U73 ( .A(i_data_alures[26]), .B(n9), .Q(n61) );
  AOI221 U74 ( .A(i_data_lwW[26]), .B(n1), .C(i_data_lwM[26]), .D(n45), .Q(n60) );
  NAND31 U75 ( .A(n51), .B(n52), .C(n53), .Q(N51) );
  NAND22 U76 ( .A(i_data_alures[29]), .B(n43), .Q(n52) );
  AOI221 U77 ( .A(i_data_lwW[29]), .B(n1), .C(i_data_lwM[29]), .D(n45), .Q(n51) );
  NAND31 U78 ( .A(n138), .B(n139), .C(n140), .Q(N22) );
  NAND22 U79 ( .A(i_data_alures[0]), .B(n9), .Q(n139) );
  AOI221 U80 ( .A(i_data_lwW[0]), .B(n44), .C(i_data_lwM[0]), .D(n3), .Q(n138)
         );
  NAND31 U81 ( .A(n135), .B(n136), .C(n137), .Q(N23) );
  NAND22 U82 ( .A(i_data_alures[1]), .B(n9), .Q(n136) );
  AOI221 U83 ( .A(i_data_lwW[1]), .B(n44), .C(i_data_lwM[1]), .D(n3), .Q(n135)
         );
  NAND31 U84 ( .A(n129), .B(n130), .C(n131), .Q(N25) );
  NAND22 U85 ( .A(i_data_alures[3]), .B(n9), .Q(n130) );
  AOI221 U86 ( .A(i_data_lwW[3]), .B(n44), .C(i_data_lwM[3]), .D(n3), .Q(n129)
         );
  NAND31 U87 ( .A(n126), .B(n127), .C(n128), .Q(N26) );
  NAND22 U88 ( .A(i_data_alures[4]), .B(n9), .Q(n127) );
  AOI221 U89 ( .A(i_data_lwW[4]), .B(n44), .C(i_data_lwM[4]), .D(n3), .Q(n126)
         );
  NAND31 U90 ( .A(n120), .B(n121), .C(n122), .Q(N28) );
  NAND22 U91 ( .A(i_data_alures[6]), .B(n9), .Q(n121) );
  AOI221 U92 ( .A(i_data_lwW[6]), .B(n44), .C(i_data_lwM[6]), .D(n3), .Q(n120)
         );
  NAND31 U93 ( .A(n117), .B(n118), .C(n119), .Q(N29) );
  NAND22 U94 ( .A(i_data_alures[7]), .B(n43), .Q(n118) );
  NAND31 U95 ( .A(n111), .B(n112), .C(n113), .Q(N31) );
  NAND22 U96 ( .A(i_data_alures[9]), .B(n43), .Q(n112) );
  AOI221 U97 ( .A(i_data_lwW[9]), .B(n44), .C(i_data_lwM[9]), .D(n3), .Q(n111)
         );
  NAND31 U98 ( .A(n108), .B(n109), .C(n110), .Q(N32) );
  NAND22 U99 ( .A(i_data_alures[10]), .B(n9), .Q(n109) );
  AOI221 U100 ( .A(i_data_lwW[10]), .B(n44), .C(i_data_lwM[10]), .D(n3), .Q(
        n108) );
  NAND31 U101 ( .A(n102), .B(n103), .C(n104), .Q(N34) );
  NAND22 U102 ( .A(i_data_alures[12]), .B(n43), .Q(n103) );
  AOI221 U103 ( .A(i_data_lwW[12]), .B(n44), .C(i_data_lwM[12]), .D(n3), .Q(
        n102) );
  NAND31 U104 ( .A(n99), .B(n100), .C(n101), .Q(N35) );
  NAND22 U105 ( .A(i_data_alures[13]), .B(n9), .Q(n100) );
  AOI221 U106 ( .A(i_data_lwW[13]), .B(n44), .C(i_data_lwM[13]), .D(n3), .Q(
        n99) );
  NAND31 U107 ( .A(n93), .B(n94), .C(n95), .Q(N37) );
  NAND22 U108 ( .A(i_data_alures[15]), .B(n43), .Q(n94) );
  AOI221 U109 ( .A(i_data_lwW[15]), .B(n1), .C(i_data_lwM[15]), .D(n45), .Q(
        n93) );
  NAND31 U110 ( .A(n90), .B(n91), .C(n92), .Q(N38) );
  NAND22 U111 ( .A(i_data_alures[16]), .B(n9), .Q(n91) );
  AOI221 U112 ( .A(i_data_lwW[16]), .B(n1), .C(i_data_lwM[16]), .D(n45), .Q(
        n90) );
  NAND31 U113 ( .A(n84), .B(n85), .C(n86), .Q(N40) );
  NAND22 U114 ( .A(i_data_alures[18]), .B(n43), .Q(n85) );
  AOI221 U115 ( .A(i_data_lwW[18]), .B(n1), .C(i_data_lwM[18]), .D(n45), .Q(
        n84) );
  NAND31 U116 ( .A(n81), .B(n82), .C(n83), .Q(N41) );
  NAND22 U117 ( .A(i_data_alures[19]), .B(n9), .Q(n82) );
  AOI221 U118 ( .A(i_data_lwW[19]), .B(n1), .C(i_data_lwM[19]), .D(n45), .Q(
        n81) );
  NAND31 U119 ( .A(n75), .B(n76), .C(n77), .Q(N43) );
  NAND22 U120 ( .A(i_data_alures[21]), .B(n9), .Q(n76) );
  AOI221 U121 ( .A(i_data_lwW[21]), .B(n1), .C(i_data_lwM[21]), .D(n45), .Q(
        n75) );
  NAND31 U122 ( .A(n72), .B(n73), .C(n74), .Q(N44) );
  NAND22 U123 ( .A(i_data_alures[22]), .B(n9), .Q(n73) );
  AOI221 U124 ( .A(i_data_lwW[22]), .B(n1), .C(i_data_lwM[22]), .D(n45), .Q(
        n72) );
  NAND31 U125 ( .A(n66), .B(n67), .C(n68), .Q(N46) );
  NAND22 U126 ( .A(i_data_alures[24]), .B(n9), .Q(n67) );
  AOI221 U127 ( .A(i_data_lwW[24]), .B(n1), .C(i_data_lwM[24]), .D(n45), .Q(
        n66) );
  NAND31 U128 ( .A(n63), .B(n64), .C(n65), .Q(N47) );
  NAND22 U129 ( .A(i_data_alures[25]), .B(n9), .Q(n64) );
  AOI221 U130 ( .A(i_data_lwW[25]), .B(n1), .C(i_data_lwM[25]), .D(n45), .Q(
        n63) );
  NAND31 U131 ( .A(n57), .B(n58), .C(n59), .Q(N49) );
  NAND22 U132 ( .A(i_data_alures[27]), .B(n9), .Q(n58) );
  AOI221 U133 ( .A(i_data_lwW[27]), .B(n1), .C(i_data_lwM[27]), .D(n45), .Q(
        n57) );
  NAND31 U134 ( .A(n54), .B(n55), .C(n56), .Q(N50) );
  NAND22 U135 ( .A(i_data_alures[28]), .B(n9), .Q(n55) );
  AOI221 U136 ( .A(i_data_lwW[28]), .B(n1), .C(i_data_lwM[28]), .D(n45), .Q(
        n54) );
  NAND31 U137 ( .A(n48), .B(n49), .C(n50), .Q(N52) );
  NAND22 U138 ( .A(i_data_alures[30]), .B(n9), .Q(n49) );
  AOI221 U139 ( .A(i_data_lwW[30]), .B(n1), .C(i_data_lwM[30]), .D(n3), .Q(n48) );
  NAND31 U140 ( .A(n38), .B(n39), .C(n40), .Q(N54) );
  NAND22 U141 ( .A(i_data_alures[31]), .B(n9), .Q(n39) );
  AOI221 U142 ( .A(i_data_lwW[31]), .B(n1), .C(i_data_lwM[31]), .D(n3), .Q(n38) );
  INV3 U143 ( .A(n42), .Q(n6) );
  NOR31 U144 ( .A(i_con_fa[1]), .B(i_con_fa[2]), .C(i_con_fa[0]), .Q(n42) );
  INV3 U145 ( .A(n41), .Q(n4) );
  NOR31 U146 ( .A(i_con_fa[1]), .B(i_con_fa[2]), .C(n13), .Q(n41) );
  INV3 U147 ( .A(i_con_fa[0]), .Q(n13) );
  INV3 U148 ( .A(i_con_fa[2]), .Q(n10) );
  LOGIC1 U149 ( .Q(n2) );
endmodule


module E_fbmux5 ( i_data_rt, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fb, o_data_alusrb );
  input [31:0] i_data_rt;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fb;
  output [31:0] o_data_alusrb;
  wire   N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N54, n2, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13;

  DLPQ3 o_data_alusrb_reg_31_ ( .SN(n2), .D(N54), .GN(n46), .Q(
        o_data_alusrb[31]) );
  DLPQ3 o_data_alusrb_reg_30_ ( .SN(n2), .D(N52), .GN(n46), .Q(
        o_data_alusrb[30]) );
  DLPQ3 o_data_alusrb_reg_29_ ( .SN(n2), .D(N51), .GN(n46), .Q(
        o_data_alusrb[29]) );
  DLPQ3 o_data_alusrb_reg_28_ ( .SN(n2), .D(N50), .GN(n46), .Q(
        o_data_alusrb[28]) );
  DLPQ3 o_data_alusrb_reg_27_ ( .SN(n2), .D(N49), .GN(n8), .Q(
        o_data_alusrb[27]) );
  DLPQ3 o_data_alusrb_reg_26_ ( .SN(n2), .D(N48), .GN(n8), .Q(
        o_data_alusrb[26]) );
  DLPQ3 o_data_alusrb_reg_25_ ( .SN(n2), .D(N47), .GN(n46), .Q(
        o_data_alusrb[25]) );
  DLPQ3 o_data_alusrb_reg_24_ ( .SN(n2), .D(N46), .GN(n46), .Q(
        o_data_alusrb[24]) );
  DLPQ3 o_data_alusrb_reg_23_ ( .SN(n2), .D(N45), .GN(n8), .Q(
        o_data_alusrb[23]) );
  DLPQ3 o_data_alusrb_reg_22_ ( .SN(n2), .D(N44), .GN(n8), .Q(
        o_data_alusrb[22]) );
  DLPQ3 o_data_alusrb_reg_21_ ( .SN(n2), .D(N43), .GN(n8), .Q(
        o_data_alusrb[21]) );
  DLPQ3 o_data_alusrb_reg_20_ ( .SN(n2), .D(N42), .GN(n8), .Q(
        o_data_alusrb[20]) );
  DLPQ3 o_data_alusrb_reg_19_ ( .SN(n2), .D(N41), .GN(n8), .Q(
        o_data_alusrb[19]) );
  DLPQ3 o_data_alusrb_reg_18_ ( .SN(n2), .D(N40), .GN(n8), .Q(
        o_data_alusrb[18]) );
  DLPQ3 o_data_alusrb_reg_17_ ( .SN(n2), .D(N39), .GN(n8), .Q(
        o_data_alusrb[17]) );
  DLPQ3 o_data_alusrb_reg_16_ ( .SN(n2), .D(N38), .GN(n46), .Q(
        o_data_alusrb[16]) );
  DLPQ3 o_data_alusrb_reg_15_ ( .SN(n2), .D(N37), .GN(n8), .Q(
        o_data_alusrb[15]) );
  DLPQ3 o_data_alusrb_reg_14_ ( .SN(n2), .D(N36), .GN(n8), .Q(
        o_data_alusrb[14]) );
  DLPQ3 o_data_alusrb_reg_13_ ( .SN(n2), .D(N35), .GN(n8), .Q(
        o_data_alusrb[13]) );
  DLPQ3 o_data_alusrb_reg_12_ ( .SN(n2), .D(N34), .GN(n8), .Q(
        o_data_alusrb[12]) );
  DLPQ3 o_data_alusrb_reg_11_ ( .SN(n2), .D(N33), .GN(n8), .Q(
        o_data_alusrb[11]) );
  DLPQ3 o_data_alusrb_reg_10_ ( .SN(n2), .D(N32), .GN(n8), .Q(
        o_data_alusrb[10]) );
  DLPQ3 o_data_alusrb_reg_9_ ( .SN(n2), .D(N31), .GN(n46), .Q(o_data_alusrb[9]) );
  DLPQ3 o_data_alusrb_reg_8_ ( .SN(n2), .D(N30), .GN(n8), .Q(o_data_alusrb[8])
         );
  DLPQ3 o_data_alusrb_reg_7_ ( .SN(n2), .D(N29), .GN(n8), .Q(o_data_alusrb[7])
         );
  DLPQ3 o_data_alusrb_reg_6_ ( .SN(n2), .D(N28), .GN(n8), .Q(o_data_alusrb[6])
         );
  DLPQ3 o_data_alusrb_reg_5_ ( .SN(n2), .D(N27), .GN(n8), .Q(o_data_alusrb[5])
         );
  DLPQ3 o_data_alusrb_reg_4_ ( .SN(n2), .D(N26), .GN(n8), .Q(o_data_alusrb[4])
         );
  DLPQ3 o_data_alusrb_reg_3_ ( .SN(n2), .D(N25), .GN(n8), .Q(o_data_alusrb[3])
         );
  DLPQ3 o_data_alusrb_reg_2_ ( .SN(n2), .D(N24), .GN(n8), .Q(o_data_alusrb[2])
         );
  DLPQ3 o_data_alusrb_reg_1_ ( .SN(n2), .D(N23), .GN(n8), .Q(o_data_alusrb[1])
         );
  DLPQ3 o_data_alusrb_reg_0_ ( .SN(n2), .D(N22), .GN(n8), .Q(o_data_alusrb[0])
         );
  AOI220 U2 ( .A(i_data_writeres[0]), .B(n41), .C(i_data_rt[0]), .D(n42), .Q(
        n140) );
  AOI220 U3 ( .A(i_data_writeres[1]), .B(n41), .C(i_data_rt[1]), .D(n7), .Q(
        n137) );
  AOI220 U4 ( .A(i_data_writeres[3]), .B(n5), .C(i_data_rt[3]), .D(n42), .Q(
        n131) );
  AOI220 U5 ( .A(i_data_writeres[4]), .B(n41), .C(i_data_rt[4]), .D(n7), .Q(
        n128) );
  AOI220 U6 ( .A(i_data_writeres[6]), .B(n41), .C(i_data_rt[6]), .D(n42), .Q(
        n122) );
  AOI220 U7 ( .A(i_data_lwW[7]), .B(n44), .C(i_data_lwM[7]), .D(n3), .Q(n117)
         );
  AOI220 U8 ( .A(i_data_writeres[7]), .B(n41), .C(i_data_rt[7]), .D(n7), .Q(
        n119) );
  AOI220 U9 ( .A(i_data_writeres[9]), .B(n5), .C(i_data_rt[9]), .D(n42), .Q(
        n113) );
  AOI220 U10 ( .A(i_data_writeres[10]), .B(n41), .C(i_data_rt[10]), .D(n7), 
        .Q(n110) );
  AOI220 U11 ( .A(i_data_writeres[12]), .B(n41), .C(i_data_rt[12]), .D(n42), 
        .Q(n104) );
  AOI220 U12 ( .A(i_data_writeres[13]), .B(n41), .C(i_data_rt[13]), .D(n7), 
        .Q(n101) );
  AOI220 U13 ( .A(i_data_writeres[15]), .B(n5), .C(i_data_rt[15]), .D(n42), 
        .Q(n95) );
  AOI220 U14 ( .A(i_data_writeres[16]), .B(n41), .C(i_data_rt[16]), .D(n7), 
        .Q(n92) );
  AOI220 U15 ( .A(i_data_writeres[18]), .B(n41), .C(i_data_rt[18]), .D(n42), 
        .Q(n86) );
  AOI220 U16 ( .A(i_data_writeres[19]), .B(n41), .C(i_data_rt[19]), .D(n7), 
        .Q(n83) );
  AOI220 U17 ( .A(i_data_writeres[21]), .B(n5), .C(i_data_rt[21]), .D(n42), 
        .Q(n77) );
  AOI220 U18 ( .A(i_data_writeres[22]), .B(n41), .C(i_data_rt[22]), .D(n7), 
        .Q(n74) );
  AOI220 U19 ( .A(i_data_writeres[24]), .B(n41), .C(i_data_rt[24]), .D(n42), 
        .Q(n68) );
  AOI220 U20 ( .A(i_data_writeres[25]), .B(n41), .C(i_data_rt[25]), .D(n7), 
        .Q(n65) );
  AOI220 U21 ( .A(i_data_writeres[27]), .B(n5), .C(i_data_rt[27]), .D(n42), 
        .Q(n59) );
  AOI220 U22 ( .A(i_data_writeres[28]), .B(n41), .C(i_data_rt[28]), .D(n7), 
        .Q(n56) );
  AOI220 U23 ( .A(i_data_writeres[30]), .B(n41), .C(i_data_rt[30]), .D(n7), 
        .Q(n50) );
  AOI220 U24 ( .A(i_data_writeres[31]), .B(n5), .C(i_data_rt[31]), .D(n7), .Q(
        n40) );
  AOI220 U25 ( .A(i_data_writeres[2]), .B(n5), .C(i_data_rt[2]), .D(n7), .Q(
        n134) );
  AOI220 U26 ( .A(i_data_writeres[5]), .B(n5), .C(i_data_rt[5]), .D(n42), .Q(
        n125) );
  AOI220 U27 ( .A(i_data_writeres[8]), .B(n5), .C(i_data_rt[8]), .D(n7), .Q(
        n116) );
  AOI220 U28 ( .A(i_data_writeres[11]), .B(n5), .C(i_data_rt[11]), .D(n42), 
        .Q(n107) );
  AOI220 U29 ( .A(i_data_writeres[14]), .B(n5), .C(i_data_rt[14]), .D(n7), .Q(
        n98) );
  AOI220 U30 ( .A(i_data_writeres[17]), .B(n5), .C(i_data_rt[17]), .D(n42), 
        .Q(n89) );
  AOI220 U31 ( .A(i_data_writeres[20]), .B(n5), .C(i_data_rt[20]), .D(n7), .Q(
        n80) );
  AOI220 U32 ( .A(i_data_writeres[23]), .B(n5), .C(i_data_rt[23]), .D(n42), 
        .Q(n71) );
  AOI220 U33 ( .A(i_data_writeres[26]), .B(n5), .C(i_data_rt[26]), .D(n7), .Q(
        n62) );
  AOI220 U34 ( .A(i_data_writeres[29]), .B(n5), .C(i_data_rt[29]), .D(n42), 
        .Q(n53) );
  BUF2 U35 ( .A(n46), .Q(n8) );
  NOR40 U36 ( .A(n44), .B(n3), .C(n11), .D(n9), .Q(n46) );
  INV3 U37 ( .A(n47), .Q(n11) );
  NOR21 U38 ( .A(n42), .B(n5), .Q(n47) );
  BUF2 U39 ( .A(n44), .Q(n1) );
  BUF2 U40 ( .A(n45), .Q(n3) );
  INV3 U41 ( .A(n4), .Q(n5) );
  INV3 U42 ( .A(n6), .Q(n7) );
  BUF2 U43 ( .A(n43), .Q(n9) );
  NOR31 U44 ( .A(i_con_fb[0]), .B(i_con_fb[2]), .C(n12), .Q(n43) );
  INV3 U45 ( .A(i_con_fb[1]), .Q(n12) );
  NOR31 U46 ( .A(i_con_fb[0]), .B(i_con_fb[1]), .C(n10), .Q(n45) );
  NOR31 U47 ( .A(n13), .B(i_con_fb[1]), .C(n10), .Q(n44) );
  NAND31 U48 ( .A(n132), .B(n133), .C(n134), .Q(N24) );
  NAND22 U49 ( .A(i_data_alures[2]), .B(n9), .Q(n133) );
  AOI221 U50 ( .A(i_data_lwW[2]), .B(n44), .C(i_data_lwM[2]), .D(n3), .Q(n132)
         );
  NAND31 U51 ( .A(n123), .B(n124), .C(n125), .Q(N27) );
  NAND22 U52 ( .A(i_data_alures[5]), .B(n9), .Q(n124) );
  AOI221 U53 ( .A(i_data_lwW[5]), .B(n44), .C(i_data_lwM[5]), .D(n3), .Q(n123)
         );
  NAND31 U54 ( .A(n114), .B(n115), .C(n116), .Q(N30) );
  NAND22 U55 ( .A(i_data_alures[8]), .B(n43), .Q(n115) );
  AOI221 U56 ( .A(i_data_lwW[8]), .B(n44), .C(i_data_lwM[8]), .D(n3), .Q(n114)
         );
  NAND31 U57 ( .A(n105), .B(n106), .C(n107), .Q(N33) );
  NAND22 U58 ( .A(i_data_alures[11]), .B(n43), .Q(n106) );
  AOI221 U59 ( .A(i_data_lwW[11]), .B(n44), .C(i_data_lwM[11]), .D(n3), .Q(
        n105) );
  NAND31 U60 ( .A(n96), .B(n97), .C(n98), .Q(N36) );
  NAND22 U61 ( .A(i_data_alures[14]), .B(n43), .Q(n97) );
  AOI221 U62 ( .A(i_data_lwW[14]), .B(n44), .C(i_data_lwM[14]), .D(n3), .Q(n96) );
  NAND31 U63 ( .A(n87), .B(n88), .C(n89), .Q(N39) );
  NAND22 U64 ( .A(i_data_alures[17]), .B(n43), .Q(n88) );
  AOI221 U65 ( .A(i_data_lwW[17]), .B(n1), .C(i_data_lwM[17]), .D(n45), .Q(n87) );
  NAND31 U66 ( .A(n78), .B(n79), .C(n80), .Q(N42) );
  NAND22 U67 ( .A(i_data_alures[20]), .B(n43), .Q(n79) );
  AOI221 U68 ( .A(i_data_lwW[20]), .B(n1), .C(i_data_lwM[20]), .D(n45), .Q(n78) );
  NAND31 U69 ( .A(n69), .B(n70), .C(n71), .Q(N45) );
  NAND22 U70 ( .A(i_data_alures[23]), .B(n43), .Q(n70) );
  AOI221 U71 ( .A(i_data_lwW[23]), .B(n1), .C(i_data_lwM[23]), .D(n45), .Q(n69) );
  NAND31 U72 ( .A(n60), .B(n61), .C(n62), .Q(N48) );
  NAND22 U73 ( .A(i_data_alures[26]), .B(n9), .Q(n61) );
  AOI221 U74 ( .A(i_data_lwW[26]), .B(n1), .C(i_data_lwM[26]), .D(n45), .Q(n60) );
  NAND31 U75 ( .A(n51), .B(n52), .C(n53), .Q(N51) );
  NAND22 U76 ( .A(i_data_alures[29]), .B(n43), .Q(n52) );
  AOI221 U77 ( .A(i_data_lwW[29]), .B(n1), .C(i_data_lwM[29]), .D(n45), .Q(n51) );
  NAND31 U78 ( .A(n138), .B(n139), .C(n140), .Q(N22) );
  NAND22 U79 ( .A(i_data_alures[0]), .B(n9), .Q(n139) );
  AOI221 U80 ( .A(i_data_lwW[0]), .B(n44), .C(i_data_lwM[0]), .D(n3), .Q(n138)
         );
  NAND31 U81 ( .A(n135), .B(n136), .C(n137), .Q(N23) );
  NAND22 U82 ( .A(i_data_alures[1]), .B(n9), .Q(n136) );
  AOI221 U83 ( .A(i_data_lwW[1]), .B(n44), .C(i_data_lwM[1]), .D(n3), .Q(n135)
         );
  NAND31 U84 ( .A(n129), .B(n130), .C(n131), .Q(N25) );
  NAND22 U85 ( .A(i_data_alures[3]), .B(n9), .Q(n130) );
  AOI221 U86 ( .A(i_data_lwW[3]), .B(n44), .C(i_data_lwM[3]), .D(n3), .Q(n129)
         );
  NAND31 U87 ( .A(n126), .B(n127), .C(n128), .Q(N26) );
  NAND22 U88 ( .A(i_data_alures[4]), .B(n9), .Q(n127) );
  AOI221 U89 ( .A(i_data_lwW[4]), .B(n44), .C(i_data_lwM[4]), .D(n3), .Q(n126)
         );
  NAND31 U90 ( .A(n120), .B(n121), .C(n122), .Q(N28) );
  NAND22 U91 ( .A(i_data_alures[6]), .B(n9), .Q(n121) );
  AOI221 U92 ( .A(i_data_lwW[6]), .B(n44), .C(i_data_lwM[6]), .D(n3), .Q(n120)
         );
  NAND31 U93 ( .A(n117), .B(n118), .C(n119), .Q(N29) );
  NAND22 U94 ( .A(i_data_alures[7]), .B(n43), .Q(n118) );
  NAND31 U95 ( .A(n111), .B(n112), .C(n113), .Q(N31) );
  NAND22 U96 ( .A(i_data_alures[9]), .B(n43), .Q(n112) );
  AOI221 U97 ( .A(i_data_lwW[9]), .B(n44), .C(i_data_lwM[9]), .D(n3), .Q(n111)
         );
  NAND31 U98 ( .A(n108), .B(n109), .C(n110), .Q(N32) );
  NAND22 U99 ( .A(i_data_alures[10]), .B(n9), .Q(n109) );
  AOI221 U100 ( .A(i_data_lwW[10]), .B(n44), .C(i_data_lwM[10]), .D(n3), .Q(
        n108) );
  NAND31 U101 ( .A(n102), .B(n103), .C(n104), .Q(N34) );
  NAND22 U102 ( .A(i_data_alures[12]), .B(n43), .Q(n103) );
  AOI221 U103 ( .A(i_data_lwW[12]), .B(n44), .C(i_data_lwM[12]), .D(n3), .Q(
        n102) );
  NAND31 U104 ( .A(n99), .B(n100), .C(n101), .Q(N35) );
  NAND22 U105 ( .A(i_data_alures[13]), .B(n9), .Q(n100) );
  AOI221 U106 ( .A(i_data_lwW[13]), .B(n44), .C(i_data_lwM[13]), .D(n3), .Q(
        n99) );
  NAND31 U107 ( .A(n93), .B(n94), .C(n95), .Q(N37) );
  NAND22 U108 ( .A(i_data_alures[15]), .B(n43), .Q(n94) );
  AOI221 U109 ( .A(i_data_lwW[15]), .B(n1), .C(i_data_lwM[15]), .D(n45), .Q(
        n93) );
  NAND31 U110 ( .A(n90), .B(n91), .C(n92), .Q(N38) );
  NAND22 U111 ( .A(i_data_alures[16]), .B(n9), .Q(n91) );
  AOI221 U112 ( .A(i_data_lwW[16]), .B(n1), .C(i_data_lwM[16]), .D(n45), .Q(
        n90) );
  NAND31 U113 ( .A(n84), .B(n85), .C(n86), .Q(N40) );
  NAND22 U114 ( .A(i_data_alures[18]), .B(n43), .Q(n85) );
  AOI221 U115 ( .A(i_data_lwW[18]), .B(n1), .C(i_data_lwM[18]), .D(n45), .Q(
        n84) );
  NAND31 U116 ( .A(n81), .B(n82), .C(n83), .Q(N41) );
  NAND22 U117 ( .A(i_data_alures[19]), .B(n9), .Q(n82) );
  AOI221 U118 ( .A(i_data_lwW[19]), .B(n1), .C(i_data_lwM[19]), .D(n45), .Q(
        n81) );
  NAND31 U119 ( .A(n75), .B(n76), .C(n77), .Q(N43) );
  NAND22 U120 ( .A(i_data_alures[21]), .B(n9), .Q(n76) );
  AOI221 U121 ( .A(i_data_lwW[21]), .B(n1), .C(i_data_lwM[21]), .D(n45), .Q(
        n75) );
  NAND31 U122 ( .A(n72), .B(n73), .C(n74), .Q(N44) );
  NAND22 U123 ( .A(i_data_alures[22]), .B(n9), .Q(n73) );
  AOI221 U124 ( .A(i_data_lwW[22]), .B(n1), .C(i_data_lwM[22]), .D(n45), .Q(
        n72) );
  NAND31 U125 ( .A(n66), .B(n67), .C(n68), .Q(N46) );
  NAND22 U126 ( .A(i_data_alures[24]), .B(n9), .Q(n67) );
  AOI221 U127 ( .A(i_data_lwW[24]), .B(n1), .C(i_data_lwM[24]), .D(n45), .Q(
        n66) );
  NAND31 U128 ( .A(n63), .B(n64), .C(n65), .Q(N47) );
  NAND22 U129 ( .A(i_data_alures[25]), .B(n9), .Q(n64) );
  AOI221 U130 ( .A(i_data_lwW[25]), .B(n1), .C(i_data_lwM[25]), .D(n45), .Q(
        n63) );
  NAND31 U131 ( .A(n57), .B(n58), .C(n59), .Q(N49) );
  NAND22 U132 ( .A(i_data_alures[27]), .B(n9), .Q(n58) );
  AOI221 U133 ( .A(i_data_lwW[27]), .B(n1), .C(i_data_lwM[27]), .D(n45), .Q(
        n57) );
  NAND31 U134 ( .A(n54), .B(n55), .C(n56), .Q(N50) );
  NAND22 U135 ( .A(i_data_alures[28]), .B(n9), .Q(n55) );
  AOI221 U136 ( .A(i_data_lwW[28]), .B(n1), .C(i_data_lwM[28]), .D(n45), .Q(
        n54) );
  NAND31 U137 ( .A(n48), .B(n49), .C(n50), .Q(N52) );
  NAND22 U138 ( .A(i_data_alures[30]), .B(n9), .Q(n49) );
  AOI221 U139 ( .A(i_data_lwW[30]), .B(n1), .C(i_data_lwM[30]), .D(n3), .Q(n48) );
  NAND31 U140 ( .A(n38), .B(n39), .C(n40), .Q(N54) );
  NAND22 U141 ( .A(i_data_alures[31]), .B(n9), .Q(n39) );
  AOI221 U142 ( .A(i_data_lwW[31]), .B(n1), .C(i_data_lwM[31]), .D(n3), .Q(n38) );
  INV3 U143 ( .A(n42), .Q(n6) );
  NOR31 U144 ( .A(i_con_fb[1]), .B(i_con_fb[2]), .C(i_con_fb[0]), .Q(n42) );
  INV3 U145 ( .A(n41), .Q(n4) );
  NOR31 U146 ( .A(i_con_fb[1]), .B(i_con_fb[2]), .C(n13), .Q(n41) );
  INV3 U147 ( .A(i_con_fb[0]), .Q(n13) );
  INV3 U148 ( .A(i_con_fb[2]), .Q(n10) );
  LOGIC1 U149 ( .Q(n2) );
endmodule


module E_alubmux ( i_data_fb, i_data_imm, i_con_imm, o_data_alub );
  input [31:0] i_data_fb;
  input [31:0] i_data_imm;
  output [31:0] o_data_alub;
  input i_con_imm;
  wire   n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  CLKIN1 U1 ( .A(i_data_imm[3]), .Q(n21) );
  NAND23 U2 ( .A(n20), .B(n19), .Q(o_data_alub[2]) );
  INV3 U3 ( .A(i_data_imm[11]), .Q(n28) );
  INV3 U4 ( .A(i_data_imm[4]), .Q(n23) );
  MUX22 U5 ( .A(i_data_fb[31]), .B(i_data_imm[31]), .S(n14), .Q(
        o_data_alub[31]) );
  CLKIN6 U6 ( .A(n10), .Q(o_data_alub[5]) );
  CLKIN8 U7 ( .A(n8), .Q(o_data_alub[6]) );
  INV3 U8 ( .A(n12), .Q(n9) );
  INV3 U9 ( .A(i_data_imm[13]), .Q(n32) );
  INV3 U10 ( .A(i_data_imm[14]), .Q(n34) );
  NAND21 U11 ( .A(i_data_imm[0]), .B(n15), .Q(n6) );
  NAND20 U12 ( .A(i_data_fb[20]), .B(n16), .Q(n47) );
  INV2 U13 ( .A(n16), .Q(n3) );
  IMUX22 U14 ( .A(n24), .B(n23), .S(n1), .Q(o_data_alub[4]) );
  INV15 U15 ( .A(n16), .Q(n1) );
  INV12 U16 ( .A(n16), .Q(n14) );
  MUX24 U17 ( .A(i_data_fb[7]), .B(i_data_imm[7]), .S(n14), .Q(o_data_alub[7])
         );
  IMUX22 U18 ( .A(n57), .B(n56), .S(n14), .Q(o_data_alub[27]) );
  CLKIN6 U19 ( .A(n16), .Q(n15) );
  IMUX22 U20 ( .A(n37), .B(n36), .S(n14), .Q(o_data_alub[15]) );
  MUX22 U21 ( .A(i_data_fb[26]), .B(i_data_imm[26]), .S(n1), .Q(
        o_data_alub[26]) );
  IMUX21 U22 ( .A(n49), .B(n48), .S(n14), .Q(o_data_alub[22]) );
  IMUX22 U23 ( .A(n31), .B(n30), .S(n14), .Q(o_data_alub[12]) );
  NAND22 U24 ( .A(i_data_fb[2]), .B(n2), .Q(n20) );
  INV2 U25 ( .A(n15), .Q(n4) );
  CLKIN2 U26 ( .A(n1), .Q(n2) );
  IMUX22 U27 ( .A(n22), .B(n21), .S(n15), .Q(o_data_alub[3]) );
  IMUX22 U28 ( .A(n35), .B(n34), .S(n1), .Q(o_data_alub[14]) );
  MUX22 U29 ( .A(i_data_fb[9]), .B(i_data_imm[9]), .S(n1), .Q(o_data_alub[9])
         );
  INV3 U30 ( .A(n27), .Q(o_data_alub[10]) );
  IMUX21 U31 ( .A(n43), .B(n42), .S(n14), .Q(o_data_alub[18]) );
  NAND21 U32 ( .A(n15), .B(i_data_imm[2]), .Q(n19) );
  NAND22 U33 ( .A(n5), .B(n6), .Q(o_data_alub[0]) );
  CLKIN15 U34 ( .A(i_con_imm), .Q(n16) );
  IMUX22 U35 ( .A(n29), .B(n28), .S(n1), .Q(o_data_alub[11]) );
  AOI221 U36 ( .A(i_data_fb[10]), .B(n16), .C(i_data_imm[10]), .D(n3), .Q(n27)
         );
  NAND22 U37 ( .A(i_data_fb[0]), .B(n4), .Q(n5) );
  CLKIN2 U38 ( .A(i_data_imm[6]), .Q(n12) );
  INV3 U39 ( .A(i_data_imm[24]), .Q(n52) );
  INV3 U40 ( .A(i_data_imm[19]), .Q(n44) );
  CLKIN2 U41 ( .A(i_data_imm[8]), .Q(n13) );
  MUX21 U42 ( .A(i_data_fb[29]), .B(i_data_imm[29]), .S(n1), .Q(
        o_data_alub[29]) );
  MUX21 U43 ( .A(i_data_fb[30]), .B(i_data_imm[30]), .S(n1), .Q(
        o_data_alub[30]) );
  MUX21 U44 ( .A(i_data_fb[28]), .B(i_data_imm[28]), .S(n14), .Q(
        o_data_alub[28]) );
  MUX21 U45 ( .A(i_data_fb[21]), .B(i_data_imm[21]), .S(i_con_imm), .Q(
        o_data_alub[21]) );
  INV3 U46 ( .A(i_data_fb[25]), .Q(n55) );
  INV3 U47 ( .A(i_data_imm[25]), .Q(n54) );
  INV3 U48 ( .A(i_data_fb[24]), .Q(n53) );
  INV3 U49 ( .A(i_data_fb[27]), .Q(n57) );
  INV3 U50 ( .A(i_data_imm[27]), .Q(n56) );
  INV3 U51 ( .A(n25), .Q(n11) );
  INV3 U52 ( .A(i_data_fb[23]), .Q(n51) );
  INV3 U53 ( .A(i_data_imm[23]), .Q(n50) );
  INV3 U54 ( .A(i_data_fb[18]), .Q(n43) );
  INV3 U55 ( .A(i_data_imm[18]), .Q(n42) );
  INV3 U56 ( .A(i_data_fb[17]), .Q(n41) );
  INV3 U57 ( .A(i_data_imm[17]), .Q(n40) );
  INV3 U58 ( .A(i_data_fb[13]), .Q(n33) );
  INV3 U59 ( .A(i_data_fb[15]), .Q(n37) );
  INV3 U60 ( .A(i_data_imm[15]), .Q(n36) );
  INV3 U61 ( .A(i_data_fb[19]), .Q(n45) );
  INV3 U62 ( .A(i_data_fb[14]), .Q(n35) );
  INV3 U63 ( .A(i_data_fb[22]), .Q(n49) );
  INV3 U64 ( .A(i_data_imm[22]), .Q(n48) );
  INV3 U65 ( .A(i_data_fb[11]), .Q(n29) );
  INV3 U66 ( .A(i_data_fb[3]), .Q(n22) );
  INV3 U67 ( .A(i_data_fb[4]), .Q(n24) );
  INV3 U68 ( .A(i_data_fb[16]), .Q(n39) );
  INV3 U69 ( .A(i_data_imm[16]), .Q(n38) );
  INV3 U70 ( .A(i_data_fb[1]), .Q(n18) );
  INV3 U71 ( .A(i_data_fb[8]), .Q(n26) );
  INV3 U72 ( .A(i_data_fb[12]), .Q(n31) );
  INV3 U73 ( .A(i_data_imm[12]), .Q(n30) );
  IMUX22 U74 ( .A(n18), .B(n17), .S(n1), .Q(o_data_alub[1]) );
  IMUX22 U75 ( .A(n45), .B(n44), .S(n1), .Q(o_data_alub[19]) );
  INV2 U76 ( .A(i_data_imm[5]), .Q(n25) );
  IMUX22 U77 ( .A(n26), .B(n13), .S(n1), .Q(o_data_alub[8]) );
  NAND22 U78 ( .A(n1), .B(i_data_imm[20]), .Q(n46) );
  NAND22 U79 ( .A(n47), .B(n46), .Q(o_data_alub[20]) );
  IMUX22 U80 ( .A(i_data_fb[6]), .B(n9), .S(n14), .Q(n8) );
  IMUX22 U81 ( .A(i_data_fb[5]), .B(n11), .S(n1), .Q(n10) );
  CLKIN2 U82 ( .A(i_data_imm[1]), .Q(n17) );
  IMUX21 U83 ( .A(n51), .B(n50), .S(n1), .Q(o_data_alub[23]) );
  IMUX21 U84 ( .A(n39), .B(n38), .S(n14), .Q(o_data_alub[16]) );
  IMUX21 U85 ( .A(n55), .B(n54), .S(n15), .Q(o_data_alub[25]) );
  IMUX21 U86 ( .A(n53), .B(n52), .S(n1), .Q(o_data_alub[24]) );
  IMUX22 U87 ( .A(n41), .B(n40), .S(n14), .Q(o_data_alub[17]) );
  IMUX22 U88 ( .A(n33), .B(n32), .S(n14), .Q(o_data_alub[13]) );
endmodule


module E_rdmux ( i_data_rtE, i_data_rdE, i_con_regdst, i_con_aluPC4, 
        o_data_writeE );
  input [4:0] i_data_rtE;
  input [4:0] i_data_rdE;
  output [4:0] o_data_writeE;
  input i_con_regdst, i_con_aluPC4;
  wire   n8, n9, n10, n11, n12, n1, n2, n3, n4, n5, n6, n7;

  OAI2112 U6 ( .A(n1), .B(n4), .C(n7), .D(n10), .Q(o_data_writeE[2]) );
  OAI2112 U8 ( .A(n1), .B(n5), .C(n7), .D(n11), .Q(o_data_writeE[1]) );
  BUF6 U2 ( .A(i_con_regdst), .Q(n1) );
  OAI2111 U3 ( .A(n1), .B(n6), .C(n7), .D(n12), .Q(o_data_writeE[0]) );
  OAI2111 U4 ( .A(n1), .B(n2), .C(n7), .D(n8), .Q(o_data_writeE[4]) );
  INV3 U5 ( .A(i_data_rtE[4]), .Q(n2) );
  NAND22 U7 ( .A(i_data_rdE[4]), .B(n1), .Q(n8) );
  INV3 U9 ( .A(i_data_rtE[2]), .Q(n4) );
  NAND22 U10 ( .A(i_data_rdE[2]), .B(n1), .Q(n10) );
  OAI2111 U11 ( .A(n1), .B(n3), .C(n7), .D(n9), .Q(o_data_writeE[3]) );
  INV3 U12 ( .A(i_data_rtE[3]), .Q(n3) );
  NAND22 U13 ( .A(i_data_rdE[3]), .B(n1), .Q(n9) );
  INV3 U14 ( .A(i_data_rtE[1]), .Q(n5) );
  NAND22 U15 ( .A(i_data_rdE[1]), .B(n1), .Q(n11) );
  INV3 U16 ( .A(i_data_rtE[0]), .Q(n6) );
  NAND22 U17 ( .A(i_data_rdE[0]), .B(n1), .Q(n12) );
  INV3 U18 ( .A(i_con_aluPC4), .Q(n7) );
endmodule


module D_compare_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48;

  INV3 U1 ( .A(NE), .Q(EQ) );
  INV3 U2 ( .A(n27), .Q(n2) );
  INV3 U3 ( .A(A[1]), .Q(n4) );
  INV3 U4 ( .A(B[0]), .Q(n3) );
  NAND20 U5 ( .A(n5), .B(n6), .Q(NE) );
  NOR40 U6 ( .A(n7), .B(n8), .C(n9), .D(n10), .Q(n6) );
  NAND40 U7 ( .A(n11), .B(n12), .C(n13), .D(n14), .Q(n10) );
  XNR20 U8 ( .A(B[11]), .B(A[11]), .Q(n14) );
  XNR20 U9 ( .A(B[12]), .B(A[12]), .Q(n13) );
  XNR20 U10 ( .A(B[13]), .B(A[13]), .Q(n12) );
  XNR20 U11 ( .A(B[14]), .B(A[14]), .Q(n11) );
  NAND40 U12 ( .A(n15), .B(n16), .C(n17), .D(n18), .Q(n9) );
  XNR20 U13 ( .A(B[7]), .B(A[7]), .Q(n18) );
  XNR20 U14 ( .A(B[8]), .B(A[8]), .Q(n17) );
  XNR20 U15 ( .A(B[9]), .B(A[9]), .Q(n16) );
  XNR20 U16 ( .A(B[10]), .B(A[10]), .Q(n15) );
  NAND40 U17 ( .A(n19), .B(n20), .C(n21), .D(n22), .Q(n8) );
  XNR20 U18 ( .A(B[3]), .B(A[3]), .Q(n22) );
  XNR20 U19 ( .A(B[4]), .B(A[4]), .Q(n21) );
  XNR20 U20 ( .A(B[5]), .B(A[5]), .Q(n20) );
  XNR20 U21 ( .A(B[6]), .B(A[6]), .Q(n19) );
  NAND40 U22 ( .A(n23), .B(n24), .C(n2), .D(n25), .Q(n7) );
  OAI220 U23 ( .A(n26), .B(n4), .C(B[1]), .D(n26), .Q(n25) );
  NOR20 U24 ( .A(n3), .B(A[0]), .Q(n26) );
  AOI220 U25 ( .A(n4), .B(n28), .C(n28), .D(B[1]), .Q(n27) );
  NAND20 U26 ( .A(A[0]), .B(n3), .Q(n28) );
  XNR20 U27 ( .A(B[31]), .B(A[31]), .Q(n24) );
  XNR20 U28 ( .A(B[2]), .B(A[2]), .Q(n23) );
  NOR40 U29 ( .A(n29), .B(n30), .C(n31), .D(n32), .Q(n5) );
  NAND40 U30 ( .A(n33), .B(n34), .C(n35), .D(n36), .Q(n32) );
  XNR20 U31 ( .A(B[27]), .B(A[27]), .Q(n36) );
  XNR20 U32 ( .A(B[28]), .B(A[28]), .Q(n35) );
  XNR20 U33 ( .A(B[29]), .B(A[29]), .Q(n34) );
  XNR20 U34 ( .A(B[30]), .B(A[30]), .Q(n33) );
  NAND40 U35 ( .A(n37), .B(n38), .C(n39), .D(n40), .Q(n31) );
  XNR20 U36 ( .A(B[23]), .B(A[23]), .Q(n40) );
  XNR20 U37 ( .A(B[24]), .B(A[24]), .Q(n39) );
  XNR20 U38 ( .A(B[25]), .B(A[25]), .Q(n38) );
  XNR20 U39 ( .A(B[26]), .B(A[26]), .Q(n37) );
  NAND40 U40 ( .A(n41), .B(n42), .C(n43), .D(n44), .Q(n30) );
  XNR20 U41 ( .A(B[19]), .B(A[19]), .Q(n44) );
  XNR20 U42 ( .A(B[20]), .B(A[20]), .Q(n43) );
  XNR20 U43 ( .A(B[21]), .B(A[21]), .Q(n42) );
  XNR20 U44 ( .A(B[22]), .B(A[22]), .Q(n41) );
  NAND40 U45 ( .A(n45), .B(n46), .C(n47), .D(n48), .Q(n29) );
  XNR20 U46 ( .A(B[15]), .B(A[15]), .Q(n48) );
  XNR20 U47 ( .A(B[16]), .B(A[16]), .Q(n47) );
  XNR20 U48 ( .A(B[17]), .B(A[17]), .Q(n46) );
  XNR20 U49 ( .A(B[18]), .B(A[18]), .Q(n45) );
endmodule


module D_compare ( o_con_ifbranch, i_data_rs, i_data_rt, i_con_bop );
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [2:0] i_con_bop;
  output o_con_ifbranch;
  wire   N34, N35, n5, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n1, n2, n3, n4;

  OAI222 U3 ( .A(n10), .B(n2), .C(i_con_bop[2]), .D(n11), .Q(o_con_ifbranch)
         );
  OAI222 U9 ( .A(n4), .B(n1), .C(i_con_bop[0]), .D(n14), .Q(n16) );
  OAI212 U10 ( .A(n17), .B(n18), .C(n1), .Q(n14) );
  D_compare_DW01_cmp6_0 r49 ( .A(i_data_rs), .B(i_data_rt), .TC(n5), .EQ(N34), 
        .NE(N35) );
  NOR21 U2 ( .A(n13), .B(n3), .Q(n12) );
  AOI221 U4 ( .A(i_con_bop[0]), .B(n14), .C(N35), .D(n4), .Q(n13) );
  INV3 U5 ( .A(i_con_bop[2]), .Q(n2) );
  AOI221 U6 ( .A(n15), .B(i_con_bop[1]), .C(n16), .D(n3), .Q(n10) );
  AOI311 U7 ( .A(N34), .B(n3), .C(i_con_bop[0]), .D(n12), .Q(n11) );
  INV3 U8 ( .A(i_con_bop[1]), .Q(n3) );
  NOR21 U11 ( .A(i_data_rs[31]), .B(i_con_bop[0]), .Q(n15) );
  INV3 U12 ( .A(i_con_bop[0]), .Q(n4) );
  NOR40 U13 ( .A(i_data_rs[15]), .B(i_data_rs[14]), .C(i_data_rs[13]), .D(
        i_data_rs[12]), .Q(n20) );
  NOR40 U14 ( .A(i_data_rs[26]), .B(i_data_rs[25]), .C(i_data_rs[24]), .D(
        i_data_rs[23]), .Q(n23) );
  NOR40 U15 ( .A(i_data_rs[9]), .B(i_data_rs[8]), .C(i_data_rs[7]), .D(
        i_data_rs[6]), .Q(n26) );
  NOR40 U16 ( .A(i_data_rs[2]), .B(i_data_rs[29]), .C(i_data_rs[28]), .D(
        i_data_rs[27]), .Q(n24) );
  NOR40 U17 ( .A(i_data_rs[22]), .B(i_data_rs[21]), .C(i_data_rs[20]), .D(
        i_data_rs[1]), .Q(n22) );
  NOR40 U18 ( .A(i_data_rs[5]), .B(i_data_rs[4]), .C(i_data_rs[3]), .D(
        i_data_rs[30]), .Q(n25) );
  NOR40 U19 ( .A(i_data_rs[19]), .B(i_data_rs[18]), .C(i_data_rs[17]), .D(
        i_data_rs[16]), .Q(n21) );
  NAND41 U20 ( .A(n19), .B(n20), .C(n21), .D(n22), .Q(n18) );
  NAND41 U21 ( .A(n23), .B(n24), .C(n25), .D(n26), .Q(n17) );
  NOR31 U22 ( .A(i_data_rs[0]), .B(i_data_rs[11]), .C(i_data_rs[10]), .Q(n19)
         );
  INV3 U23 ( .A(i_data_rs[31]), .Q(n1) );
  LOGIC0 U24 ( .Q(n5) );
endmodule


module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Ealuop, i_con_Ealusrc, 
        i_con_Eregdst, i_con_Mmemread, i_con_Mmemwrite, i_con_Wloadmux, 
        i_con_Walupc8, i_con_Wmemtoreg, i_con_Wregwrite, i_con_Efamux, 
        i_con_Efbmux, i_con_bop, o_data_pc4, o_data_alures, o_data_rt, 
        o_addr_regdst, o_con_Mmemread, o_con_Mmemwrite, o_con_Wloadmux, 
        o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_addr_Erd, 
        o_addr_Mrt, o_FaluresE, o_con_ifbranch );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [5:0] i_con_Ealuop;
  input [1:0] i_con_Wloadmux;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [2:0] i_con_bop;
  output [31:0] o_data_pc4;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [1:0] o_con_Wloadmux;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  output [31:0] o_FaluresE;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Walupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Walupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch;
  wire   n119, n1, n3, n33, n34;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;

  DFC3 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[0]) );
  DFC3 pipe_alures_reg_30_ ( .D(o_FaluresE[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[30]) );
  DFC3 pipe_alures_reg_4_ ( .D(o_FaluresE[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[4]) );
  DFC3 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC3 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC3 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC3 pipe_rt_reg_28_ ( .D(compare_i_data_rt[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[28]) );
  DFC3 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  DFC3 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC3 pipe_rt_reg_25_ ( .D(compare_i_data_rt[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[25]) );
  DFC3 pipe_rt_reg_24_ ( .D(compare_i_data_rt[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[24]) );
  DFC3 pipe_rt_reg_23_ ( .D(compare_i_data_rt[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[23]) );
  DFC3 pipe_rt_reg_22_ ( .D(compare_i_data_rt[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[22]) );
  DFC3 pipe_rt_reg_21_ ( .D(compare_i_data_rt[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[21]) );
  DFC3 pipe_rt_reg_20_ ( .D(compare_i_data_rt[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[20]) );
  DFC3 pipe_rt_reg_19_ ( .D(compare_i_data_rt[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[19]) );
  DFC3 pipe_rt_reg_18_ ( .D(compare_i_data_rt[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[18]) );
  DFC3 pipe_rt_reg_17_ ( .D(compare_i_data_rt[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[17]) );
  DFC3 pipe_rt_reg_16_ ( .D(compare_i_data_rt[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[16]) );
  DFC3 pipe_rt_reg_15_ ( .D(compare_i_data_rt[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[15]) );
  DFC3 pipe_rt_reg_14_ ( .D(compare_i_data_rt[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[14]) );
  DFC3 pipe_rt_reg_13_ ( .D(compare_i_data_rt[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[13]) );
  DFC3 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC3 pipe_rt_reg_11_ ( .D(compare_i_data_rt[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[11]) );
  DFC3 pipe_rt_reg_10_ ( .D(compare_i_data_rt[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[10]) );
  DFC3 pipe_rt_reg_9_ ( .D(compare_i_data_rt[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[9]) );
  DFC3 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC3 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC3 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC3 pipe_rt_reg_5_ ( .D(compare_i_data_rt[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[5]) );
  DFC3 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(compare_i_data_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[2]) );
  DFC3 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC3 pipe_rt_reg_0_ ( .D(compare_i_data_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[0]) );
  DFC3 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC3 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC3 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC3 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC3 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC3 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wloadmux_reg_1_ ( .D(i_con_Wloadmux[1]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[1]) );
  DFC3 pipe_con_Wloadmux_reg_0_ ( .D(i_con_Wloadmux[0]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[0]) );
  DFC3 pipe_con_Walupc8_reg ( .D(i_con_Walupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Walupc8) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  E_alu u_alu ( .o_data_AluRes(o_FaluresE), .i_data_A(compare_i_data_rs), 
        .i_data_B({alu_i_data_B[31:4], n33, alu_i_data_B[2], n34, 
        alu_i_data_B[0]}), .i_con_AluCtrl(alu_i_con_AluCtrl), .i_data_shamt({
        i_data_immext[10], n1, i_data_immext[8:6]}) );
  E_alu_control u_alu_control ( .o_con_AluCtrl(alu_i_con_AluCtrl), 
        .i_con_AluOp(i_con_Ealuop), .i_con_FuncCode(i_data_immext[5:0]) );
  E_famux5 u_famux5 ( .i_data_rs(i_data_rs), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fa(i_con_Efamux), .o_data_alusra(
        compare_i_data_rs) );
  E_fbmux5 u_fbmux ( .i_data_rt(i_data_rt), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fb(i_con_Efbmux), .o_data_alusrb(
        compare_i_data_rt) );
  E_alubmux u_alubmux ( .i_data_fb(compare_i_data_rt), .i_data_imm({
        i_data_immext[31:10], n1, i_data_immext[8:0]}), .i_con_imm(
        i_con_Ealusrc), .o_data_alub(alu_i_data_B) );
  E_rdmux u_rdmux ( .i_data_rtE(i_addr_rt), .i_data_rdE(i_addr_rd), 
        .i_con_regdst(i_con_Eregdst), .i_con_aluPC4(i_con_Walupc8), 
        .o_data_writeE({o_addr_Erd[4:1], n119}) );
  D_compare u_compare ( .o_con_ifbranch(o_con_ifbranch), .i_data_rs(
        compare_i_data_rs), .i_data_rt(compare_i_data_rt), .i_con_bop(
        i_con_bop) );
  DFC1 pipe_alures_reg_28_ ( .D(o_FaluresE[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[28]) );
  DFC1 pipe_alures_reg_1_ ( .D(o_FaluresE[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[1]) );
  DFC1 pipe_alures_reg_31_ ( .D(o_FaluresE[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[31]) );
  DFC1 pipe_alures_reg_27_ ( .D(o_FaluresE[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[27]) );
  DFC1 pipe_alures_reg_26_ ( .D(o_FaluresE[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[26]) );
  DFC1 pipe_alures_reg_25_ ( .D(o_FaluresE[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[25]) );
  DFC1 pipe_alures_reg_24_ ( .D(o_FaluresE[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[24]) );
  DFC1 pipe_alures_reg_23_ ( .D(o_FaluresE[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[23]) );
  DFC1 pipe_alures_reg_22_ ( .D(o_FaluresE[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[22]) );
  DFC1 pipe_alures_reg_21_ ( .D(o_FaluresE[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[21]) );
  DFC1 pipe_alures_reg_20_ ( .D(o_FaluresE[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[20]) );
  DFC1 pipe_alures_reg_19_ ( .D(o_FaluresE[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[19]) );
  DFC1 pipe_alures_reg_18_ ( .D(o_FaluresE[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[18]) );
  DFC1 pipe_alures_reg_17_ ( .D(o_FaluresE[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[17]) );
  DFC1 pipe_alures_reg_16_ ( .D(o_FaluresE[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[16]) );
  DFC1 pipe_alures_reg_15_ ( .D(o_FaluresE[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[15]) );
  DFC1 pipe_alures_reg_14_ ( .D(o_FaluresE[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[14]) );
  DFC1 pipe_alures_reg_13_ ( .D(o_FaluresE[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[13]) );
  DFC1 pipe_alures_reg_12_ ( .D(o_FaluresE[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[12]) );
  DFC1 pipe_alures_reg_11_ ( .D(o_FaluresE[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[11]) );
  DFC1 pipe_alures_reg_10_ ( .D(o_FaluresE[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[10]) );
  DFC1 pipe_alures_reg_9_ ( .D(o_FaluresE[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[9]) );
  DFC1 pipe_alures_reg_8_ ( .D(o_FaluresE[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[8]) );
  DFC1 pipe_alures_reg_7_ ( .D(o_FaluresE[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[7]) );
  DFC1 pipe_alures_reg_6_ ( .D(o_FaluresE[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[6]) );
  DFC1 pipe_alures_reg_5_ ( .D(o_FaluresE[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[5]) );
  DFC1 pipe_alures_reg_3_ ( .D(o_FaluresE[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[3]) );
  DFC1 pipe_alures_reg_2_ ( .D(o_FaluresE[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[2]) );
  DFC1 pipe_alures_reg_29_ ( .D(o_FaluresE[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[29]) );
  DFC1 pipe_alures_reg_0_ ( .D(o_FaluresE[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_alures[0]) );
  BUF6 U3 ( .A(i_data_immext[9]), .Q(n1) );
  INV3 U4 ( .A(n3), .Q(o_addr_Erd[0]) );
  INV3 U5 ( .A(n119), .Q(n3) );
  CLKBU15 U6 ( .A(alu_i_data_B[1]), .Q(n34) );
  CLKBU15 U7 ( .A(alu_i_data_B[3]), .Q(n33) );
endmodule


module mem_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   A_1_, A_0_, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103;
  assign SUM[1] = A_1_;
  assign A_1_ = A[1];
  assign SUM[0] = A_0_;
  assign A_0_ = A[0];

  NOR21 U2 ( .A(n67), .B(n65), .Q(n66) );
  NAND22 U3 ( .A(n50), .B(A[21]), .Q(n51) );
  NAND22 U4 ( .A(n36), .B(A[25]), .Q(n37) );
  NAND22 U5 ( .A(n16), .B(n17), .Q(n18) );
  NOR21 U6 ( .A(n67), .B(n63), .Q(n62) );
  INV3 U7 ( .A(n64), .Q(n63) );
  NOR21 U8 ( .A(n65), .B(n58), .Q(n64) );
  INV3 U9 ( .A(n67), .Q(n23) );
  NAND22 U10 ( .A(n68), .B(n69), .Q(n67) );
  NOR21 U11 ( .A(n71), .B(n72), .Q(n69) );
  NOR31 U12 ( .A(n77), .B(n78), .C(n79), .Q(n68) );
  INV3 U13 ( .A(n97), .Q(n3) );
  NAND22 U14 ( .A(n98), .B(n99), .Q(n97) );
  NOR21 U15 ( .A(SUM[2]), .B(n103), .Q(n98) );
  INV3 U16 ( .A(n22), .Q(n17) );
  NAND22 U17 ( .A(n23), .B(n24), .Q(n22) );
  NOR21 U18 ( .A(n25), .B(n26), .Q(n24) );
  NAND22 U19 ( .A(n27), .B(n28), .Q(n25) );
  NOR21 U20 ( .A(n8), .B(n10), .Q(n6) );
  XNR21 U21 ( .A(n50), .B(n44), .Q(SUM[21]) );
  XNR21 U22 ( .A(n36), .B(n31), .Q(SUM[25]) );
  XNR21 U23 ( .A(n62), .B(n59), .Q(SUM[18]) );
  XNR21 U24 ( .A(n66), .B(n58), .Q(SUM[17]) );
  XNR21 U25 ( .A(n83), .B(n76), .Q(SUM[13]) );
  XNR21 U26 ( .A(n94), .B(n92), .Q(SUM[10]) );
  XOR21 U27 ( .A(n2), .B(n1), .Q(SUM[9]) );
  NAND22 U28 ( .A(A[8]), .B(n3), .Q(n2) );
  XOR21 U29 ( .A(n84), .B(n75), .Q(SUM[14]) );
  NAND22 U30 ( .A(n83), .B(A[13]), .Q(n84) );
  XNR21 U31 ( .A(A[22]), .B(n51), .Q(SUM[22]) );
  XNR21 U32 ( .A(A[26]), .B(n37), .Q(SUM[26]) );
  NAND22 U33 ( .A(n73), .B(A[2]), .Q(n72) );
  NOR21 U34 ( .A(n75), .B(n76), .Q(n73) );
  NOR21 U35 ( .A(n30), .B(n31), .Q(n27) );
  XNR21 U36 ( .A(n6), .B(n7), .Q(SUM[6]) );
  INV3 U37 ( .A(n95), .Q(n94) );
  NAND22 U38 ( .A(n96), .B(n3), .Q(n95) );
  NOR21 U39 ( .A(n1), .B(n4), .Q(n96) );
  XNR21 U40 ( .A(n9), .B(n8), .Q(SUM[5]) );
  NOR21 U41 ( .A(n76), .B(n75), .Q(n82) );
  NOR21 U42 ( .A(n44), .B(n45), .Q(n49) );
  NOR21 U43 ( .A(n31), .B(n30), .Q(n35) );
  NAND22 U44 ( .A(n89), .B(n90), .Q(n77) );
  NOR21 U45 ( .A(n1), .B(n92), .Q(n89) );
  INV3 U46 ( .A(n91), .Q(n90) );
  NAND22 U47 ( .A(A[11]), .B(A[8]), .Q(n91) );
  NOR21 U48 ( .A(n67), .B(n52), .Q(n50) );
  NAND22 U49 ( .A(A[20]), .B(n42), .Q(n52) );
  NOR21 U50 ( .A(n67), .B(n38), .Q(n36) );
  NAND22 U51 ( .A(A[24]), .B(n39), .Q(n38) );
  XOR21 U52 ( .A(n60), .B(A[19]), .Q(SUM[19]) );
  NOR21 U53 ( .A(n59), .B(n61), .Q(n60) );
  XOR21 U54 ( .A(n46), .B(A[23]), .Q(SUM[23]) );
  NOR21 U55 ( .A(n47), .B(n48), .Q(n46) );
  INV3 U56 ( .A(n49), .Q(n48) );
  XOR21 U57 ( .A(n32), .B(A[27]), .Q(SUM[27]) );
  NOR21 U58 ( .A(n33), .B(n34), .Q(n32) );
  INV3 U59 ( .A(n35), .Q(n34) );
  INV3 U60 ( .A(A[9]), .Q(n1) );
  NAND22 U61 ( .A(n41), .B(n42), .Q(n26) );
  NOR31 U62 ( .A(n45), .B(n43), .C(n44), .Q(n41) );
  NAND22 U63 ( .A(A[23]), .B(A[20]), .Q(n43) );
  INV3 U64 ( .A(A[21]), .Q(n44) );
  INV3 U65 ( .A(A[13]), .Q(n76) );
  INV3 U66 ( .A(A[25]), .Q(n31) );
  NAND22 U67 ( .A(n100), .B(n101), .Q(n71) );
  NOR21 U68 ( .A(n70), .B(n102), .Q(n100) );
  NOR21 U69 ( .A(n8), .B(n7), .Q(n101) );
  INV3 U70 ( .A(A[7]), .Q(n102) );
  INV3 U71 ( .A(A[5]), .Q(n8) );
  INV3 U72 ( .A(A[14]), .Q(n75) );
  INV3 U73 ( .A(A[22]), .Q(n45) );
  INV3 U74 ( .A(A[10]), .Q(n92) );
  INV3 U75 ( .A(A[18]), .Q(n59) );
  INV3 U76 ( .A(A[17]), .Q(n58) );
  XOR21 U77 ( .A(n17), .B(A[28]), .Q(SUM[28]) );
  XOR21 U78 ( .A(n54), .B(A[20]), .Q(SUM[20]) );
  NOR21 U79 ( .A(n67), .B(n53), .Q(n54) );
  XOR21 U80 ( .A(n40), .B(A[24]), .Q(SUM[24]) );
  NOR21 U81 ( .A(n67), .B(n26), .Q(n40) );
  XOR21 U82 ( .A(n23), .B(A[16]), .Q(SUM[16]) );
  XOR21 U83 ( .A(n93), .B(A[11]), .Q(SUM[11]) );
  NOR21 U84 ( .A(n92), .B(n95), .Q(n93) );
  XOR21 U85 ( .A(n80), .B(A[15]), .Q(SUM[15]) );
  NOR21 U86 ( .A(n85), .B(n81), .Q(n80) );
  INV3 U87 ( .A(n82), .Q(n81) );
  XOR21 U88 ( .A(n13), .B(A[31]), .Q(SUM[31]) );
  NOR21 U89 ( .A(n14), .B(n15), .Q(n13) );
  INV3 U90 ( .A(A[30]), .Q(n14) );
  NAND22 U91 ( .A(n16), .B(n17), .Q(n15) );
  XOR21 U92 ( .A(n20), .B(n21), .Q(SUM[29]) );
  INV3 U93 ( .A(A[29]), .Q(n20) );
  NAND22 U94 ( .A(A[28]), .B(n17), .Q(n21) );
  XNR21 U95 ( .A(A[30]), .B(n18), .Q(SUM[30]) );
  INV3 U96 ( .A(A[6]), .Q(n7) );
  NAND22 U97 ( .A(A[15]), .B(A[3]), .Q(n79) );
  INV3 U98 ( .A(A[26]), .Q(n30) );
  XOR21 U99 ( .A(n78), .B(n87), .Q(SUM[12]) );
  NAND22 U100 ( .A(n88), .B(n3), .Q(n87) );
  INV3 U101 ( .A(n77), .Q(n88) );
  XOR21 U102 ( .A(n102), .B(n5), .Q(SUM[7]) );
  NAND22 U103 ( .A(n6), .B(A[6]), .Q(n5) );
  INV3 U104 ( .A(n85), .Q(n83) );
  NAND22 U105 ( .A(n86), .B(n3), .Q(n85) );
  NOR21 U106 ( .A(n77), .B(n78), .Q(n86) );
  INV3 U107 ( .A(n12), .Q(n11) );
  NAND22 U108 ( .A(A[3]), .B(A[2]), .Q(n12) );
  INV3 U109 ( .A(A[2]), .Q(SUM[2]) );
  INV3 U110 ( .A(n10), .Q(n9) );
  NAND22 U111 ( .A(A[4]), .B(n11), .Q(n10) );
  INV3 U112 ( .A(A[3]), .Q(n103) );
  INV3 U113 ( .A(A[4]), .Q(n70) );
  INV3 U114 ( .A(A[12]), .Q(n78) );
  NAND22 U115 ( .A(n55), .B(n56), .Q(n53) );
  NOR21 U116 ( .A(n58), .B(n59), .Q(n55) );
  INV3 U117 ( .A(n57), .Q(n56) );
  NAND22 U118 ( .A(A[19]), .B(A[16]), .Q(n57) );
  INV3 U119 ( .A(n29), .Q(n28) );
  NAND22 U120 ( .A(A[27]), .B(A[24]), .Q(n29) );
  XOR21 U121 ( .A(n3), .B(A[8]), .Q(SUM[8]) );
  XOR21 U122 ( .A(n11), .B(A[4]), .Q(SUM[4]) );
  NOR21 U123 ( .A(n19), .B(n20), .Q(n16) );
  INV3 U124 ( .A(A[16]), .Q(n65) );
  INV3 U125 ( .A(A[28]), .Q(n19) );
  INV3 U126 ( .A(A[8]), .Q(n4) );
  XOR21 U127 ( .A(A[3]), .B(A[2]), .Q(SUM[3]) );
  CLKIN3 U128 ( .A(n36), .Q(n33) );
  CLKIN3 U129 ( .A(n26), .Q(n39) );
  CLKIN3 U130 ( .A(n50), .Q(n47) );
  CLKIN3 U131 ( .A(n53), .Q(n42) );
  CLKIN3 U132 ( .A(n62), .Q(n61) );
  CLKIN3 U133 ( .A(n71), .Q(n99) );
endmodule


module mem ( i_clk, i_nrst, i_data_pc4, i_data_alures, i_data_memout, 
        i_addr_regdst, i_con_Wloadmux, i_con_Walupc8, i_con_Wmemtoreg, 
        i_con_Wregwrite, i_con_FWmemread, i_addr_Mrt, o_data_pc8, 
        o_data_alures, o_data_memout, o_addr_regdst, o_con_Wloadmux, 
        o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread, 
        o_addr_Wrt );
  input [31:0] i_data_pc4;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [4:0] i_addr_regdst;
  input [1:0] i_con_Wloadmux;
  input [4:0] i_addr_Mrt;
  output [31:0] o_data_pc8;
  output [31:0] o_data_alures;
  output [31:0] o_data_memout;
  output [4:0] o_addr_regdst;
  output [1:0] o_con_Wloadmux;
  output [4:0] o_addr_Wrt;
  input i_clk, i_nrst, i_con_Walupc8, i_con_Wmemtoreg, i_con_Wregwrite,
         i_con_FWmemread;
  output o_con_Walupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread;
  wire   n_Logic1_, n_Logic0_;
  wire   [31:0] pc8;

  DFC3 pipe_rt_reg_4_ ( .D(i_addr_Mrt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(i_addr_Mrt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(i_addr_Mrt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[2]) );
  DFC3 pipe_rt_reg_1_ ( .D(i_addr_Mrt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[1]) );
  DFC3 pipe_rt_reg_0_ ( .D(i_addr_Mrt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[0]) );
  DFC3 pipe_data_pc8_reg_31_ ( .D(pc8[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[31]) );
  DFC3 pipe_data_pc8_reg_30_ ( .D(pc8[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[30]) );
  DFC3 pipe_data_pc8_reg_29_ ( .D(pc8[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[29]) );
  DFC3 pipe_data_pc8_reg_28_ ( .D(pc8[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[28]) );
  DFC3 pipe_data_pc8_reg_27_ ( .D(pc8[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[27]) );
  DFC3 pipe_data_pc8_reg_26_ ( .D(pc8[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[26]) );
  DFC3 pipe_data_pc8_reg_25_ ( .D(pc8[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[25]) );
  DFC3 pipe_data_pc8_reg_24_ ( .D(pc8[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[24]) );
  DFC3 pipe_data_pc8_reg_23_ ( .D(pc8[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[23]) );
  DFC3 pipe_data_pc8_reg_22_ ( .D(pc8[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[22]) );
  DFC3 pipe_data_pc8_reg_21_ ( .D(pc8[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[21]) );
  DFC3 pipe_data_pc8_reg_20_ ( .D(pc8[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[20]) );
  DFC3 pipe_data_pc8_reg_19_ ( .D(pc8[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[19]) );
  DFC3 pipe_data_pc8_reg_18_ ( .D(pc8[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[18]) );
  DFC3 pipe_data_pc8_reg_17_ ( .D(pc8[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[17]) );
  DFC3 pipe_data_pc8_reg_16_ ( .D(pc8[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[16]) );
  DFC3 pipe_data_pc8_reg_15_ ( .D(pc8[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[15]) );
  DFC3 pipe_data_pc8_reg_14_ ( .D(pc8[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[14]) );
  DFC3 pipe_data_pc8_reg_13_ ( .D(pc8[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[13]) );
  DFC3 pipe_data_pc8_reg_12_ ( .D(pc8[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[12]) );
  DFC3 pipe_data_pc8_reg_11_ ( .D(pc8[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[11]) );
  DFC3 pipe_data_pc8_reg_10_ ( .D(pc8[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[10]) );
  DFC3 pipe_data_pc8_reg_9_ ( .D(pc8[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[9]) );
  DFC3 pipe_data_pc8_reg_8_ ( .D(pc8[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[8]) );
  DFC3 pipe_data_pc8_reg_7_ ( .D(pc8[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[7]) );
  DFC3 pipe_data_pc8_reg_6_ ( .D(pc8[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[6]) );
  DFC3 pipe_data_pc8_reg_5_ ( .D(pc8[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[5]) );
  DFC3 pipe_data_pc8_reg_4_ ( .D(pc8[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[4]) );
  DFC3 pipe_data_pc8_reg_3_ ( .D(pc8[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[3]) );
  DFC3 pipe_data_pc8_reg_2_ ( .D(pc8[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[2]) );
  DFC3 pipe_data_pc8_reg_1_ ( .D(pc8[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[1]) );
  DFC3 pipe_data_pc8_reg_0_ ( .D(pc8[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc8[0]) );
  DFC3 pipe_data_alures_reg_31_ ( .D(i_data_alures[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[31]) );
  DFC3 pipe_data_alures_reg_30_ ( .D(i_data_alures[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[30]) );
  DFC3 pipe_data_alures_reg_29_ ( .D(i_data_alures[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[29]) );
  DFC3 pipe_data_alures_reg_28_ ( .D(i_data_alures[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[28]) );
  DFC3 pipe_data_alures_reg_27_ ( .D(i_data_alures[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[27]) );
  DFC3 pipe_data_alures_reg_26_ ( .D(i_data_alures[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[26]) );
  DFC3 pipe_data_alures_reg_25_ ( .D(i_data_alures[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[25]) );
  DFC3 pipe_data_alures_reg_24_ ( .D(i_data_alures[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[24]) );
  DFC3 pipe_data_alures_reg_23_ ( .D(i_data_alures[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[23]) );
  DFC3 pipe_data_alures_reg_22_ ( .D(i_data_alures[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[22]) );
  DFC3 pipe_data_alures_reg_21_ ( .D(i_data_alures[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[21]) );
  DFC3 pipe_data_alures_reg_20_ ( .D(i_data_alures[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[20]) );
  DFC3 pipe_data_alures_reg_19_ ( .D(i_data_alures[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[19]) );
  DFC3 pipe_data_alures_reg_18_ ( .D(i_data_alures[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[18]) );
  DFC3 pipe_data_alures_reg_17_ ( .D(i_data_alures[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[17]) );
  DFC3 pipe_data_alures_reg_16_ ( .D(i_data_alures[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[16]) );
  DFC3 pipe_data_alures_reg_15_ ( .D(i_data_alures[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[15]) );
  DFC3 pipe_data_alures_reg_14_ ( .D(i_data_alures[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[14]) );
  DFC3 pipe_data_alures_reg_13_ ( .D(i_data_alures[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[13]) );
  DFC3 pipe_data_alures_reg_12_ ( .D(i_data_alures[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[12]) );
  DFC3 pipe_data_alures_reg_11_ ( .D(i_data_alures[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[11]) );
  DFC3 pipe_data_alures_reg_10_ ( .D(i_data_alures[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_alures[10]) );
  DFC3 pipe_data_alures_reg_9_ ( .D(i_data_alures[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC3 pipe_data_alures_reg_8_ ( .D(i_data_alures[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC3 pipe_data_alures_reg_7_ ( .D(i_data_alures[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC3 pipe_data_alures_reg_6_ ( .D(i_data_alures[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC3 pipe_data_alures_reg_5_ ( .D(i_data_alures[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC3 pipe_data_alures_reg_4_ ( .D(i_data_alures[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC3 pipe_data_alures_reg_3_ ( .D(i_data_alures[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC3 pipe_data_alures_reg_2_ ( .D(i_data_alures[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC3 pipe_data_alures_reg_1_ ( .D(i_data_alures[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC3 pipe_data_alures_reg_0_ ( .D(i_data_alures[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC3 pipe_data_memout_reg_31_ ( .D(i_data_memout[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[31]) );
  DFC3 pipe_data_memout_reg_30_ ( .D(i_data_memout[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[30]) );
  DFC3 pipe_data_memout_reg_29_ ( .D(i_data_memout[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[29]) );
  DFC3 pipe_data_memout_reg_28_ ( .D(i_data_memout[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[28]) );
  DFC3 pipe_data_memout_reg_27_ ( .D(i_data_memout[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[27]) );
  DFC3 pipe_data_memout_reg_26_ ( .D(i_data_memout[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[26]) );
  DFC3 pipe_data_memout_reg_25_ ( .D(i_data_memout[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[25]) );
  DFC3 pipe_data_memout_reg_24_ ( .D(i_data_memout[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[24]) );
  DFC3 pipe_data_memout_reg_23_ ( .D(i_data_memout[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[23]) );
  DFC3 pipe_data_memout_reg_22_ ( .D(i_data_memout[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[22]) );
  DFC3 pipe_data_memout_reg_21_ ( .D(i_data_memout[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[21]) );
  DFC3 pipe_data_memout_reg_20_ ( .D(i_data_memout[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[20]) );
  DFC3 pipe_data_memout_reg_19_ ( .D(i_data_memout[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[19]) );
  DFC3 pipe_data_memout_reg_18_ ( .D(i_data_memout[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[18]) );
  DFC3 pipe_data_memout_reg_17_ ( .D(i_data_memout[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[17]) );
  DFC3 pipe_data_memout_reg_16_ ( .D(i_data_memout[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[16]) );
  DFC3 pipe_data_memout_reg_15_ ( .D(i_data_memout[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[15]) );
  DFC3 pipe_data_memout_reg_14_ ( .D(i_data_memout[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[14]) );
  DFC3 pipe_data_memout_reg_13_ ( .D(i_data_memout[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[13]) );
  DFC3 pipe_data_memout_reg_12_ ( .D(i_data_memout[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[12]) );
  DFC3 pipe_data_memout_reg_11_ ( .D(i_data_memout[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[11]) );
  DFC3 pipe_data_memout_reg_10_ ( .D(i_data_memout[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[10]) );
  DFC3 pipe_data_memout_reg_9_ ( .D(i_data_memout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[9]) );
  DFC3 pipe_data_memout_reg_8_ ( .D(i_data_memout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[8]) );
  DFC3 pipe_data_memout_reg_7_ ( .D(i_data_memout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[7]) );
  DFC3 pipe_data_memout_reg_6_ ( .D(i_data_memout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[6]) );
  DFC3 pipe_data_memout_reg_5_ ( .D(i_data_memout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[5]) );
  DFC3 pipe_data_memout_reg_4_ ( .D(i_data_memout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[4]) );
  DFC3 pipe_data_memout_reg_3_ ( .D(i_data_memout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[3]) );
  DFC3 pipe_data_memout_reg_2_ ( .D(i_data_memout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[2]) );
  DFC3 pipe_data_memout_reg_1_ ( .D(i_data_memout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[1]) );
  DFC3 pipe_data_memout_reg_0_ ( .D(i_data_memout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[0]) );
  DFC3 pipe_addr_regdst_reg_4_ ( .D(i_addr_regdst[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[4]) );
  DFC3 pipe_addr_regdst_reg_3_ ( .D(i_addr_regdst[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[3]) );
  DFC3 pipe_addr_regdst_reg_2_ ( .D(i_addr_regdst[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[2]) );
  DFC3 pipe_addr_regdst_reg_1_ ( .D(i_addr_regdst[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[1]) );
  DFC3 pipe_addr_regdst_reg_0_ ( .D(i_addr_regdst[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[0]) );
  DFC3 pipe_con_Wloadmux_reg_1_ ( .D(i_con_Wloadmux[1]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[1]) );
  DFC3 pipe_con_Wloadmux_reg_0_ ( .D(i_con_Wloadmux[0]), .C(i_clk), .RN(i_nrst), .Q(o_con_Wloadmux[0]) );
  DFC3 pipe_con_Walupc8_reg ( .D(i_con_Walupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Walupc8) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_con_FWmemread_reg ( .D(i_con_FWmemread), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_FWmemread) );
  mem_DW01_add_1 add_31 ( .A(i_data_pc4), .B({n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic1_, n_Logic0_, n_Logic0_}), .CI(n_Logic0_), .SUM(pc8) );
  LOGIC0 U3 ( .Q(n_Logic0_) );
  LOGIC1 U4 ( .Q(n_Logic1_) );
endmodule


module W_resmux ( i_data_alures, i_data_pc8, i_con_pc8, o_data_alu );
  input [31:0] i_data_alures;
  input [31:0] i_data_pc8;
  output [31:0] o_data_alu;
  input i_con_pc8;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n1, n2, n3, n4, n5;

  CLKIN3 U1 ( .A(n36), .Q(o_data_alu[8]) );
  CLKIN3 U2 ( .A(n35), .Q(o_data_alu[9]) );
  CLKIN3 U3 ( .A(n37), .Q(o_data_alu[7]) );
  INV3 U4 ( .A(n5), .Q(n1) );
  BUF2 U5 ( .A(n5), .Q(n2) );
  BUF2 U6 ( .A(n5), .Q(n3) );
  BUF2 U7 ( .A(n5), .Q(n4) );
  INV3 U8 ( .A(n66), .Q(o_data_alu[0]) );
  INV3 U9 ( .A(n55), .Q(o_data_alu[1]) );
  INV3 U10 ( .A(n44), .Q(o_data_alu[2]) );
  INV3 U11 ( .A(n41), .Q(o_data_alu[3]) );
  INV3 U12 ( .A(n40), .Q(o_data_alu[4]) );
  INV3 U13 ( .A(n39), .Q(o_data_alu[5]) );
  INV3 U14 ( .A(n38), .Q(o_data_alu[6]) );
  INV3 U15 ( .A(n59), .Q(o_data_alu[16]) );
  INV3 U16 ( .A(n58), .Q(o_data_alu[17]) );
  INV3 U17 ( .A(n57), .Q(o_data_alu[18]) );
  INV3 U18 ( .A(n56), .Q(o_data_alu[19]) );
  INV3 U19 ( .A(n54), .Q(o_data_alu[20]) );
  INV3 U20 ( .A(n53), .Q(o_data_alu[21]) );
  INV3 U21 ( .A(n52), .Q(o_data_alu[22]) );
  INV3 U22 ( .A(n51), .Q(o_data_alu[23]) );
  INV3 U23 ( .A(n50), .Q(o_data_alu[24]) );
  INV3 U24 ( .A(n49), .Q(o_data_alu[25]) );
  INV3 U25 ( .A(n48), .Q(o_data_alu[26]) );
  INV3 U26 ( .A(n47), .Q(o_data_alu[27]) );
  INV3 U27 ( .A(n46), .Q(o_data_alu[28]) );
  INV3 U28 ( .A(n45), .Q(o_data_alu[29]) );
  INV3 U29 ( .A(n43), .Q(o_data_alu[30]) );
  INV3 U30 ( .A(n42), .Q(o_data_alu[31]) );
  AOI221 U31 ( .A(i_data_alures[0]), .B(n4), .C(i_data_pc8[0]), .D(n1), .Q(n66) );
  AOI221 U32 ( .A(i_data_alures[1]), .B(n2), .C(i_data_pc8[1]), .D(n1), .Q(n55) );
  AOI221 U33 ( .A(i_data_alures[2]), .B(n3), .C(i_data_pc8[2]), .D(n1), .Q(n44) );
  AOI221 U34 ( .A(i_data_alures[3]), .B(n4), .C(i_data_pc8[3]), .D(n1), .Q(n41) );
  AOI221 U35 ( .A(i_data_alures[16]), .B(n3), .C(i_data_pc8[16]), .D(i_con_pc8), .Q(n59) );
  AOI221 U36 ( .A(i_data_alures[17]), .B(n2), .C(i_data_pc8[17]), .D(i_con_pc8), .Q(n58) );
  AOI221 U37 ( .A(i_data_alures[18]), .B(n2), .C(i_data_pc8[18]), .D(i_con_pc8), .Q(n57) );
  AOI221 U38 ( .A(i_data_alures[19]), .B(n2), .C(i_data_pc8[19]), .D(i_con_pc8), .Q(n56) );
  AOI221 U39 ( .A(i_data_alures[20]), .B(n2), .C(i_data_pc8[20]), .D(i_con_pc8), .Q(n54) );
  AOI221 U40 ( .A(i_data_alures[21]), .B(n2), .C(i_data_pc8[21]), .D(n1), .Q(
        n53) );
  AOI221 U41 ( .A(i_data_alures[22]), .B(n2), .C(i_data_pc8[22]), .D(n1), .Q(
        n52) );
  AOI221 U42 ( .A(i_data_alures[23]), .B(n2), .C(i_data_pc8[23]), .D(n1), .Q(
        n51) );
  AOI221 U43 ( .A(i_data_alures[24]), .B(n3), .C(i_data_pc8[24]), .D(n1), .Q(
        n50) );
  AOI221 U44 ( .A(i_data_alures[25]), .B(n3), .C(i_data_pc8[25]), .D(n1), .Q(
        n49) );
  AOI221 U45 ( .A(i_data_alures[26]), .B(n3), .C(i_data_pc8[26]), .D(n1), .Q(
        n48) );
  AOI221 U46 ( .A(i_data_alures[27]), .B(n3), .C(i_data_pc8[27]), .D(n1), .Q(
        n47) );
  AOI221 U47 ( .A(i_data_alures[28]), .B(n3), .C(i_data_pc8[28]), .D(n1), .Q(
        n46) );
  AOI221 U48 ( .A(i_data_alures[29]), .B(n3), .C(i_data_pc8[29]), .D(n1), .Q(
        n45) );
  AOI221 U49 ( .A(i_data_alures[30]), .B(n3), .C(i_data_pc8[30]), .D(n1), .Q(
        n43) );
  AOI221 U50 ( .A(i_data_alures[31]), .B(n4), .C(i_data_pc8[31]), .D(n1), .Q(
        n42) );
  AOI221 U51 ( .A(i_data_alures[4]), .B(n4), .C(i_data_pc8[4]), .D(n1), .Q(n40) );
  AOI221 U52 ( .A(i_data_alures[5]), .B(n4), .C(i_data_pc8[5]), .D(n1), .Q(n39) );
  AOI221 U53 ( .A(i_data_alures[6]), .B(n4), .C(i_data_pc8[6]), .D(n1), .Q(n38) );
  AOI221 U54 ( .A(i_data_alures[7]), .B(n4), .C(i_data_pc8[7]), .D(n1), .Q(n37) );
  AOI221 U55 ( .A(i_data_alures[8]), .B(n4), .C(i_data_pc8[8]), .D(n1), .Q(n36) );
  AOI221 U56 ( .A(i_data_alures[9]), .B(n4), .C(i_data_pc8[9]), .D(n1), .Q(n35) );
  INV3 U57 ( .A(i_con_pc8), .Q(n5) );
  INV3 U58 ( .A(n65), .Q(o_data_alu[10]) );
  AOI221 U59 ( .A(i_data_alures[10]), .B(n2), .C(i_data_pc8[10]), .D(i_con_pc8), .Q(n65) );
  INV3 U60 ( .A(n64), .Q(o_data_alu[11]) );
  AOI221 U61 ( .A(i_data_alures[11]), .B(n4), .C(i_data_pc8[11]), .D(i_con_pc8), .Q(n64) );
  INV3 U62 ( .A(n63), .Q(o_data_alu[12]) );
  AOI221 U63 ( .A(i_data_alures[12]), .B(n3), .C(i_data_pc8[12]), .D(i_con_pc8), .Q(n63) );
  INV3 U64 ( .A(n62), .Q(o_data_alu[13]) );
  AOI221 U65 ( .A(i_data_alures[13]), .B(n2), .C(i_data_pc8[13]), .D(i_con_pc8), .Q(n62) );
  INV3 U66 ( .A(n61), .Q(o_data_alu[14]) );
  AOI221 U67 ( .A(i_data_alures[14]), .B(n4), .C(i_data_pc8[14]), .D(i_con_pc8), .Q(n61) );
  INV3 U68 ( .A(n60), .Q(o_data_alu[15]) );
  AOI221 U69 ( .A(i_data_alures[15]), .B(n3), .C(i_data_pc8[15]), .D(i_con_pc8), .Q(n60) );
endmodule


module W_loadmux3 ( i_data_Rdata, i_con_loadsig, o_data_Wdata );
  input [31:0] i_data_Rdata;
  input [1:0] i_con_loadsig;
  output [31:0] o_data_Wdata;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n1, n2, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n52;

  BUF6 U2 ( .A(n24), .Q(n2) );
  AOI211 U3 ( .A(n42), .B(i_data_Rdata[15]), .C(n22), .Q(n24) );
  NOR20 U4 ( .A(n20), .B(n11), .Q(o_data_Wdata[7]) );
  NAND22 U5 ( .A(i_con_loadsig[1]), .B(n52), .Q(n49) );
  CLKIN3 U6 ( .A(i_con_loadsig[0]), .Q(n52) );
  NAND22 U7 ( .A(n50), .B(n49), .Q(n51) );
  AOI210 U8 ( .A(n19), .B(i_data_Rdata[10]), .C(n22), .Q(n48) );
  AOI210 U9 ( .A(n19), .B(i_data_Rdata[11]), .C(n22), .Q(n47) );
  AOI210 U10 ( .A(n19), .B(i_data_Rdata[12]), .C(n22), .Q(n46) );
  AOI210 U11 ( .A(n19), .B(i_data_Rdata[13]), .C(n22), .Q(n45) );
  AOI210 U12 ( .A(n19), .B(i_data_Rdata[14]), .C(n22), .Q(n44) );
  AOI210 U13 ( .A(n19), .B(i_data_Rdata[15]), .C(n22), .Q(n43) );
  NOR20 U14 ( .A(n52), .B(i_con_loadsig[1]), .Q(n42) );
  NAND20 U15 ( .A(i_data_Rdata[16]), .B(n26), .Q(n41) );
  NAND20 U16 ( .A(i_data_Rdata[17]), .B(n26), .Q(n40) );
  NAND20 U17 ( .A(i_data_Rdata[18]), .B(n26), .Q(n39) );
  NAND20 U18 ( .A(i_data_Rdata[19]), .B(n26), .Q(n38) );
  NAND20 U19 ( .A(i_data_Rdata[20]), .B(n26), .Q(n37) );
  NAND20 U20 ( .A(i_data_Rdata[21]), .B(n26), .Q(n36) );
  NAND20 U21 ( .A(i_data_Rdata[22]), .B(n26), .Q(n35) );
  CLKIN3 U22 ( .A(n23), .Q(o_data_Wdata[8]) );
  AOI210 U23 ( .A(n19), .B(i_data_Rdata[8]), .C(n22), .Q(n23) );
  CLKIN3 U24 ( .A(n21), .Q(o_data_Wdata[9]) );
  AOI210 U25 ( .A(n19), .B(i_data_Rdata[9]), .C(n22), .Q(n21) );
  INV3 U26 ( .A(n50), .Q(n19) );
  NOR21 U27 ( .A(n11), .B(n49), .Q(n22) );
  INV3 U28 ( .A(n51), .Q(n20) );
  BUF2 U29 ( .A(n26), .Q(n1) );
  NOR21 U30 ( .A(n42), .B(n26), .Q(n50) );
  INV3 U31 ( .A(n48), .Q(o_data_Wdata[10]) );
  INV3 U32 ( .A(n47), .Q(o_data_Wdata[11]) );
  INV3 U33 ( .A(n46), .Q(o_data_Wdata[12]) );
  INV3 U34 ( .A(n45), .Q(o_data_Wdata[13]) );
  INV3 U35 ( .A(n44), .Q(o_data_Wdata[14]) );
  INV3 U36 ( .A(n43), .Q(o_data_Wdata[15]) );
  NOR21 U37 ( .A(i_con_loadsig[0]), .B(i_con_loadsig[1]), .Q(n26) );
  NOR21 U38 ( .A(n20), .B(n18), .Q(o_data_Wdata[0]) );
  INV3 U39 ( .A(i_data_Rdata[0]), .Q(n18) );
  NOR21 U40 ( .A(n20), .B(n17), .Q(o_data_Wdata[1]) );
  INV3 U41 ( .A(i_data_Rdata[1]), .Q(n17) );
  NOR21 U42 ( .A(n20), .B(n16), .Q(o_data_Wdata[2]) );
  INV3 U43 ( .A(i_data_Rdata[2]), .Q(n16) );
  NOR21 U44 ( .A(n20), .B(n15), .Q(o_data_Wdata[3]) );
  INV3 U45 ( .A(i_data_Rdata[3]), .Q(n15) );
  NOR21 U46 ( .A(n20), .B(n14), .Q(o_data_Wdata[4]) );
  INV3 U47 ( .A(i_data_Rdata[4]), .Q(n14) );
  NOR21 U48 ( .A(n20), .B(n13), .Q(o_data_Wdata[5]) );
  INV3 U49 ( .A(i_data_Rdata[5]), .Q(n13) );
  NOR21 U50 ( .A(n20), .B(n12), .Q(o_data_Wdata[6]) );
  INV3 U51 ( .A(i_data_Rdata[6]), .Q(n12) );
  INV3 U52 ( .A(i_data_Rdata[7]), .Q(n11) );
  NAND22 U53 ( .A(n2), .B(n41), .Q(o_data_Wdata[16]) );
  NAND22 U54 ( .A(n2), .B(n40), .Q(o_data_Wdata[17]) );
  NAND22 U55 ( .A(n2), .B(n39), .Q(o_data_Wdata[18]) );
  NAND22 U56 ( .A(n2), .B(n38), .Q(o_data_Wdata[19]) );
  NAND22 U57 ( .A(n2), .B(n37), .Q(o_data_Wdata[20]) );
  NAND22 U58 ( .A(n2), .B(n36), .Q(o_data_Wdata[21]) );
  NAND22 U59 ( .A(n2), .B(n35), .Q(o_data_Wdata[22]) );
  NAND22 U60 ( .A(n2), .B(n34), .Q(o_data_Wdata[23]) );
  NAND22 U61 ( .A(i_data_Rdata[23]), .B(n1), .Q(n34) );
  NAND22 U62 ( .A(n2), .B(n33), .Q(o_data_Wdata[24]) );
  NAND22 U63 ( .A(i_data_Rdata[24]), .B(n1), .Q(n33) );
  NAND22 U64 ( .A(n2), .B(n32), .Q(o_data_Wdata[25]) );
  NAND22 U65 ( .A(i_data_Rdata[25]), .B(n1), .Q(n32) );
  NAND22 U66 ( .A(n2), .B(n31), .Q(o_data_Wdata[26]) );
  NAND22 U67 ( .A(i_data_Rdata[26]), .B(n1), .Q(n31) );
  NAND22 U68 ( .A(n2), .B(n30), .Q(o_data_Wdata[27]) );
  NAND22 U69 ( .A(i_data_Rdata[27]), .B(n1), .Q(n30) );
  NAND22 U70 ( .A(n2), .B(n29), .Q(o_data_Wdata[28]) );
  NAND22 U71 ( .A(i_data_Rdata[28]), .B(n1), .Q(n29) );
  NAND22 U72 ( .A(n2), .B(n28), .Q(o_data_Wdata[29]) );
  NAND22 U73 ( .A(i_data_Rdata[29]), .B(n1), .Q(n28) );
  NAND22 U74 ( .A(n2), .B(n27), .Q(o_data_Wdata[30]) );
  NAND22 U75 ( .A(i_data_Rdata[30]), .B(n1), .Q(n27) );
  NAND22 U76 ( .A(n2), .B(n25), .Q(o_data_Wdata[31]) );
  NAND22 U77 ( .A(i_data_Rdata[31]), .B(n1), .Q(n25) );
endmodule


module W_datamux ( i_data_alu, i_data_load, i_con_memtoreg, o_data_toreg );
  input [31:0] i_data_alu;
  input [31:0] i_data_load;
  output [31:0] o_data_toreg;
  input i_con_memtoreg;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n1, n2, n3, n4, n5, n6, n7;

  CLKIN3 U1 ( .A(n59), .Q(o_data_toreg[16]) );
  CLKIN3 U2 ( .A(n58), .Q(o_data_toreg[17]) );
  CLKIN3 U3 ( .A(n57), .Q(o_data_toreg[18]) );
  CLKIN3 U4 ( .A(n56), .Q(o_data_toreg[19]) );
  CLKIN3 U5 ( .A(n54), .Q(o_data_toreg[20]) );
  CLKIN3 U6 ( .A(n53), .Q(o_data_toreg[21]) );
  CLKIN3 U7 ( .A(n52), .Q(o_data_toreg[22]) );
  CLKIN3 U8 ( .A(n51), .Q(o_data_toreg[23]) );
  CLKIN3 U9 ( .A(n50), .Q(o_data_toreg[24]) );
  CLKIN3 U10 ( .A(n49), .Q(o_data_toreg[25]) );
  CLKIN3 U11 ( .A(n48), .Q(o_data_toreg[26]) );
  CLKIN3 U12 ( .A(n47), .Q(o_data_toreg[27]) );
  CLKIN3 U13 ( .A(n46), .Q(o_data_toreg[28]) );
  CLKIN3 U14 ( .A(n45), .Q(o_data_toreg[29]) );
  CLKIN3 U15 ( .A(n43), .Q(o_data_toreg[30]) );
  CLKIN3 U16 ( .A(n42), .Q(o_data_toreg[31]) );
  CLKIN3 U17 ( .A(n36), .Q(o_data_toreg[8]) );
  CLKIN3 U18 ( .A(n35), .Q(o_data_toreg[9]) );
  CLKIN3 U19 ( .A(n65), .Q(o_data_toreg[10]) );
  CLKIN3 U20 ( .A(n64), .Q(o_data_toreg[11]) );
  CLKIN3 U21 ( .A(n63), .Q(o_data_toreg[12]) );
  CLKIN3 U22 ( .A(n62), .Q(o_data_toreg[13]) );
  CLKIN3 U23 ( .A(n61), .Q(o_data_toreg[14]) );
  CLKIN3 U24 ( .A(n60), .Q(o_data_toreg[15]) );
  CLKIN3 U25 ( .A(n66), .Q(o_data_toreg[0]) );
  CLKIN3 U26 ( .A(n55), .Q(o_data_toreg[1]) );
  CLKIN3 U27 ( .A(n44), .Q(o_data_toreg[2]) );
  CLKIN3 U28 ( .A(n41), .Q(o_data_toreg[3]) );
  CLKIN3 U29 ( .A(n40), .Q(o_data_toreg[4]) );
  CLKIN3 U30 ( .A(n39), .Q(o_data_toreg[5]) );
  CLKIN3 U31 ( .A(n38), .Q(o_data_toreg[6]) );
  CLKIN3 U32 ( .A(n37), .Q(o_data_toreg[7]) );
  INV3 U33 ( .A(n2), .Q(n1) );
  BUF2 U34 ( .A(n7), .Q(n3) );
  BUF2 U35 ( .A(n7), .Q(n4) );
  BUF2 U36 ( .A(n7), .Q(n5) );
  BUF2 U37 ( .A(n7), .Q(n6) );
  AOI221 U38 ( .A(i_data_alu[0]), .B(n3), .C(i_data_load[0]), .D(n1), .Q(n66)
         );
  AOI221 U39 ( .A(i_data_alu[1]), .B(n4), .C(i_data_load[1]), .D(n1), .Q(n55)
         );
  AOI221 U40 ( .A(i_data_alu[2]), .B(n5), .C(i_data_load[2]), .D(n1), .Q(n44)
         );
  AOI221 U41 ( .A(i_data_alu[3]), .B(n6), .C(i_data_load[3]), .D(n1), .Q(n41)
         );
  AOI221 U42 ( .A(i_data_alu[4]), .B(n6), .C(i_data_load[4]), .D(n1), .Q(n40)
         );
  AOI221 U43 ( .A(i_data_alu[5]), .B(n6), .C(i_data_load[5]), .D(n1), .Q(n39)
         );
  AOI221 U44 ( .A(i_data_alu[6]), .B(n6), .C(i_data_load[6]), .D(n1), .Q(n38)
         );
  AOI221 U45 ( .A(i_data_alu[7]), .B(n6), .C(i_data_load[7]), .D(n1), .Q(n37)
         );
  AOI221 U46 ( .A(i_data_alu[8]), .B(n6), .C(i_data_load[8]), .D(n1), .Q(n36)
         );
  AOI221 U47 ( .A(i_data_alu[9]), .B(n6), .C(i_data_load[9]), .D(n1), .Q(n35)
         );
  AOI221 U48 ( .A(i_data_alu[10]), .B(n3), .C(i_data_load[10]), .D(n1), .Q(n65) );
  AOI221 U49 ( .A(i_data_alu[11]), .B(n3), .C(i_data_load[11]), .D(n1), .Q(n64) );
  AOI221 U50 ( .A(i_data_alu[12]), .B(n3), .C(i_data_load[12]), .D(n1), .Q(n63) );
  AOI221 U51 ( .A(i_data_alu[13]), .B(n3), .C(i_data_load[13]), .D(n1), .Q(n62) );
  AOI221 U52 ( .A(i_data_alu[14]), .B(n3), .C(i_data_load[14]), .D(n1), .Q(n61) );
  AOI221 U53 ( .A(i_data_alu[15]), .B(n3), .C(i_data_load[15]), .D(n1), .Q(n60) );
  AOI221 U54 ( .A(i_data_alu[16]), .B(n3), .C(i_data_load[16]), .D(n1), .Q(n59) );
  AOI221 U55 ( .A(i_data_alu[17]), .B(n4), .C(i_data_load[17]), .D(n1), .Q(n58) );
  AOI221 U56 ( .A(i_data_alu[18]), .B(n4), .C(i_data_load[18]), .D(n1), .Q(n57) );
  AOI221 U57 ( .A(i_data_alu[19]), .B(n4), .C(i_data_load[19]), .D(n1), .Q(n56) );
  AOI221 U58 ( .A(i_data_alu[20]), .B(n4), .C(i_data_load[20]), .D(n1), .Q(n54) );
  AOI221 U59 ( .A(i_data_alu[21]), .B(n4), .C(i_data_load[21]), .D(
        i_con_memtoreg), .Q(n53) );
  AOI221 U60 ( .A(i_data_alu[22]), .B(n4), .C(i_data_load[22]), .D(
        i_con_memtoreg), .Q(n52) );
  AOI221 U61 ( .A(i_data_alu[23]), .B(n4), .C(i_data_load[23]), .D(
        i_con_memtoreg), .Q(n51) );
  AOI221 U62 ( .A(i_data_alu[24]), .B(n5), .C(i_data_load[24]), .D(
        i_con_memtoreg), .Q(n50) );
  AOI221 U63 ( .A(i_data_alu[25]), .B(n5), .C(i_data_load[25]), .D(
        i_con_memtoreg), .Q(n49) );
  AOI221 U64 ( .A(i_data_alu[26]), .B(n5), .C(i_data_load[26]), .D(
        i_con_memtoreg), .Q(n48) );
  AOI221 U65 ( .A(i_data_alu[27]), .B(n5), .C(i_data_load[27]), .D(
        i_con_memtoreg), .Q(n47) );
  AOI221 U66 ( .A(i_data_alu[28]), .B(n5), .C(i_data_load[28]), .D(
        i_con_memtoreg), .Q(n46) );
  AOI221 U67 ( .A(i_data_alu[29]), .B(n5), .C(i_data_load[29]), .D(
        i_con_memtoreg), .Q(n45) );
  AOI221 U68 ( .A(i_data_alu[30]), .B(n5), .C(i_data_load[30]), .D(
        i_con_memtoreg), .Q(n43) );
  AOI221 U69 ( .A(i_data_alu[31]), .B(n6), .C(i_data_load[31]), .D(
        i_con_memtoreg), .Q(n42) );
  BUF2 U70 ( .A(n7), .Q(n2) );
  INV3 U71 ( .A(i_con_memtoreg), .Q(n7) );
endmodule


module writeback ( i_data_pc8, i_data_alures, i_data_memout, i_con_Wloadmux, 
        i_con_Walupc8, i_con_Wmemtoreg, o_data_regwrite );
  input [31:0] i_data_pc8;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [1:0] i_con_Wloadmux;
  output [31:0] o_data_regwrite;
  input i_con_Walupc8, i_con_Wmemtoreg;

  wire   [31:0] datamux_i_data_alu;
  wire   [31:0] datamux_i_data_load;

  W_resmux u_resmux ( .i_data_alures(i_data_alures), .i_data_pc8(i_data_pc8), 
        .i_con_pc8(i_con_Walupc8), .o_data_alu(datamux_i_data_alu) );
  W_loadmux3 u_loadmux ( .i_data_Rdata(i_data_memout), .i_con_loadsig(
        i_con_Wloadmux), .o_data_Wdata(datamux_i_data_load) );
  W_datamux u_datamux ( .i_data_alu(datamux_i_data_alu), .i_data_load(
        datamux_i_data_load), .i_con_memtoreg(i_con_Wmemtoreg), .o_data_toreg(
        o_data_regwrite) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Walupc8, mem_con_Walupc8, mem_con_Wmemtoreg, wb_con_Walupc8,
         wb_con_Wmemtoreg, n1;
  wire   [31:0] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [31:0] id_addr_pc4;
  wire   [31:0] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] for_aluresE;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] wb_data_memout;
  wire   [31:0] mem_data_pc4;
  wire   [1:0] mem_con_Wloadmux;
  wire   [31:0] wb_data_pc8;
  wire   [31:0] mem_data_alures;
  wire   [1:0] wb_con_Wloadmux;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  fetch u_fetch ( .i_clk(clk), .i_nrst(rst_n), .i_addr_b(if_addr_b), 
        .i_addr_j({if_addr_j, n1, n1}), .i_addr_jr(id_data_jr), .i_con_b(
        if_con_b), .i_con_j(if_con_j), .i_data_instr(read_instruction), 
        .i_con_ifstall(if_con_ifstall), .o_addr_pc(instruction_address), 
        .o_addr_pc4(id_addr_pc4), .o_data_instr(id_data_instr) );
  decode u_decode ( .i_clk(clk), .i_nrst(rst_n), .i_addr_pc4(id_addr_pc4), 
        .i_data_instr(id_data_instr), .i_con_Wregwrite(id_con_Wregwrite), 
        .i_data_Wregwrite(id_data_Wregwrite), .i_addr_Wregwrite(
        id_addr_Wregwrite), .i_addr_Erd(for_o_addr_Erd), .i_addr_Mrd(
        mem_addr_regdst), .i_con_Eregwrite(ex_con_Wregwrite), 
        .i_con_Mregwrite(mem_con_Wregwrite), .i_addr_rtM(for_addr_rtM), 
        .i_addr_rtW(for_addr_rtW), .i_con_memreadM(mem_read), .i_con_memreadW(
        for_FWmemread), .i_data_aluresE(for_aluresE), .i_data_memoutM(
        read_data), .o_data_rs(id_data_rs), .o_data_rt(ex_data_rt), 
        .o_addr_rd(ex_addr_rd), .o_addr_rt(ex_addr_rt), .o_data_jr(id_data_jr), 
        .o_con_jump(if_con_j), .o_addr_pc4(ex_data_pc4), .o_addr_branch(
        if_addr_b), .o_addr_jump({if_addr_j, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1}), .o_con_Ealuop(ex_con_Ealuop), 
        .o_con_Ealusrc(ex_con_Ealusrc), .o_con_Eregdst(ex_con_Eregdst), 
        .o_con_Walupc8(ex_con_Walupc8), .o_con_Wregwrite(ex_con_Wregwrite), 
        .o_con_ifstall(if_con_ifstall), .o_con_Ebop(ex_con_bop), 
        .o_data_signext(ex_data_immext), .o_con_Efamux(for_o_con_Efamux), 
        .o_con_Efbmux(for_o_con_Efbmux), .o_data_Fmemout(for_memout) );
  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext(
        ex_data_immext), .i_addr_rt(ex_addr_rt), .i_addr_rd(ex_addr_rd), 
        .i_data_FEalures(data_address), .i_data_FMalures(id_data_Wregwrite), 
        .i_data_FMmemout(wb_data_memout), .i_data_FWmemout(for_memout), 
        .i_con_Ealuop(ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(n1), .i_con_Mmemwrite(
        n1), .i_con_Wloadmux({n1, n1}), .i_con_Walupc8(ex_con_Walupc8), 
        .i_con_Wmemtoreg(n1), .i_con_Wregwrite(ex_con_Wregwrite), 
        .i_con_Efamux(for_o_con_Efamux), .i_con_Efbmux(for_o_con_Efbmux), 
        .i_con_bop(ex_con_bop), .o_data_pc4(mem_data_pc4), .o_data_alures(
        data_address), .o_data_rt(write_data), .o_addr_regdst(mem_addr_regdst), 
        .o_con_Mmemread(mem_read), .o_con_Mmemwrite(mem_write), 
        .o_con_Wloadmux(mem_con_Wloadmux), .o_con_Walupc8(mem_con_Walupc8), 
        .o_con_Wmemtoreg(mem_con_Wmemtoreg), .o_con_Wregwrite(
        mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), .o_addr_Mrt(
        for_addr_rtM), .o_FaluresE(for_aluresE), .o_con_ifbranch(if_con_b) );
  mem u_mem ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(mem_data_pc4), 
        .i_data_alures(data_address), .i_data_memout(read_data), 
        .i_addr_regdst(mem_addr_regdst), .i_con_Wloadmux(mem_con_Wloadmux), 
        .i_con_Walupc8(mem_con_Walupc8), .i_con_Wmemtoreg(mem_con_Wmemtoreg), 
        .i_con_Wregwrite(mem_con_Wregwrite), .i_con_FWmemread(n1), 
        .i_addr_Mrt(for_addr_rtM), .o_data_pc8(wb_data_pc8), .o_data_alures(
        mem_data_alures), .o_data_memout(wb_data_memout), .o_addr_regdst(
        id_addr_Wregwrite), .o_con_Wloadmux(wb_con_Wloadmux), .o_con_Walupc8(
        wb_con_Walupc8), .o_con_Wmemtoreg(wb_con_Wmemtoreg), .o_con_Wregwrite(
        id_con_Wregwrite), .o_con_FWmemread(for_FWmemread), .o_addr_Wrt(
        for_addr_rtW) );
  writeback u_writeback ( .i_data_pc8(wb_data_pc8), .i_data_alures(
        mem_data_alures), .i_data_memout(wb_data_memout), .i_con_Wloadmux(
        wb_con_Wloadmux), .i_con_Walupc8(wb_con_Walupc8), .i_con_Wmemtoreg(
        wb_con_Wmemtoreg), .o_data_regwrite(id_data_Wregwrite) );
  LOGIC0 U1 ( .Q(n1) );
endmodule

