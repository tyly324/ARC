
module F_jumpmux ( i_addr_j, i_addr_jr, i_addr_pc4, i_con_jump, o_addr_jumpmux
 );
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [31:0] i_addr_pc4;
  input [1:0] i_con_jump;
  output [31:0] o_addr_jumpmux;
  wire   n3, n4, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n23,
         n24, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n1, n2, n5, n6, n19, n20,
         n21, n22, n25, n26, n27, n28, n29, n30, n31, n32, n69, n70, n71, n72;

  BUF2 U1 ( .A(n71), .Q(n1) );
  AOI221 U2 ( .A(i_addr_pc4[3]), .B(n1), .C(i_addr_jr[3]), .D(n70), .Q(n17) );
  AOI221 U3 ( .A(i_addr_pc4[4]), .B(n1), .C(i_addr_jr[4]), .D(n70), .Q(n15) );
  AOI221 U4 ( .A(i_addr_pc4[5]), .B(n1), .C(i_addr_jr[5]), .D(n70), .Q(n13) );
  AOI221 U5 ( .A(i_addr_pc4[6]), .B(n1), .C(i_addr_jr[6]), .D(n70), .Q(n11) );
  AOI221 U6 ( .A(i_addr_pc4[7]), .B(n1), .C(i_addr_jr[7]), .D(n70), .Q(n9) );
  AOI221 U7 ( .A(i_addr_pc4[8]), .B(n1), .C(i_addr_jr[8]), .D(n70), .Q(n7) );
  AOI221 U8 ( .A(i_addr_pc4[9]), .B(n1), .C(i_addr_jr[9]), .D(n70), .Q(n3) );
  AOI221 U9 ( .A(i_addr_pc4[2]), .B(n71), .C(i_addr_jr[2]), .D(n70), .Q(n23)
         );
  AOI221 U10 ( .A(i_addr_pc4[15]), .B(n1), .C(i_addr_jr[15]), .D(n70), .Q(n55)
         );
  AOI221 U11 ( .A(i_addr_pc4[16]), .B(n71), .C(i_addr_jr[16]), .D(n70), .Q(n53) );
  AOI221 U12 ( .A(i_addr_pc4[17]), .B(n71), .C(i_addr_jr[17]), .D(n70), .Q(n51) );
  AOI221 U13 ( .A(i_addr_pc4[18]), .B(n71), .C(i_addr_jr[18]), .D(n70), .Q(n49) );
  AOI221 U14 ( .A(i_addr_pc4[19]), .B(n71), .C(i_addr_jr[19]), .D(n70), .Q(n47) );
  AOI221 U15 ( .A(i_addr_pc4[20]), .B(n71), .C(i_addr_jr[20]), .D(n70), .Q(n43) );
  AOI221 U16 ( .A(i_addr_pc4[21]), .B(n71), .C(i_addr_jr[21]), .D(n70), .Q(n41) );
  AOI221 U17 ( .A(i_addr_pc4[22]), .B(n71), .C(i_addr_jr[22]), .D(n70), .Q(n39) );
  AOI221 U18 ( .A(i_addr_pc4[23]), .B(n71), .C(i_addr_jr[23]), .D(n70), .Q(n37) );
  AOI221 U19 ( .A(i_addr_pc4[24]), .B(n71), .C(i_addr_jr[24]), .D(n70), .Q(n35) );
  AOI221 U20 ( .A(i_addr_pc4[25]), .B(n1), .C(i_addr_jr[25]), .D(n70), .Q(n33)
         );
  AOI221 U21 ( .A(i_addr_pc4[10]), .B(n1), .C(i_addr_jr[10]), .D(n70), .Q(n65)
         );
  AOI221 U22 ( .A(i_addr_pc4[11]), .B(n1), .C(i_addr_jr[11]), .D(n70), .Q(n63)
         );
  AOI221 U23 ( .A(i_addr_pc4[12]), .B(n1), .C(i_addr_jr[12]), .D(n70), .Q(n61)
         );
  AOI221 U24 ( .A(i_addr_pc4[13]), .B(n1), .C(i_addr_jr[13]), .D(n70), .Q(n59)
         );
  AOI221 U25 ( .A(i_addr_pc4[14]), .B(n1), .C(i_addr_jr[14]), .D(n70), .Q(n57)
         );
  INV3 U26 ( .A(n19), .Q(n70) );
  NAND22 U27 ( .A(n67), .B(n68), .Q(o_addr_jumpmux[0]) );
  NAND22 U28 ( .A(i_addr_j[0]), .B(n72), .Q(n68) );
  NAND22 U29 ( .A(n65), .B(n66), .Q(o_addr_jumpmux[10]) );
  NAND22 U30 ( .A(i_addr_j[10]), .B(n72), .Q(n66) );
  NAND22 U31 ( .A(n63), .B(n64), .Q(o_addr_jumpmux[11]) );
  NAND22 U32 ( .A(i_addr_j[11]), .B(n72), .Q(n64) );
  NAND22 U33 ( .A(n61), .B(n62), .Q(o_addr_jumpmux[12]) );
  NAND22 U34 ( .A(i_addr_j[12]), .B(n72), .Q(n62) );
  NAND22 U35 ( .A(n59), .B(n60), .Q(o_addr_jumpmux[13]) );
  NAND22 U36 ( .A(i_addr_j[13]), .B(n72), .Q(n60) );
  NAND22 U37 ( .A(n57), .B(n58), .Q(o_addr_jumpmux[14]) );
  NAND22 U38 ( .A(i_addr_j[14]), .B(n72), .Q(n58) );
  NAND22 U39 ( .A(n55), .B(n56), .Q(o_addr_jumpmux[15]) );
  NAND22 U40 ( .A(i_addr_j[15]), .B(n72), .Q(n56) );
  NAND22 U41 ( .A(n53), .B(n54), .Q(o_addr_jumpmux[16]) );
  NAND22 U42 ( .A(i_addr_j[16]), .B(n72), .Q(n54) );
  NAND22 U43 ( .A(n51), .B(n52), .Q(o_addr_jumpmux[17]) );
  NAND22 U44 ( .A(i_addr_j[17]), .B(n72), .Q(n52) );
  NAND22 U45 ( .A(n49), .B(n50), .Q(o_addr_jumpmux[18]) );
  NAND22 U46 ( .A(i_addr_j[18]), .B(n72), .Q(n50) );
  NAND22 U47 ( .A(n47), .B(n48), .Q(o_addr_jumpmux[19]) );
  NAND22 U48 ( .A(i_addr_j[19]), .B(n72), .Q(n48) );
  NAND22 U49 ( .A(n3), .B(n4), .Q(o_addr_jumpmux[9]) );
  NAND22 U50 ( .A(i_addr_j[9]), .B(n72), .Q(n4) );
  NAND22 U51 ( .A(n45), .B(n46), .Q(o_addr_jumpmux[1]) );
  NAND22 U52 ( .A(i_addr_j[1]), .B(n72), .Q(n46) );
  NAND22 U53 ( .A(n23), .B(n24), .Q(o_addr_jumpmux[2]) );
  NAND22 U54 ( .A(i_addr_j[2]), .B(n72), .Q(n24) );
  NAND22 U55 ( .A(n17), .B(n18), .Q(o_addr_jumpmux[3]) );
  NAND22 U56 ( .A(i_addr_j[3]), .B(n72), .Q(n18) );
  NAND22 U57 ( .A(n15), .B(n16), .Q(o_addr_jumpmux[4]) );
  NAND22 U58 ( .A(i_addr_j[4]), .B(n72), .Q(n16) );
  NAND22 U59 ( .A(n13), .B(n14), .Q(o_addr_jumpmux[5]) );
  NAND22 U60 ( .A(i_addr_j[5]), .B(n72), .Q(n14) );
  NAND22 U61 ( .A(n11), .B(n12), .Q(o_addr_jumpmux[6]) );
  NAND22 U62 ( .A(i_addr_j[6]), .B(n72), .Q(n12) );
  NAND22 U63 ( .A(n9), .B(n10), .Q(o_addr_jumpmux[7]) );
  NAND22 U64 ( .A(i_addr_j[7]), .B(n72), .Q(n10) );
  NAND22 U65 ( .A(n7), .B(n8), .Q(o_addr_jumpmux[8]) );
  NAND22 U66 ( .A(i_addr_j[8]), .B(n72), .Q(n8) );
  NAND22 U67 ( .A(n43), .B(n44), .Q(o_addr_jumpmux[20]) );
  NAND22 U68 ( .A(i_addr_j[20]), .B(n72), .Q(n44) );
  NAND22 U69 ( .A(n41), .B(n42), .Q(o_addr_jumpmux[21]) );
  NAND22 U70 ( .A(i_addr_j[21]), .B(n72), .Q(n42) );
  NAND22 U71 ( .A(n39), .B(n40), .Q(o_addr_jumpmux[22]) );
  NAND22 U72 ( .A(i_addr_j[22]), .B(n72), .Q(n40) );
  NAND22 U73 ( .A(n37), .B(n38), .Q(o_addr_jumpmux[23]) );
  NAND22 U74 ( .A(i_addr_j[23]), .B(n72), .Q(n38) );
  NAND22 U75 ( .A(n35), .B(n36), .Q(o_addr_jumpmux[24]) );
  NAND22 U76 ( .A(i_addr_j[24]), .B(n72), .Q(n36) );
  NAND22 U77 ( .A(n33), .B(n34), .Q(o_addr_jumpmux[25]) );
  NAND22 U78 ( .A(i_addr_j[25]), .B(n72), .Q(n34) );
  AOI221 U79 ( .A(i_addr_j[26]), .B(n72), .C(i_addr_pc4[26]), .D(n1), .Q(n21)
         );
  AOI221 U80 ( .A(i_addr_j[27]), .B(n72), .C(i_addr_pc4[27]), .D(n1), .Q(n25)
         );
  AOI221 U81 ( .A(i_addr_j[28]), .B(n72), .C(i_addr_pc4[28]), .D(n71), .Q(n27)
         );
  AOI221 U82 ( .A(i_addr_j[29]), .B(n72), .C(i_addr_pc4[29]), .D(n71), .Q(n29)
         );
  AOI221 U83 ( .A(i_addr_j[30]), .B(n72), .C(i_addr_pc4[30]), .D(n71), .Q(n31)
         );
  AOI221 U84 ( .A(i_addr_j[31]), .B(n72), .C(i_addr_pc4[31]), .D(n71), .Q(n69)
         );
  AOI221 U85 ( .A(i_addr_pc4[1]), .B(n1), .C(i_addr_jr[1]), .D(n70), .Q(n45)
         );
  AOI221 U86 ( .A(i_addr_pc4[0]), .B(n1), .C(i_addr_jr[0]), .D(n70), .Q(n67)
         );
  CLKIN3 U87 ( .A(i_con_jump[1]), .Q(n2) );
  NAND22 U88 ( .A(i_con_jump[0]), .B(n2), .Q(n5) );
  CLKIN3 U89 ( .A(n5), .Q(n72) );
  XNR21 U90 ( .A(i_con_jump[0]), .B(i_con_jump[1]), .Q(n71) );
  CLKIN3 U91 ( .A(i_con_jump[0]), .Q(n6) );
  NAND22 U92 ( .A(i_con_jump[1]), .B(n6), .Q(n19) );
  NAND22 U93 ( .A(i_addr_jr[26]), .B(n70), .Q(n20) );
  NAND22 U94 ( .A(n21), .B(n20), .Q(o_addr_jumpmux[26]) );
  NAND22 U95 ( .A(i_addr_jr[27]), .B(n70), .Q(n22) );
  NAND22 U96 ( .A(n25), .B(n22), .Q(o_addr_jumpmux[27]) );
  NAND22 U97 ( .A(i_addr_jr[28]), .B(n70), .Q(n26) );
  NAND22 U98 ( .A(n27), .B(n26), .Q(o_addr_jumpmux[28]) );
  NAND22 U99 ( .A(i_addr_jr[29]), .B(n70), .Q(n28) );
  NAND22 U100 ( .A(n29), .B(n28), .Q(o_addr_jumpmux[29]) );
  NAND22 U101 ( .A(i_addr_jr[30]), .B(n70), .Q(n30) );
  NAND22 U102 ( .A(n31), .B(n30), .Q(o_addr_jumpmux[30]) );
  NAND22 U103 ( .A(i_addr_jr[31]), .B(n70), .Q(n32) );
  NAND22 U104 ( .A(n69), .B(n32), .Q(o_addr_jumpmux[31]) );
endmodule


module F_branchmux ( i_addr_jumpmux, i_addr_b, i_con_ifbranch, o_addr_nextpc
 );
  input [31:0] i_addr_jumpmux;
  input [31:0] i_addr_b;
  output [31:0] o_addr_nextpc;
  input i_con_ifbranch;
  wire   n34, n35, n36, n37, n38, n39, n40, n43, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n1, n2,
         n3, n4, n5;

  INV3 U1 ( .A(n5), .Q(n1) );
  INV3 U2 ( .A(n5), .Q(n2) );
  BUF2 U3 ( .A(n5), .Q(n3) );
  BUF2 U4 ( .A(n5), .Q(n4) );
  INV3 U5 ( .A(i_con_ifbranch), .Q(n5) );
  INV3 U6 ( .A(n65), .Q(o_addr_nextpc[0]) );
  AOI221 U7 ( .A(i_addr_b[0]), .B(n1), .C(i_addr_jumpmux[0]), .D(n4), .Q(n65)
         );
  INV3 U8 ( .A(n64), .Q(o_addr_nextpc[10]) );
  AOI221 U9 ( .A(i_addr_b[10]), .B(n1), .C(i_addr_jumpmux[10]), .D(n4), .Q(n64) );
  INV3 U10 ( .A(n63), .Q(o_addr_nextpc[11]) );
  AOI221 U11 ( .A(i_addr_b[11]), .B(n1), .C(i_addr_jumpmux[11]), .D(n4), .Q(
        n63) );
  INV3 U12 ( .A(n62), .Q(o_addr_nextpc[12]) );
  AOI221 U13 ( .A(i_addr_b[12]), .B(n1), .C(i_addr_jumpmux[12]), .D(n4), .Q(
        n62) );
  INV3 U14 ( .A(n61), .Q(o_addr_nextpc[13]) );
  AOI221 U15 ( .A(i_addr_b[13]), .B(n1), .C(i_addr_jumpmux[13]), .D(n4), .Q(
        n61) );
  INV3 U16 ( .A(n60), .Q(o_addr_nextpc[14]) );
  AOI221 U17 ( .A(i_addr_b[14]), .B(n1), .C(i_addr_jumpmux[14]), .D(n4), .Q(
        n60) );
  INV3 U18 ( .A(n59), .Q(o_addr_nextpc[15]) );
  AOI221 U19 ( .A(i_addr_b[15]), .B(n1), .C(i_addr_jumpmux[15]), .D(n4), .Q(
        n59) );
  INV3 U20 ( .A(n58), .Q(o_addr_nextpc[16]) );
  AOI221 U21 ( .A(i_addr_b[16]), .B(n1), .C(i_addr_jumpmux[16]), .D(n3), .Q(
        n58) );
  INV3 U22 ( .A(n57), .Q(o_addr_nextpc[17]) );
  AOI221 U23 ( .A(i_addr_b[17]), .B(n1), .C(i_addr_jumpmux[17]), .D(n3), .Q(
        n57) );
  INV3 U24 ( .A(n56), .Q(o_addr_nextpc[18]) );
  AOI221 U25 ( .A(i_addr_b[18]), .B(n1), .C(i_addr_jumpmux[18]), .D(n3), .Q(
        n56) );
  INV3 U26 ( .A(n55), .Q(o_addr_nextpc[19]) );
  AOI221 U27 ( .A(i_addr_b[19]), .B(n1), .C(i_addr_jumpmux[19]), .D(n3), .Q(
        n55) );
  INV3 U28 ( .A(n34), .Q(o_addr_nextpc[9]) );
  AOI221 U29 ( .A(n2), .B(i_addr_b[9]), .C(i_addr_jumpmux[9]), .D(n5), .Q(n34)
         );
  INV3 U30 ( .A(n54), .Q(o_addr_nextpc[1]) );
  AOI221 U31 ( .A(i_addr_b[1]), .B(n2), .C(i_addr_jumpmux[1]), .D(n3), .Q(n54)
         );
  INV3 U32 ( .A(n43), .Q(o_addr_nextpc[2]) );
  AOI221 U33 ( .A(i_addr_b[2]), .B(n2), .C(i_addr_jumpmux[2]), .D(n5), .Q(n43)
         );
  INV3 U34 ( .A(n40), .Q(o_addr_nextpc[3]) );
  AOI221 U35 ( .A(i_addr_b[3]), .B(n2), .C(i_addr_jumpmux[3]), .D(n5), .Q(n40)
         );
  INV3 U36 ( .A(n39), .Q(o_addr_nextpc[4]) );
  AOI221 U37 ( .A(i_addr_b[4]), .B(n2), .C(i_addr_jumpmux[4]), .D(n5), .Q(n39)
         );
  INV3 U38 ( .A(n38), .Q(o_addr_nextpc[5]) );
  AOI221 U39 ( .A(i_addr_b[5]), .B(n2), .C(i_addr_jumpmux[5]), .D(n5), .Q(n38)
         );
  INV3 U40 ( .A(n37), .Q(o_addr_nextpc[6]) );
  AOI221 U41 ( .A(i_addr_b[6]), .B(n2), .C(i_addr_jumpmux[6]), .D(n5), .Q(n37)
         );
  INV3 U42 ( .A(n36), .Q(o_addr_nextpc[7]) );
  AOI221 U43 ( .A(i_addr_b[7]), .B(n2), .C(i_addr_jumpmux[7]), .D(n4), .Q(n36)
         );
  INV3 U44 ( .A(n35), .Q(o_addr_nextpc[8]) );
  AOI221 U45 ( .A(i_addr_b[8]), .B(n2), .C(i_addr_jumpmux[8]), .D(n5), .Q(n35)
         );
  INV3 U46 ( .A(n53), .Q(o_addr_nextpc[20]) );
  AOI221 U47 ( .A(i_addr_b[20]), .B(n2), .C(i_addr_jumpmux[20]), .D(n3), .Q(
        n53) );
  INV3 U48 ( .A(n52), .Q(o_addr_nextpc[21]) );
  AOI221 U49 ( .A(i_addr_b[21]), .B(n2), .C(i_addr_jumpmux[21]), .D(n3), .Q(
        n52) );
  INV3 U50 ( .A(n51), .Q(o_addr_nextpc[22]) );
  AOI221 U51 ( .A(i_addr_b[22]), .B(n2), .C(i_addr_jumpmux[22]), .D(n3), .Q(
        n51) );
  INV3 U52 ( .A(n50), .Q(o_addr_nextpc[23]) );
  AOI221 U53 ( .A(i_addr_b[23]), .B(n2), .C(i_addr_jumpmux[23]), .D(n5), .Q(
        n50) );
  INV3 U54 ( .A(n49), .Q(o_addr_nextpc[24]) );
  AOI221 U55 ( .A(i_addr_b[24]), .B(n2), .C(i_addr_jumpmux[24]), .D(n5), .Q(
        n49) );
  INV3 U56 ( .A(n48), .Q(o_addr_nextpc[25]) );
  AOI221 U57 ( .A(i_addr_b[25]), .B(n2), .C(i_addr_jumpmux[25]), .D(n5), .Q(
        n48) );
  MUX22 U58 ( .A(i_addr_jumpmux[26]), .B(i_addr_b[26]), .S(n1), .Q(
        o_addr_nextpc[26]) );
  MUX22 U59 ( .A(i_addr_jumpmux[27]), .B(i_addr_b[27]), .S(n1), .Q(
        o_addr_nextpc[27]) );
  MUX22 U60 ( .A(i_addr_jumpmux[28]), .B(i_addr_b[28]), .S(n1), .Q(
        o_addr_nextpc[28]) );
  MUX22 U61 ( .A(i_addr_jumpmux[29]), .B(i_addr_b[29]), .S(n1), .Q(
        o_addr_nextpc[29]) );
  MUX22 U62 ( .A(i_addr_jumpmux[30]), .B(i_addr_b[30]), .S(n1), .Q(
        o_addr_nextpc[30]) );
  MUX22 U63 ( .A(i_addr_jumpmux[31]), .B(i_addr_b[31]), .S(n1), .Q(
        o_addr_nextpc[31]) );
endmodule


module F_pc ( i_clk, i_rst_n, i_con_stall, i_addr_next_pc, o_addr_pc );
  input [31:0] i_addr_next_pc;
  output [31:0] o_addr_pc;
  input i_clk, i_rst_n, i_con_stall;


  DFEC1 program_counter_reg_31_ ( .D(i_addr_next_pc[31]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[31]) );
  DFEC1 program_counter_reg_1_ ( .D(i_addr_next_pc[1]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[1]) );
  DFEC1 program_counter_reg_0_ ( .D(i_addr_next_pc[0]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[0]) );
  DFEC1 program_counter_reg_30_ ( .D(i_addr_next_pc[30]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[30]) );
  DFEC1 program_counter_reg_29_ ( .D(i_addr_next_pc[29]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[29]) );
  DFEC1 program_counter_reg_26_ ( .D(i_addr_next_pc[26]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[26]) );
  DFEC1 program_counter_reg_25_ ( .D(i_addr_next_pc[25]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[25]) );
  DFEC1 program_counter_reg_27_ ( .D(i_addr_next_pc[27]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[27]) );
  DFEC1 program_counter_reg_28_ ( .D(i_addr_next_pc[28]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[28]) );
  DFEC1 program_counter_reg_22_ ( .D(i_addr_next_pc[22]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[22]) );
  DFEC1 program_counter_reg_21_ ( .D(i_addr_next_pc[21]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[21]) );
  DFEC1 program_counter_reg_18_ ( .D(i_addr_next_pc[18]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[18]) );
  DFEC1 program_counter_reg_17_ ( .D(i_addr_next_pc[17]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[17]) );
  DFEC1 program_counter_reg_14_ ( .D(i_addr_next_pc[14]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[14]) );
  DFEC1 program_counter_reg_13_ ( .D(i_addr_next_pc[13]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[13]) );
  DFEC1 program_counter_reg_10_ ( .D(i_addr_next_pc[10]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[10]) );
  DFEC1 program_counter_reg_9_ ( .D(i_addr_next_pc[9]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[9]) );
  DFEC1 program_counter_reg_23_ ( .D(i_addr_next_pc[23]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[23]) );
  DFEC1 program_counter_reg_19_ ( .D(i_addr_next_pc[19]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[19]) );
  DFEC1 program_counter_reg_15_ ( .D(i_addr_next_pc[15]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[15]) );
  DFEC1 program_counter_reg_11_ ( .D(i_addr_next_pc[11]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[11]) );
  DFEC1 program_counter_reg_24_ ( .D(i_addr_next_pc[24]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[24]) );
  DFEC1 program_counter_reg_20_ ( .D(i_addr_next_pc[20]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[20]) );
  DFEC1 program_counter_reg_16_ ( .D(i_addr_next_pc[16]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[16]) );
  DFEC1 program_counter_reg_12_ ( .D(i_addr_next_pc[12]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[12]) );
  DFEC1 program_counter_reg_6_ ( .D(i_addr_next_pc[6]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[6]) );
  DFEC1 program_counter_reg_5_ ( .D(i_addr_next_pc[5]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[5]) );
  DFEC1 program_counter_reg_2_ ( .D(i_addr_next_pc[2]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[2]) );
  DFEC1 program_counter_reg_7_ ( .D(i_addr_next_pc[7]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[7]) );
  DFEC1 program_counter_reg_3_ ( .D(i_addr_next_pc[3]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[3]) );
  DFEC1 program_counter_reg_8_ ( .D(i_addr_next_pc[8]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[8]) );
  DFEC1 program_counter_reg_4_ ( .D(i_addr_next_pc[4]), .E(i_con_stall), .C(
        i_clk), .RN(i_rst_n), .Q(o_addr_pc[4]) );
endmodule


module F_add4_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  NOR21 U2 ( .A(n81), .B(n82), .Q(n80) );
  INV3 U3 ( .A(n83), .Q(n81) );
  NOR31 U4 ( .A(n10), .B(n84), .C(n7), .Q(n83) );
  NAND22 U5 ( .A(n34), .B(n35), .Q(n33) );
  NOR31 U6 ( .A(n38), .B(n36), .C(n37), .Q(n35) );
  NOR21 U7 ( .A(n22), .B(n33), .Q(n21) );
  INV3 U8 ( .A(n23), .Q(n22) );
  NOR31 U9 ( .A(n26), .B(n24), .C(n25), .Q(n23) );
  XNR21 U10 ( .A(n29), .B(n25), .Q(SUM[26]) );
  NOR21 U11 ( .A(n26), .B(n30), .Q(n29) );
  INV3 U12 ( .A(n57), .Q(n46) );
  NAND31 U13 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  NOR21 U14 ( .A(n62), .B(n63), .Q(n58) );
  INV3 U15 ( .A(n61), .Q(n59) );
  XNR21 U16 ( .A(n31), .B(n26), .Q(SUM[25]) );
  XNR21 U17 ( .A(n68), .B(n63), .Q(SUM[13]) );
  XNR21 U18 ( .A(n55), .B(n50), .Q(SUM[17]) );
  XNR21 U19 ( .A(n43), .B(n38), .Q(SUM[21]) );
  XNR21 U20 ( .A(n66), .B(n62), .Q(SUM[14]) );
  XNR21 U21 ( .A(n53), .B(n49), .Q(SUM[18]) );
  XNR21 U22 ( .A(n41), .B(n37), .Q(SUM[22]) );
  XNR21 U23 ( .A(n77), .B(n74), .Q(SUM[10]) );
  NOR21 U24 ( .A(n78), .B(n2), .Q(n77) );
  NOR21 U25 ( .A(n50), .B(n54), .Q(n53) );
  NOR21 U26 ( .A(n63), .B(n67), .Q(n66) );
  NOR21 U27 ( .A(n38), .B(n42), .Q(n41) );
  XNR21 U28 ( .A(n1), .B(n2), .Q(SUM[9]) );
  XNR21 U29 ( .A(n9), .B(n10), .Q(SUM[5]) );
  XNR21 U30 ( .A(n6), .B(n7), .Q(SUM[6]) );
  INV3 U31 ( .A(n8), .Q(n6) );
  NAND22 U32 ( .A(n9), .B(A[5]), .Q(n8) );
  NAND22 U33 ( .A(A[3]), .B(A[2]), .Q(n82) );
  XNR21 U34 ( .A(A[29]), .B(n15), .Q(SUM[29]) );
  XOR21 U35 ( .A(A[30]), .B(n14), .Q(SUM[30]) );
  XOR21 U36 ( .A(n27), .B(n28), .Q(SUM[27]) );
  INV3 U37 ( .A(A[27]), .Q(n27) );
  NAND22 U38 ( .A(n29), .B(A[26]), .Q(n28) );
  XOR21 U39 ( .A(n12), .B(n13), .Q(SUM[31]) );
  INV3 U40 ( .A(A[31]), .Q(n12) );
  NAND22 U41 ( .A(A[30]), .B(n14), .Q(n13) );
  NOR21 U42 ( .A(n19), .B(n20), .Q(n18) );
  INV3 U43 ( .A(A[28]), .Q(n20) );
  NOR21 U44 ( .A(n71), .B(n3), .Q(n60) );
  INV3 U45 ( .A(n72), .Q(n71) );
  NOR31 U46 ( .A(n2), .B(n73), .C(n74), .Q(n72) );
  NAND22 U47 ( .A(A[11]), .B(A[8]), .Q(n73) );
  NOR21 U48 ( .A(n33), .B(n32), .Q(n31) );
  INV3 U49 ( .A(A[24]), .Q(n32) );
  INV3 U50 ( .A(A[5]), .Q(n10) );
  NOR21 U51 ( .A(n15), .B(n16), .Q(n14) );
  INV3 U52 ( .A(A[29]), .Q(n16) );
  INV3 U53 ( .A(A[6]), .Q(n7) );
  NAND22 U54 ( .A(A[7]), .B(A[4]), .Q(n84) );
  INV3 U55 ( .A(A[2]), .Q(SUM[2]) );
  INV3 U56 ( .A(n45), .Q(n34) );
  NAND22 U57 ( .A(n46), .B(n47), .Q(n45) );
  NOR31 U58 ( .A(n50), .B(n48), .C(n49), .Q(n47) );
  NAND22 U59 ( .A(A[19]), .B(A[16]), .Q(n48) );
  XNR21 U60 ( .A(A[28]), .B(n19), .Q(SUM[28]) );
  XNR21 U61 ( .A(A[12]), .B(n69), .Q(SUM[12]) );
  XNR21 U62 ( .A(A[16]), .B(n57), .Q(SUM[16]) );
  XNR21 U63 ( .A(A[20]), .B(n45), .Q(SUM[20]) );
  XNR21 U64 ( .A(A[24]), .B(n33), .Q(SUM[24]) );
  XOR21 U65 ( .A(n75), .B(n76), .Q(SUM[11]) );
  INV3 U66 ( .A(A[11]), .Q(n75) );
  NAND22 U67 ( .A(n77), .B(A[10]), .Q(n76) );
  XOR21 U68 ( .A(n64), .B(n65), .Q(SUM[15]) );
  INV3 U69 ( .A(A[15]), .Q(n64) );
  NAND22 U70 ( .A(n66), .B(A[14]), .Q(n65) );
  XOR21 U71 ( .A(n51), .B(n52), .Q(SUM[19]) );
  INV3 U72 ( .A(A[19]), .Q(n51) );
  NAND22 U73 ( .A(n53), .B(A[18]), .Q(n52) );
  XOR21 U74 ( .A(n39), .B(n40), .Q(SUM[23]) );
  INV3 U75 ( .A(A[23]), .Q(n39) );
  NAND22 U76 ( .A(n41), .B(A[22]), .Q(n40) );
  INV3 U77 ( .A(A[17]), .Q(n50) );
  INV3 U78 ( .A(A[21]), .Q(n38) );
  NOR21 U79 ( .A(n3), .B(n79), .Q(n1) );
  INV3 U80 ( .A(A[8]), .Q(n79) );
  INV3 U81 ( .A(A[9]), .Q(n2) );
  INV3 U82 ( .A(A[13]), .Q(n63) );
  INV3 U83 ( .A(A[14]), .Q(n62) );
  NOR21 U84 ( .A(n69), .B(n70), .Q(n68) );
  INV3 U85 ( .A(A[12]), .Q(n70) );
  INV3 U86 ( .A(A[10]), .Q(n74) );
  INV3 U87 ( .A(A[18]), .Q(n49) );
  INV3 U88 ( .A(A[22]), .Q(n37) );
  NOR21 U89 ( .A(n57), .B(n56), .Q(n55) );
  INV3 U90 ( .A(A[16]), .Q(n56) );
  NOR21 U91 ( .A(n45), .B(n44), .Q(n43) );
  INV3 U92 ( .A(A[20]), .Q(n44) );
  NAND22 U93 ( .A(A[23]), .B(A[20]), .Q(n36) );
  NAND22 U94 ( .A(A[27]), .B(A[24]), .Q(n24) );
  NAND22 U95 ( .A(A[15]), .B(A[12]), .Q(n61) );
  XNR21 U96 ( .A(A[4]), .B(n82), .Q(SUM[4]) );
  XNR21 U97 ( .A(A[8]), .B(n3), .Q(SUM[8]) );
  XOR21 U98 ( .A(n4), .B(n5), .Q(SUM[7]) );
  INV3 U99 ( .A(A[7]), .Q(n4) );
  NAND22 U100 ( .A(n6), .B(A[6]), .Q(n5) );
  NOR21 U101 ( .A(n82), .B(n11), .Q(n9) );
  INV3 U102 ( .A(A[4]), .Q(n11) );
  INV3 U103 ( .A(A[25]), .Q(n26) );
  INV3 U104 ( .A(A[26]), .Q(n25) );
  XOR21 U105 ( .A(A[3]), .B(A[2]), .Q(SUM[3]) );
  CLKIN3 U106 ( .A(n18), .Q(n15) );
  CLKIN3 U107 ( .A(n21), .Q(n19) );
  CLKIN3 U108 ( .A(n31), .Q(n30) );
  CLKIN3 U109 ( .A(n43), .Q(n42) );
  CLKIN3 U110 ( .A(n55), .Q(n54) );
  CLKIN3 U111 ( .A(n68), .Q(n67) );
  CLKIN3 U112 ( .A(n60), .Q(n69) );
  CLKIN3 U113 ( .A(n1), .Q(n78) );
  CLKIN3 U114 ( .A(n80), .Q(n3) );
endmodule


module F_add4 ( i_addr_pc, o_addr_pcadd4 );
  input [31:0] i_addr_pc;
  output [31:0] o_addr_pcadd4;
  wire   n2, n1;

  F_add4_DW01_add_1 add_5 ( .A(i_addr_pc), .B({n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, n1, 
        n1, n1, n1, n2, n1, n1}), .CI(n1), .SUM(o_addr_pcadd4) );
  LOGIC0 U3 ( .Q(n1) );
  LOGIC1 U4 ( .Q(n2) );
endmodule


module fetch ( i_clk, i_nrst, i_addr_b, i_addr_j, i_addr_jr, i_con_b, i_con_j, 
        i_data_instr, i_con_ifstall, o_addr_pc, o_addr_pc4, o_data_instr );
  input [31:0] i_addr_b;
  input [31:0] i_addr_j;
  input [31:0] i_addr_jr;
  input [1:0] i_con_j;
  input [31:0] i_data_instr;
  output [31:0] o_addr_pc;
  output [31:0] o_addr_pc4;
  output [31:0] o_data_instr;
  input i_clk, i_nrst, i_con_b, i_con_ifstall;

  wire   [31:0] jmux_i_addr_pc4;
  wire   [31:0] bmux_i_addr_jumpmux;
  wire   [31:0] pc_i_addr_next_pc;

  DFC3 pipe_instr_reg_31_ ( .D(i_data_instr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[31]) );
  DFC3 pipe_instr_reg_30_ ( .D(i_data_instr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[30]) );
  DFC3 pipe_instr_reg_29_ ( .D(i_data_instr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[29]) );
  DFC3 pipe_instr_reg_28_ ( .D(i_data_instr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[28]) );
  DFC3 pipe_instr_reg_27_ ( .D(i_data_instr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[27]) );
  DFC3 pipe_instr_reg_26_ ( .D(i_data_instr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[26]) );
  DFC3 pipe_instr_reg_25_ ( .D(i_data_instr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[25]) );
  DFC3 pipe_instr_reg_24_ ( .D(i_data_instr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[24]) );
  DFC3 pipe_instr_reg_23_ ( .D(i_data_instr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[23]) );
  DFC3 pipe_instr_reg_22_ ( .D(i_data_instr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[22]) );
  DFC3 pipe_instr_reg_21_ ( .D(i_data_instr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[21]) );
  DFC3 pipe_instr_reg_20_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[20]) );
  DFC3 pipe_instr_reg_19_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[19]) );
  DFC3 pipe_instr_reg_18_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[18]) );
  DFC3 pipe_instr_reg_17_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[17]) );
  DFC3 pipe_instr_reg_16_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[16]) );
  DFC3 pipe_instr_reg_15_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[15]) );
  DFC3 pipe_instr_reg_14_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[14]) );
  DFC3 pipe_instr_reg_13_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[13]) );
  DFC3 pipe_instr_reg_12_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[12]) );
  DFC3 pipe_instr_reg_11_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[11]) );
  DFC3 pipe_instr_reg_10_ ( .D(i_data_instr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[10]) );
  DFC3 pipe_instr_reg_9_ ( .D(i_data_instr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[9]) );
  DFC3 pipe_instr_reg_8_ ( .D(i_data_instr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[8]) );
  DFC3 pipe_instr_reg_7_ ( .D(i_data_instr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[7]) );
  DFC3 pipe_instr_reg_6_ ( .D(i_data_instr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[6]) );
  DFC3 pipe_instr_reg_5_ ( .D(i_data_instr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[5]) );
  DFC3 pipe_instr_reg_4_ ( .D(i_data_instr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[4]) );
  DFC3 pipe_instr_reg_3_ ( .D(i_data_instr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[3]) );
  DFC3 pipe_instr_reg_2_ ( .D(i_data_instr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[2]) );
  DFC3 pipe_instr_reg_1_ ( .D(i_data_instr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[1]) );
  DFC3 pipe_instr_reg_0_ ( .D(i_data_instr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_instr[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(jmux_i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(jmux_i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(jmux_i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(jmux_i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(jmux_i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(jmux_i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(jmux_i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(jmux_i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(jmux_i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(jmux_i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(jmux_i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(jmux_i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(jmux_i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(jmux_i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(jmux_i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(jmux_i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(jmux_i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(jmux_i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(jmux_i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(jmux_i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(jmux_i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(jmux_i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(jmux_i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(jmux_i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(jmux_i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(jmux_i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(jmux_i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(jmux_i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(jmux_i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(jmux_i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(jmux_i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(jmux_i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  F_jumpmux u_jumpmux ( .i_addr_j(i_addr_j), .i_addr_jr(i_addr_jr), 
        .i_addr_pc4(jmux_i_addr_pc4), .i_con_jump(i_con_j), .o_addr_jumpmux(
        bmux_i_addr_jumpmux) );
  F_branchmux u_branchmux ( .i_addr_jumpmux(bmux_i_addr_jumpmux), .i_addr_b(
        i_addr_b), .i_con_ifbranch(i_con_b), .o_addr_nextpc(pc_i_addr_next_pc)
         );
  F_pc u_pc ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_con_stall(i_con_ifstall), 
        .i_addr_next_pc(pc_i_addr_next_pc), .o_addr_pc(o_addr_pc) );
  F_add4 u_add4 ( .i_addr_pc(o_addr_pc), .o_addr_pcadd4(jmux_i_addr_pc4) );
endmodule


module D_control ( o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite, 
        o_con_alusrc, o_con_regwrite, o_con_ifsign, o_con_aluop, i_con_instru
 );
  output [5:0] o_con_aluop;
  input [5:0] i_con_instru;
  output o_con_regdst, o_con_memread, o_con_memtoreg, o_con_memwrite,
         o_con_alusrc, o_con_regwrite, o_con_ifsign;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n1, n2, n3, n5, n6, n7, n8, n9, n10;

  OAI212 U2 ( .A(i_con_instru[3]), .B(n11), .C(n12), .Q(o_con_regwrite) );
  OAI212 U3 ( .A(n5), .B(n13), .C(n3), .Q(n12) );
  OAI222 U6 ( .A(i_con_instru[3]), .B(n15), .C(i_con_instru[4]), .D(n17), .Q(
        o_con_memread) );
  OAI212 U23 ( .A(i_con_instru[5]), .B(n20), .C(n14), .Q(o_con_aluop[1]) );
  NAND31 U4 ( .A(n24), .B(n3), .C(n13), .Q(n14) );
  NAND22 U5 ( .A(n9), .B(n13), .Q(n11) );
  AOI211 U7 ( .A(n5), .B(n8), .C(o_con_memwrite), .Q(n18) );
  INV3 U8 ( .A(n20), .Q(n5) );
  INV3 U9 ( .A(n24), .Q(n9) );
  NAND22 U10 ( .A(n20), .B(n15), .Q(o_con_alusrc) );
  NAND22 U11 ( .A(n15), .B(n16), .Q(o_con_memtoreg) );
  NOR21 U12 ( .A(n11), .B(n21), .Q(o_con_aluop[5]) );
  INV3 U13 ( .A(n16), .Q(o_con_memwrite) );
  INV3 U14 ( .A(n21), .Q(n2) );
  NOR31 U15 ( .A(i_con_instru[2]), .B(i_con_instru[4]), .C(n27), .Q(n13) );
  XNR21 U16 ( .A(i_con_instru[1]), .B(n10), .Q(n27) );
  NAND22 U17 ( .A(i_con_instru[0]), .B(i_con_instru[1]), .Q(n24) );
  NAND22 U18 ( .A(i_con_instru[3]), .B(n6), .Q(n20) );
  INV3 U19 ( .A(i_con_instru[4]), .Q(n6) );
  NAND22 U20 ( .A(i_con_instru[5]), .B(n5), .Q(n16) );
  OAI2111 U21 ( .A(n9), .B(n18), .C(n19), .D(n15), .Q(o_con_ifsign) );
  NAND31 U22 ( .A(n9), .B(n5), .C(i_con_instru[2]), .Q(n19) );
  INV3 U24 ( .A(i_con_instru[0]), .Q(n10) );
  NOR21 U25 ( .A(i_con_instru[3]), .B(n14), .Q(o_con_regdst) );
  NAND22 U26 ( .A(i_con_instru[5]), .B(n7), .Q(n15) );
  INV3 U27 ( .A(n11), .Q(n7) );
  NAND22 U28 ( .A(i_con_instru[3]), .B(n3), .Q(n21) );
  NAND31 U29 ( .A(n2), .B(n9), .C(i_con_instru[2]), .Q(n17) );
  NAND31 U30 ( .A(i_con_instru[1]), .B(n10), .C(n2), .Q(n23) );
  INV3 U31 ( .A(i_con_instru[2]), .Q(n8) );
  AOI2111 U32 ( .A(n24), .B(n26), .C(n21), .D(i_con_instru[4]), .Q(
        o_con_aluop[2]) );
  NAND22 U33 ( .A(i_con_instru[2]), .B(n10), .Q(n26) );
  NOR21 U34 ( .A(i_con_instru[4]), .B(n21), .Q(o_con_aluop[0]) );
  AOI211 U35 ( .A(n23), .B(n25), .C(i_con_instru[4]), .Q(o_con_aluop[3]) );
  NAND31 U36 ( .A(n2), .B(i_con_instru[0]), .C(i_con_instru[2]), .Q(n25) );
  AOI211 U37 ( .A(n17), .B(n22), .C(i_con_instru[4]), .Q(o_con_aluop[4]) );
  NAND22 U38 ( .A(n1), .B(n8), .Q(n22) );
  INV3 U39 ( .A(n23), .Q(n1) );
  INV3 U40 ( .A(i_con_instru[5]), .Q(n3) );
endmodule


module D_jb_control ( o_con_jump, o_con_bop, o_con_aluPC4, o_con_ifstall, 
        i_con_instru, i_con_func, i_con_rt );
  output [1:0] o_con_jump;
  output [2:0] o_con_bop;
  input [5:0] i_con_instru;
  input [5:0] i_con_func;
  input i_con_rt;
  output o_con_aluPC4, o_con_ifstall;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n2, n3, n4,
         n5, n6;

  OAI222 U13 ( .A(n5), .B(n16), .C(n14), .D(n17), .Q(o_con_bop[1]) );
  NAND31 U3 ( .A(n5), .B(n3), .C(n6), .Q(n8) );
  NAND22 U4 ( .A(n7), .B(n8), .Q(o_con_jump[1]) );
  INV3 U5 ( .A(n7), .Q(n2) );
  INV3 U6 ( .A(n13), .Q(o_con_ifstall) );
  AOI211 U7 ( .A(n3), .B(n14), .C(n2), .Q(n13) );
  NAND22 U8 ( .A(n7), .B(n4), .Q(n17) );
  OAI311 U9 ( .A(n4), .B(n2), .C(n14), .D(n16), .Q(o_con_bop[0]) );
  OAI2111 U10 ( .A(n9), .B(n8), .C(n10), .D(n7), .Q(o_con_jump[0]) );
  NOR40 U11 ( .A(n11), .B(i_con_func[2]), .C(i_con_func[5]), .D(i_con_func[4]), 
        .Q(n9) );
  NAND22 U12 ( .A(i_con_instru[1]), .B(n3), .Q(n10) );
  NAND22 U14 ( .A(n12), .B(i_con_func[3]), .Q(n11) );
  NOR31 U15 ( .A(i_con_instru[3]), .B(i_con_instru[5]), .C(i_con_instru[4]), 
        .Q(n7) );
  INV3 U16 ( .A(i_con_instru[2]), .Q(n3) );
  INV3 U17 ( .A(i_con_instru[1]), .Q(n5) );
  INV3 U18 ( .A(i_con_instru[0]), .Q(n6) );
  NOR21 U19 ( .A(i_con_func[1]), .B(i_con_func[0]), .Q(n12) );
  NAND22 U20 ( .A(i_con_instru[0]), .B(n5), .Q(n14) );
  NOR40 U21 ( .A(i_con_instru[2]), .B(n2), .C(n5), .D(n6), .Q(o_con_aluPC4) );
  NAND31 U22 ( .A(n7), .B(n6), .C(i_con_instru[2]), .Q(n16) );
  NOR31 U23 ( .A(n15), .B(n2), .C(n6), .Q(o_con_bop[2]) );
  XNR21 U24 ( .A(n5), .B(i_con_instru[2]), .Q(n15) );
  INV3 U25 ( .A(n18), .Q(n4) );
  NOR21 U26 ( .A(i_con_instru[2]), .B(i_con_rt), .Q(n18) );
endmodule


module D_pcadd_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258;

  NAND22 U2 ( .A(n30), .B(n27), .Q(n31) );
  NAND22 U3 ( .A(n204), .B(n214), .Q(n221) );
  NAND22 U4 ( .A(n169), .B(n179), .Q(n188) );
  NAND22 U5 ( .A(n133), .B(n143), .Q(n154) );
  NAND22 U6 ( .A(n100), .B(n108), .Q(n119) );
  NAND22 U7 ( .A(n79), .B(n82), .Q(n89) );
  INV3 U8 ( .A(B[23]), .Q(n6) );
  XOR21 U9 ( .A(n22), .B(n24), .Q(SUM[6]) );
  NOR21 U10 ( .A(n248), .B(n25), .Q(n24) );
  INV3 U11 ( .A(B[30]), .Q(n9) );
  NAND31 U12 ( .A(n230), .B(n231), .C(n232), .Q(n228) );
  NOR21 U13 ( .A(n244), .B(n245), .Q(n231) );
  NOR21 U14 ( .A(n25), .B(n246), .Q(n230) );
  NAND31 U15 ( .A(n71), .B(n72), .C(n73), .Q(n70) );
  NOR21 U16 ( .A(n75), .B(n76), .Q(n72) );
  NOR21 U17 ( .A(n77), .B(n78), .Q(n71) );
  INV3 U18 ( .A(n74), .Q(n73) );
  AOI211 U19 ( .A(n237), .B(n42), .C(n43), .Q(n233) );
  XNR21 U20 ( .A(n89), .B(n88), .Q(SUM[26]) );
  INV3 U21 ( .A(n211), .Q(n210) );
  AOI211 U22 ( .A(n212), .B(n204), .C(n213), .Q(n211) );
  INV3 U23 ( .A(n214), .Q(n213) );
  INV3 U24 ( .A(n176), .Q(n175) );
  AOI211 U25 ( .A(n177), .B(n169), .C(n178), .Q(n176) );
  INV3 U26 ( .A(n179), .Q(n178) );
  INV3 U27 ( .A(n140), .Q(n139) );
  AOI211 U28 ( .A(n141), .B(n133), .C(n142), .Q(n140) );
  INV3 U29 ( .A(n143), .Q(n142) );
  INV3 U30 ( .A(n26), .Q(n248) );
  AOI211 U31 ( .A(n80), .B(n79), .C(n81), .Q(n68) );
  INV3 U32 ( .A(n82), .Q(n81) );
  AOI211 U33 ( .A(n106), .B(n100), .C(n107), .Q(n103) );
  INV3 U34 ( .A(n108), .Q(n107) );
  XNR21 U35 ( .A(n188), .B(n187), .Q(SUM[14]) );
  XNR21 U36 ( .A(n221), .B(n220), .Q(SUM[10]) );
  XOR21 U37 ( .A(n193), .B(n189), .Q(SUM[13]) );
  NAND22 U38 ( .A(n190), .B(n181), .Q(n193) );
  XOR21 U39 ( .A(n158), .B(n155), .Q(SUM[17]) );
  NAND22 U40 ( .A(n156), .B(n145), .Q(n158) );
  XOR21 U41 ( .A(n123), .B(n120), .Q(SUM[21]) );
  NAND22 U42 ( .A(n121), .B(n111), .Q(n123) );
  XOR21 U43 ( .A(n93), .B(n90), .Q(SUM[25]) );
  NAND22 U44 ( .A(n91), .B(n84), .Q(n93) );
  NAND22 U45 ( .A(n144), .B(n160), .Q(n159) );
  NAND22 U46 ( .A(n161), .B(n134), .Q(n160) );
  INV3 U47 ( .A(n162), .Q(n161) );
  XNR21 U48 ( .A(n154), .B(n153), .Q(SUM[18]) );
  XNR21 U49 ( .A(n119), .B(n118), .Q(SUM[22]) );
  INV3 U50 ( .A(n79), .Q(n78) );
  XNR21 U51 ( .A(n31), .B(n29), .Q(SUM[5]) );
  XOR21 U52 ( .A(n10), .B(n11), .Q(SUM[9]) );
  NAND22 U53 ( .A(n12), .B(n13), .Q(n10) );
  NAND22 U54 ( .A(n27), .B(n28), .Q(n22) );
  NAND22 U55 ( .A(n29), .B(n30), .Q(n28) );
  XOR21 U56 ( .A(n41), .B(n54), .Q(SUM[2]) );
  NOR21 U57 ( .A(n43), .B(n55), .Q(n54) );
  XNR21 U58 ( .A(n58), .B(n149), .Q(SUM[1]) );
  NAND22 U59 ( .A(n59), .B(n56), .Q(n149) );
  INV3 U60 ( .A(n144), .Q(n184) );
  NAND22 U61 ( .A(n56), .B(n57), .Q(n41) );
  NAND22 U62 ( .A(n58), .B(n59), .Q(n57) );
  INV3 U63 ( .A(n150), .Q(n58) );
  AOI311 U64 ( .A(n99), .B(n100), .C(n101), .D(n102), .Q(n74) );
  NOR31 U65 ( .A(n109), .B(n112), .C(n113), .Q(n99) );
  NOR21 U66 ( .A(B[20]), .B(A[20]), .Q(n112) );
  OAI2111 U67 ( .A(n226), .B(n227), .C(n228), .D(n229), .Q(n205) );
  NOR21 U68 ( .A(A[7]), .B(B[7]), .Q(n227) );
  NAND22 U69 ( .A(B[7]), .B(A[7]), .Q(n229) );
  AOI211 U70 ( .A(n247), .B(n23), .C(n248), .Q(n226) );
  NAND22 U71 ( .A(B[29]), .B(A[29]), .Q(n53) );
  NOR21 U72 ( .A(A[29]), .B(B[29]), .Q(n52) );
  NAND22 U73 ( .A(n253), .B(n254), .Q(n204) );
  INV3 U74 ( .A(A[10]), .Q(n254) );
  INV3 U75 ( .A(B[10]), .Q(n253) );
  NOR21 U76 ( .A(n66), .B(n67), .Q(n62) );
  INV3 U77 ( .A(n85), .Q(n66) );
  NAND22 U78 ( .A(B[27]), .B(A[27]), .Q(n85) );
  NAND22 U79 ( .A(B[2]), .B(A[2]), .Q(n238) );
  NAND22 U80 ( .A(B[10]), .B(A[10]), .Q(n214) );
  XOR21 U81 ( .A(n44), .B(n45), .Q(SUM[31]) );
  XNR21 U82 ( .A(B[31]), .B(A[31]), .Q(n44) );
  AOI211 U83 ( .A(n46), .B(n47), .C(n48), .Q(n45) );
  NOR21 U84 ( .A(n49), .B(n9), .Q(n48) );
  XOR21 U85 ( .A(n86), .B(n87), .Q(SUM[27]) );
  XNR21 U86 ( .A(B[27]), .B(A[27]), .Q(n86) );
  AOI211 U87 ( .A(n88), .B(n79), .C(n81), .Q(n87) );
  XOR21 U88 ( .A(n116), .B(n117), .Q(SUM[23]) );
  XNR21 U89 ( .A(B[23]), .B(A[23]), .Q(n116) );
  AOI211 U90 ( .A(n118), .B(n100), .C(n107), .Q(n117) );
  NAND22 U91 ( .A(n130), .B(n131), .Q(n101) );
  AOI221 U92 ( .A(A[19]), .B(B[19]), .C(n138), .D(n139), .Q(n130) );
  NAND31 U93 ( .A(n132), .B(n133), .C(n134), .Q(n131) );
  INV3 U94 ( .A(n146), .Q(n138) );
  NAND22 U95 ( .A(n166), .B(n167), .Q(n134) );
  AOI221 U96 ( .A(A[15]), .B(B[15]), .C(n174), .D(n175), .Q(n166) );
  NAND31 U97 ( .A(n168), .B(n169), .C(n170), .Q(n167) );
  INV3 U98 ( .A(n182), .Q(n174) );
  NAND22 U99 ( .A(B[5]), .B(A[5]), .Q(n27) );
  NAND22 U100 ( .A(B[4]), .B(A[4]), .Q(n34) );
  NAND22 U101 ( .A(B[8]), .B(A[8]), .Q(n19) );
  NAND22 U102 ( .A(B[12]), .B(A[12]), .Q(n180) );
  NOR21 U103 ( .A(A[24]), .B(B[24]), .Q(n95) );
  NOR21 U104 ( .A(B[4]), .B(A[4]), .Q(n244) );
  NAND22 U105 ( .A(B[9]), .B(A[9]), .Q(n13) );
  NAND22 U106 ( .A(B[17]), .B(A[17]), .Q(n145) );
  NAND22 U107 ( .A(n249), .B(n250), .Q(n23) );
  INV3 U108 ( .A(A[6]), .Q(n250) );
  INV3 U109 ( .A(B[6]), .Q(n249) );
  NOR21 U110 ( .A(A[20]), .B(B[20]), .Q(n126) );
  NAND22 U111 ( .A(B[28]), .B(A[28]), .Q(n64) );
  NOR21 U112 ( .A(A[28]), .B(B[28]), .Q(n63) );
  NOR21 U113 ( .A(B[7]), .B(A[7]), .Q(n245) );
  NAND22 U114 ( .A(B[6]), .B(A[6]), .Q(n26) );
  NAND22 U115 ( .A(n201), .B(n202), .Q(n170) );
  AOI221 U116 ( .A(A[11]), .B(B[11]), .C(n209), .D(n210), .Q(n201) );
  NAND31 U117 ( .A(n203), .B(n204), .C(n205), .Q(n202) );
  INV3 U118 ( .A(n215), .Q(n209) );
  INV3 U119 ( .A(n232), .Q(n32) );
  INV3 U120 ( .A(A[3]), .Q(n235) );
  INV3 U121 ( .A(B[3]), .Q(n236) );
  NOR31 U122 ( .A(n135), .B(n136), .C(n137), .Q(n132) );
  NOR21 U123 ( .A(B[16]), .B(A[16]), .Q(n136) );
  NOR21 U124 ( .A(B[19]), .B(A[19]), .Q(n137) );
  NOR31 U125 ( .A(n206), .B(n207), .C(n208), .Q(n203) );
  NOR21 U126 ( .A(B[11]), .B(A[11]), .Q(n207) );
  NOR21 U127 ( .A(B[8]), .B(A[8]), .Q(n208) );
  NAND22 U128 ( .A(n222), .B(n223), .Q(n12) );
  INV3 U129 ( .A(A[9]), .Q(n223) );
  INV3 U130 ( .A(B[9]), .Q(n222) );
  NAND22 U131 ( .A(n197), .B(n198), .Q(n190) );
  INV3 U132 ( .A(A[13]), .Q(n198) );
  INV3 U133 ( .A(B[13]), .Q(n197) );
  XOR21 U134 ( .A(n65), .B(n62), .Q(SUM[28]) );
  XNR21 U135 ( .A(B[28]), .B(A[28]), .Q(n65) );
  XOR21 U136 ( .A(n60), .B(n51), .Q(SUM[29]) );
  XNR21 U137 ( .A(B[29]), .B(A[29]), .Q(n60) );
  XOR21 U138 ( .A(n1), .B(n47), .Q(SUM[30]) );
  XOR21 U139 ( .A(B[30]), .B(A[30]), .Q(n1) );
  NOR21 U140 ( .A(A[3]), .B(B[3]), .Q(n234) );
  NAND22 U141 ( .A(n251), .B(n252), .Q(n30) );
  INV3 U142 ( .A(A[5]), .Q(n252) );
  INV3 U143 ( .A(B[5]), .Q(n251) );
  NAND22 U144 ( .A(n2), .B(n163), .Q(n156) );
  INV3 U145 ( .A(A[17]), .Q(n163) );
  INV3 U146 ( .A(B[17]), .Q(n2) );
  NAND22 U147 ( .A(n191), .B(n192), .Q(n169) );
  INV3 U148 ( .A(A[14]), .Q(n192) );
  INV3 U149 ( .A(B[14]), .Q(n191) );
  NAND22 U150 ( .A(B[16]), .B(A[16]), .Q(n144) );
  NAND22 U151 ( .A(B[14]), .B(A[14]), .Q(n179) );
  NAND22 U152 ( .A(B[18]), .B(A[18]), .Q(n143) );
  NAND22 U153 ( .A(B[22]), .B(A[22]), .Q(n108) );
  NAND22 U154 ( .A(B[26]), .B(A[26]), .Q(n82) );
  XOR21 U155 ( .A(n185), .B(n186), .Q(SUM[15]) );
  XNR21 U156 ( .A(B[15]), .B(A[15]), .Q(n185) );
  AOI211 U157 ( .A(n187), .B(n169), .C(n178), .Q(n186) );
  XOR21 U158 ( .A(n151), .B(n152), .Q(SUM[19]) );
  XNR21 U159 ( .A(B[19]), .B(A[19]), .Q(n151) );
  AOI211 U160 ( .A(n153), .B(n133), .C(n142), .Q(n152) );
  NAND22 U161 ( .A(B[20]), .B(A[20]), .Q(n110) );
  NAND22 U162 ( .A(B[24]), .B(A[24]), .Q(n83) );
  NAND22 U163 ( .A(B[13]), .B(A[13]), .Q(n181) );
  NAND22 U164 ( .A(B[21]), .B(A[21]), .Q(n111) );
  NAND22 U165 ( .A(B[25]), .B(A[25]), .Q(n84) );
  NOR21 U166 ( .A(A[8]), .B(B[8]), .Q(n225) );
  NOR21 U167 ( .A(A[12]), .B(B[12]), .Q(n196) );
  NOR31 U168 ( .A(n171), .B(n172), .C(n173), .Q(n168) );
  NOR21 U169 ( .A(B[15]), .B(A[15]), .Q(n173) );
  NOR21 U170 ( .A(B[12]), .B(A[12]), .Q(n172) );
  NAND22 U171 ( .A(n4), .B(n127), .Q(n121) );
  INV3 U172 ( .A(A[21]), .Q(n127) );
  INV3 U173 ( .A(B[21]), .Q(n4) );
  XOR21 U174 ( .A(n218), .B(n219), .Q(SUM[11]) );
  XNR21 U175 ( .A(B[11]), .B(A[11]), .Q(n218) );
  AOI211 U176 ( .A(n220), .B(n204), .C(n213), .Q(n219) );
  NOR21 U177 ( .A(B[23]), .B(A[23]), .Q(n113) );
  NOR21 U178 ( .A(A[15]), .B(B[15]), .Q(n182) );
  NOR21 U179 ( .A(A[11]), .B(B[11]), .Q(n215) );
  NOR21 U180 ( .A(A[19]), .B(B[19]), .Q(n146) );
  NOR21 U181 ( .A(A[23]), .B(B[23]), .Q(n104) );
  IMUX21 U182 ( .A(n97), .B(n98), .S(n74), .Q(SUM[24]) );
  XNR21 U183 ( .A(B[24]), .B(A[24]), .Q(n98) );
  NOR21 U184 ( .A(n114), .B(n115), .Q(n97) );
  NOR21 U185 ( .A(B[24]), .B(A[24]), .Q(n114) );
  IMUX21 U186 ( .A(n128), .B(n129), .S(n125), .Q(SUM[20]) );
  XNR21 U187 ( .A(B[20]), .B(A[20]), .Q(n129) );
  NOR21 U188 ( .A(n147), .B(n148), .Q(n128) );
  NOR21 U189 ( .A(B[20]), .B(A[20]), .Q(n147) );
  NAND22 U190 ( .A(n5), .B(n122), .Q(n100) );
  INV3 U191 ( .A(A[22]), .Q(n122) );
  INV3 U192 ( .A(B[22]), .Q(n5) );
  NAND22 U193 ( .A(n8), .B(n92), .Q(n79) );
  INV3 U194 ( .A(A[26]), .Q(n92) );
  INV3 U195 ( .A(B[26]), .Q(n8) );
  NAND22 U196 ( .A(n3), .B(n157), .Q(n133) );
  INV3 U197 ( .A(A[18]), .Q(n157) );
  INV3 U198 ( .A(B[18]), .Q(n3) );
  NAND22 U199 ( .A(n7), .B(n96), .Q(n91) );
  INV3 U200 ( .A(A[25]), .Q(n96) );
  INV3 U201 ( .A(B[25]), .Q(n7) );
  NOR21 U202 ( .A(A[4]), .B(B[4]), .Q(n33) );
  NOR21 U203 ( .A(A[16]), .B(B[16]), .Q(n162) );
  NOR21 U204 ( .A(B[24]), .B(A[24]), .Q(n75) );
  XOR21 U205 ( .A(n20), .B(n21), .Q(SUM[7]) );
  XNR21 U206 ( .A(B[7]), .B(A[7]), .Q(n20) );
  AOI211 U207 ( .A(n22), .B(n23), .C(n248), .Q(n21) );
  NOR21 U208 ( .A(B[27]), .B(A[27]), .Q(n76) );
  NOR21 U209 ( .A(A[27]), .B(B[27]), .Q(n69) );
  IMUX21 U210 ( .A(n164), .B(n165), .S(n134), .Q(SUM[16]) );
  NOR21 U211 ( .A(n183), .B(n184), .Q(n165) );
  XNR21 U212 ( .A(B[16]), .B(A[16]), .Q(n164) );
  NOR21 U213 ( .A(B[16]), .B(A[16]), .Q(n183) );
  IMUX21 U214 ( .A(n14), .B(n15), .S(n16), .Q(SUM[8]) );
  NOR21 U215 ( .A(n17), .B(n18), .Q(n14) );
  XNR21 U216 ( .A(B[8]), .B(A[8]), .Q(n15) );
  NOR21 U217 ( .A(B[8]), .B(A[8]), .Q(n17) );
  IMUX21 U218 ( .A(n199), .B(n200), .S(n195), .Q(SUM[12]) );
  NOR21 U219 ( .A(n216), .B(n217), .Q(n199) );
  XNR21 U220 ( .A(B[12]), .B(A[12]), .Q(n200) );
  NOR21 U221 ( .A(B[12]), .B(A[12]), .Q(n216) );
  INV3 U222 ( .A(A[23]), .Q(n105) );
  INV3 U223 ( .A(n50), .Q(n46) );
  NOR21 U224 ( .A(A[30]), .B(B[30]), .Q(n50) );
  NAND22 U225 ( .A(n242), .B(n243), .Q(n42) );
  INV3 U226 ( .A(A[2]), .Q(n243) );
  INV3 U227 ( .A(B[2]), .Q(n242) );
  XOR21 U228 ( .A(n39), .B(n40), .Q(SUM[3]) );
  XNR21 U229 ( .A(B[3]), .B(A[3]), .Q(n39) );
  AOI211 U230 ( .A(n41), .B(n42), .C(n43), .Q(n40) );
  IMUX21 U231 ( .A(n35), .B(n36), .S(n32), .Q(SUM[4]) );
  NOR21 U232 ( .A(n37), .B(n38), .Q(n35) );
  XNR21 U233 ( .A(B[4]), .B(A[4]), .Q(n36) );
  NOR21 U234 ( .A(B[4]), .B(A[4]), .Q(n37) );
  INV3 U235 ( .A(B[0]), .Q(n255) );
  INV3 U236 ( .A(n257), .Q(n256) );
  NOR21 U237 ( .A(B[0]), .B(n258), .Q(n257) );
  INV3 U238 ( .A(A[30]), .Q(n49) );
  INV3 U239 ( .A(A[0]), .Q(n258) );
  NAND22 U240 ( .A(n240), .B(n241), .Q(n59) );
  INV3 U241 ( .A(B[1]), .Q(n240) );
  INV3 U242 ( .A(A[1]), .Q(n241) );
  NAND22 U243 ( .A(B[1]), .B(A[1]), .Q(n56) );
  NAND22 U244 ( .A(B[0]), .B(A[0]), .Q(n150) );
  CLKIN3 U245 ( .A(n19), .Q(n18) );
  OAI212 U246 ( .A(n32), .B(n33), .C(n34), .Q(n29) );
  CLKIN3 U247 ( .A(n34), .Q(n38) );
  OAI212 U248 ( .A(n51), .B(n52), .C(n53), .Q(n47) );
  CLKIN3 U249 ( .A(n42), .Q(n55) );
  CLKIN3 U250 ( .A(n61), .Q(n51) );
  OAI212 U251 ( .A(n62), .B(n63), .C(n64), .Q(n61) );
  OAI212 U252 ( .A(n68), .B(n69), .C(n70), .Q(n67) );
  OAI212 U253 ( .A(n77), .B(n83), .C(n84), .Q(n80) );
  OAI212 U254 ( .A(n77), .B(n90), .C(n84), .Q(n88) );
  CLKIN3 U255 ( .A(n91), .Q(n77) );
  CLKIN3 U256 ( .A(n94), .Q(n90) );
  OAI212 U257 ( .A(n74), .B(n95), .C(n83), .Q(n94) );
  OAI222 U258 ( .A(n103), .B(n104), .C(n6), .D(n105), .Q(n102) );
  OAI212 U259 ( .A(n109), .B(n110), .C(n111), .Q(n106) );
  CLKIN3 U260 ( .A(n83), .Q(n115) );
  OAI212 U261 ( .A(n109), .B(n120), .C(n111), .Q(n118) );
  CLKIN3 U262 ( .A(n121), .Q(n109) );
  CLKIN3 U263 ( .A(n124), .Q(n120) );
  OAI212 U264 ( .A(n125), .B(n126), .C(n110), .Q(n124) );
  CLKIN3 U265 ( .A(n101), .Q(n125) );
  OAI212 U266 ( .A(n135), .B(n144), .C(n145), .Q(n141) );
  CLKIN3 U267 ( .A(n110), .Q(n148) );
  OAI212 U268 ( .A(n135), .B(n155), .C(n145), .Q(n153) );
  CLKIN3 U269 ( .A(n156), .Q(n135) );
  CLKIN3 U270 ( .A(n159), .Q(n155) );
  OAI212 U271 ( .A(n171), .B(n180), .C(n181), .Q(n177) );
  OAI212 U272 ( .A(n171), .B(n189), .C(n181), .Q(n187) );
  CLKIN3 U273 ( .A(n190), .Q(n171) );
  CLKIN3 U274 ( .A(n194), .Q(n189) );
  OAI212 U275 ( .A(n195), .B(n196), .C(n180), .Q(n194) );
  CLKIN3 U276 ( .A(n170), .Q(n195) );
  OAI212 U277 ( .A(n206), .B(n19), .C(n13), .Q(n212) );
  CLKIN3 U278 ( .A(n180), .Q(n217) );
  OAI212 U279 ( .A(n11), .B(n206), .C(n13), .Q(n220) );
  CLKIN3 U280 ( .A(n12), .Q(n206) );
  CLKIN3 U281 ( .A(n224), .Q(n11) );
  OAI212 U282 ( .A(n16), .B(n225), .C(n19), .Q(n224) );
  CLKIN3 U283 ( .A(n205), .Q(n16) );
  OAI222 U284 ( .A(n233), .B(n234), .C(n235), .D(n236), .Q(n232) );
  CLKIN3 U285 ( .A(n238), .Q(n43) );
  OAI212 U286 ( .A(n239), .B(n150), .C(n56), .Q(n237) );
  CLKIN3 U287 ( .A(n59), .Q(n239) );
  CLKIN3 U288 ( .A(n23), .Q(n25) );
  OAI212 U289 ( .A(n246), .B(n34), .C(n27), .Q(n247) );
  CLKIN3 U290 ( .A(n30), .Q(n246) );
  OAI212 U291 ( .A(A[0]), .B(n255), .C(n256), .Q(SUM[0]) );
endmodule


module D_pcadd ( i_addr_pcadd4E, i_data_immshiftl, o_addr_pcbranchE );
  input [31:0] i_addr_pcadd4E;
  input [31:0] i_data_immshiftl;
  output [31:0] o_addr_pcbranchE;
  wire   n1;

  D_pcadd_DW01_add_1 add_5 ( .A(i_addr_pcadd4E), .B(i_data_immshiftl), .CI(n1), 
        .SUM(o_addr_pcbranchE) );
  LOGIC0 U1 ( .Q(n1) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_addr_Rt, i_con_RegWr, 
        i_addr_Rd, i_data_Rd, o_data_Rs, o_data_Rt );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rt;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr;
  wire   n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777;
  wire   [1023:0] regs;

  DFEC1 regs_reg_15__31_ ( .D(i_data_Rd[31]), .E(n757), .C(i_clk), .RN(n735), 
        .Q(regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(i_data_Rd[30]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(i_data_Rd[29]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(i_data_Rd[28]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[508]) );
  DFEC1 regs_reg_14__31_ ( .D(i_data_Rd[31]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(i_data_Rd[30]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(i_data_Rd[29]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(i_data_Rd[28]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[476]) );
  DFEC1 regs_reg_13__31_ ( .D(i_data_Rd[31]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(i_data_Rd[30]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(i_data_Rd[29]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(i_data_Rd[28]), .E(n759), .C(i_clk), .RN(n732), 
        .Q(regs[444]) );
  DFEC1 regs_reg_12__31_ ( .D(i_data_Rd[31]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(i_data_Rd[30]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(i_data_Rd[29]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(i_data_Rd[28]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[412]) );
  DFEC1 regs_reg_11__31_ ( .D(i_data_Rd[31]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(i_data_Rd[30]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(i_data_Rd[29]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(i_data_Rd[28]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[380]) );
  DFEC1 regs_reg_10__31_ ( .D(i_data_Rd[31]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(i_data_Rd[30]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(i_data_Rd[29]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(i_data_Rd[28]), .E(n762), .C(i_clk), .RN(n733), 
        .Q(regs[348]) );
  DFEC1 regs_reg_9__31_ ( .D(i_data_Rd[31]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(i_data_Rd[30]), .E(n763), .C(i_clk), .RN(n737), 
        .Q(regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(i_data_Rd[29]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(i_data_Rd[28]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[316]) );
  DFEC1 regs_reg_8__31_ ( .D(i_data_Rd[31]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(i_data_Rd[30]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(i_data_Rd[29]), .E(n764), .C(i_clk), .RN(n732), 
        .Q(regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(i_data_Rd[28]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[284]) );
  DFEC1 regs_reg_7__31_ ( .D(i_data_Rd[31]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(i_data_Rd[30]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(i_data_Rd[29]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(i_data_Rd[28]), .E(n765), .C(i_clk), .RN(n734), 
        .Q(regs[252]) );
  DFEC1 regs_reg_6__31_ ( .D(i_data_Rd[31]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(i_data_Rd[30]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(i_data_Rd[29]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(i_data_Rd[28]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[220]) );
  DFEC1 regs_reg_5__31_ ( .D(i_data_Rd[31]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(i_data_Rd[30]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(i_data_Rd[29]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(i_data_Rd[28]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[188]) );
  DFEC1 regs_reg_4__31_ ( .D(i_data_Rd[31]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(i_data_Rd[30]), .E(n768), .C(i_clk), .RN(n737), 
        .Q(regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(i_data_Rd[29]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(i_data_Rd[28]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[156]) );
  DFEC1 regs_reg_3__31_ ( .D(i_data_Rd[31]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(i_data_Rd[30]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(i_data_Rd[29]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(i_data_Rd[28]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[124]) );
  DFEC1 regs_reg_2__31_ ( .D(i_data_Rd[31]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(i_data_Rd[30]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(i_data_Rd[29]), .E(n770), .C(i_clk), .RN(n731), 
        .Q(regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(i_data_Rd[28]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[92]) );
  DFEC1 regs_reg_1__31_ ( .D(i_data_Rd[31]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(i_data_Rd[30]), .E(n771), .C(i_clk), .RN(n737), 
        .Q(regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(i_data_Rd[29]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(i_data_Rd[28]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[60]) );
  DFEC1 regs_reg_0__31_ ( .D(i_data_Rd[31]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(i_data_Rd[30]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(i_data_Rd[29]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(i_data_Rd[28]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[28]) );
  DFEC1 regs_reg_15__27_ ( .D(i_data_Rd[27]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(i_data_Rd[26]), .E(n757), .C(i_clk), .RN(n732), 
        .Q(regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(i_data_Rd[25]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(i_data_Rd[24]), .E(n757), .C(i_clk), .RN(n737), 
        .Q(regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(i_data_Rd[23]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(i_data_Rd[22]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(i_data_Rd[21]), .E(n757), .C(i_clk), .RN(n736), 
        .Q(regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(i_data_Rd[20]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(i_data_Rd[19]), .E(n757), .C(i_clk), .RN(n734), 
        .Q(regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(i_data_Rd[18]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(i_data_Rd[17]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(i_data_Rd[16]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(i_data_Rd[15]), .E(n757), .C(i_clk), .RN(n736), 
        .Q(regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(i_data_Rd[13]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(i_data_Rd[12]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(i_data_Rd[11]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n757), .C(i_clk), .RN(i_rst_n), .Q(regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(i_data_Rd[9]), .E(n757), .C(i_clk), .RN(n734), 
        .Q(regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(i_data_Rd[8]), .E(n757), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(i_data_Rd[7]), .E(n757), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(i_data_Rd[6]), .E(n757), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(i_data_Rd[5]), .E(n757), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(i_data_Rd[4]), .E(n757), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(i_data_Rd[3]), .E(n757), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(i_data_Rd[2]), .E(n757), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(i_data_Rd[1]), .E(n757), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(i_data_Rd[0]), .E(n757), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[480]) );
  DFEC1 regs_reg_14__27_ ( .D(i_data_Rd[27]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(i_data_Rd[26]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(i_data_Rd[25]), .E(n758), .C(i_clk), .RN(n737), 
        .Q(regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(i_data_Rd[24]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(i_data_Rd[23]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(i_data_Rd[22]), .E(n758), .C(i_clk), .RN(n733), 
        .Q(regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(i_data_Rd[21]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(i_data_Rd[20]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(i_data_Rd[19]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(i_data_Rd[18]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(i_data_Rd[17]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(i_data_Rd[16]), .E(n758), .C(i_clk), .RN(n738), 
        .Q(regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(i_data_Rd[15]), .E(n758), .C(i_clk), .RN(n733), 
        .Q(regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n758), .C(i_clk), .RN(n734), 
        .Q(regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(i_data_Rd[13]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(i_data_Rd[12]), .E(n758), .C(i_clk), .RN(n734), 
        .Q(regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(i_data_Rd[11]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n758), .C(i_clk), .RN(i_rst_n), .Q(regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(i_data_Rd[9]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(i_data_Rd[8]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(i_data_Rd[7]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(i_data_Rd[6]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(i_data_Rd[5]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(i_data_Rd[4]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(i_data_Rd[3]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(i_data_Rd[2]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(i_data_Rd[1]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(i_data_Rd[0]), .E(n758), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[448]) );
  DFEC1 regs_reg_13__27_ ( .D(i_data_Rd[27]), .E(n759), .C(i_clk), .RN(n733), 
        .Q(regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(i_data_Rd[26]), .E(n759), .C(i_clk), .RN(n734), 
        .Q(regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(i_data_Rd[25]), .E(n759), .C(i_clk), .RN(n735), 
        .Q(regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(i_data_Rd[24]), .E(n759), .C(i_clk), .RN(n736), 
        .Q(regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(i_data_Rd[23]), .E(n759), .C(i_clk), .RN(n737), 
        .Q(regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(i_data_Rd[22]), .E(n759), .C(i_clk), .RN(n735), 
        .Q(regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(i_data_Rd[21]), .E(n759), .C(i_clk), .RN(n733), 
        .Q(regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(i_data_Rd[20]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(i_data_Rd[19]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(i_data_Rd[18]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(i_data_Rd[17]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(i_data_Rd[16]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(i_data_Rd[15]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(i_data_Rd[13]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(i_data_Rd[12]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(i_data_Rd[11]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n759), .C(i_clk), .RN(i_rst_n), .Q(regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(i_data_Rd[9]), .E(n759), .C(i_clk), .RN(n739), 
        .Q(regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(i_data_Rd[8]), .E(n759), .C(i_clk), .RN(n738), 
        .Q(regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(i_data_Rd[7]), .E(n759), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(i_data_Rd[6]), .E(n759), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(i_data_Rd[5]), .E(n759), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(i_data_Rd[4]), .E(n759), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(i_data_Rd[3]), .E(n759), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(i_data_Rd[2]), .E(n759), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(i_data_Rd[1]), .E(n759), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(i_data_Rd[0]), .E(n759), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[416]) );
  DFEC1 regs_reg_12__27_ ( .D(i_data_Rd[27]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(i_data_Rd[26]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(i_data_Rd[25]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(i_data_Rd[24]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(i_data_Rd[23]), .E(n760), .C(i_clk), .RN(n737), 
        .Q(regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(i_data_Rd[22]), .E(n760), .C(i_clk), .RN(n735), 
        .Q(regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(i_data_Rd[21]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(i_data_Rd[20]), .E(n760), .C(i_clk), .RN(n734), 
        .Q(regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(i_data_Rd[19]), .E(n760), .C(i_clk), .RN(n735), 
        .Q(regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(i_data_Rd[18]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(i_data_Rd[17]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(i_data_Rd[16]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(i_data_Rd[15]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(i_data_Rd[13]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(i_data_Rd[12]), .E(n760), .C(i_clk), .RN(n738), 
        .Q(regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(i_data_Rd[11]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n760), .C(i_clk), .RN(i_rst_n), .Q(regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(i_data_Rd[9]), .E(n760), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(i_data_Rd[8]), .E(n760), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(i_data_Rd[7]), .E(n760), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(i_data_Rd[6]), .E(n760), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(i_data_Rd[5]), .E(n760), .C(i_clk), .RN(n739), 
        .Q(regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(i_data_Rd[4]), .E(n760), .C(i_clk), .RN(n735), 
        .Q(regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(i_data_Rd[3]), .E(n760), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(i_data_Rd[2]), .E(n760), .C(i_clk), .RN(n738), 
        .Q(regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(i_data_Rd[1]), .E(n760), .C(i_clk), .RN(n732), 
        .Q(regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(i_data_Rd[0]), .E(n760), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[384]) );
  DFEC1 regs_reg_11__27_ ( .D(i_data_Rd[27]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(i_data_Rd[26]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(i_data_Rd[25]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(i_data_Rd[24]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(i_data_Rd[23]), .E(n761), .C(i_clk), .RN(n737), 
        .Q(regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(i_data_Rd[22]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(i_data_Rd[21]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(i_data_Rd[20]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(i_data_Rd[19]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(i_data_Rd[18]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(i_data_Rd[17]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(i_data_Rd[16]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(i_data_Rd[15]), .E(n761), .C(i_clk), .RN(n731), 
        .Q(regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(i_data_Rd[13]), .E(n761), .C(i_clk), .RN(n732), 
        .Q(regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(i_data_Rd[12]), .E(n761), .C(i_clk), .RN(n739), 
        .Q(regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(i_data_Rd[11]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(i_data_Rd[10]), .E(n761), .C(i_clk), .RN(i_rst_n), .Q(regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(i_data_Rd[9]), .E(n761), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(i_data_Rd[8]), .E(n761), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(i_data_Rd[7]), .E(n761), .C(i_clk), .RN(n733), 
        .Q(regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(i_data_Rd[6]), .E(n761), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(i_data_Rd[5]), .E(n761), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(i_data_Rd[4]), .E(n761), .C(i_clk), .RN(n736), 
        .Q(regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(i_data_Rd[3]), .E(n761), .C(i_clk), .RN(n734), 
        .Q(regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(i_data_Rd[2]), .E(n761), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(i_data_Rd[1]), .E(n761), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(i_data_Rd[0]), .E(n761), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[352]) );
  DFEC1 regs_reg_10__27_ ( .D(i_data_Rd[27]), .E(n762), .C(i_clk), .RN(n734), 
        .Q(regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(i_data_Rd[26]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(i_data_Rd[25]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(i_data_Rd[24]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(i_data_Rd[23]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(i_data_Rd[22]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(i_data_Rd[21]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(i_data_Rd[20]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(i_data_Rd[19]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(i_data_Rd[18]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(i_data_Rd[17]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(i_data_Rd[16]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(i_data_Rd[15]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(i_data_Rd[13]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(i_data_Rd[12]), .E(n762), .C(i_clk), .RN(n735), 
        .Q(regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(i_data_Rd[11]), .E(n762), .C(i_clk), .RN(i_rst_n), .Q(regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n762), .C(i_clk), .RN(n731), 
        .Q(regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(i_data_Rd[9]), .E(n762), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(i_data_Rd[8]), .E(n762), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(i_data_Rd[7]), .E(n762), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(i_data_Rd[6]), .E(n762), .C(i_clk), .RN(n739), 
        .Q(regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(i_data_Rd[5]), .E(n762), .C(i_clk), .RN(n738), 
        .Q(regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(i_data_Rd[4]), .E(n762), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(i_data_Rd[3]), .E(n762), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(i_data_Rd[2]), .E(n762), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(i_data_Rd[1]), .E(n762), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(i_data_Rd[0]), .E(n762), .C(i_clk), .RN(n731), 
        .Q(regs[320]) );
  DFEC1 regs_reg_9__27_ ( .D(i_data_Rd[27]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(i_data_Rd[26]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(i_data_Rd[25]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(i_data_Rd[24]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(i_data_Rd[23]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(i_data_Rd[22]), .E(n763), .C(i_clk), .RN(n734), 
        .Q(regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(i_data_Rd[21]), .E(n763), .C(i_clk), .RN(n732), 
        .Q(regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(i_data_Rd[20]), .E(n763), .C(i_clk), .RN(n733), 
        .Q(regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(i_data_Rd[19]), .E(n763), .C(i_clk), .RN(n731), 
        .Q(regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(i_data_Rd[18]), .E(n763), .C(i_clk), .RN(n732), 
        .Q(regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(i_data_Rd[17]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(i_data_Rd[16]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(i_data_Rd[15]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(i_data_Rd[14]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(i_data_Rd[13]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(i_data_Rd[12]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(i_data_Rd[11]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(i_data_Rd[10]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(i_data_Rd[9]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(i_data_Rd[8]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(i_data_Rd[7]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(i_data_Rd[6]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(i_data_Rd[5]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(i_data_Rd[4]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(i_data_Rd[3]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(i_data_Rd[2]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(i_data_Rd[1]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(i_data_Rd[0]), .E(n763), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[288]) );
  DFEC1 regs_reg_8__27_ ( .D(i_data_Rd[27]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(i_data_Rd[26]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(i_data_Rd[25]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(i_data_Rd[24]), .E(n764), .C(i_clk), .RN(n736), 
        .Q(regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(i_data_Rd[23]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(i_data_Rd[22]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(i_data_Rd[21]), .E(n764), .C(i_clk), .RN(n731), 
        .Q(regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(i_data_Rd[20]), .E(n764), .C(i_clk), .RN(n731), 
        .Q(regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(i_data_Rd[19]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(i_data_Rd[18]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(i_data_Rd[17]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(i_data_Rd[16]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(i_data_Rd[15]), .E(n764), .C(i_clk), .RN(n731), 
        .Q(regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(i_data_Rd[14]), .E(n764), .C(i_clk), .RN(n733), 
        .Q(regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(i_data_Rd[13]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(i_data_Rd[12]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(i_data_Rd[11]), .E(n764), .C(i_clk), .RN(n739), 
        .Q(regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(i_data_Rd[10]), .E(n764), .C(i_clk), .RN(n736), 
        .Q(regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(i_data_Rd[9]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(i_data_Rd[8]), .E(n764), .C(i_clk), .RN(n732), .Q(
        regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(i_data_Rd[7]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(i_data_Rd[6]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(i_data_Rd[5]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(i_data_Rd[4]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(i_data_Rd[3]), .E(n764), .C(i_clk), .RN(n731), .Q(
        regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(i_data_Rd[2]), .E(n764), .C(i_clk), .RN(n738), .Q(
        regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(i_data_Rd[1]), .E(n764), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(i_data_Rd[0]), .E(n764), .C(i_clk), .RN(n738), .Q(
        regs[256]) );
  DFEC1 regs_reg_7__27_ ( .D(i_data_Rd[27]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(i_data_Rd[26]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(i_data_Rd[25]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(i_data_Rd[24]), .E(n765), .C(i_clk), .RN(n739), 
        .Q(regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(i_data_Rd[23]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(i_data_Rd[22]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(i_data_Rd[21]), .E(n765), .C(i_clk), .RN(n737), 
        .Q(regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(i_data_Rd[20]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(i_data_Rd[19]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(i_data_Rd[18]), .E(n765), .C(i_clk), .RN(n739), 
        .Q(regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(i_data_Rd[17]), .E(n765), .C(i_clk), .RN(n738), 
        .Q(regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(i_data_Rd[16]), .E(n765), .C(i_clk), .RN(n732), 
        .Q(regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(i_data_Rd[15]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(i_data_Rd[14]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(i_data_Rd[13]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(i_data_Rd[12]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(i_data_Rd[11]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(i_data_Rd[10]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(i_data_Rd[9]), .E(n765), .C(i_clk), .RN(n735), .Q(
        regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(i_data_Rd[8]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(i_data_Rd[7]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(i_data_Rd[6]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(i_data_Rd[5]), .E(n765), .C(i_clk), .RN(n735), .Q(
        regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(i_data_Rd[4]), .E(n765), .C(i_clk), .RN(n739), .Q(
        regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(i_data_Rd[3]), .E(n765), .C(i_clk), .RN(n738), .Q(
        regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(i_data_Rd[2]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(i_data_Rd[1]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(i_data_Rd[0]), .E(n765), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[224]) );
  DFEC1 regs_reg_6__27_ ( .D(i_data_Rd[27]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(i_data_Rd[26]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(i_data_Rd[25]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(i_data_Rd[24]), .E(n766), .C(i_clk), .RN(n731), 
        .Q(regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(i_data_Rd[23]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(i_data_Rd[22]), .E(n766), .C(i_clk), .RN(n733), 
        .Q(regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(i_data_Rd[21]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(i_data_Rd[20]), .E(n766), .C(i_clk), .RN(n738), 
        .Q(regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(i_data_Rd[19]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(i_data_Rd[18]), .E(n766), .C(i_clk), .RN(n733), 
        .Q(regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(i_data_Rd[17]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(i_data_Rd[16]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(i_data_Rd[15]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(i_data_Rd[14]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(i_data_Rd[13]), .E(n766), .C(i_clk), .RN(n739), 
        .Q(regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(i_data_Rd[12]), .E(n766), .C(i_clk), .RN(n731), 
        .Q(regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(i_data_Rd[11]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(i_data_Rd[10]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(i_data_Rd[9]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(i_data_Rd[8]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(i_data_Rd[7]), .E(n766), .C(i_clk), .RN(n737), .Q(
        regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(i_data_Rd[6]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(i_data_Rd[5]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(i_data_Rd[4]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(i_data_Rd[3]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(i_data_Rd[2]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(i_data_Rd[1]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(i_data_Rd[0]), .E(n766), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[192]) );
  DFEC1 regs_reg_5__27_ ( .D(i_data_Rd[27]), .E(n767), .C(i_clk), .RN(n735), 
        .Q(regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(i_data_Rd[26]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(i_data_Rd[25]), .E(n767), .C(i_clk), .RN(n739), 
        .Q(regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(i_data_Rd[24]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(i_data_Rd[23]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(i_data_Rd[22]), .E(n767), .C(i_clk), .RN(n733), 
        .Q(regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(i_data_Rd[21]), .E(n767), .C(i_clk), .RN(n739), 
        .Q(regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(i_data_Rd[20]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(i_data_Rd[19]), .E(n767), .C(i_clk), .RN(n739), 
        .Q(regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(i_data_Rd[18]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(i_data_Rd[17]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(i_data_Rd[16]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(i_data_Rd[15]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(i_data_Rd[14]), .E(n767), .C(i_clk), .RN(n733), 
        .Q(regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(i_data_Rd[13]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(i_data_Rd[12]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(i_data_Rd[11]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(i_data_Rd[10]), .E(n767), .C(i_clk), .RN(n734), 
        .Q(regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(i_data_Rd[9]), .E(n767), .C(i_clk), .RN(n731), .Q(
        regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(i_data_Rd[8]), .E(n767), .C(i_clk), .RN(n738), .Q(
        regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(i_data_Rd[7]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(i_data_Rd[6]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(i_data_Rd[5]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(i_data_Rd[4]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(i_data_Rd[3]), .E(n767), .C(i_clk), .RN(n737), .Q(
        regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(i_data_Rd[2]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(i_data_Rd[1]), .E(n767), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(i_data_Rd[0]), .E(n767), .C(i_clk), .RN(n735), .Q(
        regs[160]) );
  DFEC1 regs_reg_4__27_ ( .D(i_data_Rd[27]), .E(n768), .C(i_clk), .RN(n735), 
        .Q(regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(i_data_Rd[26]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(i_data_Rd[25]), .E(n768), .C(i_clk), .RN(n731), 
        .Q(regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(i_data_Rd[24]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(i_data_Rd[23]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(i_data_Rd[22]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(i_data_Rd[21]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(i_data_Rd[20]), .E(n768), .C(i_clk), .RN(n736), 
        .Q(regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(i_data_Rd[19]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(i_data_Rd[18]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(i_data_Rd[17]), .E(n768), .C(i_clk), .RN(n733), 
        .Q(regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(i_data_Rd[16]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(i_data_Rd[15]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(i_data_Rd[14]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(i_data_Rd[13]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(i_data_Rd[12]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(i_data_Rd[11]), .E(n768), .C(i_clk), .RN(n739), 
        .Q(regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(i_data_Rd[10]), .E(n768), .C(i_clk), .RN(n738), 
        .Q(regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(i_data_Rd[9]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(i_data_Rd[8]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(i_data_Rd[7]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(i_data_Rd[6]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(i_data_Rd[5]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(i_data_Rd[4]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(i_data_Rd[3]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(i_data_Rd[2]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(i_data_Rd[1]), .E(n768), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(i_data_Rd[0]), .E(n768), .C(i_clk), .RN(n732), .Q(
        regs[128]) );
  DFEC1 regs_reg_3__27_ ( .D(i_data_Rd[27]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(i_data_Rd[26]), .E(n769), .C(i_clk), .RN(n733), 
        .Q(regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(i_data_Rd[25]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(i_data_Rd[24]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(i_data_Rd[23]), .E(n769), .C(i_clk), .RN(n734), 
        .Q(regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(i_data_Rd[22]), .E(n769), .C(i_clk), .RN(n732), 
        .Q(regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(i_data_Rd[21]), .E(n769), .C(i_clk), .RN(n736), 
        .Q(regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(i_data_Rd[20]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(i_data_Rd[19]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(i_data_Rd[18]), .E(n769), .C(i_clk), .RN(n738), 
        .Q(regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(i_data_Rd[17]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(i_data_Rd[16]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(i_data_Rd[15]), .E(n769), .C(i_clk), .RN(n731), 
        .Q(regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(i_data_Rd[14]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(i_data_Rd[13]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(i_data_Rd[12]), .E(n769), .C(i_clk), .RN(n738), 
        .Q(regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(i_data_Rd[11]), .E(n769), .C(i_clk), .RN(n736), 
        .Q(regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(i_data_Rd[10]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(i_data_Rd[9]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(i_data_Rd[8]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(i_data_Rd[7]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(i_data_Rd[6]), .E(n769), .C(i_clk), .RN(n732), .Q(
        regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(i_data_Rd[5]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(i_data_Rd[4]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(i_data_Rd[3]), .E(n769), .C(i_clk), .RN(n734), .Q(
        regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(i_data_Rd[2]), .E(n769), .C(i_clk), .RN(n739), .Q(
        regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(i_data_Rd[1]), .E(n769), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(i_data_Rd[0]), .E(n769), .C(i_clk), .RN(n737), .Q(
        regs[96]) );
  DFEC1 regs_reg_2__27_ ( .D(i_data_Rd[27]), .E(n770), .C(i_clk), .RN(n731), 
        .Q(regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(i_data_Rd[26]), .E(n770), .C(i_clk), .RN(n735), 
        .Q(regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(i_data_Rd[25]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(i_data_Rd[24]), .E(n770), .C(i_clk), .RN(n731), 
        .Q(regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(i_data_Rd[23]), .E(n770), .C(i_clk), .RN(n736), 
        .Q(regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(i_data_Rd[22]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(i_data_Rd[21]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(i_data_Rd[20]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(i_data_Rd[19]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(i_data_Rd[18]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(i_data_Rd[17]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(i_data_Rd[16]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(i_data_Rd[15]), .E(n770), .C(i_clk), .RN(n739), 
        .Q(regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(i_data_Rd[14]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(i_data_Rd[13]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(i_data_Rd[12]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(i_data_Rd[11]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(i_data_Rd[10]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(i_data_Rd[9]), .E(n770), .C(i_clk), .RN(n732), .Q(
        regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(i_data_Rd[8]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(i_data_Rd[7]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(i_data_Rd[6]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(i_data_Rd[5]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(i_data_Rd[4]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(i_data_Rd[3]), .E(n770), .C(i_clk), .RN(n739), .Q(
        regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(i_data_Rd[2]), .E(n770), .C(i_clk), .RN(n738), .Q(
        regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(i_data_Rd[1]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(i_data_Rd[0]), .E(n770), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[64]) );
  DFEC1 regs_reg_1__27_ ( .D(i_data_Rd[27]), .E(n771), .C(i_clk), .RN(n736), 
        .Q(regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(i_data_Rd[26]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(i_data_Rd[25]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(i_data_Rd[24]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(i_data_Rd[23]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(i_data_Rd[22]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(i_data_Rd[21]), .E(n771), .C(i_clk), .RN(n738), 
        .Q(regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(i_data_Rd[20]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(i_data_Rd[19]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(i_data_Rd[18]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(i_data_Rd[17]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(i_data_Rd[16]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(i_data_Rd[15]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(i_data_Rd[14]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(i_data_Rd[13]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(i_data_Rd[12]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(i_data_Rd[11]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(i_data_Rd[10]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(i_data_Rd[9]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(i_data_Rd[8]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(i_data_Rd[7]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(i_data_Rd[6]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(i_data_Rd[5]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(i_data_Rd[4]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(i_data_Rd[3]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(i_data_Rd[2]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(i_data_Rd[1]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(i_data_Rd[0]), .E(n771), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[32]) );
  DFEC1 regs_reg_0__27_ ( .D(i_data_Rd[27]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(i_data_Rd[26]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(i_data_Rd[25]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(i_data_Rd[24]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(i_data_Rd[23]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(i_data_Rd[22]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(i_data_Rd[21]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(i_data_Rd[20]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(i_data_Rd[19]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(i_data_Rd[18]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(i_data_Rd[17]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(i_data_Rd[16]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(i_data_Rd[15]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(i_data_Rd[14]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(i_data_Rd[13]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(i_data_Rd[12]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(i_data_Rd[11]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(i_data_Rd[10]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(i_data_Rd[9]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(i_data_Rd[8]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(i_data_Rd[7]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(i_data_Rd[6]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(i_data_Rd[5]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(i_data_Rd[4]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(i_data_Rd[3]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(i_data_Rd[2]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(i_data_Rd[1]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(i_data_Rd[0]), .E(n772), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[0]) );
  DFEC1 regs_reg_31__31_ ( .D(i_data_Rd[31]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1023]) );
  DFEC1 regs_reg_31__30_ ( .D(i_data_Rd[30]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(i_data_Rd[29]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(i_data_Rd[28]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1020]) );
  DFEC1 regs_reg_24__31_ ( .D(i_data_Rd[31]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(i_data_Rd[30]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(i_data_Rd[29]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(i_data_Rd[28]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[796]) );
  DFEC1 regs_reg_23__31_ ( .D(i_data_Rd[31]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(i_data_Rd[30]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(i_data_Rd[29]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(i_data_Rd[28]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[764]) );
  DFEC1 regs_reg_30__31_ ( .D(i_data_Rd[31]), .E(n741), .C(i_clk), .RN(n732), 
        .Q(regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(i_data_Rd[30]), .E(n741), .C(i_clk), .RN(n732), 
        .Q(regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(i_data_Rd[29]), .E(n741), .C(i_clk), .RN(n732), 
        .Q(regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(i_data_Rd[28]), .E(n741), .C(i_clk), .RN(n732), 
        .Q(regs[988]) );
  DFEC1 regs_reg_29__31_ ( .D(i_data_Rd[31]), .E(n742), .C(i_clk), .RN(n736), 
        .Q(regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(i_data_Rd[30]), .E(n742), .C(i_clk), .RN(n736), 
        .Q(regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(i_data_Rd[29]), .E(n742), .C(i_clk), .RN(n736), 
        .Q(regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(i_data_Rd[28]), .E(n742), .C(i_clk), .RN(n736), 
        .Q(regs[956]) );
  DFEC1 regs_reg_28__31_ ( .D(i_data_Rd[31]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(i_data_Rd[30]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(i_data_Rd[29]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(i_data_Rd[28]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[924]) );
  DFEC1 regs_reg_27__31_ ( .D(i_data_Rd[31]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(i_data_Rd[30]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(i_data_Rd[29]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(i_data_Rd[28]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[892]) );
  DFEC1 regs_reg_26__31_ ( .D(i_data_Rd[31]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(i_data_Rd[30]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(i_data_Rd[29]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(i_data_Rd[28]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[860]) );
  DFEC1 regs_reg_25__31_ ( .D(i_data_Rd[31]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(i_data_Rd[30]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(i_data_Rd[29]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(i_data_Rd[28]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[828]) );
  DFEC1 regs_reg_31__27_ ( .D(i_data_Rd[27]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(i_data_Rd[26]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(i_data_Rd[25]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(i_data_Rd[24]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(i_data_Rd[23]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(i_data_Rd[22]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(i_data_Rd[21]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(i_data_Rd[20]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(i_data_Rd[18]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(i_data_Rd[17]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(i_data_Rd[16]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(i_data_Rd[15]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(i_data_Rd[14]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(i_data_Rd[13]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(i_data_Rd[12]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(i_data_Rd[11]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(i_data_Rd[10]), .E(n740), .C(i_clk), .RN(i_rst_n), .Q(regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(i_data_Rd[9]), .E(n740), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(i_data_Rd[8]), .E(n740), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(i_data_Rd[7]), .E(n740), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n740), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(i_data_Rd[5]), .E(n740), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(i_data_Rd[4]), .E(n740), .C(i_clk), .RN(n732), 
        .Q(regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(i_data_Rd[3]), .E(n740), .C(i_clk), .RN(n732), 
        .Q(regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(i_data_Rd[2]), .E(n740), .C(i_clk), .RN(n732), 
        .Q(regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n740), .C(i_clk), .RN(n732), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(i_data_Rd[0]), .E(n740), .C(i_clk), .RN(n732), 
        .Q(regs[992]) );
  DFEC1 regs_reg_24__27_ ( .D(i_data_Rd[27]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(i_data_Rd[26]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(i_data_Rd[25]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(i_data_Rd[24]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(i_data_Rd[23]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(i_data_Rd[22]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(i_data_Rd[21]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(i_data_Rd[20]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(i_data_Rd[19]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(i_data_Rd[18]), .E(n747), .C(i_clk), .RN(n739), 
        .Q(regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(i_data_Rd[17]), .E(n747), .C(i_clk), .RN(n737), 
        .Q(regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(i_data_Rd[16]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(i_data_Rd[15]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(i_data_Rd[14]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(i_data_Rd[13]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(i_data_Rd[12]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(i_data_Rd[11]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(i_data_Rd[10]), .E(n747), .C(i_clk), .RN(i_rst_n), .Q(regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(i_data_Rd[9]), .E(n747), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(i_data_Rd[8]), .E(n747), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(i_data_Rd[7]), .E(n747), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(i_data_Rd[6]), .E(n747), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(i_data_Rd[5]), .E(n747), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(i_data_Rd[4]), .E(n747), .C(i_clk), .RN(n739), 
        .Q(regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(i_data_Rd[3]), .E(n747), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(i_data_Rd[2]), .E(n747), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(i_data_Rd[1]), .E(n747), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(i_data_Rd[0]), .E(n747), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[768]) );
  DFEC1 regs_reg_22__31_ ( .D(i_data_Rd[31]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(i_data_Rd[30]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(i_data_Rd[29]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(i_data_Rd[28]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[732]) );
  DFEC1 regs_reg_21__31_ ( .D(i_data_Rd[31]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(i_data_Rd[30]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(i_data_Rd[29]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(i_data_Rd[28]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[700]) );
  DFEC1 regs_reg_20__31_ ( .D(i_data_Rd[31]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(i_data_Rd[30]), .E(n751), .C(i_clk), .RN(n732), 
        .Q(regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(i_data_Rd[29]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(i_data_Rd[28]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[668]) );
  DFEC1 regs_reg_19__31_ ( .D(i_data_Rd[31]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(i_data_Rd[30]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(i_data_Rd[29]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(i_data_Rd[28]), .E(n752), .C(i_clk), .RN(n732), 
        .Q(regs[636]) );
  DFEC1 regs_reg_18__31_ ( .D(i_data_Rd[31]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(i_data_Rd[30]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(i_data_Rd[29]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(i_data_Rd[28]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[604]) );
  DFEC1 regs_reg_17__31_ ( .D(i_data_Rd[31]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(i_data_Rd[30]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(i_data_Rd[29]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(i_data_Rd[28]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[572]) );
  DFEC1 regs_reg_16__31_ ( .D(i_data_Rd[31]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(i_data_Rd[30]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(i_data_Rd[29]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(i_data_Rd[28]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[540]) );
  DFEC1 regs_reg_23__27_ ( .D(i_data_Rd[27]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(i_data_Rd[26]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(i_data_Rd[25]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(i_data_Rd[24]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(i_data_Rd[23]), .E(n748), .C(i_clk), .RN(n731), 
        .Q(regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(i_data_Rd[22]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(i_data_Rd[21]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(i_data_Rd[20]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(i_data_Rd[19]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(i_data_Rd[18]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(i_data_Rd[17]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(i_data_Rd[16]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(i_data_Rd[15]), .E(n748), .C(i_clk), .RN(n739), 
        .Q(regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(i_data_Rd[14]), .E(n748), .C(i_clk), .RN(n738), 
        .Q(regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(i_data_Rd[13]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(i_data_Rd[12]), .E(n748), .C(i_clk), .RN(n738), 
        .Q(regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(i_data_Rd[11]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(i_data_Rd[10]), .E(n748), .C(i_clk), .RN(i_rst_n), .Q(regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(i_data_Rd[9]), .E(n748), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(i_data_Rd[8]), .E(n748), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(i_data_Rd[7]), .E(n748), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(i_data_Rd[6]), .E(n748), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(i_data_Rd[5]), .E(n748), .C(i_clk), .RN(n732), 
        .Q(regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(i_data_Rd[4]), .E(n748), .C(i_clk), .RN(n733), 
        .Q(regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(i_data_Rd[3]), .E(n748), .C(i_clk), .RN(n734), 
        .Q(regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(i_data_Rd[2]), .E(n748), .C(i_clk), .RN(n735), 
        .Q(regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(i_data_Rd[1]), .E(n748), .C(i_clk), .RN(n736), 
        .Q(regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(i_data_Rd[0]), .E(n748), .C(i_clk), .RN(n737), 
        .Q(regs[736]) );
  DFEC1 regs_reg_30__27_ ( .D(i_data_Rd[27]), .E(n741), .C(i_clk), .RN(n733), 
        .Q(regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(i_data_Rd[26]), .E(n741), .C(i_clk), .RN(n733), 
        .Q(regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(i_data_Rd[25]), .E(n741), .C(i_clk), .RN(n733), 
        .Q(regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(i_data_Rd[24]), .E(n741), .C(i_clk), .RN(n733), 
        .Q(regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(i_data_Rd[23]), .E(n741), .C(i_clk), .RN(n733), 
        .Q(regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(i_data_Rd[22]), .E(n741), .C(i_clk), .RN(n733), 
        .Q(regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(i_data_Rd[21]), .E(n741), .C(i_clk), .RN(n733), 
        .Q(regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(i_data_Rd[20]), .E(n741), .C(i_clk), .RN(n733), 
        .Q(regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n741), .C(i_clk), .RN(n733), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(i_data_Rd[18]), .E(n741), .C(i_clk), .RN(n734), 
        .Q(regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(i_data_Rd[17]), .E(n741), .C(i_clk), .RN(n734), 
        .Q(regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(i_data_Rd[16]), .E(n741), .C(i_clk), .RN(n734), 
        .Q(regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(i_data_Rd[15]), .E(n741), .C(i_clk), .RN(n734), 
        .Q(regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(i_data_Rd[14]), .E(n741), .C(i_clk), .RN(n734), 
        .Q(regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(i_data_Rd[13]), .E(n741), .C(i_clk), .RN(n734), 
        .Q(regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(i_data_Rd[12]), .E(n741), .C(i_clk), .RN(n734), 
        .Q(regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(i_data_Rd[11]), .E(n741), .C(i_clk), .RN(n734), 
        .Q(regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(i_data_Rd[10]), .E(n741), .C(i_clk), .RN(n734), 
        .Q(regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(i_data_Rd[9]), .E(n741), .C(i_clk), .RN(n735), 
        .Q(regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(i_data_Rd[8]), .E(n741), .C(i_clk), .RN(n735), 
        .Q(regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(i_data_Rd[7]), .E(n741), .C(i_clk), .RN(n735), 
        .Q(regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n741), .C(i_clk), .RN(n735), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(i_data_Rd[5]), .E(n741), .C(i_clk), .RN(n735), 
        .Q(regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(i_data_Rd[4]), .E(n741), .C(i_clk), .RN(n735), 
        .Q(regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(i_data_Rd[3]), .E(n741), .C(i_clk), .RN(n735), 
        .Q(regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(i_data_Rd[2]), .E(n741), .C(i_clk), .RN(n735), 
        .Q(regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n741), .C(i_clk), .RN(n735), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(i_data_Rd[0]), .E(n741), .C(i_clk), .RN(n736), 
        .Q(regs[960]) );
  DFEC1 regs_reg_29__27_ ( .D(i_data_Rd[27]), .E(n742), .C(i_clk), .RN(n736), 
        .Q(regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(i_data_Rd[26]), .E(n742), .C(i_clk), .RN(n736), 
        .Q(regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(i_data_Rd[25]), .E(n742), .C(i_clk), .RN(n736), 
        .Q(regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(i_data_Rd[24]), .E(n742), .C(i_clk), .RN(n736), 
        .Q(regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(i_data_Rd[23]), .E(n742), .C(i_clk), .RN(n737), 
        .Q(regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(i_data_Rd[22]), .E(n742), .C(i_clk), .RN(n737), 
        .Q(regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(i_data_Rd[21]), .E(n742), .C(i_clk), .RN(n737), 
        .Q(regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(i_data_Rd[20]), .E(n742), .C(i_clk), .RN(n737), 
        .Q(regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n742), .C(i_clk), .RN(n737), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(i_data_Rd[18]), .E(n742), .C(i_clk), .RN(n737), 
        .Q(regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(i_data_Rd[17]), .E(n742), .C(i_clk), .RN(n737), 
        .Q(regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(i_data_Rd[16]), .E(n742), .C(i_clk), .RN(n737), 
        .Q(regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(i_data_Rd[15]), .E(n742), .C(i_clk), .RN(n737), 
        .Q(regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(i_data_Rd[14]), .E(n742), .C(i_clk), .RN(i_rst_n), .Q(regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(i_data_Rd[13]), .E(n742), .C(i_clk), .RN(i_rst_n), .Q(regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(i_data_Rd[12]), .E(n742), .C(i_clk), .RN(i_rst_n), .Q(regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(i_data_Rd[11]), .E(n742), .C(i_clk), .RN(i_rst_n), .Q(regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(i_data_Rd[10]), .E(n742), .C(i_clk), .RN(i_rst_n), .Q(regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(i_data_Rd[9]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(i_data_Rd[8]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(i_data_Rd[7]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(i_data_Rd[5]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(i_data_Rd[4]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(i_data_Rd[3]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(i_data_Rd[2]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(i_data_Rd[0]), .E(n742), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[928]) );
  DFEC1 regs_reg_28__27_ ( .D(i_data_Rd[27]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(i_data_Rd[26]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(i_data_Rd[25]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(i_data_Rd[24]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(i_data_Rd[23]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(i_data_Rd[22]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(i_data_Rd[21]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(i_data_Rd[20]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(i_data_Rd[18]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(i_data_Rd[17]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(i_data_Rd[16]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(i_data_Rd[15]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(i_data_Rd[14]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(i_data_Rd[13]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(i_data_Rd[12]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(i_data_Rd[11]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(i_data_Rd[10]), .E(n743), .C(i_clk), .RN(i_rst_n), .Q(regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(i_data_Rd[9]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(i_data_Rd[8]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(i_data_Rd[7]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(i_data_Rd[5]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(i_data_Rd[4]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(i_data_Rd[3]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(i_data_Rd[2]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(i_data_Rd[0]), .E(n743), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[896]) );
  DFEC1 regs_reg_27__27_ ( .D(i_data_Rd[27]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(i_data_Rd[26]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(i_data_Rd[25]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(i_data_Rd[24]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(i_data_Rd[23]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(i_data_Rd[22]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(i_data_Rd[21]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(i_data_Rd[20]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(i_data_Rd[18]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(i_data_Rd[17]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(i_data_Rd[16]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(i_data_Rd[15]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(i_data_Rd[14]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(i_data_Rd[13]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(i_data_Rd[12]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(i_data_Rd[11]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(i_data_Rd[10]), .E(n744), .C(i_clk), .RN(i_rst_n), .Q(regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(i_data_Rd[9]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(i_data_Rd[8]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(i_data_Rd[7]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(i_data_Rd[5]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(i_data_Rd[4]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(i_data_Rd[3]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(i_data_Rd[2]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(i_data_Rd[1]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(i_data_Rd[0]), .E(n744), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[864]) );
  DFEC1 regs_reg_26__27_ ( .D(i_data_Rd[27]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(i_data_Rd[26]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(i_data_Rd[25]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(i_data_Rd[24]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(i_data_Rd[23]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(i_data_Rd[22]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(i_data_Rd[21]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(i_data_Rd[20]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(i_data_Rd[18]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(i_data_Rd[17]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(i_data_Rd[16]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(i_data_Rd[15]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(i_data_Rd[14]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(i_data_Rd[13]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(i_data_Rd[12]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(i_data_Rd[11]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(i_data_Rd[10]), .E(n745), .C(i_clk), .RN(i_rst_n), .Q(regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(i_data_Rd[9]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(i_data_Rd[8]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(i_data_Rd[7]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(i_data_Rd[5]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(i_data_Rd[4]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(i_data_Rd[3]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(i_data_Rd[2]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(i_data_Rd[0]), .E(n745), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[832]) );
  DFEC1 regs_reg_25__27_ ( .D(i_data_Rd[27]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(i_data_Rd[26]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(i_data_Rd[25]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(i_data_Rd[24]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(i_data_Rd[23]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(i_data_Rd[22]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(i_data_Rd[21]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(i_data_Rd[20]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(i_data_Rd[19]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(i_data_Rd[18]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(i_data_Rd[17]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(i_data_Rd[16]), .E(n746), .C(i_clk), .RN(n733), 
        .Q(regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(i_data_Rd[15]), .E(n746), .C(i_clk), .RN(n734), 
        .Q(regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(i_data_Rd[14]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(i_data_Rd[13]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(i_data_Rd[12]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(i_data_Rd[11]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(i_data_Rd[10]), .E(n746), .C(i_clk), .RN(i_rst_n), .Q(regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(i_data_Rd[9]), .E(n746), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(i_data_Rd[8]), .E(n746), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(i_data_Rd[7]), .E(n746), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(i_data_Rd[6]), .E(n746), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(i_data_Rd[5]), .E(n746), .C(i_clk), .RN(n738), 
        .Q(regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(i_data_Rd[4]), .E(n746), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(i_data_Rd[3]), .E(n746), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(i_data_Rd[2]), .E(n746), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(i_data_Rd[1]), .E(n746), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(i_data_Rd[0]), .E(n746), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[800]) );
  DFEC1 regs_reg_22__27_ ( .D(i_data_Rd[27]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(i_data_Rd[26]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(i_data_Rd[25]), .E(n749), .C(i_clk), .RN(n739), 
        .Q(regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(i_data_Rd[24]), .E(n749), .C(i_clk), .RN(n734), 
        .Q(regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(i_data_Rd[23]), .E(n749), .C(i_clk), .RN(n731), 
        .Q(regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(i_data_Rd[22]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(i_data_Rd[21]), .E(n749), .C(i_clk), .RN(n737), 
        .Q(regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(i_data_Rd[20]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(i_data_Rd[19]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(i_data_Rd[18]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(i_data_Rd[17]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(i_data_Rd[16]), .E(n749), .C(i_clk), .RN(n736), 
        .Q(regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(i_data_Rd[15]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(i_data_Rd[14]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(i_data_Rd[13]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(i_data_Rd[12]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(i_data_Rd[11]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(i_data_Rd[10]), .E(n749), .C(i_clk), .RN(i_rst_n), .Q(regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(i_data_Rd[9]), .E(n749), .C(i_clk), .RN(n739), 
        .Q(regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(i_data_Rd[8]), .E(n749), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(i_data_Rd[7]), .E(n749), .C(i_clk), .RN(n731), 
        .Q(regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(i_data_Rd[6]), .E(n749), .C(i_clk), .RN(n732), 
        .Q(regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(i_data_Rd[5]), .E(n749), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(i_data_Rd[4]), .E(n749), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(i_data_Rd[3]), .E(n749), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(i_data_Rd[2]), .E(n749), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(i_data_Rd[1]), .E(n749), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(i_data_Rd[0]), .E(n749), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[704]) );
  DFEC1 regs_reg_21__27_ ( .D(i_data_Rd[27]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(i_data_Rd[26]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(i_data_Rd[25]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(i_data_Rd[24]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(i_data_Rd[23]), .E(n750), .C(i_clk), .RN(n731), 
        .Q(regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(i_data_Rd[22]), .E(n750), .C(i_clk), .RN(n739), 
        .Q(regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(i_data_Rd[21]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(i_data_Rd[20]), .E(n750), .C(i_clk), .RN(n731), 
        .Q(regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(i_data_Rd[19]), .E(n750), .C(i_clk), .RN(n732), 
        .Q(regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(i_data_Rd[18]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(i_data_Rd[17]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(i_data_Rd[16]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(i_data_Rd[15]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(i_data_Rd[14]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(i_data_Rd[13]), .E(n750), .C(i_clk), .RN(n736), 
        .Q(regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(i_data_Rd[12]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(i_data_Rd[11]), .E(n750), .C(i_clk), .RN(n738), 
        .Q(regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(i_data_Rd[10]), .E(n750), .C(i_clk), .RN(i_rst_n), .Q(regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(i_data_Rd[9]), .E(n750), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(i_data_Rd[8]), .E(n750), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(i_data_Rd[7]), .E(n750), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(i_data_Rd[6]), .E(n750), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(i_data_Rd[5]), .E(n750), .C(i_clk), .RN(n734), 
        .Q(regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(i_data_Rd[4]), .E(n750), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(i_data_Rd[3]), .E(n750), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(i_data_Rd[2]), .E(n750), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(i_data_Rd[1]), .E(n750), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(i_data_Rd[0]), .E(n750), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[672]) );
  DFEC1 regs_reg_20__27_ ( .D(i_data_Rd[27]), .E(n751), .C(i_clk), .RN(n738), 
        .Q(regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(i_data_Rd[26]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(i_data_Rd[25]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(i_data_Rd[24]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(i_data_Rd[23]), .E(n751), .C(i_clk), .RN(n731), 
        .Q(regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(i_data_Rd[22]), .E(n751), .C(i_clk), .RN(n737), 
        .Q(regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(i_data_Rd[21]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(i_data_Rd[20]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(i_data_Rd[19]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(i_data_Rd[18]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(i_data_Rd[17]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(i_data_Rd[16]), .E(n751), .C(i_clk), .RN(n739), 
        .Q(regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(i_data_Rd[15]), .E(n751), .C(i_clk), .RN(n738), 
        .Q(regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(i_data_Rd[14]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(i_data_Rd[13]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(i_data_Rd[12]), .E(n751), .C(i_clk), .RN(n733), 
        .Q(regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(i_data_Rd[11]), .E(n751), .C(i_clk), .RN(n731), 
        .Q(regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(i_data_Rd[10]), .E(n751), .C(i_clk), .RN(i_rst_n), .Q(regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(i_data_Rd[9]), .E(n751), .C(i_clk), .RN(n738), 
        .Q(regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(i_data_Rd[8]), .E(n751), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(i_data_Rd[7]), .E(n751), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(i_data_Rd[6]), .E(n751), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(i_data_Rd[5]), .E(n751), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(i_data_Rd[4]), .E(n751), .C(i_clk), .RN(n737), 
        .Q(regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(i_data_Rd[3]), .E(n751), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(i_data_Rd[2]), .E(n751), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(i_data_Rd[1]), .E(n751), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(i_data_Rd[0]), .E(n751), .C(i_clk), .RN(n734), 
        .Q(regs[640]) );
  DFEC1 regs_reg_19__27_ ( .D(i_data_Rd[27]), .E(n752), .C(i_clk), .RN(n731), 
        .Q(regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(i_data_Rd[26]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(i_data_Rd[25]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(i_data_Rd[24]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(i_data_Rd[23]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(i_data_Rd[22]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(i_data_Rd[21]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(i_data_Rd[20]), .E(n752), .C(i_clk), .RN(n731), 
        .Q(regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(i_data_Rd[19]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(i_data_Rd[18]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(i_data_Rd[17]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(i_data_Rd[16]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(i_data_Rd[15]), .E(n752), .C(i_clk), .RN(n739), 
        .Q(regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(i_data_Rd[14]), .E(n752), .C(i_clk), .RN(n738), 
        .Q(regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(i_data_Rd[13]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(i_data_Rd[12]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(i_data_Rd[11]), .E(n752), .C(i_clk), .RN(i_rst_n), .Q(regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(i_data_Rd[10]), .E(n752), .C(i_clk), .RN(n734), 
        .Q(regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(i_data_Rd[9]), .E(n752), .C(i_clk), .RN(n735), 
        .Q(regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(i_data_Rd[8]), .E(n752), .C(i_clk), .RN(n736), 
        .Q(regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(i_data_Rd[7]), .E(n752), .C(i_clk), .RN(n737), 
        .Q(regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(i_data_Rd[6]), .E(n752), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(i_data_Rd[5]), .E(n752), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(i_data_Rd[4]), .E(n752), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(i_data_Rd[3]), .E(n752), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(i_data_Rd[2]), .E(n752), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(i_data_Rd[1]), .E(n752), .C(i_clk), .RN(n733), 
        .Q(regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(i_data_Rd[0]), .E(n752), .C(i_clk), .RN(n738), 
        .Q(regs[608]) );
  DFEC1 regs_reg_18__27_ ( .D(i_data_Rd[27]), .E(n753), .C(i_clk), .RN(n731), 
        .Q(regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(i_data_Rd[26]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(i_data_Rd[25]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(i_data_Rd[24]), .E(n753), .C(i_clk), .RN(n733), 
        .Q(regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(i_data_Rd[23]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(i_data_Rd[22]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(i_data_Rd[21]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(i_data_Rd[20]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(i_data_Rd[19]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(i_data_Rd[18]), .E(n753), .C(i_clk), .RN(n735), 
        .Q(regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(i_data_Rd[17]), .E(n753), .C(i_clk), .RN(n736), 
        .Q(regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(i_data_Rd[16]), .E(n753), .C(i_clk), .RN(n732), 
        .Q(regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(i_data_Rd[15]), .E(n753), .C(i_clk), .RN(n739), 
        .Q(regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(i_data_Rd[14]), .E(n753), .C(i_clk), .RN(n735), 
        .Q(regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(i_data_Rd[13]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(i_data_Rd[12]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(i_data_Rd[11]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(i_data_Rd[10]), .E(n753), .C(i_clk), .RN(i_rst_n), .Q(regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(i_data_Rd[9]), .E(n753), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(i_data_Rd[8]), .E(n753), .C(i_clk), .RN(n735), 
        .Q(regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(i_data_Rd[7]), .E(n753), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(i_data_Rd[6]), .E(n753), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(i_data_Rd[5]), .E(n753), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(i_data_Rd[4]), .E(n753), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(i_data_Rd[3]), .E(n753), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(i_data_Rd[2]), .E(n753), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(i_data_Rd[1]), .E(n753), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(i_data_Rd[0]), .E(n753), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[576]) );
  DFEC1 regs_reg_17__27_ ( .D(i_data_Rd[27]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(i_data_Rd[26]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(i_data_Rd[25]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(i_data_Rd[24]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(i_data_Rd[23]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(i_data_Rd[22]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(i_data_Rd[21]), .E(n754), .C(i_clk), .RN(n739), 
        .Q(regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(i_data_Rd[20]), .E(n754), .C(i_clk), .RN(n731), 
        .Q(regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(i_data_Rd[19]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(i_data_Rd[18]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(i_data_Rd[17]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(i_data_Rd[16]), .E(n754), .C(i_clk), .RN(n736), 
        .Q(regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(i_data_Rd[15]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(i_data_Rd[14]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(i_data_Rd[13]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(i_data_Rd[12]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(i_data_Rd[11]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(i_data_Rd[10]), .E(n754), .C(i_clk), .RN(i_rst_n), .Q(regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(i_data_Rd[9]), .E(n754), .C(i_clk), .RN(n736), 
        .Q(regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(i_data_Rd[8]), .E(n754), .C(i_clk), .RN(n735), 
        .Q(regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(i_data_Rd[7]), .E(n754), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(i_data_Rd[6]), .E(n754), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(i_data_Rd[5]), .E(n754), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(i_data_Rd[4]), .E(n754), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(i_data_Rd[3]), .E(n754), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(i_data_Rd[2]), .E(n754), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(i_data_Rd[1]), .E(n754), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(i_data_Rd[0]), .E(n754), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[544]) );
  DFEC1 regs_reg_16__27_ ( .D(i_data_Rd[27]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(i_data_Rd[26]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(i_data_Rd[25]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(i_data_Rd[24]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(i_data_Rd[23]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(i_data_Rd[22]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(i_data_Rd[21]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(i_data_Rd[20]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(i_data_Rd[19]), .E(n755), .C(i_clk), .RN(n739), 
        .Q(regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(i_data_Rd[18]), .E(n755), .C(i_clk), .RN(n738), 
        .Q(regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(i_data_Rd[17]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(i_data_Rd[16]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(i_data_Rd[15]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(i_data_Rd[14]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(i_data_Rd[13]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(i_data_Rd[12]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(i_data_Rd[11]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(i_data_Rd[10]), .E(n755), .C(i_clk), .RN(i_rst_n), .Q(regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(i_data_Rd[9]), .E(n755), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(i_data_Rd[8]), .E(n755), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(i_data_Rd[7]), .E(n755), .C(i_clk), .RN(n736), 
        .Q(regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(i_data_Rd[6]), .E(n755), .C(i_clk), .RN(n737), 
        .Q(regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(i_data_Rd[5]), .E(n755), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(i_data_Rd[4]), .E(n755), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(i_data_Rd[3]), .E(n755), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(i_data_Rd[2]), .E(n755), .C(i_clk), .RN(n738), 
        .Q(regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(i_data_Rd[1]), .E(n755), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(i_data_Rd[0]), .E(n755), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[512]) );
  BUF2 U2 ( .A(n738), .Q(n737) );
  BUF2 U3 ( .A(n738), .Q(n736) );
  BUF2 U4 ( .A(n738), .Q(n735) );
  BUF2 U5 ( .A(n739), .Q(n734) );
  BUF2 U6 ( .A(n739), .Q(n733) );
  BUF2 U7 ( .A(n739), .Q(n732) );
  BUF2 U8 ( .A(n731), .Q(n738) );
  BUF2 U9 ( .A(n731), .Q(n739) );
  BUF2 U10 ( .A(i_addr_Rt[0]), .Q(n376) );
  BUF2 U11 ( .A(i_addr_Rt[0]), .Q(n377) );
  BUF2 U12 ( .A(i_addr_Rt[0]), .Q(n378) );
  BUF2 U13 ( .A(n385), .Q(n379) );
  BUF2 U14 ( .A(n385), .Q(n380) );
  BUF2 U15 ( .A(n386), .Q(n381) );
  BUF2 U16 ( .A(n386), .Q(n382) );
  BUF2 U17 ( .A(n387), .Q(n383) );
  BUF2 U18 ( .A(n387), .Q(n384) );
  BUF2 U19 ( .A(n728), .Q(n719) );
  BUF2 U20 ( .A(n729), .Q(n720) );
  BUF2 U21 ( .A(n727), .Q(n721) );
  BUF2 U22 ( .A(n727), .Q(n722) );
  BUF2 U23 ( .A(n727), .Q(n723) );
  BUF2 U24 ( .A(n729), .Q(n724) );
  BUF2 U25 ( .A(n730), .Q(n725) );
  BUF2 U26 ( .A(n730), .Q(n726) );
  INV3 U27 ( .A(n55), .Q(n740) );
  NAND22 U28 ( .A(n41), .B(n56), .Q(n55) );
  BUF2 U29 ( .A(i_addr_Rt[1]), .Q(n371) );
  BUF2 U30 ( .A(n370), .Q(n372) );
  BUF2 U31 ( .A(n714), .Q(n715) );
  BUF2 U32 ( .A(n713), .Q(n716) );
  BUF2 U33 ( .A(i_rst_n), .Q(n731) );
  NOR31 U34 ( .A(n777), .B(n756), .C(n773), .Q(n41) );
  NOR31 U35 ( .A(n775), .B(n776), .C(n774), .Q(n56) );
  INV3 U36 ( .A(n39), .Q(n748) );
  NAND22 U37 ( .A(n76), .B(n56), .Q(n39) );
  INV3 U38 ( .A(n75), .Q(n755) );
  NAND22 U39 ( .A(n42), .B(n76), .Q(n75) );
  INV3 U40 ( .A(n77), .Q(n754) );
  NAND22 U41 ( .A(n44), .B(n76), .Q(n77) );
  INV3 U42 ( .A(n78), .Q(n753) );
  NAND22 U43 ( .A(n46), .B(n76), .Q(n78) );
  INV3 U44 ( .A(n79), .Q(n752) );
  NAND22 U45 ( .A(n48), .B(n76), .Q(n79) );
  INV3 U46 ( .A(n80), .Q(n751) );
  NAND22 U47 ( .A(n50), .B(n76), .Q(n80) );
  INV3 U48 ( .A(n81), .Q(n750) );
  NAND22 U49 ( .A(n52), .B(n76), .Q(n81) );
  INV3 U50 ( .A(n82), .Q(n749) );
  NAND22 U51 ( .A(n54), .B(n76), .Q(n82) );
  INV3 U52 ( .A(n43), .Q(n746) );
  NAND22 U53 ( .A(n44), .B(n41), .Q(n43) );
  INV3 U54 ( .A(n45), .Q(n745) );
  NAND22 U55 ( .A(n46), .B(n41), .Q(n45) );
  INV3 U56 ( .A(n47), .Q(n744) );
  NAND22 U57 ( .A(n48), .B(n41), .Q(n47) );
  INV3 U58 ( .A(n49), .Q(n743) );
  NAND22 U59 ( .A(n50), .B(n41), .Q(n49) );
  INV3 U60 ( .A(n51), .Q(n742) );
  NAND22 U61 ( .A(n52), .B(n41), .Q(n51) );
  INV3 U62 ( .A(n53), .Q(n741) );
  NAND22 U63 ( .A(n54), .B(n41), .Q(n53) );
  INV3 U64 ( .A(n57), .Q(n772) );
  NAND22 U65 ( .A(n58), .B(n42), .Q(n57) );
  INV3 U66 ( .A(n60), .Q(n770) );
  NAND22 U67 ( .A(n58), .B(n46), .Q(n60) );
  INV3 U68 ( .A(n62), .Q(n768) );
  NAND22 U69 ( .A(n58), .B(n50), .Q(n62) );
  INV3 U70 ( .A(n63), .Q(n767) );
  NAND22 U71 ( .A(n58), .B(n52), .Q(n63) );
  INV3 U72 ( .A(n65), .Q(n765) );
  NAND22 U73 ( .A(n58), .B(n56), .Q(n65) );
  INV3 U74 ( .A(n69), .Q(n762) );
  NAND22 U75 ( .A(n67), .B(n46), .Q(n69) );
  INV3 U76 ( .A(n71), .Q(n760) );
  NAND22 U77 ( .A(n67), .B(n50), .Q(n71) );
  INV3 U78 ( .A(n72), .Q(n759) );
  NAND22 U79 ( .A(n67), .B(n52), .Q(n72) );
  INV3 U80 ( .A(n74), .Q(n757) );
  NAND22 U81 ( .A(n67), .B(n56), .Q(n74) );
  INV3 U82 ( .A(n40), .Q(n747) );
  NAND22 U83 ( .A(n41), .B(n42), .Q(n40) );
  INV3 U84 ( .A(n66), .Q(n764) );
  NAND22 U85 ( .A(n67), .B(n42), .Q(n66) );
  INV3 U86 ( .A(n59), .Q(n771) );
  NAND22 U87 ( .A(n58), .B(n44), .Q(n59) );
  INV3 U88 ( .A(n68), .Q(n763) );
  NAND22 U89 ( .A(n67), .B(n44), .Q(n68) );
  INV3 U90 ( .A(n61), .Q(n769) );
  NAND22 U91 ( .A(n58), .B(n48), .Q(n61) );
  INV3 U92 ( .A(n64), .Q(n766) );
  NAND22 U93 ( .A(n58), .B(n54), .Q(n64) );
  INV3 U94 ( .A(n70), .Q(n761) );
  NAND22 U95 ( .A(n67), .B(n48), .Q(n70) );
  INV3 U96 ( .A(n73), .Q(n758) );
  NAND22 U97 ( .A(n67), .B(n54), .Q(n73) );
  BUF2 U98 ( .A(n369), .Q(n373) );
  BUF2 U99 ( .A(n369), .Q(n374) );
  BUF2 U100 ( .A(n712), .Q(n717) );
  BUF2 U101 ( .A(n712), .Q(n718) );
  BUF2 U102 ( .A(i_addr_Rt[0]), .Q(n385) );
  BUF2 U103 ( .A(i_addr_Rt[0]), .Q(n386) );
  BUF2 U104 ( .A(i_addr_Rt[0]), .Q(n387) );
  BUF2 U105 ( .A(i_addr_Rs[0]), .Q(n727) );
  BUF2 U106 ( .A(i_addr_Rs[0]), .Q(n728) );
  BUF2 U107 ( .A(i_addr_Rs[0]), .Q(n729) );
  BUF2 U108 ( .A(i_addr_Rs[0]), .Q(n730) );
  BUF2 U109 ( .A(i_addr_Rt[1]), .Q(n370) );
  BUF2 U110 ( .A(i_addr_Rs[1]), .Q(n714) );
  BUF2 U111 ( .A(i_addr_Rs[1]), .Q(n713) );
  NOR31 U112 ( .A(n756), .B(i_addr_Rd[3]), .C(n777), .Q(n76) );
  NOR31 U113 ( .A(i_addr_Rd[3]), .B(i_addr_Rd[4]), .C(n777), .Q(n58) );
  NOR31 U114 ( .A(n777), .B(i_addr_Rd[4]), .C(n773), .Q(n67) );
  MUX22 U115 ( .A(n393), .B(n388), .S(n708), .Q(o_data_Rs[0]) );
  IMUX40 U116 ( .A(n389), .B(n390), .C(n391), .D(n392), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n388) );
  IMUX40 U117 ( .A(n394), .B(n395), .C(n396), .D(n397), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n393) );
  NOR31 U118 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(i_addr_Rd[0]), .Q(n42)
         );
  NOR31 U119 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n774), .Q(n50) );
  NOR31 U120 ( .A(n776), .B(i_addr_Rd[1]), .C(n774), .Q(n52) );
  NOR31 U121 ( .A(n775), .B(i_addr_Rd[0]), .C(n774), .Q(n54) );
  NOR31 U122 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[2]), .C(n776), .Q(n44) );
  NOR31 U123 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[2]), .C(n775), .Q(n46) );
  NOR31 U124 ( .A(n776), .B(i_addr_Rd[2]), .C(n775), .Q(n48) );
  IMUX40 U125 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n386), .S1(n372), .Q(n10) );
  IMUX40 U126 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n8) );
  IMUX40 U127 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n387), .S1(i_addr_Rt[1]), .Q(n7) );
  IMUX40 U128 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(i_addr_Rt[0]), .S1(n375), .Q(n5) );
  IMUX40 U129 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(i_addr_Rt[0]), .S1(n371), .Q(n3) );
  IMUX40 U130 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n2) );
  IMUX40 U131 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n386), .S1(n369), .Q(n15) );
  IMUX40 U132 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n387), .S1(i_addr_Rt[1]), .Q(n13) );
  IMUX40 U133 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n383), .S1(i_addr_Rt[1]), .Q(n12) );
  IMUX40 U134 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n387), .S1(n375), .Q(n20) );
  IMUX40 U135 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n382), .S1(i_addr_Rt[1]), .Q(n18) );
  IMUX40 U136 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(i_addr_Rt[0]), .S1(n369), .Q(n25) );
  IMUX40 U137 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n387), .S1(n374), .Q(n23) );
  IMUX40 U138 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n387), .S1(i_addr_Rt[1]), .Q(n22) );
  IMUX40 U139 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n380), .S1(n375), .Q(n30) );
  IMUX40 U140 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n28) );
  IMUX40 U141 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(n378), .S1(n371), .Q(n35) );
  IMUX40 U142 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(n376), .S1(i_addr_Rt[1]), .Q(n33) );
  IMUX40 U143 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n32) );
  IMUX40 U144 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(n383), .S1(n369), .Q(n84) );
  IMUX40 U145 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n386), .S1(i_addr_Rt[1]), .Q(n38) );
  IMUX40 U146 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(i_addr_Rt[0]), .S1(n375), .Q(n89) );
  IMUX40 U147 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n385), .S1(n370), .Q(n87) );
  IMUX40 U148 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(n381), .S1(i_addr_Rt[1]), .Q(n86) );
  IMUX40 U149 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(i_addr_Rt[0]), .S1(n371), .Q(n94) );
  IMUX40 U150 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n380), .S1(i_addr_Rt[1]), .Q(n92) );
  IMUX40 U151 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(n376), .S1(n375), .Q(n99) );
  IMUX40 U152 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n97) );
  IMUX40 U153 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(n386), .S1(n373), .Q(n96) );
  IMUX40 U154 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(n387), .S1(n375), .Q(n104) );
  IMUX40 U155 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n102) );
  IMUX40 U156 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n386), .S1(n373), .Q(n109) );
  IMUX40 U157 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n376), .S1(n372), .Q(n107) );
  IMUX40 U158 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(n382), .S1(i_addr_Rt[1]), .Q(n106) );
  IMUX40 U159 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(i_addr_Rt[0]), .S1(i_addr_Rt[1]), .Q(n114) );
  IMUX40 U160 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n385), .S1(i_addr_Rt[1]), .Q(n112) );
  IMUX40 U161 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n387), .S1(n375), .Q(n119) );
  IMUX40 U162 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n117) );
  IMUX40 U163 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n379), .S1(n370), .Q(n116) );
  IMUX40 U164 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n385), .S1(n375), .Q(n124) );
  IMUX40 U165 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n386), .S1(n372), .Q(n122) );
  IMUX40 U166 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n386), .S1(n375), .Q(n129) );
  IMUX40 U167 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n386), .S1(n371), .Q(n127) );
  IMUX40 U168 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n378), .S1(i_addr_Rt[1]), .Q(n126) );
  IMUX40 U169 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(n387), .S1(n369), .Q(n134) );
  IMUX40 U170 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n386), .S1(n375), .Q(n132) );
  IMUX40 U171 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n384), .S1(n375), .Q(n139) );
  IMUX40 U172 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n387), .S1(n369), .Q(n137) );
  IMUX40 U173 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n380), .S1(i_addr_Rt[1]), .Q(n136) );
  IMUX40 U174 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n376), .S1(i_addr_Rt[1]), .Q(n144) );
  IMUX40 U175 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n386), .S1(i_addr_Rt[1]), .Q(n142) );
  IMUX40 U176 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n383), .S1(n370), .Q(n149) );
  IMUX40 U177 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n386), .S1(n374), .Q(n147) );
  IMUX40 U178 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n387), .S1(i_addr_Rt[1]), .Q(n146) );
  IMUX40 U179 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(n377), .S1(n371), .Q(n154) );
  IMUX40 U180 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n378), .S1(n375), .Q(n152) );
  IMUX40 U181 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n376), .S1(n369), .Q(n159) );
  IMUX40 U182 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n376), .S1(n369), .Q(n157) );
  IMUX40 U183 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n376), .S1(i_addr_Rt[1]), .Q(n156) );
  IMUX40 U184 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n376), .S1(i_addr_Rt[1]), .Q(n164) );
  IMUX40 U185 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n376), .S1(n369), .Q(n162) );
  IMUX40 U186 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n376), .S1(n371), .Q(n169) );
  IMUX40 U187 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n376), .S1(n375), .Q(n167) );
  IMUX40 U188 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n376), .S1(n374), .Q(n166) );
  IMUX40 U189 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n377), .S1(i_addr_Rt[1]), .Q(n174) );
  IMUX40 U190 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n377), .S1(n372), .Q(n172) );
  IMUX40 U191 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n377), .S1(n375), .Q(n179) );
  IMUX40 U192 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n377), .S1(n369), .Q(n177) );
  IMUX40 U193 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n377), .S1(i_addr_Rt[1]), .Q(n176) );
  IMUX40 U194 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n377), .S1(n375), .Q(n184) );
  IMUX40 U195 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n377), .S1(i_addr_Rt[1]), .Q(n182) );
  IMUX40 U196 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n378), .S1(n371), .Q(n189) );
  IMUX40 U197 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n378), .S1(n371), .Q(n187) );
  IMUX40 U198 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n378), .S1(n371), .Q(n186) );
  IMUX40 U199 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n378), .S1(n371), .Q(n194) );
  IMUX40 U200 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n378), .S1(n371), .Q(n192) );
  IMUX40 U201 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n378), .S1(n371), .Q(n199) );
  IMUX40 U202 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n378), .S1(i_addr_Rt[1]), .Q(n197) );
  IMUX40 U203 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n378), .S1(i_addr_Rt[1]), .Q(n196) );
  IMUX40 U204 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n380), .S1(i_addr_Rt[1]), .Q(n204) );
  IMUX40 U205 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n382), .S1(i_addr_Rt[1]), .Q(n202) );
  IMUX40 U206 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n384), .S1(n371), .Q(n209) );
  IMUX40 U207 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n384), .S1(i_addr_Rt[1]), .Q(n207) );
  IMUX40 U208 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n384), .S1(n372), .Q(n206) );
  IMUX40 U209 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n379), .S1(n373), .Q(n214) );
  IMUX40 U210 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n380), .S1(n369), .Q(n212) );
  IMUX40 U211 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n383), .S1(n372), .Q(n219) );
  IMUX40 U212 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(i_addr_Rt[0]), .S1(n372), .Q(n217) );
  IMUX40 U213 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n379), .S1(n370), .Q(n216) );
  IMUX40 U214 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n382), .S1(n370), .Q(n224) );
  IMUX40 U215 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n378), .S1(n370), .Q(n222) );
  IMUX40 U216 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n229) );
  IMUX40 U217 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n227) );
  IMUX40 U218 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n385), .S1(n370), .Q(n226) );
  IMUX40 U219 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n379), .S1(n370), .Q(n234) );
  IMUX40 U220 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n379), .S1(n370), .Q(n232) );
  IMUX40 U221 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n379), .S1(n370), .Q(n239) );
  IMUX40 U222 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n379), .S1(n370), .Q(n237) );
  IMUX40 U223 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n379), .S1(n370), .Q(n236) );
  IMUX40 U224 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n379), .S1(n370), .Q(n244) );
  IMUX40 U225 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n379), .S1(n372), .Q(n242) );
  IMUX40 U226 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n380), .S1(n369), .Q(n249) );
  IMUX40 U227 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n380), .S1(n375), .Q(n247) );
  IMUX40 U228 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n380), .S1(n375), .Q(n246) );
  IMUX40 U229 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n380), .S1(n375), .Q(n254) );
  IMUX40 U230 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n380), .S1(n370), .Q(n252) );
  IMUX40 U231 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n380), .S1(n369), .Q(n259) );
  IMUX40 U232 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n380), .S1(n370), .Q(n257) );
  IMUX40 U233 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n380), .S1(n372), .Q(n256) );
  IMUX40 U234 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n379), .S1(n370), .Q(n264) );
  IMUX40 U235 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n385), .S1(n370), .Q(n262) );
  IMUX40 U236 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n380), .S1(n371), .Q(n269) );
  IMUX40 U237 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n385), .S1(n371), .Q(n267) );
  IMUX40 U238 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n376), .S1(n371), .Q(n266) );
  IMUX40 U239 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n387), .S1(n371), .Q(n274) );
  IMUX40 U240 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n379), .S1(n371), .Q(n272) );
  IMUX40 U241 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n381), .S1(n369), .Q(n279) );
  IMUX40 U242 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n381), .S1(n369), .Q(n277) );
  IMUX40 U243 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n381), .S1(n369), .Q(n276) );
  IMUX40 U244 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n381), .S1(n373), .Q(n284) );
  IMUX40 U245 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n381), .S1(n373), .Q(n282) );
  IMUX40 U246 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n381), .S1(n372), .Q(n289) );
  IMUX40 U247 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n381), .S1(n369), .Q(n287) );
  IMUX40 U248 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n381), .S1(n373), .Q(n286) );
  IMUX40 U249 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n382), .S1(n372), .Q(n294) );
  IMUX40 U250 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n382), .S1(n372), .Q(n292) );
  IMUX40 U251 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(n382), .S1(n373), .Q(n299) );
  IMUX40 U252 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n382), .S1(n372), .Q(n297) );
  IMUX40 U253 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(n382), .S1(n374), .Q(n296) );
  IMUX40 U254 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(n382), .S1(n374), .Q(n304) );
  IMUX40 U255 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n382), .S1(n372), .Q(n302) );
  IMUX40 U256 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n386), .S1(n371), .Q(n309) );
  IMUX40 U257 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n385), .S1(n372), .Q(n307) );
  IMUX40 U258 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n378), .S1(n372), .Q(n306) );
  IMUX40 U259 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n376), .S1(n372), .Q(n314) );
  IMUX40 U260 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n377), .S1(n372), .Q(n312) );
  IMUX40 U261 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n377), .S1(n372), .Q(n319) );
  IMUX40 U262 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n384), .S1(n372), .Q(n317) );
  IMUX40 U263 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n381), .S1(n372), .Q(n316) );
  IMUX40 U264 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n383), .S1(n374), .Q(n324) );
  IMUX40 U265 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n383), .S1(n373), .Q(n322) );
  IMUX40 U266 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n383), .S1(n370), .Q(n329) );
  IMUX40 U267 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n383), .S1(n369), .Q(n327) );
  IMUX40 U268 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n383), .S1(n374), .Q(n326) );
  IMUX40 U269 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n383), .S1(n373), .Q(n334) );
  IMUX40 U270 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n383), .S1(n374), .Q(n332) );
  IMUX40 U271 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n384), .S1(n372), .Q(n339) );
  IMUX40 U272 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n384), .S1(n372), .Q(n337) );
  IMUX40 U273 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n384), .S1(n369), .Q(n336) );
  IMUX40 U274 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n384), .S1(n374), .Q(n344) );
  IMUX40 U275 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n384), .S1(n369), .Q(n342) );
  IMUX40 U276 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n384), .S1(n373), .Q(n349) );
  IMUX40 U277 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n384), .S1(n373), .Q(n347) );
  IMUX40 U278 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n384), .S1(n373), .Q(n346) );
  IMUX40 U279 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(i_addr_Rt[0]), .S1(n373), .Q(n354) );
  IMUX40 U280 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(i_addr_Rt[0]), .S1(n373), .Q(n352) );
  IMUX40 U281 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n384), .S1(n374), .Q(n359) );
  IMUX40 U282 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n387), .S1(n374), .Q(n357) );
  IMUX40 U283 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n356) );
  IMUX40 U284 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n364) );
  IMUX40 U285 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n362) );
  IMUX40 U286 ( .A(regs[384]), .B(regs[416]), .C(regs[448]), .D(regs[480]), 
        .S0(n728), .S1(n712), .Q(n397) );
  IMUX40 U287 ( .A(regs[256]), .B(regs[288]), .C(regs[320]), .D(regs[352]), 
        .S0(n727), .S1(n713), .Q(n395) );
  IMUX40 U288 ( .A(regs[0]), .B(regs[32]), .C(regs[64]), .D(regs[96]), .S0(
        n725), .S1(i_addr_Rs[1]), .Q(n394) );
  IMUX40 U289 ( .A(regs[896]), .B(regs[928]), .C(regs[960]), .D(regs[992]), 
        .S0(n725), .S1(n713), .Q(n392) );
  IMUX40 U290 ( .A(regs[768]), .B(regs[800]), .C(regs[832]), .D(regs[864]), 
        .S0(n726), .S1(n714), .Q(n390) );
  IMUX40 U291 ( .A(regs[512]), .B(regs[544]), .C(regs[576]), .D(regs[608]), 
        .S0(n726), .S1(n714), .Q(n389) );
  IMUX40 U292 ( .A(regs[897]), .B(regs[929]), .C(regs[961]), .D(regs[993]), 
        .S0(n727), .S1(n714), .Q(n402) );
  IMUX40 U293 ( .A(regs[769]), .B(regs[801]), .C(regs[833]), .D(regs[865]), 
        .S0(n729), .S1(n714), .Q(n400) );
  IMUX40 U294 ( .A(regs[513]), .B(regs[545]), .C(regs[577]), .D(regs[609]), 
        .S0(n730), .S1(i_addr_Rs[1]), .Q(n399) );
  IMUX40 U295 ( .A(regs[385]), .B(regs[417]), .C(regs[449]), .D(regs[481]), 
        .S0(n728), .S1(n715), .Q(n407) );
  IMUX40 U296 ( .A(regs[257]), .B(regs[289]), .C(regs[321]), .D(regs[353]), 
        .S0(n729), .S1(n712), .Q(n405) );
  IMUX40 U297 ( .A(regs[898]), .B(regs[930]), .C(regs[962]), .D(regs[994]), 
        .S0(n730), .S1(n713), .Q(n412) );
  IMUX40 U298 ( .A(regs[770]), .B(regs[802]), .C(regs[834]), .D(regs[866]), 
        .S0(n726), .S1(n713), .Q(n410) );
  IMUX40 U299 ( .A(regs[514]), .B(regs[546]), .C(regs[578]), .D(regs[610]), 
        .S0(n727), .S1(n712), .Q(n409) );
  IMUX40 U300 ( .A(regs[386]), .B(regs[418]), .C(regs[450]), .D(regs[482]), 
        .S0(n728), .S1(n712), .Q(n417) );
  IMUX40 U301 ( .A(regs[258]), .B(regs[290]), .C(regs[322]), .D(regs[354]), 
        .S0(n728), .S1(n716), .Q(n415) );
  IMUX40 U302 ( .A(regs[899]), .B(regs[931]), .C(regs[963]), .D(regs[995]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n422) );
  IMUX40 U303 ( .A(regs[771]), .B(regs[803]), .C(regs[835]), .D(regs[867]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n420) );
  IMUX40 U304 ( .A(regs[515]), .B(regs[547]), .C(regs[579]), .D(regs[611]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n419) );
  IMUX40 U305 ( .A(regs[387]), .B(regs[419]), .C(regs[451]), .D(regs[483]), 
        .S0(i_addr_Rs[0]), .S1(n716), .Q(n427) );
  IMUX40 U306 ( .A(regs[259]), .B(regs[291]), .C(regs[323]), .D(regs[355]), 
        .S0(n724), .S1(i_addr_Rs[1]), .Q(n425) );
  IMUX40 U307 ( .A(regs[900]), .B(regs[932]), .C(regs[964]), .D(regs[996]), 
        .S0(n725), .S1(n713), .Q(n432) );
  IMUX40 U308 ( .A(regs[772]), .B(regs[804]), .C(regs[836]), .D(regs[868]), 
        .S0(n727), .S1(n713), .Q(n430) );
  IMUX40 U309 ( .A(regs[516]), .B(regs[548]), .C(regs[580]), .D(regs[612]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n429) );
  IMUX40 U310 ( .A(regs[388]), .B(regs[420]), .C(regs[452]), .D(regs[484]), 
        .S0(n730), .S1(n714), .Q(n437) );
  IMUX40 U311 ( .A(regs[260]), .B(regs[292]), .C(regs[324]), .D(regs[356]), 
        .S0(n719), .S1(n713), .Q(n435) );
  IMUX40 U312 ( .A(regs[901]), .B(regs[933]), .C(regs[965]), .D(regs[997]), 
        .S0(i_addr_Rs[0]), .S1(n716), .Q(n442) );
  IMUX40 U313 ( .A(regs[773]), .B(regs[805]), .C(regs[837]), .D(regs[869]), 
        .S0(n727), .S1(n714), .Q(n440) );
  IMUX40 U314 ( .A(regs[517]), .B(regs[549]), .C(regs[581]), .D(regs[613]), 
        .S0(i_addr_Rs[0]), .S1(n715), .Q(n439) );
  IMUX40 U315 ( .A(regs[389]), .B(regs[421]), .C(regs[453]), .D(regs[485]), 
        .S0(i_addr_Rs[0]), .S1(n713), .Q(n447) );
  IMUX40 U316 ( .A(regs[261]), .B(regs[293]), .C(regs[325]), .D(regs[357]), 
        .S0(i_addr_Rs[0]), .S1(n713), .Q(n445) );
  IMUX40 U317 ( .A(regs[902]), .B(regs[934]), .C(regs[966]), .D(regs[998]), 
        .S0(n729), .S1(n715), .Q(n452) );
  IMUX40 U318 ( .A(regs[774]), .B(regs[806]), .C(regs[838]), .D(regs[870]), 
        .S0(n723), .S1(n714), .Q(n450) );
  IMUX40 U319 ( .A(regs[518]), .B(regs[550]), .C(regs[582]), .D(regs[614]), 
        .S0(i_addr_Rs[0]), .S1(n714), .Q(n449) );
  IMUX40 U320 ( .A(regs[390]), .B(regs[422]), .C(regs[454]), .D(regs[486]), 
        .S0(n728), .S1(n714), .Q(n457) );
  IMUX40 U321 ( .A(regs[262]), .B(regs[294]), .C(regs[326]), .D(regs[358]), 
        .S0(n729), .S1(i_addr_Rs[1]), .Q(n455) );
  IMUX40 U322 ( .A(regs[903]), .B(regs[935]), .C(regs[967]), .D(regs[999]), 
        .S0(n727), .S1(n713), .Q(n462) );
  IMUX40 U323 ( .A(regs[775]), .B(regs[807]), .C(regs[839]), .D(regs[871]), 
        .S0(n726), .S1(n713), .Q(n460) );
  IMUX40 U324 ( .A(regs[519]), .B(regs[551]), .C(regs[583]), .D(regs[615]), 
        .S0(n730), .S1(n716), .Q(n459) );
  IMUX40 U325 ( .A(regs[391]), .B(regs[423]), .C(regs[455]), .D(regs[487]), 
        .S0(n724), .S1(n716), .Q(n467) );
  IMUX40 U326 ( .A(regs[263]), .B(regs[295]), .C(regs[327]), .D(regs[359]), 
        .S0(n727), .S1(n713), .Q(n465) );
  IMUX40 U327 ( .A(regs[904]), .B(regs[936]), .C(regs[968]), .D(regs[1000]), 
        .S0(n720), .S1(n714), .Q(n472) );
  IMUX40 U328 ( .A(regs[776]), .B(regs[808]), .C(regs[840]), .D(regs[872]), 
        .S0(n723), .S1(n716), .Q(n470) );
  IMUX40 U329 ( .A(regs[520]), .B(regs[552]), .C(regs[584]), .D(regs[616]), 
        .S0(n729), .S1(n713), .Q(n469) );
  IMUX40 U330 ( .A(regs[392]), .B(regs[424]), .C(regs[456]), .D(regs[488]), 
        .S0(i_addr_Rs[0]), .S1(n717), .Q(n477) );
  IMUX40 U331 ( .A(regs[264]), .B(regs[296]), .C(regs[328]), .D(regs[360]), 
        .S0(n725), .S1(n714), .Q(n475) );
  IMUX40 U332 ( .A(regs[905]), .B(regs[937]), .C(regs[969]), .D(regs[1001]), 
        .S0(n720), .S1(i_addr_Rs[1]), .Q(n482) );
  IMUX40 U333 ( .A(regs[777]), .B(regs[809]), .C(regs[841]), .D(regs[873]), 
        .S0(n719), .S1(n713), .Q(n480) );
  IMUX40 U334 ( .A(regs[521]), .B(regs[553]), .C(regs[585]), .D(regs[617]), 
        .S0(n722), .S1(n712), .Q(n479) );
  IMUX40 U335 ( .A(regs[393]), .B(regs[425]), .C(regs[457]), .D(regs[489]), 
        .S0(n727), .S1(i_addr_Rs[1]), .Q(n487) );
  IMUX40 U336 ( .A(regs[265]), .B(regs[297]), .C(regs[329]), .D(regs[361]), 
        .S0(n730), .S1(i_addr_Rs[1]), .Q(n485) );
  IMUX40 U337 ( .A(regs[906]), .B(regs[938]), .C(regs[970]), .D(regs[1002]), 
        .S0(n723), .S1(i_addr_Rs[1]), .Q(n492) );
  IMUX40 U338 ( .A(regs[778]), .B(regs[810]), .C(regs[842]), .D(regs[874]), 
        .S0(n727), .S1(n716), .Q(n490) );
  IMUX40 U339 ( .A(regs[522]), .B(regs[554]), .C(regs[586]), .D(regs[618]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n489) );
  IMUX40 U340 ( .A(regs[394]), .B(regs[426]), .C(regs[458]), .D(regs[490]), 
        .S0(i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n497) );
  IMUX40 U341 ( .A(regs[266]), .B(regs[298]), .C(regs[330]), .D(regs[362]), 
        .S0(n725), .S1(n713), .Q(n495) );
  IMUX40 U342 ( .A(regs[907]), .B(regs[939]), .C(regs[971]), .D(regs[1003]), 
        .S0(n719), .S1(n716), .Q(n502) );
  IMUX40 U343 ( .A(regs[779]), .B(regs[811]), .C(regs[843]), .D(regs[875]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n500) );
  IMUX40 U344 ( .A(regs[523]), .B(regs[555]), .C(regs[587]), .D(regs[619]), 
        .S0(n719), .S1(n717), .Q(n499) );
  IMUX40 U345 ( .A(regs[395]), .B(regs[427]), .C(regs[459]), .D(regs[491]), 
        .S0(n719), .S1(n715), .Q(n507) );
  IMUX40 U346 ( .A(regs[267]), .B(regs[299]), .C(regs[331]), .D(regs[363]), 
        .S0(n719), .S1(n712), .Q(n505) );
  IMUX40 U347 ( .A(regs[908]), .B(regs[940]), .C(regs[972]), .D(regs[1004]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n512) );
  IMUX40 U348 ( .A(regs[780]), .B(regs[812]), .C(regs[844]), .D(regs[876]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n510) );
  IMUX40 U349 ( .A(regs[524]), .B(regs[556]), .C(regs[588]), .D(regs[620]), 
        .S0(n719), .S1(n718), .Q(n509) );
  IMUX40 U350 ( .A(regs[396]), .B(regs[428]), .C(regs[460]), .D(regs[492]), 
        .S0(n720), .S1(i_addr_Rs[1]), .Q(n517) );
  IMUX40 U351 ( .A(regs[268]), .B(regs[300]), .C(regs[332]), .D(regs[364]), 
        .S0(n720), .S1(n712), .Q(n515) );
  IMUX40 U352 ( .A(regs[909]), .B(regs[941]), .C(regs[973]), .D(regs[1005]), 
        .S0(n720), .S1(n718), .Q(n522) );
  IMUX40 U353 ( .A(regs[781]), .B(regs[813]), .C(regs[845]), .D(regs[877]), 
        .S0(n720), .S1(n712), .Q(n520) );
  IMUX40 U354 ( .A(regs[525]), .B(regs[557]), .C(regs[589]), .D(regs[621]), 
        .S0(n720), .S1(n714), .Q(n519) );
  IMUX40 U355 ( .A(regs[397]), .B(regs[429]), .C(regs[461]), .D(regs[493]), 
        .S0(n720), .S1(n718), .Q(n527) );
  IMUX40 U356 ( .A(regs[269]), .B(regs[301]), .C(regs[333]), .D(regs[365]), 
        .S0(n720), .S1(n714), .Q(n525) );
  IMUX40 U357 ( .A(regs[910]), .B(regs[942]), .C(regs[974]), .D(regs[1006]), 
        .S0(n721), .S1(n715), .Q(n532) );
  IMUX40 U358 ( .A(regs[782]), .B(regs[814]), .C(regs[846]), .D(regs[878]), 
        .S0(n721), .S1(n717), .Q(n530) );
  IMUX40 U359 ( .A(regs[526]), .B(regs[558]), .C(regs[590]), .D(regs[622]), 
        .S0(n721), .S1(n714), .Q(n529) );
  IMUX40 U360 ( .A(regs[398]), .B(regs[430]), .C(regs[462]), .D(regs[494]), 
        .S0(n721), .S1(n717), .Q(n537) );
  IMUX40 U361 ( .A(regs[270]), .B(regs[302]), .C(regs[334]), .D(regs[366]), 
        .S0(n721), .S1(n715), .Q(n535) );
  IMUX40 U362 ( .A(regs[911]), .B(regs[943]), .C(regs[975]), .D(regs[1007]), 
        .S0(n721), .S1(n712), .Q(n542) );
  IMUX40 U363 ( .A(regs[783]), .B(regs[815]), .C(regs[847]), .D(regs[879]), 
        .S0(n721), .S1(i_addr_Rs[1]), .Q(n540) );
  IMUX40 U364 ( .A(regs[527]), .B(regs[559]), .C(regs[591]), .D(regs[623]), 
        .S0(n721), .S1(i_addr_Rs[1]), .Q(n539) );
  IMUX40 U365 ( .A(regs[399]), .B(regs[431]), .C(regs[463]), .D(regs[495]), 
        .S0(n722), .S1(i_addr_Rs[1]), .Q(n547) );
  IMUX40 U366 ( .A(regs[271]), .B(regs[303]), .C(regs[335]), .D(regs[367]), 
        .S0(n722), .S1(i_addr_Rs[1]), .Q(n545) );
  IMUX40 U367 ( .A(regs[912]), .B(regs[944]), .C(regs[976]), .D(regs[1008]), 
        .S0(n722), .S1(n712), .Q(n552) );
  IMUX40 U368 ( .A(regs[784]), .B(regs[816]), .C(regs[848]), .D(regs[880]), 
        .S0(n722), .S1(n713), .Q(n550) );
  IMUX40 U369 ( .A(regs[528]), .B(regs[560]), .C(regs[592]), .D(regs[624]), 
        .S0(n722), .S1(i_addr_Rs[1]), .Q(n549) );
  IMUX40 U370 ( .A(regs[400]), .B(regs[432]), .C(regs[464]), .D(regs[496]), 
        .S0(n722), .S1(i_addr_Rs[1]), .Q(n557) );
  IMUX40 U371 ( .A(regs[272]), .B(regs[304]), .C(regs[336]), .D(regs[368]), 
        .S0(n722), .S1(i_addr_Rs[1]), .Q(n555) );
  IMUX40 U372 ( .A(regs[913]), .B(regs[945]), .C(regs[977]), .D(regs[1009]), 
        .S0(n723), .S1(n714), .Q(n562) );
  IMUX40 U373 ( .A(regs[785]), .B(regs[817]), .C(regs[849]), .D(regs[881]), 
        .S0(n723), .S1(n713), .Q(n560) );
  IMUX40 U374 ( .A(regs[529]), .B(regs[561]), .C(regs[593]), .D(regs[625]), 
        .S0(n723), .S1(n714), .Q(n559) );
  IMUX40 U375 ( .A(regs[401]), .B(regs[433]), .C(regs[465]), .D(regs[497]), 
        .S0(n723), .S1(n714), .Q(n567) );
  IMUX40 U376 ( .A(regs[273]), .B(regs[305]), .C(regs[337]), .D(regs[369]), 
        .S0(n723), .S1(n712), .Q(n565) );
  IMUX40 U377 ( .A(regs[914]), .B(regs[946]), .C(regs[978]), .D(regs[1010]), 
        .S0(n723), .S1(n713), .Q(n572) );
  IMUX40 U378 ( .A(regs[786]), .B(regs[818]), .C(regs[850]), .D(regs[882]), 
        .S0(n723), .S1(n717), .Q(n570) );
  IMUX40 U379 ( .A(regs[530]), .B(regs[562]), .C(regs[594]), .D(regs[626]), 
        .S0(n723), .S1(n713), .Q(n569) );
  IMUX40 U380 ( .A(regs[402]), .B(regs[434]), .C(regs[466]), .D(regs[498]), 
        .S0(n727), .S1(n715), .Q(n577) );
  IMUX40 U381 ( .A(regs[274]), .B(regs[306]), .C(regs[338]), .D(regs[370]), 
        .S0(n730), .S1(n715), .Q(n575) );
  IMUX40 U382 ( .A(regs[915]), .B(regs[947]), .C(regs[979]), .D(regs[1011]), 
        .S0(n719), .S1(n715), .Q(n582) );
  IMUX40 U383 ( .A(regs[787]), .B(regs[819]), .C(regs[851]), .D(regs[883]), 
        .S0(n720), .S1(n715), .Q(n580) );
  IMUX40 U384 ( .A(regs[531]), .B(regs[563]), .C(regs[595]), .D(regs[627]), 
        .S0(n724), .S1(n714), .Q(n579) );
  IMUX40 U385 ( .A(regs[403]), .B(regs[435]), .C(regs[467]), .D(regs[499]), 
        .S0(n724), .S1(n712), .Q(n587) );
  IMUX40 U386 ( .A(regs[275]), .B(regs[307]), .C(regs[339]), .D(regs[371]), 
        .S0(n726), .S1(n715), .Q(n585) );
  IMUX40 U387 ( .A(regs[916]), .B(regs[948]), .C(regs[980]), .D(regs[1012]), 
        .S0(n729), .S1(n715), .Q(n592) );
  IMUX40 U388 ( .A(regs[788]), .B(regs[820]), .C(regs[852]), .D(regs[884]), 
        .S0(n730), .S1(n713), .Q(n590) );
  IMUX40 U389 ( .A(regs[532]), .B(regs[564]), .C(regs[596]), .D(regs[628]), 
        .S0(n723), .S1(i_addr_Rs[1]), .Q(n589) );
  IMUX40 U390 ( .A(regs[404]), .B(regs[436]), .C(regs[468]), .D(regs[500]), 
        .S0(n728), .S1(n712), .Q(n597) );
  IMUX40 U391 ( .A(regs[276]), .B(regs[308]), .C(regs[340]), .D(regs[372]), 
        .S0(n728), .S1(n718), .Q(n595) );
  IMUX40 U392 ( .A(regs[917]), .B(regs[949]), .C(regs[981]), .D(regs[1013]), 
        .S0(n728), .S1(n712), .Q(n602) );
  IMUX40 U393 ( .A(regs[789]), .B(regs[821]), .C(regs[853]), .D(regs[885]), 
        .S0(n728), .S1(n712), .Q(n600) );
  IMUX40 U394 ( .A(regs[533]), .B(regs[565]), .C(regs[597]), .D(regs[629]), 
        .S0(n721), .S1(n713), .Q(n599) );
  IMUX40 U395 ( .A(regs[405]), .B(regs[437]), .C(regs[469]), .D(regs[501]), 
        .S0(n729), .S1(n713), .Q(n607) );
  IMUX40 U396 ( .A(regs[277]), .B(regs[309]), .C(regs[341]), .D(regs[373]), 
        .S0(n727), .S1(i_addr_Rs[1]), .Q(n605) );
  IMUX40 U397 ( .A(regs[918]), .B(regs[950]), .C(regs[982]), .D(regs[1014]), 
        .S0(n728), .S1(n715), .Q(n612) );
  IMUX40 U398 ( .A(regs[790]), .B(regs[822]), .C(regs[854]), .D(regs[886]), 
        .S0(n728), .S1(n715), .Q(n610) );
  IMUX40 U399 ( .A(regs[534]), .B(regs[566]), .C(regs[598]), .D(regs[630]), 
        .S0(n727), .S1(n715), .Q(n609) );
  IMUX40 U400 ( .A(regs[406]), .B(regs[438]), .C(regs[470]), .D(regs[502]), 
        .S0(n730), .S1(n715), .Q(n617) );
  IMUX40 U401 ( .A(regs[278]), .B(regs[310]), .C(regs[342]), .D(regs[374]), 
        .S0(n729), .S1(n715), .Q(n615) );
  IMUX40 U402 ( .A(regs[919]), .B(regs[951]), .C(regs[983]), .D(regs[1015]), 
        .S0(n724), .S1(n714), .Q(n622) );
  IMUX40 U403 ( .A(regs[791]), .B(regs[823]), .C(regs[855]), .D(regs[887]), 
        .S0(n724), .S1(n717), .Q(n620) );
  IMUX40 U404 ( .A(regs[535]), .B(regs[567]), .C(regs[599]), .D(regs[631]), 
        .S0(n724), .S1(n714), .Q(n619) );
  IMUX40 U405 ( .A(regs[407]), .B(regs[439]), .C(regs[471]), .D(regs[503]), 
        .S0(n724), .S1(n712), .Q(n627) );
  IMUX40 U406 ( .A(regs[279]), .B(regs[311]), .C(regs[343]), .D(regs[375]), 
        .S0(n724), .S1(n712), .Q(n625) );
  IMUX40 U407 ( .A(regs[920]), .B(regs[952]), .C(regs[984]), .D(regs[1016]), 
        .S0(n724), .S1(n712), .Q(n632) );
  IMUX40 U408 ( .A(regs[792]), .B(regs[824]), .C(regs[856]), .D(regs[888]), 
        .S0(n724), .S1(n712), .Q(n630) );
  IMUX40 U409 ( .A(regs[536]), .B(regs[568]), .C(regs[600]), .D(regs[632]), 
        .S0(n724), .S1(n714), .Q(n629) );
  IMUX40 U410 ( .A(regs[408]), .B(regs[440]), .C(regs[472]), .D(regs[504]), 
        .S0(n730), .S1(n717), .Q(n637) );
  IMUX40 U411 ( .A(regs[280]), .B(regs[312]), .C(regs[344]), .D(regs[376]), 
        .S0(n722), .S1(n712), .Q(n635) );
  IMUX40 U412 ( .A(regs[921]), .B(regs[953]), .C(regs[985]), .D(regs[1017]), 
        .S0(i_addr_Rs[0]), .S1(n716), .Q(n642) );
  IMUX40 U413 ( .A(regs[793]), .B(regs[825]), .C(regs[857]), .D(regs[889]), 
        .S0(n728), .S1(n714), .Q(n640) );
  IMUX40 U414 ( .A(regs[537]), .B(regs[569]), .C(regs[601]), .D(regs[633]), 
        .S0(i_addr_Rs[0]), .S1(n714), .Q(n639) );
  IMUX40 U415 ( .A(regs[409]), .B(regs[441]), .C(regs[473]), .D(regs[505]), 
        .S0(i_addr_Rs[0]), .S1(n716), .Q(n647) );
  IMUX40 U416 ( .A(regs[281]), .B(regs[313]), .C(regs[345]), .D(regs[377]), 
        .S0(n729), .S1(n712), .Q(n645) );
  IMUX40 U417 ( .A(regs[922]), .B(regs[954]), .C(regs[986]), .D(regs[1018]), 
        .S0(n722), .S1(n718), .Q(n652) );
  IMUX40 U418 ( .A(regs[794]), .B(regs[826]), .C(regs[858]), .D(regs[890]), 
        .S0(n721), .S1(n714), .Q(n650) );
  IMUX40 U419 ( .A(regs[538]), .B(regs[570]), .C(regs[602]), .D(regs[634]), 
        .S0(n729), .S1(n716), .Q(n649) );
  IMUX40 U420 ( .A(regs[410]), .B(regs[442]), .C(regs[474]), .D(regs[506]), 
        .S0(n721), .S1(n716), .Q(n657) );
  IMUX40 U421 ( .A(regs[282]), .B(regs[314]), .C(regs[346]), .D(regs[378]), 
        .S0(n722), .S1(n716), .Q(n655) );
  IMUX40 U422 ( .A(regs[923]), .B(regs[955]), .C(regs[987]), .D(regs[1019]), 
        .S0(n723), .S1(n716), .Q(n662) );
  IMUX40 U423 ( .A(regs[795]), .B(regs[827]), .C(regs[859]), .D(regs[891]), 
        .S0(n729), .S1(n716), .Q(n660) );
  IMUX40 U424 ( .A(regs[539]), .B(regs[571]), .C(regs[603]), .D(regs[635]), 
        .S0(n719), .S1(n716), .Q(n659) );
  IMUX40 U425 ( .A(regs[411]), .B(regs[443]), .C(regs[475]), .D(regs[507]), 
        .S0(n725), .S1(n717), .Q(n667) );
  IMUX40 U426 ( .A(regs[283]), .B(regs[315]), .C(regs[347]), .D(regs[379]), 
        .S0(n725), .S1(n717), .Q(n665) );
  IMUX40 U427 ( .A(regs[924]), .B(regs[956]), .C(regs[988]), .D(regs[1020]), 
        .S0(n725), .S1(n718), .Q(n672) );
  IMUX40 U428 ( .A(regs[796]), .B(regs[828]), .C(regs[860]), .D(regs[892]), 
        .S0(n725), .S1(n717), .Q(n670) );
  IMUX40 U429 ( .A(regs[540]), .B(regs[572]), .C(regs[604]), .D(regs[636]), 
        .S0(n725), .S1(n716), .Q(n669) );
  IMUX40 U430 ( .A(regs[412]), .B(regs[444]), .C(regs[476]), .D(regs[508]), 
        .S0(n725), .S1(n718), .Q(n677) );
  IMUX40 U431 ( .A(regs[284]), .B(regs[316]), .C(regs[348]), .D(regs[380]), 
        .S0(n725), .S1(n717), .Q(n675) );
  IMUX40 U432 ( .A(regs[925]), .B(regs[957]), .C(regs[989]), .D(regs[1021]), 
        .S0(n726), .S1(n717), .Q(n682) );
  IMUX40 U433 ( .A(regs[797]), .B(regs[829]), .C(regs[861]), .D(regs[893]), 
        .S0(n726), .S1(n718), .Q(n680) );
  IMUX40 U434 ( .A(regs[541]), .B(regs[573]), .C(regs[605]), .D(regs[637]), 
        .S0(n726), .S1(n717), .Q(n679) );
  IMUX40 U435 ( .A(regs[413]), .B(regs[445]), .C(regs[477]), .D(regs[509]), 
        .S0(n726), .S1(n718), .Q(n687) );
  IMUX40 U436 ( .A(regs[285]), .B(regs[317]), .C(regs[349]), .D(regs[381]), 
        .S0(n726), .S1(n718), .Q(n685) );
  IMUX40 U437 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n726), .S1(n717), .Q(n684) );
  IMUX40 U438 ( .A(regs[926]), .B(regs[958]), .C(regs[990]), .D(regs[1022]), 
        .S0(n726), .S1(n717), .Q(n692) );
  IMUX40 U439 ( .A(regs[798]), .B(regs[830]), .C(regs[862]), .D(regs[894]), 
        .S0(n726), .S1(n717), .Q(n690) );
  IMUX40 U440 ( .A(regs[542]), .B(regs[574]), .C(regs[606]), .D(regs[638]), 
        .S0(n726), .S1(n717), .Q(n689) );
  IMUX40 U441 ( .A(regs[414]), .B(regs[446]), .C(regs[478]), .D(regs[510]), 
        .S0(n723), .S1(n717), .Q(n697) );
  IMUX40 U442 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        n729), .S1(n718), .Q(n694) );
  IMUX40 U443 ( .A(regs[286]), .B(regs[318]), .C(regs[350]), .D(regs[382]), 
        .S0(n725), .S1(n717), .Q(n695) );
  IMUX40 U444 ( .A(regs[927]), .B(regs[959]), .C(regs[991]), .D(regs[1023]), 
        .S0(n724), .S1(n718), .Q(n702) );
  IMUX40 U445 ( .A(regs[799]), .B(regs[831]), .C(regs[863]), .D(regs[895]), 
        .S0(n720), .S1(n718), .Q(n700) );
  IMUX40 U446 ( .A(regs[543]), .B(regs[575]), .C(regs[607]), .D(regs[639]), 
        .S0(n728), .S1(n718), .Q(n699) );
  IMUX40 U447 ( .A(regs[415]), .B(regs[447]), .C(regs[479]), .D(regs[511]), 
        .S0(n726), .S1(n718), .Q(n707) );
  IMUX40 U448 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        i_addr_Rs[0]), .S1(n718), .Q(n704) );
  IMUX40 U449 ( .A(regs[287]), .B(regs[319]), .C(regs[351]), .D(regs[383]), 
        .S0(n724), .S1(n718), .Q(n705) );
  IMUX40 U450 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n386), .S1(n371), .Q(n9) );
  IMUX40 U451 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(i_addr_Rt[0]), .S1(n375), .Q(n4) );
  IMUX40 U452 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n386), .S1(n375), .Q(n14) );
  IMUX40 U453 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n387), .S1(n370), .Q(n19) );
  IMUX40 U454 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n386), .S1(n371), .Q(n24) );
  IMUX40 U455 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n386), .S1(n375), .Q(n29) );
  IMUX40 U456 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n385), .S1(n375), .Q(n34) );
  IMUX40 U457 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n386), .S1(n375), .Q(n83) );
  IMUX40 U458 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n376), .S1(n375), .Q(n88) );
  IMUX40 U459 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n387), .S1(n369), .Q(n93) );
  IMUX40 U460 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n377), .S1(n369), .Q(n98) );
  IMUX40 U461 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(n385), .S1(n369), .Q(n103) );
  IMUX40 U462 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n377), .S1(n369), .Q(n108) );
  IMUX40 U463 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n380), .S1(n369), .Q(n113) );
  IMUX40 U464 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n386), .S1(n375), .Q(n118) );
  IMUX40 U465 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n379), .S1(n373), .Q(n123) );
  IMUX40 U466 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n387), .S1(n375), .Q(n128) );
  IMUX40 U467 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n385), .S1(n370), .Q(n133) );
  IMUX40 U468 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n385), .S1(n375), .Q(n138) );
  IMUX40 U469 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n387), .S1(n372), .Q(n143) );
  IMUX40 U470 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n377), .S1(n372), .Q(n148) );
  IMUX40 U471 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n385), .S1(n369), .Q(n153) );
  IMUX40 U472 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n376), .S1(n372), .Q(n158) );
  IMUX40 U473 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n376), .S1(i_addr_Rt[1]), .Q(n163) );
  IMUX40 U474 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n376), .S1(n371), .Q(n168) );
  IMUX40 U475 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n377), .S1(n371), .Q(n173) );
  IMUX40 U476 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n377), .S1(n375), .Q(n178) );
  IMUX40 U477 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n377), .S1(n369), .Q(n183) );
  IMUX40 U478 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n378), .S1(n371), .Q(n188) );
  IMUX40 U479 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n378), .S1(n371), .Q(n193) );
  IMUX40 U480 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n378), .S1(n369), .Q(n198) );
  IMUX40 U481 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n381), .S1(i_addr_Rt[1]), .Q(n203) );
  IMUX40 U482 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n383), .S1(n370), .Q(n208) );
  IMUX40 U483 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n381), .S1(n374), .Q(n213) );
  IMUX40 U484 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n377), .S1(n375), .Q(n218) );
  IMUX40 U485 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(i_addr_Rt[0]), .S1(n370), .Q(n223) );
  IMUX40 U486 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n386), .S1(n370), .Q(n228) );
  IMUX40 U487 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n379), .S1(n370), .Q(n233) );
  IMUX40 U488 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n379), .S1(n370), .Q(n238) );
  IMUX40 U489 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n379), .S1(n371), .Q(n243) );
  IMUX40 U490 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n380), .S1(n375), .Q(n248) );
  IMUX40 U491 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n380), .S1(n372), .Q(n253) );
  IMUX40 U492 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n380), .S1(n370), .Q(n258) );
  IMUX40 U493 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n385), .S1(n372), .Q(n263) );
  IMUX40 U494 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n379), .S1(n371), .Q(n268) );
  IMUX40 U495 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n383), .S1(n371), .Q(n273) );
  IMUX40 U496 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n381), .S1(n369), .Q(n278) );
  IMUX40 U497 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n381), .S1(n372), .Q(n283) );
  IMUX40 U498 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n381), .S1(n372), .Q(n288) );
  IMUX40 U499 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n382), .S1(n373), .Q(n293) );
  IMUX40 U500 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n382), .S1(n371), .Q(n298) );
  IMUX40 U501 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(n382), .S1(n374), .Q(n303) );
  IMUX40 U502 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n381), .S1(n371), .Q(n308) );
  IMUX40 U503 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n378), .S1(n372), .Q(n313) );
  IMUX40 U504 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n382), .S1(n372), .Q(n318) );
  IMUX40 U505 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n383), .S1(n373), .Q(n323) );
  IMUX40 U506 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n383), .S1(n369), .Q(n328) );
  IMUX40 U507 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n383), .S1(n374), .Q(n333) );
  IMUX40 U508 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n384), .S1(n369), .Q(n338) );
  IMUX40 U509 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n384), .S1(n373), .Q(n343) );
  IMUX40 U510 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n384), .S1(n373), .Q(n348) );
  IMUX40 U511 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(i_addr_Rt[0]), .S1(n373), .Q(n353) );
  IMUX40 U512 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n383), .S1(n374), .Q(n358) );
  IMUX40 U513 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(i_addr_Rt[0]), .S1(n374), .Q(n363) );
  IMUX40 U514 ( .A(regs[128]), .B(regs[160]), .C(regs[192]), .D(regs[224]), 
        .S0(n729), .S1(i_addr_Rs[1]), .Q(n396) );
  IMUX40 U515 ( .A(regs[640]), .B(regs[672]), .C(regs[704]), .D(regs[736]), 
        .S0(n721), .S1(n716), .Q(n391) );
  IMUX40 U516 ( .A(regs[641]), .B(regs[673]), .C(regs[705]), .D(regs[737]), 
        .S0(n730), .S1(n718), .Q(n401) );
  IMUX40 U517 ( .A(regs[129]), .B(regs[161]), .C(regs[193]), .D(regs[225]), 
        .S0(n730), .S1(n717), .Q(n406) );
  IMUX40 U518 ( .A(regs[642]), .B(regs[674]), .C(regs[706]), .D(regs[738]), 
        .S0(n727), .S1(n716), .Q(n411) );
  IMUX40 U519 ( .A(regs[130]), .B(regs[162]), .C(regs[194]), .D(regs[226]), 
        .S0(n720), .S1(n714), .Q(n416) );
  IMUX40 U520 ( .A(regs[643]), .B(regs[675]), .C(regs[707]), .D(regs[739]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n421) );
  IMUX40 U521 ( .A(regs[131]), .B(regs[163]), .C(regs[195]), .D(regs[227]), 
        .S0(n728), .S1(n716), .Q(n426) );
  IMUX40 U522 ( .A(regs[644]), .B(regs[676]), .C(regs[708]), .D(regs[740]), 
        .S0(n722), .S1(n713), .Q(n431) );
  IMUX40 U523 ( .A(regs[132]), .B(regs[164]), .C(regs[196]), .D(regs[228]), 
        .S0(n722), .S1(n718), .Q(n436) );
  IMUX40 U524 ( .A(regs[645]), .B(regs[677]), .C(regs[709]), .D(regs[741]), 
        .S0(n722), .S1(n712), .Q(n441) );
  IMUX40 U525 ( .A(regs[133]), .B(regs[165]), .C(regs[197]), .D(regs[229]), 
        .S0(i_addr_Rs[0]), .S1(n712), .Q(n446) );
  IMUX40 U526 ( .A(regs[646]), .B(regs[678]), .C(regs[710]), .D(regs[742]), 
        .S0(n724), .S1(n712), .Q(n451) );
  IMUX40 U527 ( .A(regs[134]), .B(regs[166]), .C(regs[198]), .D(regs[230]), 
        .S0(n719), .S1(n716), .Q(n456) );
  IMUX40 U528 ( .A(regs[647]), .B(regs[679]), .C(regs[711]), .D(regs[743]), 
        .S0(n720), .S1(n714), .Q(n461) );
  IMUX40 U529 ( .A(regs[135]), .B(regs[167]), .C(regs[199]), .D(regs[231]), 
        .S0(n728), .S1(n714), .Q(n466) );
  IMUX40 U530 ( .A(regs[648]), .B(regs[680]), .C(regs[712]), .D(regs[744]), 
        .S0(n721), .S1(i_addr_Rs[1]), .Q(n471) );
  IMUX40 U531 ( .A(regs[136]), .B(regs[168]), .C(regs[200]), .D(regs[232]), 
        .S0(n730), .S1(n715), .Q(n476) );
  IMUX40 U532 ( .A(regs[649]), .B(regs[681]), .C(regs[713]), .D(regs[745]), 
        .S0(n719), .S1(n713), .Q(n481) );
  IMUX40 U533 ( .A(regs[137]), .B(regs[169]), .C(regs[201]), .D(regs[233]), 
        .S0(n721), .S1(i_addr_Rs[1]), .Q(n486) );
  IMUX40 U534 ( .A(regs[650]), .B(regs[682]), .C(regs[714]), .D(regs[746]), 
        .S0(n720), .S1(n715), .Q(n491) );
  IMUX40 U535 ( .A(regs[138]), .B(regs[170]), .C(regs[202]), .D(regs[234]), 
        .S0(n723), .S1(n714), .Q(n496) );
  IMUX40 U536 ( .A(regs[651]), .B(regs[683]), .C(regs[715]), .D(regs[747]), 
        .S0(n719), .S1(n713), .Q(n501) );
  IMUX40 U537 ( .A(regs[139]), .B(regs[171]), .C(regs[203]), .D(regs[235]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n506) );
  IMUX40 U538 ( .A(regs[652]), .B(regs[684]), .C(regs[716]), .D(regs[748]), 
        .S0(n719), .S1(i_addr_Rs[1]), .Q(n511) );
  IMUX40 U539 ( .A(regs[140]), .B(regs[172]), .C(regs[204]), .D(regs[236]), 
        .S0(n720), .S1(i_addr_Rs[1]), .Q(n516) );
  IMUX40 U540 ( .A(regs[653]), .B(regs[685]), .C(regs[717]), .D(regs[749]), 
        .S0(n720), .S1(n713), .Q(n521) );
  IMUX40 U541 ( .A(regs[141]), .B(regs[173]), .C(regs[205]), .D(regs[237]), 
        .S0(n720), .S1(n715), .Q(n526) );
  IMUX40 U542 ( .A(regs[654]), .B(regs[686]), .C(regs[718]), .D(regs[750]), 
        .S0(n721), .S1(n712), .Q(n531) );
  IMUX40 U543 ( .A(regs[142]), .B(regs[174]), .C(regs[206]), .D(regs[238]), 
        .S0(n721), .S1(n712), .Q(n536) );
  IMUX40 U544 ( .A(regs[655]), .B(regs[687]), .C(regs[719]), .D(regs[751]), 
        .S0(n721), .S1(n715), .Q(n541) );
  IMUX40 U545 ( .A(regs[143]), .B(regs[175]), .C(regs[207]), .D(regs[239]), 
        .S0(n722), .S1(i_addr_Rs[1]), .Q(n546) );
  IMUX40 U546 ( .A(regs[656]), .B(regs[688]), .C(regs[720]), .D(regs[752]), 
        .S0(n722), .S1(n713), .Q(n551) );
  IMUX40 U547 ( .A(regs[144]), .B(regs[176]), .C(regs[208]), .D(regs[240]), 
        .S0(n722), .S1(n718), .Q(n556) );
  IMUX40 U548 ( .A(regs[657]), .B(regs[689]), .C(regs[721]), .D(regs[753]), 
        .S0(n723), .S1(n712), .Q(n561) );
  IMUX40 U549 ( .A(regs[145]), .B(regs[177]), .C(regs[209]), .D(regs[241]), 
        .S0(n723), .S1(n713), .Q(n566) );
  IMUX40 U550 ( .A(regs[658]), .B(regs[690]), .C(regs[722]), .D(regs[754]), 
        .S0(n723), .S1(n716), .Q(n571) );
  IMUX40 U551 ( .A(regs[146]), .B(regs[178]), .C(regs[210]), .D(regs[242]), 
        .S0(n721), .S1(n715), .Q(n576) );
  IMUX40 U552 ( .A(regs[659]), .B(regs[691]), .C(regs[723]), .D(regs[755]), 
        .S0(n722), .S1(n715), .Q(n581) );
  IMUX40 U553 ( .A(regs[147]), .B(regs[179]), .C(regs[211]), .D(regs[243]), 
        .S0(n723), .S1(n713), .Q(n586) );
  IMUX40 U554 ( .A(regs[660]), .B(regs[692]), .C(regs[724]), .D(regs[756]), 
        .S0(n727), .S1(n715), .Q(n591) );
  IMUX40 U555 ( .A(regs[148]), .B(regs[180]), .C(regs[212]), .D(regs[244]), 
        .S0(n729), .S1(i_addr_Rs[1]), .Q(n596) );
  IMUX40 U556 ( .A(regs[661]), .B(regs[693]), .C(regs[725]), .D(regs[757]), 
        .S0(n728), .S1(n713), .Q(n601) );
  IMUX40 U557 ( .A(regs[149]), .B(regs[181]), .C(regs[213]), .D(regs[245]), 
        .S0(n727), .S1(n714), .Q(n606) );
  IMUX40 U558 ( .A(regs[662]), .B(regs[694]), .C(regs[726]), .D(regs[758]), 
        .S0(n729), .S1(n715), .Q(n611) );
  IMUX40 U559 ( .A(regs[150]), .B(regs[182]), .C(regs[214]), .D(regs[246]), 
        .S0(n730), .S1(n715), .Q(n616) );
  IMUX40 U560 ( .A(regs[663]), .B(regs[695]), .C(regs[727]), .D(regs[759]), 
        .S0(n724), .S1(n712), .Q(n621) );
  IMUX40 U561 ( .A(regs[151]), .B(regs[183]), .C(regs[215]), .D(regs[247]), 
        .S0(n724), .S1(n716), .Q(n626) );
  IMUX40 U562 ( .A(regs[664]), .B(regs[696]), .C(regs[728]), .D(regs[760]), 
        .S0(n724), .S1(n715), .Q(n631) );
  IMUX40 U563 ( .A(regs[152]), .B(regs[184]), .C(regs[216]), .D(regs[248]), 
        .S0(n730), .S1(n716), .Q(n636) );
  IMUX40 U564 ( .A(regs[665]), .B(regs[697]), .C(regs[729]), .D(regs[761]), 
        .S0(n724), .S1(n712), .Q(n641) );
  IMUX40 U565 ( .A(regs[153]), .B(regs[185]), .C(regs[217]), .D(regs[249]), 
        .S0(i_addr_Rs[0]), .S1(n712), .Q(n646) );
  IMUX40 U566 ( .A(regs[666]), .B(regs[698]), .C(regs[730]), .D(regs[762]), 
        .S0(n726), .S1(n716), .Q(n651) );
  IMUX40 U567 ( .A(regs[154]), .B(regs[186]), .C(regs[218]), .D(regs[250]), 
        .S0(n728), .S1(n716), .Q(n656) );
  IMUX40 U568 ( .A(regs[667]), .B(regs[699]), .C(regs[731]), .D(regs[763]), 
        .S0(n728), .S1(n716), .Q(n661) );
  IMUX40 U569 ( .A(regs[155]), .B(regs[187]), .C(regs[219]), .D(regs[251]), 
        .S0(n725), .S1(n718), .Q(n666) );
  IMUX40 U570 ( .A(regs[668]), .B(regs[700]), .C(regs[732]), .D(regs[764]), 
        .S0(n725), .S1(n717), .Q(n671) );
  IMUX40 U571 ( .A(regs[156]), .B(regs[188]), .C(regs[220]), .D(regs[252]), 
        .S0(n725), .S1(n717), .Q(n676) );
  IMUX40 U572 ( .A(regs[669]), .B(regs[701]), .C(regs[733]), .D(regs[765]), 
        .S0(n726), .S1(n718), .Q(n681) );
  IMUX40 U573 ( .A(regs[670]), .B(regs[702]), .C(regs[734]), .D(regs[766]), 
        .S0(n726), .S1(n717), .Q(n691) );
  IMUX40 U574 ( .A(regs[671]), .B(regs[703]), .C(regs[735]), .D(regs[767]), 
        .S0(n730), .S1(n718), .Q(n701) );
  BUF2 U575 ( .A(i_addr_Rt[3]), .Q(n366) );
  BUF2 U576 ( .A(i_addr_Rt[3]), .Q(n367) );
  BUF2 U577 ( .A(i_addr_Rs[3]), .Q(n709) );
  BUF2 U578 ( .A(i_addr_Rs[3]), .Q(n710) );
  INV3 U579 ( .A(i_addr_Rd[0]), .Q(n776) );
  INV3 U580 ( .A(i_addr_Rd[1]), .Q(n775) );
  INV3 U581 ( .A(i_addr_Rd[2]), .Q(n774) );
  INV3 U582 ( .A(i_con_RegWr), .Q(n777) );
  BUF2 U583 ( .A(i_addr_Rs[4]), .Q(n708) );
  BUF2 U584 ( .A(i_addr_Rs[2]), .Q(n711) );
  INV3 U585 ( .A(i_addr_Rd[4]), .Q(n756) );
  INV3 U586 ( .A(i_addr_Rd[3]), .Q(n773) );
  MUX22 U587 ( .A(n403), .B(n398), .S(n708), .Q(o_data_Rs[1]) );
  IMUX40 U588 ( .A(n404), .B(n405), .C(n406), .D(n407), .S0(i_addr_Rs[3]), 
        .S1(n711), .Q(n403) );
  IMUX40 U589 ( .A(n399), .B(n400), .C(n401), .D(n402), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n398) );
  IMUX40 U590 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n727), .S1(n714), .Q(n404) );
  MUX22 U591 ( .A(n413), .B(n408), .S(n708), .Q(o_data_Rs[2]) );
  IMUX40 U592 ( .A(n414), .B(n415), .C(n416), .D(n417), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n413) );
  IMUX40 U593 ( .A(n409), .B(n410), .C(n411), .D(n412), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n408) );
  IMUX40 U594 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n730), .S1(n713), .Q(n414) );
  MUX22 U595 ( .A(n423), .B(n418), .S(n708), .Q(o_data_Rs[3]) );
  IMUX40 U596 ( .A(n424), .B(n425), .C(n426), .D(n427), .S0(n709), .S1(n711), 
        .Q(n423) );
  IMUX40 U597 ( .A(n419), .B(n420), .C(n421), .D(n422), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n418) );
  IMUX40 U598 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n424) );
  MUX22 U599 ( .A(n433), .B(n428), .S(n708), .Q(o_data_Rs[4]) );
  IMUX40 U600 ( .A(n434), .B(n435), .C(n436), .D(n437), .S0(n709), .S1(n711), 
        .Q(n433) );
  IMUX40 U601 ( .A(n429), .B(n430), .C(n431), .D(n432), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n428) );
  IMUX40 U602 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        i_addr_Rs[0]), .S1(n714), .Q(n434) );
  MUX22 U603 ( .A(n443), .B(n438), .S(n708), .Q(o_data_Rs[5]) );
  IMUX40 U604 ( .A(n444), .B(n445), .C(n446), .D(n447), .S0(n709), .S1(n711), 
        .Q(n443) );
  IMUX40 U605 ( .A(n439), .B(n440), .C(n441), .D(n442), .S0(n709), .S1(n711), 
        .Q(n438) );
  IMUX40 U606 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n444) );
  MUX22 U607 ( .A(n453), .B(n448), .S(i_addr_Rs[4]), .Q(o_data_Rs[6]) );
  IMUX40 U608 ( .A(n454), .B(n455), .C(n456), .D(n457), .S0(n709), .S1(n711), 
        .Q(n453) );
  IMUX40 U609 ( .A(n449), .B(n450), .C(n451), .D(n452), .S0(n709), .S1(n711), 
        .Q(n448) );
  IMUX40 U610 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        i_addr_Rs[0]), .S1(n717), .Q(n454) );
  MUX22 U611 ( .A(n463), .B(n458), .S(i_addr_Rs[4]), .Q(o_data_Rs[7]) );
  IMUX40 U612 ( .A(n464), .B(n465), .C(n466), .D(n467), .S0(n709), .S1(n711), 
        .Q(n463) );
  IMUX40 U613 ( .A(n459), .B(n460), .C(n461), .D(n462), .S0(n709), .S1(n711), 
        .Q(n458) );
  IMUX40 U614 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n727), .S1(n714), .Q(n464) );
  MUX22 U615 ( .A(n473), .B(n468), .S(i_addr_Rs[4]), .Q(o_data_Rs[8]) );
  IMUX40 U616 ( .A(n474), .B(n475), .C(n476), .D(n477), .S0(n710), .S1(n711), 
        .Q(n473) );
  IMUX40 U617 ( .A(n469), .B(n470), .C(n471), .D(n472), .S0(n710), .S1(n711), 
        .Q(n468) );
  IMUX40 U618 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n729), .S1(n718), .Q(n474) );
  MUX22 U619 ( .A(n483), .B(n478), .S(i_addr_Rs[4]), .Q(o_data_Rs[9]) );
  IMUX40 U620 ( .A(n484), .B(n485), .C(n486), .D(n487), .S0(n710), .S1(n711), 
        .Q(n483) );
  IMUX40 U621 ( .A(n479), .B(n480), .C(n481), .D(n482), .S0(n710), .S1(n711), 
        .Q(n478) );
  IMUX40 U622 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        i_addr_Rs[0]), .S1(i_addr_Rs[1]), .Q(n484) );
  MUX22 U623 ( .A(n493), .B(n488), .S(i_addr_Rs[4]), .Q(o_data_Rs[10]) );
  IMUX40 U624 ( .A(n494), .B(n495), .C(n496), .D(n497), .S0(n710), .S1(n711), 
        .Q(n493) );
  IMUX40 U625 ( .A(n489), .B(n490), .C(n491), .D(n492), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n488) );
  IMUX40 U626 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        i_addr_Rs[0]), .S1(n714), .Q(n494) );
  MUX22 U627 ( .A(n503), .B(n498), .S(i_addr_Rs[4]), .Q(o_data_Rs[11]) );
  IMUX40 U628 ( .A(n504), .B(n505), .C(n506), .D(n507), .S0(n710), .S1(n711), 
        .Q(n503) );
  IMUX40 U629 ( .A(n499), .B(n500), .C(n501), .D(n502), .S0(n710), .S1(n711), 
        .Q(n498) );
  IMUX40 U630 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n719), .S1(n712), .Q(n504) );
  MUX22 U631 ( .A(n513), .B(n508), .S(i_addr_Rs[4]), .Q(o_data_Rs[12]) );
  IMUX40 U632 ( .A(n514), .B(n515), .C(n516), .D(n517), .S0(n710), .S1(n711), 
        .Q(n513) );
  IMUX40 U633 ( .A(n509), .B(n510), .C(n511), .D(n512), .S0(n710), .S1(n711), 
        .Q(n508) );
  IMUX40 U634 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n720), .S1(i_addr_Rs[1]), .Q(n514) );
  MUX22 U635 ( .A(n523), .B(n518), .S(i_addr_Rs[4]), .Q(o_data_Rs[13]) );
  IMUX40 U636 ( .A(n524), .B(n525), .C(n526), .D(n527), .S0(n710), .S1(n711), 
        .Q(n523) );
  IMUX40 U637 ( .A(n519), .B(n520), .C(n521), .D(n522), .S0(n710), .S1(n711), 
        .Q(n518) );
  IMUX40 U638 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n720), .S1(n716), .Q(n524) );
  MUX22 U639 ( .A(n533), .B(n528), .S(i_addr_Rs[4]), .Q(o_data_Rs[14]) );
  IMUX40 U640 ( .A(n534), .B(n535), .C(n536), .D(n537), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n533) );
  IMUX40 U641 ( .A(n529), .B(n530), .C(n531), .D(n532), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n528) );
  IMUX40 U642 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n721), .S1(n718), .Q(n534) );
  MUX22 U643 ( .A(n543), .B(n538), .S(i_addr_Rs[4]), .Q(o_data_Rs[15]) );
  IMUX40 U644 ( .A(n544), .B(n545), .C(n546), .D(n547), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n543) );
  IMUX40 U645 ( .A(n539), .B(n540), .C(n541), .D(n542), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n538) );
  IMUX40 U646 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n722), .S1(i_addr_Rs[1]), .Q(n544) );
  MUX22 U647 ( .A(n553), .B(n548), .S(i_addr_Rs[4]), .Q(o_data_Rs[16]) );
  IMUX40 U648 ( .A(n554), .B(n555), .C(n556), .D(n557), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n553) );
  IMUX40 U649 ( .A(n549), .B(n550), .C(n551), .D(n552), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n548) );
  IMUX40 U650 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n722), .S1(i_addr_Rs[1]), .Q(n554) );
  MUX22 U651 ( .A(n563), .B(n558), .S(i_addr_Rs[4]), .Q(o_data_Rs[17]) );
  IMUX40 U652 ( .A(n564), .B(n565), .C(n566), .D(n567), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n563) );
  IMUX40 U653 ( .A(n559), .B(n560), .C(n561), .D(n562), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n558) );
  IMUX40 U654 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n723), .S1(n713), .Q(n564) );
  MUX22 U655 ( .A(n573), .B(n568), .S(i_addr_Rs[4]), .Q(o_data_Rs[18]) );
  IMUX40 U656 ( .A(n574), .B(n575), .C(n576), .D(n577), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n573) );
  IMUX40 U657 ( .A(n569), .B(n570), .C(n571), .D(n572), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n568) );
  IMUX40 U658 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n729), .S1(n714), .Q(n574) );
  MUX22 U659 ( .A(n583), .B(n578), .S(n708), .Q(o_data_Rs[19]) );
  IMUX40 U660 ( .A(n584), .B(n585), .C(n586), .D(n587), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n583) );
  IMUX40 U661 ( .A(n579), .B(n580), .C(n581), .D(n582), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n578) );
  IMUX40 U662 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n728), .S1(n712), .Q(n584) );
  MUX22 U663 ( .A(n593), .B(n588), .S(n708), .Q(o_data_Rs[20]) );
  IMUX40 U664 ( .A(n594), .B(n595), .C(n596), .D(n597), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n593) );
  IMUX40 U665 ( .A(n589), .B(n590), .C(n591), .D(n592), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n588) );
  IMUX40 U666 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n721), .S1(i_addr_Rs[1]), .Q(n594) );
  MUX22 U667 ( .A(n603), .B(n598), .S(n708), .Q(o_data_Rs[21]) );
  IMUX40 U668 ( .A(n604), .B(n605), .C(n606), .D(n607), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n603) );
  IMUX40 U669 ( .A(n599), .B(n600), .C(n601), .D(n602), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n598) );
  IMUX40 U670 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n730), .S1(n715), .Q(n604) );
  MUX22 U671 ( .A(n613), .B(n608), .S(n708), .Q(o_data_Rs[22]) );
  IMUX40 U672 ( .A(n614), .B(n615), .C(n616), .D(n617), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n613) );
  IMUX40 U673 ( .A(n609), .B(n610), .C(n611), .D(n612), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n608) );
  IMUX40 U674 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n729), .S1(n715), .Q(n614) );
  MUX22 U675 ( .A(n623), .B(n618), .S(n708), .Q(o_data_Rs[23]) );
  IMUX40 U676 ( .A(n624), .B(n625), .C(n626), .D(n627), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n623) );
  IMUX40 U677 ( .A(n619), .B(n620), .C(n621), .D(n622), .S0(n709), .S1(
        i_addr_Rs[2]), .Q(n618) );
  IMUX40 U678 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n724), .S1(n718), .Q(n624) );
  MUX22 U679 ( .A(n633), .B(n628), .S(n708), .Q(o_data_Rs[24]) );
  IMUX40 U680 ( .A(n634), .B(n635), .C(n636), .D(n637), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n633) );
  IMUX40 U681 ( .A(n629), .B(n630), .C(n631), .D(n632), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n628) );
  IMUX40 U682 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n730), .S1(n717), .Q(n634) );
  MUX22 U683 ( .A(n643), .B(n638), .S(n708), .Q(o_data_Rs[25]) );
  IMUX40 U684 ( .A(n644), .B(n645), .C(n646), .D(n647), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n643) );
  IMUX40 U685 ( .A(n639), .B(n640), .C(n641), .D(n642), .S0(n710), .S1(
        i_addr_Rs[2]), .Q(n638) );
  IMUX40 U686 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n727), .S1(n717), .Q(n644) );
  MUX22 U687 ( .A(n653), .B(n648), .S(i_addr_Rs[4]), .Q(o_data_Rs[26]) );
  IMUX40 U688 ( .A(n654), .B(n655), .C(n656), .D(n657), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n653) );
  IMUX40 U689 ( .A(n649), .B(n650), .C(n651), .D(n652), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n648) );
  IMUX40 U690 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n720), .S1(n716), .Q(n654) );
  MUX22 U691 ( .A(n663), .B(n658), .S(i_addr_Rs[4]), .Q(o_data_Rs[27]) );
  IMUX40 U692 ( .A(n664), .B(n665), .C(n666), .D(n667), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n663) );
  IMUX40 U693 ( .A(n659), .B(n660), .C(n661), .D(n662), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n658) );
  IMUX40 U694 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n725), .S1(n713), .Q(n664) );
  MUX22 U695 ( .A(n673), .B(n668), .S(i_addr_Rs[4]), .Q(o_data_Rs[28]) );
  IMUX40 U696 ( .A(n674), .B(n675), .C(n676), .D(n677), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n673) );
  IMUX40 U697 ( .A(n669), .B(n670), .C(n671), .D(n672), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n668) );
  IMUX40 U698 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n725), .S1(n718), .Q(n674) );
  MUX22 U699 ( .A(n683), .B(n678), .S(i_addr_Rs[4]), .Q(o_data_Rs[29]) );
  IMUX40 U700 ( .A(n684), .B(n685), .C(n686), .D(n687), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n683) );
  IMUX40 U701 ( .A(n679), .B(n680), .C(n681), .D(n682), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n678) );
  IMUX40 U702 ( .A(regs[157]), .B(regs[189]), .C(regs[221]), .D(regs[253]), 
        .S0(n726), .S1(n717), .Q(n686) );
  MUX22 U703 ( .A(n693), .B(n688), .S(i_addr_Rs[4]), .Q(o_data_Rs[30]) );
  IMUX40 U704 ( .A(n694), .B(n695), .C(n696), .D(n697), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n693) );
  IMUX40 U705 ( .A(n689), .B(n690), .C(n691), .D(n692), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n688) );
  IMUX40 U706 ( .A(regs[158]), .B(regs[190]), .C(regs[222]), .D(regs[254]), 
        .S0(n729), .S1(n717), .Q(n696) );
  MUX22 U707 ( .A(n703), .B(n698), .S(i_addr_Rs[4]), .Q(o_data_Rs[31]) );
  IMUX40 U708 ( .A(n704), .B(n705), .C(n706), .D(n707), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n703) );
  IMUX40 U709 ( .A(n699), .B(n700), .C(n701), .D(n702), .S0(i_addr_Rs[3]), 
        .S1(i_addr_Rs[2]), .Q(n698) );
  IMUX40 U710 ( .A(regs[159]), .B(regs[191]), .C(regs[223]), .D(regs[255]), 
        .S0(n725), .S1(n718), .Q(n706) );
  BUF2 U711 ( .A(n375), .Q(n369) );
  BUF2 U712 ( .A(i_addr_Rt[1]), .Q(n375) );
  BUF2 U713 ( .A(i_addr_Rs[1]), .Q(n712) );
  MUX22 U714 ( .A(n6), .B(n1), .S(i_addr_Rt[4]), .Q(o_data_Rt[0]) );
  IMUX40 U715 ( .A(n2), .B(n3), .C(n4), .D(n5), .S0(n365), .S1(i_addr_Rt[2]), 
        .Q(n1) );
  IMUX40 U716 ( .A(n7), .B(n8), .C(n9), .D(n10), .S0(n365), .S1(i_addr_Rt[2]), 
        .Q(n6) );
  MUX22 U717 ( .A(n16), .B(n11), .S(i_addr_Rt[4]), .Q(o_data_Rt[1]) );
  IMUX40 U718 ( .A(n17), .B(n18), .C(n19), .D(n20), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n16) );
  IMUX40 U719 ( .A(n12), .B(n13), .C(n14), .D(n15), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n11) );
  IMUX40 U720 ( .A(regs[1]), .B(regs[33]), .C(regs[65]), .D(regs[97]), .S0(
        n379), .S1(n370), .Q(n17) );
  MUX22 U721 ( .A(n26), .B(n21), .S(i_addr_Rt[4]), .Q(o_data_Rt[2]) );
  IMUX40 U722 ( .A(n27), .B(n28), .C(n29), .D(n30), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n26) );
  IMUX40 U723 ( .A(n22), .B(n23), .C(n24), .D(n25), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n21) );
  IMUX40 U724 ( .A(regs[2]), .B(regs[34]), .C(regs[66]), .D(regs[98]), .S0(
        n378), .S1(i_addr_Rt[1]), .Q(n27) );
  MUX22 U725 ( .A(n36), .B(n31), .S(i_addr_Rt[4]), .Q(o_data_Rt[3]) );
  IMUX40 U726 ( .A(n37), .B(n38), .C(n83), .D(n84), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n36) );
  IMUX40 U727 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n31) );
  IMUX40 U728 ( .A(regs[3]), .B(regs[35]), .C(regs[67]), .D(regs[99]), .S0(
        n381), .S1(n369), .Q(n37) );
  MUX22 U729 ( .A(n90), .B(n85), .S(i_addr_Rt[4]), .Q(o_data_Rt[4]) );
  IMUX40 U730 ( .A(n91), .B(n92), .C(n93), .D(n94), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n90) );
  IMUX40 U731 ( .A(n86), .B(n87), .C(n88), .D(n89), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n85) );
  IMUX40 U732 ( .A(regs[4]), .B(regs[36]), .C(regs[68]), .D(regs[100]), .S0(
        n376), .S1(i_addr_Rt[1]), .Q(n91) );
  MUX22 U733 ( .A(n100), .B(n95), .S(i_addr_Rt[4]), .Q(o_data_Rt[5]) );
  IMUX40 U734 ( .A(n101), .B(n102), .C(n103), .D(n104), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n100) );
  IMUX40 U735 ( .A(n96), .B(n97), .C(n98), .D(n99), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n95) );
  IMUX40 U736 ( .A(regs[5]), .B(regs[37]), .C(regs[69]), .D(regs[101]), .S0(
        n387), .S1(n375), .Q(n101) );
  MUX22 U737 ( .A(n110), .B(n105), .S(i_addr_Rt[4]), .Q(o_data_Rt[6]) );
  IMUX40 U738 ( .A(n111), .B(n112), .C(n113), .D(n114), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n110) );
  IMUX40 U739 ( .A(n106), .B(n107), .C(n108), .D(n109), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n105) );
  IMUX40 U740 ( .A(regs[6]), .B(regs[38]), .C(regs[70]), .D(regs[102]), .S0(
        n385), .S1(i_addr_Rt[1]), .Q(n111) );
  MUX22 U741 ( .A(n120), .B(n115), .S(i_addr_Rt[4]), .Q(o_data_Rt[7]) );
  IMUX40 U742 ( .A(n121), .B(n122), .C(n123), .D(n124), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n120) );
  IMUX40 U743 ( .A(n116), .B(n117), .C(n118), .D(n119), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n115) );
  IMUX40 U744 ( .A(regs[7]), .B(regs[39]), .C(regs[71]), .D(regs[103]), .S0(
        n385), .S1(n373), .Q(n121) );
  MUX22 U745 ( .A(n130), .B(n125), .S(i_addr_Rt[4]), .Q(o_data_Rt[8]) );
  IMUX40 U746 ( .A(n131), .B(n132), .C(n133), .D(n134), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n130) );
  IMUX40 U747 ( .A(n126), .B(n127), .C(n128), .D(n129), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n125) );
  IMUX40 U748 ( .A(regs[8]), .B(regs[40]), .C(regs[72]), .D(regs[104]), .S0(
        n382), .S1(n375), .Q(n131) );
  MUX22 U749 ( .A(n140), .B(n135), .S(i_addr_Rt[4]), .Q(o_data_Rt[9]) );
  IMUX40 U750 ( .A(n141), .B(n142), .C(n143), .D(n144), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n140) );
  IMUX40 U751 ( .A(n136), .B(n137), .C(n138), .D(n139), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n135) );
  IMUX40 U752 ( .A(regs[9]), .B(regs[41]), .C(regs[73]), .D(regs[105]), .S0(
        n387), .S1(i_addr_Rt[1]), .Q(n141) );
  MUX22 U753 ( .A(n150), .B(n145), .S(i_addr_Rt[4]), .Q(o_data_Rt[10]) );
  IMUX40 U754 ( .A(n151), .B(n152), .C(n153), .D(n154), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n150) );
  IMUX40 U755 ( .A(n146), .B(n147), .C(n148), .D(n149), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n145) );
  IMUX40 U756 ( .A(regs[10]), .B(regs[42]), .C(regs[74]), .D(regs[106]), .S0(
        n381), .S1(i_addr_Rt[1]), .Q(n151) );
  MUX22 U757 ( .A(n160), .B(n155), .S(i_addr_Rt[4]), .Q(o_data_Rt[11]) );
  IMUX40 U758 ( .A(n161), .B(n162), .C(n163), .D(n164), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n160) );
  IMUX40 U759 ( .A(n156), .B(n157), .C(n158), .D(n159), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n155) );
  IMUX40 U760 ( .A(regs[11]), .B(regs[43]), .C(regs[75]), .D(regs[107]), .S0(
        n376), .S1(n371), .Q(n161) );
  MUX22 U761 ( .A(n170), .B(n165), .S(i_addr_Rt[4]), .Q(o_data_Rt[12]) );
  IMUX40 U762 ( .A(n171), .B(n172), .C(n173), .D(n174), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n170) );
  IMUX40 U763 ( .A(n166), .B(n167), .C(n168), .D(n169), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n165) );
  IMUX40 U764 ( .A(regs[12]), .B(regs[44]), .C(regs[76]), .D(regs[108]), .S0(
        n377), .S1(i_addr_Rt[1]), .Q(n171) );
  MUX22 U765 ( .A(n180), .B(n175), .S(i_addr_Rt[4]), .Q(o_data_Rt[13]) );
  IMUX40 U766 ( .A(n181), .B(n182), .C(n183), .D(n184), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n180) );
  IMUX40 U767 ( .A(n176), .B(n177), .C(n178), .D(n179), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n175) );
  IMUX40 U768 ( .A(regs[13]), .B(regs[45]), .C(regs[77]), .D(regs[109]), .S0(
        n377), .S1(n375), .Q(n181) );
  MUX22 U769 ( .A(n190), .B(n185), .S(i_addr_Rt[4]), .Q(o_data_Rt[14]) );
  IMUX40 U770 ( .A(n191), .B(n192), .C(n193), .D(n194), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n190) );
  IMUX40 U771 ( .A(n186), .B(n187), .C(n188), .D(n189), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n185) );
  IMUX40 U772 ( .A(regs[14]), .B(regs[46]), .C(regs[78]), .D(regs[110]), .S0(
        n378), .S1(n371), .Q(n191) );
  MUX22 U773 ( .A(n200), .B(n195), .S(i_addr_Rt[4]), .Q(o_data_Rt[15]) );
  IMUX40 U774 ( .A(n201), .B(n202), .C(n203), .D(n204), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n200) );
  IMUX40 U775 ( .A(n196), .B(n197), .C(n198), .D(n199), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n195) );
  IMUX40 U776 ( .A(regs[15]), .B(regs[47]), .C(regs[79]), .D(regs[111]), .S0(
        n380), .S1(i_addr_Rt[1]), .Q(n201) );
  MUX22 U777 ( .A(n210), .B(n205), .S(i_addr_Rt[4]), .Q(o_data_Rt[16]) );
  IMUX40 U778 ( .A(n211), .B(n212), .C(n213), .D(n214), .S0(n366), .S1(
        i_addr_Rt[2]), .Q(n210) );
  IMUX40 U779 ( .A(n206), .B(n207), .C(n208), .D(n209), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n205) );
  IMUX40 U780 ( .A(regs[16]), .B(regs[48]), .C(regs[80]), .D(regs[112]), .S0(
        n382), .S1(n372), .Q(n211) );
  MUX22 U781 ( .A(n220), .B(n215), .S(i_addr_Rt[4]), .Q(o_data_Rt[17]) );
  IMUX40 U782 ( .A(n221), .B(n222), .C(n223), .D(n224), .S0(n367), .S1(
        i_addr_Rt[2]), .Q(n220) );
  IMUX40 U783 ( .A(n216), .B(n217), .C(n218), .D(n219), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n215) );
  IMUX40 U784 ( .A(regs[17]), .B(regs[49]), .C(regs[81]), .D(regs[113]), .S0(
        n384), .S1(n370), .Q(n221) );
  MUX22 U785 ( .A(n230), .B(n225), .S(i_addr_Rt[4]), .Q(o_data_Rt[18]) );
  IMUX40 U786 ( .A(n231), .B(n232), .C(n233), .D(n234), .S0(n365), .S1(n368), 
        .Q(n230) );
  IMUX40 U787 ( .A(n226), .B(n227), .C(n228), .D(n229), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n225) );
  IMUX40 U788 ( .A(regs[18]), .B(regs[50]), .C(regs[82]), .D(regs[114]), .S0(
        n379), .S1(n370), .Q(n231) );
  MUX22 U789 ( .A(n240), .B(n235), .S(i_addr_Rt[4]), .Q(o_data_Rt[19]) );
  IMUX40 U790 ( .A(n241), .B(n242), .C(n243), .D(n244), .S0(n366), .S1(n368), 
        .Q(n240) );
  IMUX40 U791 ( .A(n236), .B(n237), .C(n238), .D(n239), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n235) );
  IMUX40 U792 ( .A(regs[19]), .B(regs[51]), .C(regs[83]), .D(regs[115]), .S0(
        n379), .S1(i_addr_Rt[1]), .Q(n241) );
  MUX22 U793 ( .A(n250), .B(n245), .S(i_addr_Rt[4]), .Q(o_data_Rt[20]) );
  IMUX40 U794 ( .A(n251), .B(n252), .C(n253), .D(n254), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n250) );
  IMUX40 U795 ( .A(n246), .B(n247), .C(n248), .D(n249), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n245) );
  IMUX40 U796 ( .A(regs[20]), .B(regs[52]), .C(regs[84]), .D(regs[116]), .S0(
        n380), .S1(i_addr_Rt[1]), .Q(n251) );
  MUX22 U797 ( .A(n260), .B(n255), .S(i_addr_Rt[4]), .Q(o_data_Rt[21]) );
  IMUX40 U798 ( .A(n261), .B(n262), .C(n263), .D(n264), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n260) );
  IMUX40 U799 ( .A(n256), .B(n257), .C(n258), .D(n259), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n255) );
  IMUX40 U800 ( .A(regs[21]), .B(regs[53]), .C(regs[85]), .D(regs[117]), .S0(
        n377), .S1(n371), .Q(n261) );
  MUX22 U801 ( .A(n270), .B(n265), .S(i_addr_Rt[4]), .Q(o_data_Rt[22]) );
  IMUX40 U802 ( .A(n271), .B(n272), .C(n273), .D(n274), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n270) );
  IMUX40 U803 ( .A(n266), .B(n267), .C(n268), .D(n269), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n265) );
  IMUX40 U804 ( .A(regs[22]), .B(regs[54]), .C(regs[86]), .D(regs[118]), .S0(
        n378), .S1(n371), .Q(n271) );
  MUX22 U805 ( .A(n280), .B(n275), .S(i_addr_Rt[4]), .Q(o_data_Rt[23]) );
  IMUX40 U806 ( .A(n281), .B(n282), .C(n283), .D(n284), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n280) );
  IMUX40 U807 ( .A(n276), .B(n277), .C(n278), .D(n279), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n275) );
  IMUX40 U808 ( .A(regs[23]), .B(regs[55]), .C(regs[87]), .D(regs[119]), .S0(
        n381), .S1(n373), .Q(n281) );
  MUX22 U809 ( .A(n290), .B(n285), .S(i_addr_Rt[4]), .Q(o_data_Rt[24]) );
  IMUX40 U810 ( .A(n291), .B(n292), .C(n293), .D(n294), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n290) );
  IMUX40 U811 ( .A(n286), .B(n287), .C(n288), .D(n289), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n285) );
  IMUX40 U812 ( .A(regs[24]), .B(regs[56]), .C(regs[88]), .D(regs[120]), .S0(
        n382), .S1(n374), .Q(n291) );
  MUX22 U813 ( .A(n300), .B(n295), .S(i_addr_Rt[4]), .Q(o_data_Rt[25]) );
  IMUX40 U814 ( .A(n301), .B(n302), .C(n303), .D(n304), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n300) );
  IMUX40 U815 ( .A(n296), .B(n297), .C(n298), .D(n299), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n295) );
  IMUX40 U816 ( .A(regs[25]), .B(regs[57]), .C(regs[89]), .D(regs[121]), .S0(
        n382), .S1(n369), .Q(n301) );
  MUX22 U817 ( .A(n310), .B(n305), .S(i_addr_Rt[4]), .Q(o_data_Rt[26]) );
  IMUX40 U818 ( .A(n311), .B(n312), .C(n313), .D(n314), .S0(n365), .S1(n368), 
        .Q(n310) );
  IMUX40 U819 ( .A(n306), .B(n307), .C(n308), .D(n309), .S0(n365), .S1(n368), 
        .Q(n305) );
  IMUX40 U820 ( .A(regs[26]), .B(regs[58]), .C(regs[90]), .D(regs[122]), .S0(
        n382), .S1(n372), .Q(n311) );
  MUX22 U821 ( .A(n320), .B(n315), .S(i_addr_Rt[4]), .Q(o_data_Rt[27]) );
  IMUX40 U822 ( .A(n321), .B(n322), .C(n323), .D(n324), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n320) );
  IMUX40 U823 ( .A(n316), .B(n317), .C(n318), .D(n319), .S0(n365), .S1(n368), 
        .Q(n315) );
  IMUX40 U824 ( .A(regs[27]), .B(regs[59]), .C(regs[91]), .D(regs[123]), .S0(
        n383), .S1(n374), .Q(n321) );
  MUX22 U825 ( .A(n330), .B(n325), .S(i_addr_Rt[4]), .Q(o_data_Rt[28]) );
  IMUX40 U826 ( .A(n331), .B(n332), .C(n333), .D(n334), .S0(i_addr_Rt[3]), 
        .S1(i_addr_Rt[2]), .Q(n330) );
  IMUX40 U827 ( .A(n326), .B(n327), .C(n328), .D(n329), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n325) );
  IMUX40 U828 ( .A(regs[28]), .B(regs[60]), .C(regs[92]), .D(regs[124]), .S0(
        n383), .S1(n372), .Q(n331) );
  MUX22 U829 ( .A(n340), .B(n335), .S(i_addr_Rt[4]), .Q(o_data_Rt[29]) );
  IMUX40 U830 ( .A(n341), .B(n342), .C(n343), .D(n344), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n340) );
  IMUX40 U831 ( .A(n336), .B(n337), .C(n338), .D(n339), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n335) );
  IMUX40 U832 ( .A(regs[29]), .B(regs[61]), .C(regs[93]), .D(regs[125]), .S0(
        n384), .S1(n373), .Q(n341) );
  MUX22 U833 ( .A(n350), .B(n345), .S(i_addr_Rt[4]), .Q(o_data_Rt[30]) );
  IMUX40 U834 ( .A(n351), .B(n352), .C(n353), .D(n354), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n350) );
  IMUX40 U835 ( .A(n346), .B(n347), .C(n348), .D(n349), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n345) );
  IMUX40 U836 ( .A(regs[30]), .B(regs[62]), .C(regs[94]), .D(regs[126]), .S0(
        i_addr_Rt[0]), .S1(n374), .Q(n351) );
  MUX22 U837 ( .A(n360), .B(n355), .S(i_addr_Rt[4]), .Q(o_data_Rt[31]) );
  IMUX40 U838 ( .A(n361), .B(n362), .C(n363), .D(n364), .S0(i_addr_Rt[3]), 
        .S1(n368), .Q(n360) );
  IMUX40 U839 ( .A(n356), .B(n357), .C(n358), .D(n359), .S0(n365), .S1(
        i_addr_Rt[2]), .Q(n355) );
  IMUX40 U840 ( .A(regs[31]), .B(regs[63]), .C(regs[95]), .D(regs[127]), .S0(
        n381), .S1(n374), .Q(n361) );
  BUF2 U841 ( .A(i_addr_Rt[2]), .Q(n368) );
  BUF2 U842 ( .A(i_addr_Rt[3]), .Q(n365) );
endmodule


module D_shiftleft ( i_data_immE, o_data_immshiftl );
  input [15:0] i_data_immE;
  output [31:0] o_data_immshiftl;
  wire   n1;
  assign o_data_immshiftl[0] = o_data_immshiftl[1];
  assign o_data_immshiftl[19] = o_data_immshiftl[30];
  assign o_data_immshiftl[29] = o_data_immshiftl[30];
  assign o_data_immshiftl[25] = o_data_immshiftl[30];
  assign o_data_immshiftl[21] = o_data_immshiftl[30];
  assign o_data_immshiftl[31] = o_data_immshiftl[30];
  assign o_data_immshiftl[20] = o_data_immshiftl[30];
  assign o_data_immshiftl[27] = o_data_immshiftl[30];
  assign o_data_immshiftl[26] = o_data_immshiftl[30];
  assign o_data_immshiftl[22] = o_data_immshiftl[30];
  assign o_data_immshiftl[24] = i_data_immE[15];
  assign o_data_immshiftl[28] = i_data_immE[15];
  assign o_data_immshiftl[17] = i_data_immE[15];
  assign o_data_immshiftl[18] = i_data_immE[15];
  assign o_data_immshiftl[23] = i_data_immE[15];
  assign o_data_immshiftl[16] = i_data_immE[14];
  assign o_data_immshiftl[15] = i_data_immE[13];
  assign o_data_immshiftl[14] = i_data_immE[12];
  assign o_data_immshiftl[13] = i_data_immE[11];
  assign o_data_immshiftl[12] = i_data_immE[10];
  assign o_data_immshiftl[11] = i_data_immE[9];
  assign o_data_immshiftl[10] = i_data_immE[8];
  assign o_data_immshiftl[9] = i_data_immE[7];
  assign o_data_immshiftl[8] = i_data_immE[6];
  assign o_data_immshiftl[7] = i_data_immE[5];
  assign o_data_immshiftl[6] = i_data_immE[4];
  assign o_data_immshiftl[5] = i_data_immE[3];
  assign o_data_immshiftl[4] = i_data_immE[2];
  assign o_data_immshiftl[3] = i_data_immE[1];
  assign o_data_immshiftl[2] = i_data_immE[0];

  INV3 U2 ( .A(n1), .Q(o_data_immshiftl[30]) );
  INV3 U3 ( .A(i_data_immE[15]), .Q(n1) );
  LOGIC0 U4 ( .Q(o_data_immshiftl[1]) );
endmodule


module D_sign_extend ( i_data_immD, i_con_signext, o_data_immD );
  input [15:0] i_data_immD;
  output [31:0] o_data_immD;
  input i_con_signext;
  wire   n2;
  assign o_data_immD[15] = i_data_immD[15];
  assign o_data_immD[14] = i_data_immD[14];
  assign o_data_immD[13] = i_data_immD[13];
  assign o_data_immD[12] = i_data_immD[12];
  assign o_data_immD[11] = i_data_immD[11];
  assign o_data_immD[10] = i_data_immD[10];
  assign o_data_immD[9] = i_data_immD[9];
  assign o_data_immD[8] = i_data_immD[8];
  assign o_data_immD[7] = i_data_immD[7];
  assign o_data_immD[6] = i_data_immD[6];
  assign o_data_immD[5] = i_data_immD[5];
  assign o_data_immD[4] = i_data_immD[4];
  assign o_data_immD[3] = i_data_immD[3];
  assign o_data_immD[2] = i_data_immD[2];
  assign o_data_immD[1] = i_data_immD[1];
  assign o_data_immD[0] = i_data_immD[0];
  assign o_data_immD[16] = o_data_immD[31];
  assign o_data_immD[17] = o_data_immD[31];
  assign o_data_immD[18] = o_data_immD[31];
  assign o_data_immD[19] = o_data_immD[31];
  assign o_data_immD[20] = o_data_immD[31];
  assign o_data_immD[21] = o_data_immD[31];
  assign o_data_immD[22] = o_data_immD[31];
  assign o_data_immD[23] = o_data_immD[31];
  assign o_data_immD[24] = o_data_immD[31];
  assign o_data_immD[25] = o_data_immD[31];
  assign o_data_immD[26] = o_data_immD[31];
  assign o_data_immD[27] = o_data_immD[31];
  assign o_data_immD[28] = o_data_immD[31];
  assign o_data_immD[29] = o_data_immD[31];
  assign o_data_immD[30] = o_data_immD[31];

  INV3 U2 ( .A(n2), .Q(o_data_immD[31]) );
  NAND22 U3 ( .A(i_con_signext), .B(i_data_immD[15]), .Q(n2) );
endmodule


module D_jump_ext ( i_addr_j, i_PC4_j, o_addr_j );
  input [25:0] i_addr_j;
  input [3:0] i_PC4_j;
  output [31:0] o_addr_j;

  assign o_addr_j[0] = o_addr_j[1];
  assign o_addr_j[31] = i_PC4_j[3];
  assign o_addr_j[30] = i_PC4_j[2];
  assign o_addr_j[29] = i_PC4_j[1];
  assign o_addr_j[28] = i_PC4_j[0];
  assign o_addr_j[27] = i_addr_j[25];
  assign o_addr_j[26] = i_addr_j[24];
  assign o_addr_j[25] = i_addr_j[23];
  assign o_addr_j[24] = i_addr_j[22];
  assign o_addr_j[23] = i_addr_j[21];
  assign o_addr_j[22] = i_addr_j[20];
  assign o_addr_j[21] = i_addr_j[19];
  assign o_addr_j[20] = i_addr_j[18];
  assign o_addr_j[19] = i_addr_j[17];
  assign o_addr_j[18] = i_addr_j[16];
  assign o_addr_j[17] = i_addr_j[15];
  assign o_addr_j[16] = i_addr_j[14];
  assign o_addr_j[15] = i_addr_j[13];
  assign o_addr_j[14] = i_addr_j[12];
  assign o_addr_j[13] = i_addr_j[11];
  assign o_addr_j[12] = i_addr_j[10];
  assign o_addr_j[11] = i_addr_j[9];
  assign o_addr_j[10] = i_addr_j[8];
  assign o_addr_j[9] = i_addr_j[7];
  assign o_addr_j[8] = i_addr_j[6];
  assign o_addr_j[7] = i_addr_j[5];
  assign o_addr_j[6] = i_addr_j[4];
  assign o_addr_j[5] = i_addr_j[3];
  assign o_addr_j[4] = i_addr_j[2];
  assign o_addr_j[3] = i_addr_j[1];
  assign o_addr_j[2] = i_addr_j[0];

  LOGIC0 U2 ( .Q(o_addr_j[1]) );
endmodule


module D_forward ( i_addr_rs, i_addr_rt, i_addr_rdE, i_addr_rdM, i_addr_rtM, 
        i_addr_rtW, i_con_regwriteE, i_con_regwriteM, i_con_memreadM, 
        i_con_memreadW, o_con_fa, o_con_fb );
  input [4:0] i_addr_rs;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rdE;
  input [4:0] i_addr_rdM;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  output [2:0] o_con_fa;
  output [2:0] o_con_fb;
  input i_con_regwriteE, i_con_regwriteM, i_con_memreadM, i_con_memreadW;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;

  OAI310 U1 ( .A(n1), .B(n2), .C(n3), .D(n4), .Q(o_con_fb[2]) );
  NOR40 U2 ( .A(n5), .B(n6), .C(n7), .D(n8), .Q(o_con_fb[1]) );
  CLKIN0 U3 ( .A(n9), .Q(n6) );
  NAND20 U4 ( .A(n4), .B(n10), .Q(o_con_fb[0]) );
  NAND40 U5 ( .A(n11), .B(i_con_regwriteM), .C(n12), .D(n13), .Q(n10) );
  NOR40 U6 ( .A(n14), .B(n15), .C(n16), .D(n17), .Q(n13) );
  XOR20 U7 ( .A(i_addr_rdM[4]), .B(i_addr_rt[4]), .Q(n17) );
  XNR20 U8 ( .A(n18), .B(i_addr_rt[2]), .Q(n16) );
  XNR20 U9 ( .A(n19), .B(i_addr_rt[1]), .Q(n15) );
  XNR20 U10 ( .A(n20), .B(i_addr_rt[0]), .Q(n14) );
  CLKIN0 U11 ( .A(n21), .Q(n12) );
  OAI210 U12 ( .A(n8), .B(n7), .C(n9), .Q(n21) );
  NAND40 U13 ( .A(n22), .B(n23), .C(n24), .D(n25), .Q(n7) );
  XNR20 U14 ( .A(i_addr_rt[0]), .B(i_addr_rdE[0]), .Q(n25) );
  NOR20 U15 ( .A(n26), .B(n27), .Q(n24) );
  XNR20 U16 ( .A(n28), .B(i_addr_rt[3]), .Q(n27) );
  XOR20 U17 ( .A(i_addr_rdE[1]), .B(i_addr_rt[1]), .Q(n26) );
  XNR20 U18 ( .A(i_addr_rt[2]), .B(i_addr_rdE[2]), .Q(n23) );
  XNR20 U19 ( .A(i_addr_rt[4]), .B(i_addr_rdE[4]), .Q(n22) );
  CLKIN0 U20 ( .A(i_con_regwriteE), .Q(n8) );
  XNR20 U21 ( .A(i_addr_rt[3]), .B(i_addr_rdM[3]), .Q(n11) );
  NAND20 U22 ( .A(n9), .B(n5), .Q(n4) );
  CLKIN0 U23 ( .A(n29), .Q(n5) );
  NAND40 U24 ( .A(n30), .B(i_con_memreadW), .C(n31), .D(n32), .Q(n29) );
  NOR30 U25 ( .A(n33), .B(n34), .C(n35), .Q(n32) );
  XOR20 U26 ( .A(i_addr_rtW[2]), .B(i_addr_rt[2]), .Q(n35) );
  XOR20 U27 ( .A(i_addr_rtW[4]), .B(i_addr_rt[4]), .Q(n34) );
  XOR20 U28 ( .A(i_addr_rtW[3]), .B(i_addr_rt[3]), .Q(n33) );
  XNR20 U29 ( .A(i_addr_rt[0]), .B(i_addr_rtW[0]), .Q(n31) );
  XNR20 U30 ( .A(i_addr_rt[1]), .B(i_addr_rtW[1]), .Q(n30) );
  AOI210 U31 ( .A(n36), .B(i_con_memreadM), .C(n2), .Q(n9) );
  NOR30 U32 ( .A(i_addr_rt[0]), .B(i_addr_rt[1]), .C(n37), .Q(n2) );
  CLKIN0 U33 ( .A(n38), .Q(n37) );
  NOR30 U34 ( .A(i_addr_rt[2]), .B(i_addr_rt[4]), .C(i_addr_rt[3]), .Q(n38) );
  CLKIN0 U35 ( .A(n3), .Q(n36) );
  NAND40 U36 ( .A(n39), .B(n40), .C(n41), .D(n42), .Q(n3) );
  XNR20 U37 ( .A(i_addr_rt[0]), .B(i_addr_rtM[0]), .Q(n42) );
  NOR20 U38 ( .A(n43), .B(n44), .Q(n41) );
  XOR20 U39 ( .A(i_addr_rtM[3]), .B(i_addr_rt[3]), .Q(n44) );
  XNR20 U40 ( .A(n45), .B(i_addr_rt[1]), .Q(n43) );
  XNR20 U41 ( .A(i_addr_rt[2]), .B(i_addr_rtM[2]), .Q(n40) );
  XNR20 U42 ( .A(i_addr_rt[4]), .B(i_addr_rtM[4]), .Q(n39) );
  NOR20 U43 ( .A(o_con_fa[2]), .B(n46), .Q(o_con_fa[1]) );
  OAI210 U44 ( .A(n47), .B(n48), .C(n49), .Q(o_con_fa[0]) );
  NAND20 U45 ( .A(n50), .B(n51), .Q(n49) );
  NOR40 U46 ( .A(o_con_fa[2]), .B(n52), .C(n53), .D(n54), .Q(n51) );
  XNR20 U47 ( .A(n20), .B(i_addr_rs[0]), .Q(n54) );
  CLKIN0 U48 ( .A(i_addr_rdM[0]), .Q(n20) );
  CLKIN0 U49 ( .A(i_con_regwriteM), .Q(n53) );
  CLKIN0 U50 ( .A(n46), .Q(n52) );
  NAND40 U51 ( .A(n55), .B(i_con_regwriteE), .C(n56), .D(n57), .Q(n46) );
  NOR30 U52 ( .A(n58), .B(n59), .C(n60), .Q(n57) );
  XNR20 U53 ( .A(n28), .B(i_addr_rs[3]), .Q(n60) );
  CLKIN0 U54 ( .A(i_addr_rdE[3]), .Q(n28) );
  XOR20 U55 ( .A(i_addr_rdE[2]), .B(i_addr_rs[2]), .Q(n59) );
  IMUX20 U56 ( .A(n61), .B(i_addr_rs[4]), .S(i_addr_rdE[4]), .Q(n58) );
  NOR20 U57 ( .A(n62), .B(i_addr_rs[4]), .Q(n61) );
  NOR40 U58 ( .A(i_addr_rdE[3]), .B(i_addr_rdE[2]), .C(i_addr_rdE[1]), .D(
        i_addr_rdE[0]), .Q(n62) );
  XNR20 U59 ( .A(i_addr_rs[0]), .B(i_addr_rdE[0]), .Q(n56) );
  XNR20 U60 ( .A(i_addr_rs[1]), .B(i_addr_rdE[1]), .Q(n55) );
  NAND20 U61 ( .A(n63), .B(n48), .Q(o_con_fa[2]) );
  NOR40 U62 ( .A(n64), .B(n65), .C(n66), .D(n67), .Q(n50) );
  IMUX20 U63 ( .A(n68), .B(i_addr_rs[4]), .S(i_addr_rdM[4]), .Q(n67) );
  NOR20 U64 ( .A(n69), .B(i_addr_rs[4]), .Q(n68) );
  NOR40 U65 ( .A(i_addr_rdM[3]), .B(i_addr_rdM[2]), .C(i_addr_rdM[1]), .D(
        i_addr_rdM[0]), .Q(n69) );
  XOR20 U66 ( .A(i_addr_rdM[3]), .B(i_addr_rs[3]), .Q(n66) );
  XNR20 U67 ( .A(n18), .B(i_addr_rs[2]), .Q(n65) );
  CLKIN0 U68 ( .A(i_addr_rdM[2]), .Q(n18) );
  XNR20 U69 ( .A(n19), .B(i_addr_rs[1]), .Q(n64) );
  CLKIN0 U70 ( .A(i_addr_rdM[1]), .Q(n19) );
  NAND40 U71 ( .A(n70), .B(n71), .C(n72), .D(n73), .Q(n48) );
  NOR40 U72 ( .A(n74), .B(n75), .C(n76), .D(n77), .Q(n73) );
  XOR20 U73 ( .A(i_addr_rtW[1]), .B(i_addr_rs[1]), .Q(n77) );
  XOR20 U74 ( .A(i_addr_rtW[0]), .B(i_addr_rs[0]), .Q(n76) );
  CLKIN0 U75 ( .A(i_con_memreadW), .Q(n75) );
  XNR20 U76 ( .A(i_addr_rtW[3]), .B(i_addr_rs[3]), .Q(n72) );
  XNR20 U77 ( .A(i_addr_rtW[4]), .B(i_addr_rs[4]), .Q(n71) );
  XNR20 U78 ( .A(i_addr_rtW[2]), .B(i_addr_rs[2]), .Q(n70) );
  CLKIN0 U79 ( .A(n63), .Q(n47) );
  NAND40 U80 ( .A(n78), .B(n79), .C(n80), .D(n81), .Q(n63) );
  NOR40 U81 ( .A(n74), .B(n1), .C(n82), .D(n83), .Q(n81) );
  XNR20 U82 ( .A(n45), .B(i_addr_rs[1]), .Q(n83) );
  CLKIN0 U83 ( .A(i_addr_rtM[1]), .Q(n45) );
  XOR20 U84 ( .A(i_addr_rtM[0]), .B(i_addr_rs[0]), .Q(n82) );
  CLKIN0 U85 ( .A(i_con_memreadM), .Q(n1) );
  NOR30 U86 ( .A(i_addr_rs[0]), .B(i_addr_rs[1]), .C(n84), .Q(n74) );
  CLKIN0 U87 ( .A(n85), .Q(n84) );
  NOR30 U88 ( .A(i_addr_rs[2]), .B(i_addr_rs[4]), .C(i_addr_rs[3]), .Q(n85) );
  XNR20 U89 ( .A(i_addr_rtM[3]), .B(i_addr_rs[3]), .Q(n80) );
  XNR20 U90 ( .A(i_addr_rtM[4]), .B(i_addr_rs[4]), .Q(n79) );
  XNR20 U91 ( .A(i_addr_rtM[2]), .B(i_addr_rs[2]), .Q(n78) );
endmodule


module decode ( i_clk, i_nrst, i_addr_pc4, i_data_instr, i_con_Wregwrite, 
        i_data_Wregwrite, i_addr_Wregwrite, i_addr_Erd, i_addr_Mrd, 
        i_con_Eregwrite, i_con_Mregwrite, i_addr_rtM, i_addr_rtW, 
        i_con_memreadM, i_con_memreadW, i_data_Wmemout, o_data_rs, o_data_rt, 
        o_addr_rd, o_addr_rt, o_data_jr, o_con_jump, o_addr_pc4, o_addr_branch, 
        o_addr_jump, o_con_Ealuop, o_con_Ealusrc, o_con_Eregdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_con_ifstall, o_con_Ebop, o_data_signext, 
        o_con_Efamux, o_con_Efbmux, o_data_Fmemout );
  input [31:0] i_addr_pc4;
  input [31:0] i_data_instr;
  input [31:0] i_data_Wregwrite;
  input [4:0] i_addr_Wregwrite;
  input [4:0] i_addr_Erd;
  input [4:0] i_addr_Mrd;
  input [4:0] i_addr_rtM;
  input [4:0] i_addr_rtW;
  input [31:0] i_data_Wmemout;
  output [31:0] o_data_rs;
  output [31:0] o_data_rt;
  output [4:0] o_addr_rd;
  output [4:0] o_addr_rt;
  output [31:0] o_data_jr;
  output [1:0] o_con_jump;
  output [31:0] o_addr_pc4;
  output [31:0] o_addr_branch;
  output [31:0] o_addr_jump;
  output [5:0] o_con_Ealuop;
  output [2:0] o_con_Ebop;
  output [31:0] o_data_signext;
  output [2:0] o_con_Efamux;
  output [2:0] o_con_Efbmux;
  output [31:0] o_data_Fmemout;
  input i_clk, i_nrst, i_con_Wregwrite, i_con_Eregwrite, i_con_Mregwrite,
         i_con_memreadM, i_con_memreadW;
  output o_con_Ealusrc, o_con_Eregdst, o_con_Mmemread, o_con_Mmemwrite,
         o_con_Malupc8, o_con_Wmemtoreg, o_con_Wregwrite, o_con_ifstall;
  wire   control_o_con_alusrc, control_o_con_regdst, jbcon_o_con_aluPC4,
         control_o_con_memread, control_o_con_memwrite, control_o_con_memtoreg,
         control_o_con_regwrite, signext_i_con_signext, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4;
  wire   [31:0] regbank_o_data_Rt;
  wire   [5:0] control_o_con_aluop;
  wire   [31:0] signext_o_data_immD;
  wire   [2:0] for_o_con_fa;
  wire   [2:0] for_o_con_fb;
  wire   [31:0] pcadd_o_addr_pcbranchE;
  wire   [2:0] jbcon_o_con_bop;
  wire   [31:2] pcadd_i_data_immshiftl;
  assign o_addr_jump[1] = o_addr_jump[0];

  DFC3 pipe_bop_reg_2_ ( .D(jbcon_o_con_bop[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[2]) );
  DFC3 pipe_bop_reg_1_ ( .D(jbcon_o_con_bop[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[1]) );
  DFC3 pipe_bop_reg_0_ ( .D(jbcon_o_con_bop[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Ebop[0]) );
  DFC3 pipe_data_rs_reg_31_ ( .D(o_data_jr[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[31]) );
  DFC3 pipe_data_rs_reg_30_ ( .D(o_data_jr[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[30]) );
  DFC3 pipe_data_rs_reg_29_ ( .D(o_data_jr[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[29]) );
  DFC3 pipe_data_rs_reg_28_ ( .D(o_data_jr[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[28]) );
  DFC3 pipe_data_rs_reg_27_ ( .D(o_data_jr[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[27]) );
  DFC3 pipe_data_rs_reg_26_ ( .D(o_data_jr[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[26]) );
  DFC3 pipe_data_rs_reg_25_ ( .D(o_data_jr[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[25]) );
  DFC3 pipe_data_rs_reg_24_ ( .D(o_data_jr[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[24]) );
  DFC3 pipe_data_rs_reg_23_ ( .D(o_data_jr[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[23]) );
  DFC3 pipe_data_rs_reg_22_ ( .D(o_data_jr[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[22]) );
  DFC3 pipe_data_rs_reg_21_ ( .D(o_data_jr[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[21]) );
  DFC3 pipe_data_rs_reg_20_ ( .D(o_data_jr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[20]) );
  DFC3 pipe_data_rs_reg_19_ ( .D(o_data_jr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[19]) );
  DFC3 pipe_data_rs_reg_18_ ( .D(o_data_jr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[18]) );
  DFC3 pipe_data_rs_reg_17_ ( .D(o_data_jr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[17]) );
  DFC3 pipe_data_rs_reg_16_ ( .D(o_data_jr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[16]) );
  DFC3 pipe_data_rs_reg_15_ ( .D(o_data_jr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[15]) );
  DFC3 pipe_data_rs_reg_14_ ( .D(o_data_jr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[14]) );
  DFC3 pipe_data_rs_reg_13_ ( .D(o_data_jr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[13]) );
  DFC3 pipe_data_rs_reg_12_ ( .D(o_data_jr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[12]) );
  DFC3 pipe_data_rs_reg_11_ ( .D(o_data_jr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[11]) );
  DFC3 pipe_data_rs_reg_10_ ( .D(o_data_jr[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[10]) );
  DFC3 pipe_data_rs_reg_9_ ( .D(o_data_jr[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[9]) );
  DFC3 pipe_data_rs_reg_8_ ( .D(o_data_jr[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[8]) );
  DFC3 pipe_data_rs_reg_7_ ( .D(o_data_jr[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[7]) );
  DFC3 pipe_data_rs_reg_6_ ( .D(o_data_jr[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[6]) );
  DFC3 pipe_data_rs_reg_5_ ( .D(o_data_jr[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[5]) );
  DFC3 pipe_data_rs_reg_4_ ( .D(o_data_jr[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[4]) );
  DFC3 pipe_data_rs_reg_3_ ( .D(o_data_jr[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[3]) );
  DFC3 pipe_data_rs_reg_2_ ( .D(o_data_jr[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[2]) );
  DFC3 pipe_data_rs_reg_1_ ( .D(o_data_jr[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[1]) );
  DFC3 pipe_data_rs_reg_0_ ( .D(o_data_jr[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rs[0]) );
  DFC3 pipe_data_rt_reg_31_ ( .D(regbank_o_data_Rt[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[31]) );
  DFC3 pipe_data_rt_reg_30_ ( .D(regbank_o_data_Rt[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[30]) );
  DFC3 pipe_data_rt_reg_29_ ( .D(regbank_o_data_Rt[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[29]) );
  DFC3 pipe_data_rt_reg_28_ ( .D(regbank_o_data_Rt[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[28]) );
  DFC3 pipe_data_rt_reg_27_ ( .D(regbank_o_data_Rt[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[27]) );
  DFC3 pipe_data_rt_reg_26_ ( .D(regbank_o_data_Rt[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[26]) );
  DFC3 pipe_data_rt_reg_25_ ( .D(regbank_o_data_Rt[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[25]) );
  DFC3 pipe_data_rt_reg_24_ ( .D(regbank_o_data_Rt[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[24]) );
  DFC3 pipe_data_rt_reg_23_ ( .D(regbank_o_data_Rt[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[23]) );
  DFC3 pipe_data_rt_reg_22_ ( .D(regbank_o_data_Rt[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[22]) );
  DFC3 pipe_data_rt_reg_21_ ( .D(regbank_o_data_Rt[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[21]) );
  DFC3 pipe_data_rt_reg_20_ ( .D(regbank_o_data_Rt[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[20]) );
  DFC3 pipe_data_rt_reg_19_ ( .D(regbank_o_data_Rt[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[19]) );
  DFC3 pipe_data_rt_reg_18_ ( .D(regbank_o_data_Rt[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[18]) );
  DFC3 pipe_data_rt_reg_17_ ( .D(regbank_o_data_Rt[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[17]) );
  DFC3 pipe_data_rt_reg_16_ ( .D(regbank_o_data_Rt[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC3 pipe_data_rt_reg_15_ ( .D(regbank_o_data_Rt[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[15]) );
  DFC3 pipe_data_rt_reg_14_ ( .D(regbank_o_data_Rt[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[14]) );
  DFC3 pipe_data_rt_reg_13_ ( .D(regbank_o_data_Rt[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[13]) );
  DFC3 pipe_data_rt_reg_12_ ( .D(regbank_o_data_Rt[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[12]) );
  DFC3 pipe_data_rt_reg_11_ ( .D(regbank_o_data_Rt[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[11]) );
  DFC3 pipe_data_rt_reg_10_ ( .D(regbank_o_data_Rt[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[10]) );
  DFC3 pipe_data_rt_reg_9_ ( .D(regbank_o_data_Rt[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[9]) );
  DFC3 pipe_data_rt_reg_8_ ( .D(regbank_o_data_Rt[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[8]) );
  DFC3 pipe_data_rt_reg_7_ ( .D(regbank_o_data_Rt[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[7]) );
  DFC3 pipe_data_rt_reg_6_ ( .D(regbank_o_data_Rt[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[6]) );
  DFC3 pipe_data_rt_reg_5_ ( .D(regbank_o_data_Rt[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[5]) );
  DFC3 pipe_data_rt_reg_4_ ( .D(regbank_o_data_Rt[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[4]) );
  DFC3 pipe_data_rt_reg_3_ ( .D(regbank_o_data_Rt[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[3]) );
  DFC3 pipe_data_rt_reg_2_ ( .D(regbank_o_data_Rt[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[2]) );
  DFC3 pipe_data_rt_reg_1_ ( .D(regbank_o_data_Rt[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[1]) );
  DFC3 pipe_data_rt_reg_0_ ( .D(regbank_o_data_Rt[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[0]) );
  DFC3 pipe_addr_rd_reg_4_ ( .D(i_data_instr[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[4]) );
  DFC3 pipe_addr_rd_reg_3_ ( .D(i_data_instr[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[3]) );
  DFC3 pipe_addr_rd_reg_2_ ( .D(i_data_instr[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[2]) );
  DFC3 pipe_addr_rd_reg_1_ ( .D(i_data_instr[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[1]) );
  DFC3 pipe_addr_rd_reg_0_ ( .D(i_data_instr[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rd[0]) );
  DFC3 pipe_addr_rt_reg_4_ ( .D(i_data_instr[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_data_instr[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_data_instr[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_data_instr[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_data_instr[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_rt[0]) );
  DFC3 pipe_addr_pc4_reg_31_ ( .D(i_addr_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[31]) );
  DFC3 pipe_addr_pc4_reg_30_ ( .D(i_addr_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[30]) );
  DFC3 pipe_addr_pc4_reg_29_ ( .D(i_addr_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[29]) );
  DFC3 pipe_addr_pc4_reg_28_ ( .D(i_addr_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[28]) );
  DFC3 pipe_addr_pc4_reg_27_ ( .D(i_addr_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[27]) );
  DFC3 pipe_addr_pc4_reg_26_ ( .D(i_addr_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[26]) );
  DFC3 pipe_addr_pc4_reg_25_ ( .D(i_addr_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[25]) );
  DFC3 pipe_addr_pc4_reg_24_ ( .D(i_addr_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[24]) );
  DFC3 pipe_addr_pc4_reg_23_ ( .D(i_addr_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[23]) );
  DFC3 pipe_addr_pc4_reg_22_ ( .D(i_addr_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[22]) );
  DFC3 pipe_addr_pc4_reg_21_ ( .D(i_addr_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[21]) );
  DFC3 pipe_addr_pc4_reg_20_ ( .D(i_addr_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[20]) );
  DFC3 pipe_addr_pc4_reg_19_ ( .D(i_addr_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[19]) );
  DFC3 pipe_addr_pc4_reg_18_ ( .D(i_addr_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[18]) );
  DFC3 pipe_addr_pc4_reg_17_ ( .D(i_addr_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[17]) );
  DFC3 pipe_addr_pc4_reg_16_ ( .D(i_addr_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[16]) );
  DFC3 pipe_addr_pc4_reg_15_ ( .D(i_addr_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[15]) );
  DFC3 pipe_addr_pc4_reg_14_ ( .D(i_addr_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[14]) );
  DFC3 pipe_addr_pc4_reg_13_ ( .D(i_addr_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[13]) );
  DFC3 pipe_addr_pc4_reg_12_ ( .D(i_addr_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[12]) );
  DFC3 pipe_addr_pc4_reg_11_ ( .D(i_addr_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[11]) );
  DFC3 pipe_addr_pc4_reg_10_ ( .D(i_addr_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[10]) );
  DFC3 pipe_addr_pc4_reg_9_ ( .D(i_addr_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[9]) );
  DFC3 pipe_addr_pc4_reg_8_ ( .D(i_addr_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[8]) );
  DFC3 pipe_addr_pc4_reg_7_ ( .D(i_addr_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[7]) );
  DFC3 pipe_addr_pc4_reg_6_ ( .D(i_addr_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[6]) );
  DFC3 pipe_addr_pc4_reg_5_ ( .D(i_addr_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[5]) );
  DFC3 pipe_addr_pc4_reg_4_ ( .D(i_addr_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[4]) );
  DFC3 pipe_addr_pc4_reg_3_ ( .D(i_addr_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[3]) );
  DFC3 pipe_addr_pc4_reg_2_ ( .D(i_addr_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[2]) );
  DFC3 pipe_addr_pc4_reg_1_ ( .D(i_addr_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[1]) );
  DFC3 pipe_addr_pc4_reg_0_ ( .D(i_addr_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_pc4[0]) );
  DFC3 pipe_con_Ealuop_reg_5_ ( .D(control_o_con_aluop[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[5]) );
  DFC3 pipe_con_Ealuop_reg_4_ ( .D(control_o_con_aluop[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[4]) );
  DFC3 pipe_con_Ealuop_reg_3_ ( .D(control_o_con_aluop[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[3]) );
  DFC3 pipe_con_Ealuop_reg_2_ ( .D(control_o_con_aluop[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[2]) );
  DFC3 pipe_con_Ealuop_reg_1_ ( .D(control_o_con_aluop[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[1]) );
  DFC3 pipe_con_Ealuop_reg_0_ ( .D(control_o_con_aluop[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Ealuop[0]) );
  DFC3 pipe_con_Ealusrc_reg ( .D(control_o_con_alusrc), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Ealusrc) );
  DFC3 pipe_con_Eregdst_reg ( .D(control_o_con_regdst), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Eregdst) );
  DFC3 pipe_con_MaluPC4_reg ( .D(jbcon_o_con_aluPC4), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Malupc8) );
  DFC3 pipe_con_Mmemread_reg ( .D(control_o_con_memread), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(control_o_con_memwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(control_o_con_memtoreg), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(control_o_con_regwrite), .C(i_clk), .RN(
        i_nrst), .Q(o_con_Wregwrite) );
  DFC3 pipe_signext_o_data_immD_reg_31_ ( .D(signext_o_data_immD[31]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[31]) );
  DFC3 pipe_signext_o_data_immD_reg_30_ ( .D(signext_o_data_immD[30]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[30]) );
  DFC3 pipe_signext_o_data_immD_reg_29_ ( .D(signext_o_data_immD[29]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[29]) );
  DFC3 pipe_signext_o_data_immD_reg_28_ ( .D(signext_o_data_immD[28]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[28]) );
  DFC3 pipe_signext_o_data_immD_reg_27_ ( .D(signext_o_data_immD[27]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[27]) );
  DFC3 pipe_signext_o_data_immD_reg_26_ ( .D(signext_o_data_immD[26]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[26]) );
  DFC3 pipe_signext_o_data_immD_reg_25_ ( .D(signext_o_data_immD[25]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[25]) );
  DFC3 pipe_signext_o_data_immD_reg_24_ ( .D(signext_o_data_immD[24]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[24]) );
  DFC3 pipe_signext_o_data_immD_reg_23_ ( .D(signext_o_data_immD[23]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[23]) );
  DFC3 pipe_signext_o_data_immD_reg_22_ ( .D(signext_o_data_immD[22]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[22]) );
  DFC3 pipe_signext_o_data_immD_reg_21_ ( .D(signext_o_data_immD[21]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[21]) );
  DFC3 pipe_signext_o_data_immD_reg_20_ ( .D(signext_o_data_immD[20]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[20]) );
  DFC3 pipe_signext_o_data_immD_reg_19_ ( .D(signext_o_data_immD[19]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[19]) );
  DFC3 pipe_signext_o_data_immD_reg_18_ ( .D(signext_o_data_immD[18]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[18]) );
  DFC3 pipe_signext_o_data_immD_reg_17_ ( .D(signext_o_data_immD[17]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[17]) );
  DFC3 pipe_signext_o_data_immD_reg_16_ ( .D(signext_o_data_immD[16]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[16]) );
  DFC3 pipe_signext_o_data_immD_reg_15_ ( .D(signext_o_data_immD[15]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[15]) );
  DFC3 pipe_signext_o_data_immD_reg_14_ ( .D(signext_o_data_immD[14]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[14]) );
  DFC3 pipe_signext_o_data_immD_reg_13_ ( .D(signext_o_data_immD[13]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[13]) );
  DFC3 pipe_signext_o_data_immD_reg_12_ ( .D(signext_o_data_immD[12]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[12]) );
  DFC3 pipe_signext_o_data_immD_reg_11_ ( .D(signext_o_data_immD[11]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[11]) );
  DFC3 pipe_signext_o_data_immD_reg_10_ ( .D(signext_o_data_immD[10]), .C(
        i_clk), .RN(i_nrst), .Q(o_data_signext[10]) );
  DFC3 pipe_signext_o_data_immD_reg_9_ ( .D(signext_o_data_immD[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[9]) );
  DFC3 pipe_signext_o_data_immD_reg_8_ ( .D(signext_o_data_immD[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[8]) );
  DFC3 pipe_signext_o_data_immD_reg_7_ ( .D(signext_o_data_immD[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[7]) );
  DFC3 pipe_signext_o_data_immD_reg_6_ ( .D(signext_o_data_immD[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[6]) );
  DFC3 pipe_signext_o_data_immD_reg_5_ ( .D(signext_o_data_immD[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[5]) );
  DFC3 pipe_signext_o_data_immD_reg_4_ ( .D(signext_o_data_immD[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[4]) );
  DFC3 pipe_signext_o_data_immD_reg_3_ ( .D(signext_o_data_immD[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[3]) );
  DFC3 pipe_signext_o_data_immD_reg_2_ ( .D(signext_o_data_immD[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[2]) );
  DFC3 pipe_signext_o_data_immD_reg_1_ ( .D(signext_o_data_immD[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[1]) );
  DFC3 pipe_signext_o_data_immD_reg_0_ ( .D(signext_o_data_immD[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_data_signext[0]) );
  DFC3 pipe_con_Efamux_reg_2_ ( .D(for_o_con_fa[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[2]) );
  DFC3 pipe_con_Efamux_reg_1_ ( .D(for_o_con_fa[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[1]) );
  DFC3 pipe_con_Efamux_reg_0_ ( .D(for_o_con_fa[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efamux[0]) );
  DFC3 pipe_con_Efbmux_reg_2_ ( .D(for_o_con_fb[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[2]) );
  DFC3 pipe_con_Efbmux_reg_1_ ( .D(for_o_con_fb[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[1]) );
  DFC3 pipe_con_Efbmux_reg_0_ ( .D(for_o_con_fb[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Efbmux[0]) );
  DFC3 pipe_FWmemout_reg_31_ ( .D(i_data_Wmemout[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[31]) );
  DFC3 pipe_FWmemout_reg_30_ ( .D(i_data_Wmemout[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[30]) );
  DFC3 pipe_FWmemout_reg_29_ ( .D(i_data_Wmemout[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[29]) );
  DFC3 pipe_FWmemout_reg_28_ ( .D(i_data_Wmemout[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[28]) );
  DFC3 pipe_FWmemout_reg_27_ ( .D(i_data_Wmemout[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[27]) );
  DFC3 pipe_FWmemout_reg_26_ ( .D(i_data_Wmemout[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[26]) );
  DFC3 pipe_FWmemout_reg_25_ ( .D(i_data_Wmemout[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[25]) );
  DFC3 pipe_FWmemout_reg_24_ ( .D(i_data_Wmemout[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[24]) );
  DFC3 pipe_FWmemout_reg_23_ ( .D(i_data_Wmemout[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[23]) );
  DFC3 pipe_FWmemout_reg_22_ ( .D(i_data_Wmemout[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[22]) );
  DFC3 pipe_FWmemout_reg_21_ ( .D(i_data_Wmemout[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[21]) );
  DFC3 pipe_FWmemout_reg_20_ ( .D(i_data_Wmemout[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[20]) );
  DFC3 pipe_FWmemout_reg_19_ ( .D(i_data_Wmemout[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[19]) );
  DFC3 pipe_FWmemout_reg_18_ ( .D(i_data_Wmemout[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[18]) );
  DFC3 pipe_FWmemout_reg_17_ ( .D(i_data_Wmemout[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[17]) );
  DFC3 pipe_FWmemout_reg_16_ ( .D(i_data_Wmemout[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[16]) );
  DFC3 pipe_FWmemout_reg_15_ ( .D(i_data_Wmemout[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[15]) );
  DFC3 pipe_FWmemout_reg_14_ ( .D(i_data_Wmemout[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[14]) );
  DFC3 pipe_FWmemout_reg_13_ ( .D(i_data_Wmemout[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[13]) );
  DFC3 pipe_FWmemout_reg_12_ ( .D(i_data_Wmemout[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[12]) );
  DFC3 pipe_FWmemout_reg_11_ ( .D(i_data_Wmemout[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[11]) );
  DFC3 pipe_FWmemout_reg_10_ ( .D(i_data_Wmemout[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[10]) );
  DFC3 pipe_FWmemout_reg_9_ ( .D(i_data_Wmemout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[9]) );
  DFC3 pipe_FWmemout_reg_8_ ( .D(i_data_Wmemout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[8]) );
  DFC3 pipe_FWmemout_reg_7_ ( .D(i_data_Wmemout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[7]) );
  DFC3 pipe_FWmemout_reg_6_ ( .D(i_data_Wmemout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[6]) );
  DFC3 pipe_FWmemout_reg_5_ ( .D(i_data_Wmemout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[5]) );
  DFC3 pipe_FWmemout_reg_4_ ( .D(i_data_Wmemout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[4]) );
  DFC3 pipe_FWmemout_reg_3_ ( .D(i_data_Wmemout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[3]) );
  DFC3 pipe_FWmemout_reg_2_ ( .D(i_data_Wmemout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[2]) );
  DFC3 pipe_FWmemout_reg_1_ ( .D(i_data_Wmemout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[1]) );
  DFC3 pipe_FWmemout_reg_0_ ( .D(i_data_Wmemout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_Fmemout[0]) );
  DFC3 pipe_addr_branch_reg_31_ ( .D(pcadd_o_addr_pcbranchE[31]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[31]) );
  DFC3 pipe_addr_branch_reg_30_ ( .D(pcadd_o_addr_pcbranchE[30]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[30]) );
  DFC3 pipe_addr_branch_reg_29_ ( .D(pcadd_o_addr_pcbranchE[29]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[29]) );
  DFC3 pipe_addr_branch_reg_28_ ( .D(pcadd_o_addr_pcbranchE[28]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[28]) );
  DFC3 pipe_addr_branch_reg_27_ ( .D(pcadd_o_addr_pcbranchE[27]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[27]) );
  DFC3 pipe_addr_branch_reg_26_ ( .D(pcadd_o_addr_pcbranchE[26]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[26]) );
  DFC3 pipe_addr_branch_reg_25_ ( .D(pcadd_o_addr_pcbranchE[25]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[25]) );
  DFC3 pipe_addr_branch_reg_24_ ( .D(pcadd_o_addr_pcbranchE[24]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[24]) );
  DFC3 pipe_addr_branch_reg_23_ ( .D(pcadd_o_addr_pcbranchE[23]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[23]) );
  DFC3 pipe_addr_branch_reg_22_ ( .D(pcadd_o_addr_pcbranchE[22]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[22]) );
  DFC3 pipe_addr_branch_reg_21_ ( .D(pcadd_o_addr_pcbranchE[21]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[21]) );
  DFC3 pipe_addr_branch_reg_20_ ( .D(pcadd_o_addr_pcbranchE[20]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[20]) );
  DFC3 pipe_addr_branch_reg_19_ ( .D(pcadd_o_addr_pcbranchE[19]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[19]) );
  DFC3 pipe_addr_branch_reg_18_ ( .D(pcadd_o_addr_pcbranchE[18]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[18]) );
  DFC3 pipe_addr_branch_reg_17_ ( .D(pcadd_o_addr_pcbranchE[17]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[17]) );
  DFC3 pipe_addr_branch_reg_16_ ( .D(pcadd_o_addr_pcbranchE[16]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[16]) );
  DFC3 pipe_addr_branch_reg_15_ ( .D(pcadd_o_addr_pcbranchE[15]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[15]) );
  DFC3 pipe_addr_branch_reg_14_ ( .D(pcadd_o_addr_pcbranchE[14]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[14]) );
  DFC3 pipe_addr_branch_reg_13_ ( .D(pcadd_o_addr_pcbranchE[13]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[13]) );
  DFC3 pipe_addr_branch_reg_12_ ( .D(pcadd_o_addr_pcbranchE[12]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[12]) );
  DFC3 pipe_addr_branch_reg_11_ ( .D(pcadd_o_addr_pcbranchE[11]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[11]) );
  DFC3 pipe_addr_branch_reg_10_ ( .D(pcadd_o_addr_pcbranchE[10]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[10]) );
  DFC3 pipe_addr_branch_reg_9_ ( .D(pcadd_o_addr_pcbranchE[9]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[9]) );
  DFC3 pipe_addr_branch_reg_8_ ( .D(pcadd_o_addr_pcbranchE[8]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[8]) );
  DFC3 pipe_addr_branch_reg_7_ ( .D(pcadd_o_addr_pcbranchE[7]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[7]) );
  DFC3 pipe_addr_branch_reg_6_ ( .D(pcadd_o_addr_pcbranchE[6]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[6]) );
  DFC3 pipe_addr_branch_reg_5_ ( .D(pcadd_o_addr_pcbranchE[5]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[5]) );
  DFC3 pipe_addr_branch_reg_4_ ( .D(pcadd_o_addr_pcbranchE[4]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[4]) );
  DFC3 pipe_addr_branch_reg_3_ ( .D(pcadd_o_addr_pcbranchE[3]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[3]) );
  DFC3 pipe_addr_branch_reg_2_ ( .D(pcadd_o_addr_pcbranchE[2]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[2]) );
  DFC3 pipe_addr_branch_reg_1_ ( .D(pcadd_o_addr_pcbranchE[1]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[1]) );
  DFC3 pipe_addr_branch_reg_0_ ( .D(pcadd_o_addr_pcbranchE[0]), .C(i_clk), 
        .RN(i_nrst), .Q(o_addr_branch[0]) );
  D_control u_control ( .o_con_regdst(control_o_con_regdst), .o_con_memread(
        control_o_con_memread), .o_con_memtoreg(control_o_con_memtoreg), 
        .o_con_memwrite(control_o_con_memwrite), .o_con_alusrc(
        control_o_con_alusrc), .o_con_regwrite(control_o_con_regwrite), 
        .o_con_ifsign(signext_i_con_signext), .o_con_aluop(control_o_con_aluop), .i_con_instru(i_data_instr[31:26]) );
  D_jb_control u_jb_control ( .o_con_jump(o_con_jump), .o_con_bop(
        jbcon_o_con_bop), .o_con_aluPC4(jbcon_o_con_aluPC4), .o_con_ifstall(
        o_con_ifstall), .i_con_instru(i_data_instr[31:26]), .i_con_func(
        i_data_instr[5:0]), .i_con_rt(i_data_instr[16]) );
  D_pcadd u_pcadd ( .i_addr_pcadd4E(i_addr_pc4), .i_data_immshiftl({
        pcadd_i_data_immshiftl, o_addr_jump[0], o_addr_jump[0]}), 
        .o_addr_pcbranchE(pcadd_o_addr_pcbranchE) );
  D_register_bank u_regbank ( .i_clk(i_clk), .i_rst_n(i_nrst), .i_addr_Rs(
        i_data_instr[25:21]), .i_addr_Rt(i_data_instr[20:16]), .i_con_RegWr(
        i_con_Wregwrite), .i_addr_Rd(i_addr_Wregwrite), .i_data_Rd(
        i_data_Wregwrite), .o_data_Rs(o_data_jr), .o_data_Rt(regbank_o_data_Rt) );
  D_shiftleft u_sl ( .i_data_immE(i_data_instr[15:0]), .o_data_immshiftl({
        pcadd_i_data_immshiftl, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2}) );
  D_sign_extend u_signext ( .i_data_immD(i_data_instr[15:0]), .i_con_signext(
        signext_i_con_signext), .o_data_immD(signext_o_data_immD) );
  D_jump_ext u_jump_ext ( .i_addr_j(i_data_instr[25:0]), .i_PC4_j(
        i_addr_pc4[31:28]), .o_addr_j({o_addr_jump[31:2], 
        SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4}) );
  D_forward u_forward ( .i_addr_rs(i_data_instr[25:21]), .i_addr_rt(
        i_data_instr[20:16]), .i_addr_rdE(i_addr_Erd), .i_addr_rdM(i_addr_Mrd), 
        .i_addr_rtM(i_addr_rtM), .i_addr_rtW(i_addr_rtW), .i_con_regwriteE(
        i_con_Eregwrite), .i_con_regwriteM(i_con_Mregwrite), .i_con_memreadM(
        i_con_memreadM), .i_con_memreadW(i_con_memreadW), .o_con_fa(
        for_o_con_fa), .o_con_fb(for_o_con_fb) );
  LOGIC0 U3 ( .Q(o_addr_jump[0]) );
endmodule


module E_alu_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   ML_int_1__31_, ML_int_1__30_, ML_int_1__29_, ML_int_1__28_,
         ML_int_1__27_, ML_int_1__26_, ML_int_1__25_, ML_int_1__24_,
         ML_int_1__23_, ML_int_1__22_, ML_int_1__21_, ML_int_1__20_,
         ML_int_1__19_, ML_int_1__18_, ML_int_1__17_, ML_int_1__16_,
         ML_int_1__15_, ML_int_1__14_, ML_int_1__13_, ML_int_1__12_,
         ML_int_1__11_, ML_int_1__10_, ML_int_1__9_, ML_int_1__8_,
         ML_int_1__7_, ML_int_1__6_, ML_int_1__5_, ML_int_1__4_, ML_int_1__3_,
         ML_int_1__2_, ML_int_1__1_, ML_int_1__0_, ML_int_2__31_,
         ML_int_2__30_, ML_int_2__29_, ML_int_2__28_, ML_int_2__27_,
         ML_int_2__26_, ML_int_2__25_, ML_int_2__24_, ML_int_2__23_,
         ML_int_2__22_, ML_int_2__21_, ML_int_2__20_, ML_int_2__19_,
         ML_int_2__18_, ML_int_2__17_, ML_int_2__16_, ML_int_2__15_,
         ML_int_2__14_, ML_int_2__13_, ML_int_2__12_, ML_int_2__11_,
         ML_int_2__10_, ML_int_2__9_, ML_int_2__8_, ML_int_2__7_, ML_int_2__6_,
         ML_int_2__5_, ML_int_2__4_, ML_int_2__3_, ML_int_2__2_, ML_int_3__31_,
         ML_int_3__30_, ML_int_3__29_, ML_int_3__28_, ML_int_3__27_,
         ML_int_3__26_, ML_int_3__25_, ML_int_3__24_, ML_int_3__23_,
         ML_int_3__22_, ML_int_3__21_, ML_int_3__20_, ML_int_3__19_,
         ML_int_3__18_, ML_int_3__17_, ML_int_3__16_, ML_int_3__15_,
         ML_int_3__14_, ML_int_3__13_, ML_int_3__12_, ML_int_3__11_,
         ML_int_3__10_, ML_int_3__9_, ML_int_3__8_, ML_int_3__7_, ML_int_3__6_,
         ML_int_3__5_, ML_int_3__4_, ML_int_3__1_, ML_int_3__0_, ML_int_4__31_,
         ML_int_4__30_, ML_int_4__29_, ML_int_4__28_, ML_int_4__27_,
         ML_int_4__26_, ML_int_4__25_, ML_int_4__24_, ML_int_4__15_,
         ML_int_4__14_, ML_int_4__13_, ML_int_4__12_, ML_int_4__11_,
         ML_int_4__10_, ML_int_4__9_, ML_int_4__8_, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36;

  MUX21 U3 ( .A(A[4]), .B(A[3]), .S(SH[0]), .Q(ML_int_1__4_) );
  MUX21 U4 ( .A(A[3]), .B(A[2]), .S(SH[0]), .Q(ML_int_1__3_) );
  MUX21 U5 ( .A(A[20]), .B(A[19]), .S(SH[0]), .Q(ML_int_1__20_) );
  MUX21 U6 ( .A(A[21]), .B(A[20]), .S(SH[0]), .Q(ML_int_1__21_) );
  INV0 U7 ( .A(A[0]), .Q(n24) );
  MUX21 U8 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Q(ML_int_1__1_) );
  MUX21 U9 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Q(ML_int_1__8_) );
  MUX21 U10 ( .A(A[9]), .B(A[8]), .S(SH[0]), .Q(ML_int_1__9_) );
  MUX21 U11 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Q(ML_int_1__10_) );
  MUX21 U12 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Q(ML_int_1__2_) );
  MUX21 U13 ( .A(A[17]), .B(A[16]), .S(SH[0]), .Q(ML_int_1__17_) );
  MUX21 U14 ( .A(A[16]), .B(A[15]), .S(SH[0]), .Q(ML_int_1__16_) );
  MUX21 U15 ( .A(A[18]), .B(A[17]), .S(SH[0]), .Q(ML_int_1__18_) );
  MUX22 U16 ( .A(ML_int_3__8_), .B(ML_int_3__0_), .S(SH[3]), .Q(ML_int_4__8_)
         );
  MUX22 U17 ( .A(ML_int_1__2_), .B(ML_int_1__0_), .S(SH[1]), .Q(ML_int_2__2_)
         );
  MUX22 U18 ( .A(ML_int_2__4_), .B(n23), .S(SH[2]), .Q(ML_int_3__4_) );
  INV3 U19 ( .A(n36), .Q(n23) );
  MUX22 U20 ( .A(ML_int_3__9_), .B(ML_int_3__1_), .S(SH[3]), .Q(ML_int_4__9_)
         );
  MUX22 U21 ( .A(ML_int_1__8_), .B(ML_int_1__6_), .S(SH[1]), .Q(ML_int_2__8_)
         );
  MUX22 U22 ( .A(ML_int_1__11_), .B(ML_int_1__9_), .S(SH[1]), .Q(ML_int_2__11_) );
  MUX22 U23 ( .A(ML_int_1__7_), .B(ML_int_1__5_), .S(SH[1]), .Q(ML_int_2__7_)
         );
  MUX22 U24 ( .A(ML_int_1__9_), .B(ML_int_1__7_), .S(SH[1]), .Q(ML_int_2__9_)
         );
  MUX22 U25 ( .A(ML_int_1__10_), .B(ML_int_1__8_), .S(SH[1]), .Q(ML_int_2__10_) );
  MUX22 U26 ( .A(ML_int_1__12_), .B(ML_int_1__10_), .S(SH[1]), .Q(
        ML_int_2__12_) );
  MUX22 U27 ( .A(ML_int_1__13_), .B(ML_int_1__11_), .S(SH[1]), .Q(
        ML_int_2__13_) );
  MUX22 U28 ( .A(ML_int_1__14_), .B(ML_int_1__12_), .S(SH[1]), .Q(
        ML_int_2__14_) );
  MUX22 U29 ( .A(ML_int_1__4_), .B(ML_int_1__2_), .S(SH[1]), .Q(ML_int_2__4_)
         );
  MUX22 U30 ( .A(ML_int_1__5_), .B(ML_int_1__3_), .S(SH[1]), .Q(ML_int_2__5_)
         );
  MUX22 U31 ( .A(ML_int_1__6_), .B(ML_int_1__4_), .S(SH[1]), .Q(ML_int_2__6_)
         );
  MUX22 U32 ( .A(ML_int_1__15_), .B(ML_int_1__13_), .S(SH[1]), .Q(
        ML_int_2__15_) );
  MUX22 U33 ( .A(ML_int_2__8_), .B(ML_int_2__4_), .S(SH[2]), .Q(ML_int_3__8_)
         );
  MUX22 U34 ( .A(ML_int_2__9_), .B(ML_int_2__5_), .S(SH[2]), .Q(ML_int_3__9_)
         );
  MUX22 U35 ( .A(ML_int_2__10_), .B(ML_int_2__6_), .S(SH[2]), .Q(ML_int_3__10_) );
  MUX22 U36 ( .A(ML_int_2__15_), .B(ML_int_2__11_), .S(SH[2]), .Q(
        ML_int_3__15_) );
  MUX22 U37 ( .A(ML_int_2__18_), .B(ML_int_2__14_), .S(SH[2]), .Q(
        ML_int_3__18_) );
  MUX22 U38 ( .A(ML_int_2__11_), .B(ML_int_2__7_), .S(SH[2]), .Q(ML_int_3__11_) );
  MUX22 U39 ( .A(ML_int_2__12_), .B(ML_int_2__8_), .S(SH[2]), .Q(ML_int_3__12_) );
  MUX22 U40 ( .A(ML_int_2__13_), .B(ML_int_2__9_), .S(SH[2]), .Q(ML_int_3__13_) );
  MUX22 U41 ( .A(ML_int_2__14_), .B(ML_int_2__10_), .S(SH[2]), .Q(
        ML_int_3__14_) );
  MUX22 U42 ( .A(ML_int_3__10_), .B(n21), .S(SH[3]), .Q(ML_int_4__10_) );
  MUX22 U43 ( .A(ML_int_3__15_), .B(ML_int_3__7_), .S(SH[3]), .Q(ML_int_4__15_) );
  MUX22 U44 ( .A(ML_int_3__11_), .B(n20), .S(SH[3]), .Q(ML_int_4__11_) );
  MUX22 U45 ( .A(ML_int_3__12_), .B(ML_int_3__4_), .S(SH[3]), .Q(ML_int_4__12_) );
  MUX22 U46 ( .A(ML_int_3__13_), .B(ML_int_3__5_), .S(SH[3]), .Q(ML_int_4__13_) );
  MUX22 U47 ( .A(ML_int_3__14_), .B(ML_int_3__6_), .S(SH[3]), .Q(ML_int_4__14_) );
  MUX22 U48 ( .A(ML_int_1__3_), .B(ML_int_1__1_), .S(SH[1]), .Q(ML_int_2__3_)
         );
  MUX22 U49 ( .A(ML_int_2__7_), .B(ML_int_2__3_), .S(SH[2]), .Q(ML_int_3__7_)
         );
  MUX22 U50 ( .A(ML_int_2__5_), .B(n22), .S(SH[2]), .Q(ML_int_3__5_) );
  INV3 U51 ( .A(n35), .Q(n22) );
  MUX22 U52 ( .A(ML_int_2__6_), .B(ML_int_2__2_), .S(SH[2]), .Q(ML_int_3__6_)
         );
  MUX22 U53 ( .A(ML_int_1__16_), .B(ML_int_1__14_), .S(SH[1]), .Q(
        ML_int_2__16_) );
  MUX22 U54 ( .A(ML_int_1__24_), .B(ML_int_1__22_), .S(SH[1]), .Q(
        ML_int_2__24_) );
  MUX22 U55 ( .A(ML_int_1__20_), .B(ML_int_1__18_), .S(SH[1]), .Q(
        ML_int_2__20_) );
  MUX22 U56 ( .A(ML_int_1__17_), .B(ML_int_1__15_), .S(SH[1]), .Q(
        ML_int_2__17_) );
  MUX22 U57 ( .A(ML_int_1__21_), .B(ML_int_1__19_), .S(SH[1]), .Q(
        ML_int_2__21_) );
  MUX22 U58 ( .A(ML_int_1__25_), .B(ML_int_1__23_), .S(SH[1]), .Q(
        ML_int_2__25_) );
  MUX22 U59 ( .A(ML_int_1__18_), .B(ML_int_1__16_), .S(SH[1]), .Q(
        ML_int_2__18_) );
  MUX22 U60 ( .A(ML_int_1__22_), .B(ML_int_1__20_), .S(SH[1]), .Q(
        ML_int_2__22_) );
  MUX22 U61 ( .A(ML_int_1__26_), .B(ML_int_1__24_), .S(SH[1]), .Q(
        ML_int_2__26_) );
  MUX22 U62 ( .A(ML_int_1__19_), .B(ML_int_1__17_), .S(SH[1]), .Q(
        ML_int_2__19_) );
  MUX22 U63 ( .A(ML_int_1__23_), .B(ML_int_1__21_), .S(SH[1]), .Q(
        ML_int_2__23_) );
  MUX22 U64 ( .A(ML_int_1__27_), .B(ML_int_1__25_), .S(SH[1]), .Q(
        ML_int_2__27_) );
  MUX22 U65 ( .A(ML_int_2__16_), .B(ML_int_2__12_), .S(SH[2]), .Q(
        ML_int_3__16_) );
  MUX22 U66 ( .A(ML_int_2__17_), .B(ML_int_2__13_), .S(SH[2]), .Q(
        ML_int_3__17_) );
  MUX22 U67 ( .A(ML_int_2__19_), .B(ML_int_2__15_), .S(SH[2]), .Q(
        ML_int_3__19_) );
  MUX22 U68 ( .A(ML_int_2__20_), .B(ML_int_2__16_), .S(SH[2]), .Q(
        ML_int_3__20_) );
  MUX22 U69 ( .A(ML_int_2__21_), .B(ML_int_2__17_), .S(SH[2]), .Q(
        ML_int_3__21_) );
  MUX22 U70 ( .A(ML_int_2__22_), .B(ML_int_2__18_), .S(SH[2]), .Q(
        ML_int_3__22_) );
  MUX22 U71 ( .A(ML_int_2__23_), .B(ML_int_2__19_), .S(SH[2]), .Q(
        ML_int_3__23_) );
  MUX22 U72 ( .A(ML_int_3__27_), .B(ML_int_3__19_), .S(SH[3]), .Q(
        ML_int_4__27_) );
  MUX22 U73 ( .A(ML_int_2__27_), .B(ML_int_2__23_), .S(SH[2]), .Q(
        ML_int_3__27_) );
  MUX22 U74 ( .A(ML_int_3__28_), .B(ML_int_3__20_), .S(SH[3]), .Q(
        ML_int_4__28_) );
  MUX22 U75 ( .A(ML_int_2__28_), .B(ML_int_2__24_), .S(SH[2]), .Q(
        ML_int_3__28_) );
  MUX22 U76 ( .A(ML_int_1__28_), .B(ML_int_1__26_), .S(SH[1]), .Q(
        ML_int_2__28_) );
  MUX22 U77 ( .A(ML_int_3__29_), .B(ML_int_3__21_), .S(SH[3]), .Q(
        ML_int_4__29_) );
  MUX22 U78 ( .A(ML_int_2__29_), .B(ML_int_2__25_), .S(SH[2]), .Q(
        ML_int_3__29_) );
  MUX22 U79 ( .A(ML_int_1__29_), .B(ML_int_1__27_), .S(SH[1]), .Q(
        ML_int_2__29_) );
  MUX22 U80 ( .A(ML_int_4__29_), .B(ML_int_4__13_), .S(SH[4]), .Q(B[29]) );
  MUX22 U81 ( .A(ML_int_4__30_), .B(ML_int_4__14_), .S(SH[4]), .Q(B[30]) );
  MUX22 U82 ( .A(ML_int_4__27_), .B(ML_int_4__11_), .S(SH[4]), .Q(B[27]) );
  MUX22 U83 ( .A(ML_int_4__28_), .B(ML_int_4__12_), .S(SH[4]), .Q(B[28]) );
  INV3 U84 ( .A(ML_int_4__8_), .Q(n19) );
  INV3 U85 ( .A(n34), .Q(n21) );
  IMUX21 U86 ( .A(n1), .B(n32), .S(SH[4]), .Q(B[16]) );
  IMUX21 U87 ( .A(ML_int_3__16_), .B(ML_int_3__8_), .S(SH[3]), .Q(n1) );
  IMUX21 U88 ( .A(n2), .B(n31), .S(SH[4]), .Q(B[17]) );
  IMUX21 U89 ( .A(ML_int_3__17_), .B(ML_int_3__9_), .S(SH[3]), .Q(n2) );
  IMUX21 U90 ( .A(n3), .B(n28), .S(SH[4]), .Q(B[20]) );
  IMUX21 U91 ( .A(ML_int_3__20_), .B(ML_int_3__12_), .S(SH[3]), .Q(n3) );
  INV3 U92 ( .A(ML_int_4__10_), .Q(n17) );
  INV3 U93 ( .A(ML_int_4__11_), .Q(n16) );
  INV3 U94 ( .A(ML_int_4__12_), .Q(n15) );
  INV3 U95 ( .A(ML_int_4__13_), .Q(n14) );
  INV3 U96 ( .A(ML_int_4__14_), .Q(n13) );
  INV3 U97 ( .A(ML_int_4__15_), .Q(n12) );
  INV3 U98 ( .A(n33), .Q(n20) );
  MUX22 U99 ( .A(A[11]), .B(A[10]), .S(SH[0]), .Q(ML_int_1__11_) );
  MUX22 U100 ( .A(A[7]), .B(A[6]), .S(SH[0]), .Q(ML_int_1__7_) );
  MUX22 U101 ( .A(A[12]), .B(A[11]), .S(SH[0]), .Q(ML_int_1__12_) );
  MUX22 U102 ( .A(A[14]), .B(A[13]), .S(SH[0]), .Q(ML_int_1__14_) );
  MUX22 U103 ( .A(A[13]), .B(A[12]), .S(SH[0]), .Q(ML_int_1__13_) );
  MUX22 U104 ( .A(A[6]), .B(A[5]), .S(SH[0]), .Q(ML_int_1__6_) );
  MUX22 U105 ( .A(A[5]), .B(A[4]), .S(SH[0]), .Q(ML_int_1__5_) );
  MUX22 U106 ( .A(A[15]), .B(A[14]), .S(SH[0]), .Q(ML_int_1__15_) );
  MUX22 U107 ( .A(ML_int_4__24_), .B(ML_int_4__8_), .S(SH[4]), .Q(B[24]) );
  MUX22 U108 ( .A(ML_int_3__24_), .B(ML_int_3__16_), .S(SH[3]), .Q(
        ML_int_4__24_) );
  MUX22 U109 ( .A(ML_int_2__24_), .B(ML_int_2__20_), .S(SH[2]), .Q(
        ML_int_3__24_) );
  MUX22 U110 ( .A(ML_int_4__25_), .B(ML_int_4__9_), .S(SH[4]), .Q(B[25]) );
  MUX22 U111 ( .A(ML_int_3__25_), .B(ML_int_3__17_), .S(SH[3]), .Q(
        ML_int_4__25_) );
  MUX22 U112 ( .A(ML_int_2__25_), .B(ML_int_2__21_), .S(SH[2]), .Q(
        ML_int_3__25_) );
  IMUX21 U113 ( .A(n4), .B(n30), .S(SH[4]), .Q(B[18]) );
  IMUX21 U114 ( .A(ML_int_3__18_), .B(ML_int_3__10_), .S(SH[3]), .Q(n4) );
  IMUX21 U115 ( .A(n5), .B(n29), .S(SH[4]), .Q(B[19]) );
  IMUX21 U116 ( .A(ML_int_3__19_), .B(ML_int_3__11_), .S(SH[3]), .Q(n5) );
  IMUX21 U117 ( .A(n6), .B(n27), .S(SH[4]), .Q(B[21]) );
  IMUX21 U118 ( .A(ML_int_3__21_), .B(ML_int_3__13_), .S(SH[3]), .Q(n6) );
  IMUX21 U119 ( .A(n7), .B(n26), .S(SH[4]), .Q(B[22]) );
  IMUX21 U120 ( .A(ML_int_3__22_), .B(ML_int_3__14_), .S(SH[3]), .Q(n7) );
  IMUX21 U121 ( .A(n8), .B(n25), .S(SH[4]), .Q(B[23]) );
  IMUX21 U122 ( .A(ML_int_3__23_), .B(ML_int_3__15_), .S(SH[3]), .Q(n8) );
  MUX22 U123 ( .A(ML_int_4__26_), .B(ML_int_4__10_), .S(SH[4]), .Q(B[26]) );
  MUX22 U124 ( .A(ML_int_3__26_), .B(ML_int_3__18_), .S(SH[3]), .Q(
        ML_int_4__26_) );
  MUX22 U125 ( .A(ML_int_2__26_), .B(ML_int_2__22_), .S(SH[2]), .Q(
        ML_int_3__26_) );
  MUX22 U126 ( .A(ML_int_4__31_), .B(ML_int_4__15_), .S(SH[4]), .Q(B[31]) );
  MUX22 U127 ( .A(ML_int_3__31_), .B(ML_int_3__23_), .S(SH[3]), .Q(
        ML_int_4__31_) );
  MUX22 U128 ( .A(ML_int_2__31_), .B(ML_int_2__27_), .S(SH[2]), .Q(
        ML_int_3__31_) );
  MUX22 U129 ( .A(ML_int_1__31_), .B(ML_int_1__29_), .S(SH[1]), .Q(
        ML_int_2__31_) );
  INV3 U130 ( .A(ML_int_4__9_), .Q(n18) );
  MUX22 U131 ( .A(A[24]), .B(A[23]), .S(SH[0]), .Q(ML_int_1__24_) );
  MUX22 U132 ( .A(A[19]), .B(A[18]), .S(SH[0]), .Q(ML_int_1__19_) );
  MUX22 U133 ( .A(A[22]), .B(A[21]), .S(SH[0]), .Q(ML_int_1__22_) );
  MUX22 U134 ( .A(A[26]), .B(A[25]), .S(SH[0]), .Q(ML_int_1__26_) );
  MUX22 U135 ( .A(A[28]), .B(A[27]), .S(SH[0]), .Q(ML_int_1__28_) );
  MUX22 U136 ( .A(A[27]), .B(A[26]), .S(SH[0]), .Q(ML_int_1__27_) );
  MUX22 U137 ( .A(A[25]), .B(A[24]), .S(SH[0]), .Q(ML_int_1__25_) );
  MUX22 U138 ( .A(A[29]), .B(A[28]), .S(SH[0]), .Q(ML_int_1__29_) );
  MUX22 U139 ( .A(A[23]), .B(A[22]), .S(SH[0]), .Q(ML_int_1__23_) );
  MUX22 U140 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Q(ML_int_1__31_) );
  MUX22 U141 ( .A(ML_int_3__30_), .B(ML_int_3__22_), .S(SH[3]), .Q(
        ML_int_4__30_) );
  MUX22 U142 ( .A(ML_int_2__30_), .B(ML_int_2__26_), .S(SH[2]), .Q(
        ML_int_3__30_) );
  MUX22 U143 ( .A(ML_int_1__30_), .B(ML_int_1__28_), .S(SH[1]), .Q(
        ML_int_2__30_) );
  MUX22 U144 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Q(ML_int_1__30_) );
  INV3 U145 ( .A(SH[2]), .Q(n10) );
  INV3 U146 ( .A(SH[1]), .Q(n9) );
  INV3 U147 ( .A(SH[3]), .Q(n11) );
  NOR20 U148 ( .A(SH[4]), .B(n18), .Q(B[9]) );
  NOR20 U149 ( .A(SH[4]), .B(n19), .Q(B[8]) );
  NOR20 U150 ( .A(SH[4]), .B(n25), .Q(B[7]) );
  NOR20 U151 ( .A(SH[4]), .B(n26), .Q(B[6]) );
  NOR20 U152 ( .A(SH[4]), .B(n27), .Q(B[5]) );
  NOR20 U153 ( .A(SH[4]), .B(n28), .Q(B[4]) );
  NOR20 U154 ( .A(SH[4]), .B(n29), .Q(B[3]) );
  NOR20 U155 ( .A(SH[4]), .B(n30), .Q(B[2]) );
  NOR20 U156 ( .A(SH[4]), .B(n31), .Q(B[1]) );
  NOR20 U157 ( .A(SH[4]), .B(n12), .Q(B[15]) );
  NOR20 U158 ( .A(SH[4]), .B(n13), .Q(B[14]) );
  NOR20 U159 ( .A(SH[4]), .B(n14), .Q(B[13]) );
  NOR20 U160 ( .A(SH[4]), .B(n15), .Q(B[12]) );
  NOR20 U161 ( .A(SH[4]), .B(n16), .Q(B[11]) );
  NOR20 U162 ( .A(SH[4]), .B(n17), .Q(B[10]) );
  NOR20 U163 ( .A(SH[4]), .B(n32), .Q(B[0]) );
  NAND20 U164 ( .A(ML_int_3__7_), .B(n11), .Q(n25) );
  NAND20 U165 ( .A(ML_int_3__6_), .B(n11), .Q(n26) );
  NAND20 U166 ( .A(ML_int_3__5_), .B(n11), .Q(n27) );
  NAND20 U167 ( .A(ML_int_3__4_), .B(n11), .Q(n28) );
  NAND20 U168 ( .A(n20), .B(n11), .Q(n29) );
  NAND20 U169 ( .A(n21), .B(n11), .Q(n30) );
  NAND20 U170 ( .A(ML_int_3__1_), .B(n11), .Q(n31) );
  NAND20 U171 ( .A(ML_int_3__0_), .B(n11), .Q(n32) );
  NAND20 U172 ( .A(ML_int_2__3_), .B(n10), .Q(n33) );
  NAND20 U173 ( .A(ML_int_2__2_), .B(n10), .Q(n34) );
  NOR20 U174 ( .A(n35), .B(SH[2]), .Q(ML_int_3__1_) );
  NOR20 U175 ( .A(n36), .B(SH[2]), .Q(ML_int_3__0_) );
  NAND20 U176 ( .A(ML_int_1__1_), .B(n9), .Q(n35) );
  NAND20 U177 ( .A(ML_int_1__0_), .B(n9), .Q(n36) );
  NOR20 U178 ( .A(n24), .B(SH[0]), .Q(ML_int_1__0_) );
endmodule


module E_alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [15:1] carry;

  ADD32 U2_14 ( .A(A[14]), .B(n10), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADD32 U2_12 ( .A(A[12]), .B(n12), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADD32 U2_11 ( .A(A[11]), .B(n13), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADD32 U2_10 ( .A(A[10]), .B(n14), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADD32 U2_9 ( .A(A[9]), .B(n15), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADD32 U2_8 ( .A(A[8]), .B(n16), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADD32 U2_6 ( .A(A[6]), .B(n18), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADD32 U2_5 ( .A(A[5]), .B(n19), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADD32 U2_4 ( .A(A[4]), .B(n20), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADD32 U2_3 ( .A(A[3]), .B(n21), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADD32 U2_2 ( .A(A[2]), .B(n22), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADD32 U2_1 ( .A(A[1]), .B(n23), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  CLKIN3 U1 ( .A(n1), .Q(n2) );
  NAND22 U2 ( .A(n5), .B(n2), .Q(carry[14]) );
  NAND22 U3 ( .A(A[0]), .B(n24), .Q(n3) );
  NAND22 U4 ( .A(carry[7]), .B(A[7]), .Q(n8) );
  NAND21 U5 ( .A(carry[13]), .B(A[13]), .Q(n5) );
  NAND22 U6 ( .A(carry[13]), .B(n11), .Q(n4) );
  NAND33 U7 ( .A(n7), .B(n8), .C(n9), .Q(carry[8]) );
  NAND22 U8 ( .A(n11), .B(A[13]), .Q(n6) );
  NAND22 U9 ( .A(n4), .B(n6), .Q(n1) );
  XNR31 U10 ( .A(A[15]), .B(B[15]), .C(carry[15]), .Q(DIFF[15]) );
  XOR20 U11 ( .A(A[0]), .B(n24), .Q(DIFF[0]) );
  INV3 U12 ( .A(B[6]), .Q(n18) );
  INV3 U13 ( .A(B[12]), .Q(n12) );
  INV3 U14 ( .A(B[8]), .Q(n16) );
  INV3 U15 ( .A(B[2]), .Q(n22) );
  INV3 U16 ( .A(B[3]), .Q(n21) );
  INV3 U17 ( .A(B[9]), .Q(n15) );
  INV3 U18 ( .A(B[10]), .Q(n14) );
  INV3 U19 ( .A(B[11]), .Q(n13) );
  INV3 U20 ( .A(B[4]), .Q(n20) );
  INV3 U21 ( .A(B[5]), .Q(n19) );
  INV3 U22 ( .A(B[14]), .Q(n10) );
  INV3 U23 ( .A(B[0]), .Q(n24) );
  INV3 U24 ( .A(B[1]), .Q(n23) );
  INV3 U25 ( .A(n3), .Q(carry[1]) );
  XOR31 U26 ( .A(carry[13]), .B(n11), .C(A[13]), .Q(DIFF[13]) );
  XOR31 U27 ( .A(carry[7]), .B(n17), .C(A[7]), .Q(DIFF[7]) );
  NAND22 U28 ( .A(carry[7]), .B(n17), .Q(n7) );
  NAND22 U29 ( .A(n17), .B(A[7]), .Q(n9) );
  INV3 U30 ( .A(B[13]), .Q(n11) );
  INV3 U31 ( .A(B[7]), .Q(n17) );
endmodule


module E_alu_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  ADD32 U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(DIFF[14]) );
  ADD32 U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(DIFF[13]) );
  ADD32 U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(DIFF[12]) );
  ADD32 U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(DIFF[11]) );
  ADD32 U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(DIFF[10]) );
  ADD32 U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9]) );
  ADD32 U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  ADD32 U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  ADD32 U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADD32 U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADD32 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADD32 U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADD32 U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADD32 U1 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  NOR21 U2 ( .A(n17), .B(A[0]), .Q(n1) );
  XNR20 U3 ( .A(A[0]), .B(n17), .Q(DIFF[0]) );
  INV3 U4 ( .A(B[15]), .Q(n2) );
  INV3 U5 ( .A(B[7]), .Q(n10) );
  INV3 U6 ( .A(B[13]), .Q(n4) );
  INV3 U7 ( .A(B[8]), .Q(n9) );
  INV3 U8 ( .A(B[1]), .Q(n16) );
  INV3 U9 ( .A(n1), .Q(carry[1]) );
  INV3 U10 ( .A(B[2]), .Q(n15) );
  INV3 U11 ( .A(B[3]), .Q(n14) );
  INV3 U12 ( .A(B[6]), .Q(n11) );
  INV3 U13 ( .A(B[4]), .Q(n13) );
  INV3 U14 ( .A(B[5]), .Q(n12) );
  INV3 U15 ( .A(B[9]), .Q(n8) );
  INV3 U16 ( .A(B[10]), .Q(n7) );
  INV3 U17 ( .A(B[11]), .Q(n6) );
  INV3 U18 ( .A(B[12]), .Q(n5) );
  INV3 U19 ( .A(B[14]), .Q(n3) );
  INV3 U20 ( .A(B[0]), .Q(n17) );
  XOR31 U21 ( .A(A[15]), .B(n2), .C(carry[15]), .Q(DIFF[15]) );
endmodule


module E_alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR31 U1 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Q(SUM[7]) );
  INV3 U2 ( .A(n1), .Q(carry[1]) );
  NOR21 U3 ( .A(B[0]), .B(A[0]), .Q(n1) );
  XNR21 U4 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
endmodule


module E_alu_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR31 U1 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Q(SUM[7]) );
  XOR21 U2 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  INV3 U3 ( .A(n1), .Q(carry[1]) );
  NAND22 U4 ( .A(A[0]), .B(B[0]), .Q(n1) );
endmodule


module E_alu_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  ADD31 U1 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD31 U2 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  NOR20 U3 ( .A(B[0]), .B(A[0]), .Q(n1) );
  ADD31 U4 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XNR20 U5 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  INV3 U6 ( .A(n1), .Q(carry[1]) );
endmodule


module E_alu_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  XOR20 U1 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  NAND20 U2 ( .A(A[0]), .B(B[0]), .Q(n1) );
  ADD31 U3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  INV3 U4 ( .A(n1), .Q(carry[1]) );
endmodule


module E_alu_DW01_add_4 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKIN3 U1 ( .A(n1), .Q(carry[1]) );
  XNR20 U2 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  NOR21 U3 ( .A(B[0]), .B(A[0]), .Q(n1) );
endmodule


module E_alu_DW01_add_5 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND21 U1 ( .A(A[0]), .B(B[0]), .Q(n1) );
  XOR20 U2 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  INV3 U3 ( .A(n1), .Q(carry[1]) );
endmodule


module E_alu_DW01_add_6 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  ADD31 U1 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  XOR20 U2 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  INV3 U3 ( .A(n1), .Q(carry[1]) );
  NAND22 U4 ( .A(A[0]), .B(B[0]), .Q(n1) );
endmodule


module E_alu_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211;

  INV3 U3 ( .A(n126), .Q(n29) );
  INV3 U4 ( .A(n103), .Q(n24) );
  INV3 U5 ( .A(n113), .Q(n15) );
  INV3 U6 ( .A(n138), .Q(n34) );
  INV3 U7 ( .A(n116), .Q(n32) );
  INV3 U8 ( .A(n142), .Q(n31) );
  INV3 U9 ( .A(n102), .Q(n21) );
  INV3 U10 ( .A(n164), .Q(n33) );
  INV3 U11 ( .A(n69), .Q(n20) );
  BUF2 U12 ( .A(n97), .Q(n4) );
  INV3 U13 ( .A(n70), .Q(n37) );
  INV3 U14 ( .A(n91), .Q(n46) );
  INV3 U15 ( .A(n63), .Q(n28) );
  INV3 U16 ( .A(A[18]), .Q(n38) );
  INV3 U17 ( .A(A[19]), .Q(n36) );
  INV3 U18 ( .A(n78), .Q(n35) );
  INV3 U19 ( .A(n159), .Q(n17) );
  INV3 U20 ( .A(n118), .Q(n49) );
  INV3 U21 ( .A(n145), .Q(n26) );
  INV3 U22 ( .A(n87), .Q(n27) );
  INV3 U23 ( .A(n82), .Q(n16) );
  INV3 U24 ( .A(n76), .Q(n25) );
  INV3 U25 ( .A(n92), .Q(n19) );
  INV3 U26 ( .A(n129), .Q(n13) );
  INV3 U27 ( .A(n106), .Q(n23) );
  INV3 U28 ( .A(n110), .Q(n43) );
  BUF2 U29 ( .A(n96), .Q(n3) );
  BUF2 U30 ( .A(n95), .Q(n2) );
  INV3 U31 ( .A(n58), .Q(n47) );
  NOR21 U32 ( .A(n49), .B(n11), .Q(n91) );
  INV3 U33 ( .A(n123), .Q(n48) );
  INV3 U34 ( .A(n88), .Q(n41) );
  INV3 U35 ( .A(n83), .Q(n40) );
  INV3 U36 ( .A(n77), .Q(n39) );
  INV3 U37 ( .A(n62), .Q(n45) );
  INV3 U38 ( .A(n54), .Q(n44) );
  INV3 U39 ( .A(n6), .Q(n5) );
  INV3 U40 ( .A(n53), .Q(n1) );
  NOR21 U41 ( .A(n50), .B(n11), .Q(n53) );
  INV3 U42 ( .A(n170), .Q(n18) );
  INV3 U43 ( .A(n120), .Q(n30) );
  INV3 U44 ( .A(n55), .Q(n14) );
  INV3 U45 ( .A(n72), .Q(n42) );
  INV3 U46 ( .A(n179), .Q(n22) );
  INV3 U47 ( .A(n117), .Q(n50) );
  INV3 U48 ( .A(n12), .Q(n11) );
  INV3 U49 ( .A(n98), .Q(n6) );
  INV3 U50 ( .A(SH[2]), .Q(n9) );
  INV3 U51 ( .A(SH[1]), .Q(n8) );
  INV3 U52 ( .A(SH[0]), .Q(n7) );
  INV3 U53 ( .A(SH[3]), .Q(n10) );
  NOR21 U54 ( .A(SH[2]), .B(SH[3]), .Q(n117) );
  INV3 U55 ( .A(SH[4]), .Q(n12) );
  NOR21 U56 ( .A(n207), .B(SH[2]), .Q(n56) );
  OAI2110 U57 ( .A(n40), .B(n46), .C(n51), .D(n52), .Q(B[9]) );
  AOI220 U58 ( .A(n53), .B(n54), .C(n11), .D(n14), .Q(n52) );
  AOI220 U59 ( .A(n56), .B(n57), .C(n58), .D(n59), .Q(n51) );
  OAI2110 U60 ( .A(n41), .B(n46), .C(n60), .D(n61), .Q(B[8]) );
  AOI220 U61 ( .A(n53), .B(n62), .C(n11), .D(n63), .Q(n61) );
  AOI220 U62 ( .A(n56), .B(n64), .C(n58), .D(n65), .Q(n60) );
  OAI2110 U63 ( .A(n42), .B(n46), .C(n66), .D(n67), .Q(B[7]) );
  AOI220 U64 ( .A(n53), .B(n68), .C(n11), .D(n69), .Q(n67) );
  AOI220 U65 ( .A(n56), .B(n70), .C(n58), .D(n71), .Q(n66) );
  OAI2110 U66 ( .A(n43), .B(n46), .C(n73), .D(n74), .Q(B[6]) );
  AOI220 U67 ( .A(n53), .B(n75), .C(n11), .D(n25), .Q(n74) );
  AOI220 U68 ( .A(n56), .B(n77), .C(n58), .D(n78), .Q(n73) );
  OAI2110 U69 ( .A(n44), .B(n46), .C(n79), .D(n80), .Q(B[5]) );
  AOI220 U70 ( .A(n53), .B(n81), .C(n11), .D(n16), .Q(n80) );
  AOI220 U71 ( .A(n56), .B(n83), .C(n58), .D(n57), .Q(n79) );
  OAI2110 U72 ( .A(n45), .B(n46), .C(n84), .D(n85), .Q(B[4]) );
  AOI220 U73 ( .A(n53), .B(n86), .C(n11), .D(n27), .Q(n85) );
  AOI220 U74 ( .A(n56), .B(n88), .C(n58), .D(n64), .Q(n84) );
  OAI2110 U75 ( .A(n37), .B(n47), .C(n89), .D(n90), .Q(B[3]) );
  AOI220 U76 ( .A(n91), .B(n68), .C(n11), .D(n92), .Q(n90) );
  NAND20 U77 ( .A(n93), .B(n94), .Q(n68) );
  AOI220 U78 ( .A(A[10]), .B(n2), .C(A[9]), .D(n3), .Q(n94) );
  AOI220 U79 ( .A(A[8]), .B(n4), .C(A[7]), .D(n5), .Q(n93) );
  AOI220 U80 ( .A(n53), .B(n99), .C(n56), .D(n72), .Q(n89) );
  NAND20 U81 ( .A(n100), .B(n101), .Q(n99) );
  AOI220 U82 ( .A(A[6]), .B(n2), .C(A[5]), .D(n3), .Q(n101) );
  AOI220 U83 ( .A(A[4]), .B(n4), .C(A[3]), .D(n5), .Q(n100) );
  NOR20 U84 ( .A(n1), .B(n102), .Q(B[31]) );
  NOR20 U85 ( .A(n103), .B(n1), .Q(B[30]) );
  OAI2110 U86 ( .A(n39), .B(n47), .C(n104), .D(n105), .Q(B[2]) );
  AOI220 U87 ( .A(n91), .B(n75), .C(n11), .D(n106), .Q(n105) );
  NAND20 U88 ( .A(n107), .B(n108), .Q(n75) );
  AOI220 U89 ( .A(A[9]), .B(n95), .C(A[8]), .D(n96), .Q(n108) );
  AOI220 U90 ( .A(A[7]), .B(n4), .C(A[6]), .D(n5), .Q(n107) );
  AOI220 U91 ( .A(n53), .B(n109), .C(n56), .D(n110), .Q(n104) );
  NAND20 U92 ( .A(n111), .B(n112), .Q(n109) );
  AOI220 U93 ( .A(A[5]), .B(n2), .C(A[4]), .D(n3), .Q(n112) );
  AOI220 U94 ( .A(A[3]), .B(n4), .C(A[2]), .D(n5), .Q(n111) );
  NOR20 U95 ( .A(n113), .B(n1), .Q(B[29]) );
  NOR20 U96 ( .A(n29), .B(n1), .Q(B[28]) );
  NOR30 U97 ( .A(n114), .B(n11), .C(SH[3]), .Q(B[27]) );
  NOR20 U98 ( .A(n11), .B(n115), .Q(B[26]) );
  NOR20 U99 ( .A(n11), .B(n55), .Q(B[25]) );
  AOI220 U100 ( .A(n116), .B(n117), .C(n15), .D(n118), .Q(n55) );
  NOR20 U101 ( .A(n11), .B(n28), .Q(B[24]) );
  OAI220 U102 ( .A(n33), .B(n50), .C(n29), .D(n49), .Q(n63) );
  NOR20 U103 ( .A(n11), .B(n20), .Q(B[23]) );
  OAI210 U104 ( .A(n34), .B(n50), .C(n119), .Q(n69) );
  AOI220 U105 ( .A(n48), .B(n21), .C(n118), .D(n120), .Q(n119) );
  NOR20 U106 ( .A(n11), .B(n76), .Q(B[22]) );
  AOI210 U107 ( .A(n121), .B(n117), .C(n122), .Q(n76) );
  OAI220 U108 ( .A(n123), .B(n103), .C(n49), .D(n31), .Q(n122) );
  NOR20 U109 ( .A(n11), .B(n82), .Q(B[21]) );
  AOI210 U110 ( .A(n59), .B(n117), .C(n124), .Q(n82) );
  OAI220 U111 ( .A(n123), .B(n113), .C(n49), .D(n32), .Q(n124) );
  NOR20 U112 ( .A(n11), .B(n87), .Q(B[20]) );
  AOI210 U113 ( .A(n65), .B(n117), .C(n125), .Q(n87) );
  OAI220 U114 ( .A(n123), .B(n29), .C(n49), .D(n33), .Q(n125) );
  OAI2110 U115 ( .A(n40), .B(n47), .C(n127), .D(n128), .Q(B[1]) );
  AOI220 U116 ( .A(n91), .B(n81), .C(n11), .D(n129), .Q(n128) );
  NAND20 U117 ( .A(n130), .B(n131), .Q(n81) );
  AOI220 U118 ( .A(A[8]), .B(n2), .C(A[7]), .D(n96), .Q(n131) );
  AOI220 U119 ( .A(A[6]), .B(n4), .C(A[5]), .D(n5), .Q(n130) );
  AOI220 U120 ( .A(n53), .B(n132), .C(n56), .D(n54), .Q(n127) );
  NAND20 U121 ( .A(n133), .B(n134), .Q(n54) );
  AOI220 U122 ( .A(A[12]), .B(n2), .C(A[11]), .D(n3), .Q(n134) );
  AOI220 U123 ( .A(A[10]), .B(n4), .C(A[9]), .D(n5), .Q(n133) );
  NAND20 U124 ( .A(n135), .B(n136), .Q(n132) );
  AOI220 U125 ( .A(A[4]), .B(n2), .C(A[3]), .D(n96), .Q(n136) );
  AOI220 U126 ( .A(A[2]), .B(n4), .C(A[1]), .D(n5), .Q(n135) );
  NOR20 U127 ( .A(n11), .B(n19), .Q(B[19]) );
  OAI210 U128 ( .A(n114), .B(n10), .C(n137), .Q(n92) );
  AOI220 U129 ( .A(n118), .B(n138), .C(n117), .D(n71), .Q(n137) );
  NOR20 U130 ( .A(n11), .B(n23), .Q(B[18]) );
  OAI2110 U131 ( .A(n35), .B(n50), .C(n139), .D(n140), .Q(n106) );
  AOI220 U132 ( .A(n141), .B(n24), .C(n48), .D(n142), .Q(n140) );
  NAND20 U133 ( .A(n118), .B(n121), .Q(n139) );
  NOR20 U134 ( .A(n11), .B(n13), .Q(B[17]) );
  NAND20 U135 ( .A(n143), .B(n144), .Q(n129) );
  AOI220 U136 ( .A(n141), .B(n15), .C(n48), .D(n116), .Q(n144) );
  AOI220 U137 ( .A(n118), .B(n59), .C(n117), .D(n57), .Q(n143) );
  NOR20 U138 ( .A(n11), .B(n26), .Q(B[16]) );
  OAI2110 U139 ( .A(n30), .B(n47), .C(n146), .D(n147), .Q(B[15]) );
  AOI220 U140 ( .A(n91), .B(n71), .C(n53), .D(n70), .Q(n147) );
  AOI220 U141 ( .A(n148), .B(n21), .C(n56), .D(n138), .Q(n146) );
  OAI2110 U142 ( .A(n31), .B(n47), .C(n149), .D(n150), .Q(B[14]) );
  AOI220 U143 ( .A(n91), .B(n78), .C(n53), .D(n77), .Q(n150) );
  AOI220 U144 ( .A(n148), .B(n24), .C(n56), .D(n121), .Q(n149) );
  OAI2110 U145 ( .A(n32), .B(n47), .C(n151), .D(n152), .Q(B[13]) );
  AOI220 U146 ( .A(n91), .B(n57), .C(n53), .D(n83), .Q(n152) );
  NAND20 U147 ( .A(n153), .B(n154), .Q(n83) );
  AOI220 U148 ( .A(A[16]), .B(n95), .C(A[15]), .D(n3), .Q(n154) );
  AOI220 U149 ( .A(A[14]), .B(n97), .C(A[13]), .D(n5), .Q(n153) );
  NAND20 U150 ( .A(n155), .B(n156), .Q(n57) );
  AOI220 U151 ( .A(A[20]), .B(n2), .C(A[19]), .D(n3), .Q(n156) );
  AOI220 U152 ( .A(A[18]), .B(n97), .C(A[17]), .D(n5), .Q(n155) );
  AOI220 U153 ( .A(n148), .B(n15), .C(n56), .D(n59), .Q(n151) );
  NAND20 U154 ( .A(n157), .B(n158), .Q(n59) );
  AOI220 U155 ( .A(A[24]), .B(n95), .C(A[23]), .D(n3), .Q(n158) );
  AOI220 U156 ( .A(A[22]), .B(n97), .C(A[21]), .D(n5), .Q(n157) );
  AOI210 U157 ( .A(n98), .B(A[29]), .C(n17), .Q(n113) );
  AOI220 U158 ( .A(A[31]), .B(n3), .C(A[30]), .D(n97), .Q(n159) );
  NAND20 U159 ( .A(n160), .B(n161), .Q(n116) );
  AOI220 U160 ( .A(A[28]), .B(n2), .C(A[27]), .D(n3), .Q(n161) );
  AOI220 U161 ( .A(A[26]), .B(n4), .C(A[25]), .D(n5), .Q(n160) );
  OAI2110 U162 ( .A(n33), .B(n47), .C(n162), .D(n163), .Q(B[12]) );
  AOI220 U163 ( .A(n91), .B(n64), .C(n53), .D(n88), .Q(n163) );
  AOI220 U164 ( .A(n148), .B(n126), .C(n56), .D(n65), .Q(n162) );
  NOR20 U165 ( .A(n12), .B(n50), .Q(n148) );
  OAI2110 U166 ( .A(n34), .B(n47), .C(n18), .D(n165), .Q(B[11]) );
  AOI220 U167 ( .A(n91), .B(n70), .C(n53), .D(n72), .Q(n165) );
  NAND20 U168 ( .A(n166), .B(n167), .Q(n72) );
  AOI220 U169 ( .A(A[14]), .B(n95), .C(A[13]), .D(n3), .Q(n167) );
  AOI220 U170 ( .A(A[12]), .B(n97), .C(A[11]), .D(n5), .Q(n166) );
  NAND20 U171 ( .A(n168), .B(n169), .Q(n70) );
  AOI220 U172 ( .A(A[18]), .B(n95), .C(A[17]), .D(n3), .Q(n169) );
  AOI220 U173 ( .A(A[16]), .B(n97), .C(A[15]), .D(n98), .Q(n168) );
  OAI310 U174 ( .A(n114), .B(SH[3]), .C(n12), .D(n171), .Q(n170) );
  NAND20 U175 ( .A(n71), .B(n56), .Q(n171) );
  OAI2110 U176 ( .A(n36), .B(n6), .C(n172), .D(n173), .Q(n71) );
  AOI220 U177 ( .A(A[22]), .B(n2), .C(A[21]), .D(n3), .Q(n173) );
  NAND20 U178 ( .A(n4), .B(A[20]), .Q(n172) );
  IMUX20 U179 ( .A(n21), .B(n120), .S(n9), .Q(n114) );
  NAND20 U180 ( .A(n174), .B(n175), .Q(n120) );
  AOI220 U181 ( .A(A[30]), .B(n2), .C(A[29]), .D(n3), .Q(n175) );
  AOI220 U182 ( .A(A[28]), .B(n4), .C(A[27]), .D(n5), .Q(n174) );
  NAND20 U183 ( .A(A[31]), .B(n98), .Q(n102) );
  NAND20 U184 ( .A(n176), .B(n177), .Q(n138) );
  AOI220 U185 ( .A(A[26]), .B(n2), .C(A[25]), .D(n3), .Q(n177) );
  AOI220 U186 ( .A(A[24]), .B(n4), .C(A[23]), .D(n5), .Q(n176) );
  OAI2110 U187 ( .A(n39), .B(n46), .C(n178), .D(n22), .Q(B[10]) );
  OAI220 U188 ( .A(n1), .B(n43), .C(n12), .D(n115), .Q(n179) );
  AOI220 U189 ( .A(n142), .B(n117), .C(n24), .D(n118), .Q(n115) );
  AOI220 U190 ( .A(n5), .B(A[30]), .C(n4), .D(A[31]), .Q(n103) );
  NAND20 U191 ( .A(n180), .B(n181), .Q(n142) );
  AOI220 U192 ( .A(A[29]), .B(n2), .C(A[28]), .D(n3), .Q(n181) );
  AOI220 U193 ( .A(A[27]), .B(n4), .C(A[26]), .D(n98), .Q(n180) );
  NAND20 U194 ( .A(n182), .B(n183), .Q(n110) );
  AOI220 U195 ( .A(A[13]), .B(n95), .C(A[12]), .D(n3), .Q(n183) );
  AOI220 U196 ( .A(A[11]), .B(n4), .C(A[10]), .D(n5), .Q(n182) );
  AOI220 U197 ( .A(n56), .B(n78), .C(n58), .D(n121), .Q(n178) );
  NAND20 U198 ( .A(n184), .B(n185), .Q(n121) );
  AOI220 U199 ( .A(A[25]), .B(n2), .C(A[24]), .D(n3), .Q(n185) );
  AOI220 U200 ( .A(A[23]), .B(n4), .C(A[22]), .D(n98), .Q(n184) );
  OAI2110 U201 ( .A(n38), .B(n6), .C(n186), .D(n187), .Q(n78) );
  AOI220 U202 ( .A(A[21]), .B(n95), .C(n3), .D(A[20]), .Q(n187) );
  NAND20 U203 ( .A(n97), .B(A[19]), .Q(n186) );
  NAND20 U204 ( .A(n188), .B(n189), .Q(n77) );
  AOI220 U205 ( .A(A[17]), .B(n95), .C(A[16]), .D(n96), .Q(n189) );
  AOI220 U206 ( .A(A[15]), .B(n4), .C(A[14]), .D(n5), .Q(n188) );
  OAI2110 U207 ( .A(n41), .B(n47), .C(n190), .D(n191), .Q(B[0]) );
  AOI220 U208 ( .A(n91), .B(n86), .C(n11), .D(n145), .Q(n191) );
  NAND20 U209 ( .A(n192), .B(n193), .Q(n145) );
  AOI220 U210 ( .A(n141), .B(n126), .C(n48), .D(n164), .Q(n193) );
  NAND20 U211 ( .A(n194), .B(n195), .Q(n164) );
  AOI220 U212 ( .A(A[27]), .B(n95), .C(A[26]), .D(n96), .Q(n195) );
  AOI220 U213 ( .A(A[25]), .B(n4), .C(A[24]), .D(n5), .Q(n194) );
  NAND20 U214 ( .A(SH[3]), .B(n9), .Q(n123) );
  NAND20 U215 ( .A(n196), .B(n197), .Q(n126) );
  AOI220 U216 ( .A(A[31]), .B(n2), .C(A[30]), .D(n96), .Q(n197) );
  AOI220 U217 ( .A(A[29]), .B(n97), .C(A[28]), .D(n98), .Q(n196) );
  NOR20 U218 ( .A(n9), .B(n10), .Q(n141) );
  AOI220 U219 ( .A(n118), .B(n65), .C(n117), .D(n64), .Q(n192) );
  NAND20 U220 ( .A(n198), .B(n199), .Q(n64) );
  AOI220 U221 ( .A(A[19]), .B(n2), .C(A[18]), .D(n3), .Q(n199) );
  AOI220 U222 ( .A(A[17]), .B(n97), .C(A[16]), .D(n5), .Q(n198) );
  NAND20 U223 ( .A(n200), .B(n201), .Q(n65) );
  AOI220 U224 ( .A(A[23]), .B(n2), .C(A[22]), .D(n3), .Q(n201) );
  AOI220 U225 ( .A(A[21]), .B(n4), .C(n98), .D(A[20]), .Q(n200) );
  NAND20 U226 ( .A(n202), .B(n203), .Q(n86) );
  AOI220 U227 ( .A(A[7]), .B(n2), .C(A[6]), .D(n96), .Q(n203) );
  AOI220 U228 ( .A(A[5]), .B(n4), .C(A[4]), .D(n5), .Q(n202) );
  NOR20 U229 ( .A(n9), .B(SH[3]), .Q(n118) );
  AOI220 U230 ( .A(n53), .B(n204), .C(n56), .D(n62), .Q(n190) );
  NAND20 U231 ( .A(n205), .B(n206), .Q(n62) );
  AOI220 U232 ( .A(A[11]), .B(n2), .C(A[10]), .D(n96), .Q(n206) );
  AOI220 U233 ( .A(A[9]), .B(n4), .C(A[8]), .D(n98), .Q(n205) );
  NAND20 U234 ( .A(n208), .B(n209), .Q(n204) );
  AOI220 U235 ( .A(A[3]), .B(n2), .C(A[2]), .D(n96), .Q(n209) );
  AOI220 U236 ( .A(A[1]), .B(n4), .C(A[0]), .D(n5), .Q(n208) );
  NOR20 U237 ( .A(n9), .B(n207), .Q(n58) );
  NAND20 U238 ( .A(SH[3]), .B(n12), .Q(n207) );
  NAND20 U239 ( .A(n210), .B(n211), .Q(n88) );
  AOI220 U240 ( .A(A[15]), .B(n2), .C(A[14]), .D(n3), .Q(n211) );
  NOR20 U241 ( .A(n8), .B(SH[0]), .Q(n96) );
  NOR20 U242 ( .A(n8), .B(n7), .Q(n95) );
  AOI220 U243 ( .A(A[13]), .B(n4), .C(A[12]), .D(n5), .Q(n210) );
  NOR20 U244 ( .A(SH[0]), .B(SH[1]), .Q(n98) );
  NOR20 U245 ( .A(n7), .B(SH[1]), .Q(n97) );
endmodule


module E_alu_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151;

  INV2 U1 ( .A(A[5]), .Q(n89) );
  NAND20 U2 ( .A(A[2]), .B(n119), .Q(n111) );
  INV0 U3 ( .A(A[2]), .Q(n101) );
  AOI220 U4 ( .A(B[22]), .B(n37), .C(B[21]), .D(n51), .Q(n32) );
  INV0 U5 ( .A(A[19]), .Q(n34) );
  NOR20 U6 ( .A(B[16]), .B(n47), .Q(n45) );
  INV0 U7 ( .A(B[16]), .Q(n67) );
  INV0 U8 ( .A(B[9]), .Q(n96) );
  INV0 U9 ( .A(B[8]), .Q(n95) );
  AOI2110 U10 ( .A(n71), .B(B[8]), .C(n72), .D(n73), .Q(n70) );
  INV0 U11 ( .A(B[0]), .Q(n108) );
  NOR20 U12 ( .A(B[0]), .B(n110), .Q(n109) );
  INV0 U13 ( .A(B[1]), .Q(n107) );
  NAND20 U14 ( .A(B[9]), .B(n77), .Q(n74) );
  NAND30 U15 ( .A(n102), .B(n117), .C(B[1]), .Q(n112) );
  INV3 U16 ( .A(A[23]), .Q(n143) );
  NAND41 U17 ( .A(n120), .B(n121), .C(n122), .D(n123), .Q(n56) );
  NAND22 U18 ( .A(A[12]), .B(n135), .Q(n121) );
  NAND22 U19 ( .A(A[13]), .B(n136), .Q(n120) );
  INV3 U20 ( .A(n63), .Q(n122) );
  NAND41 U21 ( .A(n137), .B(n138), .C(n26), .D(n139), .Q(n17) );
  NAND22 U22 ( .A(A[24]), .B(n151), .Q(n138) );
  NAND22 U23 ( .A(A[25]), .B(n27), .Q(n137) );
  AOI311 U24 ( .A(n34), .B(n35), .C(B[19]), .D(n36), .Q(n33) );
  AOI221 U25 ( .A(n140), .B(n141), .C(n142), .D(n141), .Q(n139) );
  NOR21 U26 ( .A(B[22]), .B(n37), .Q(n140) );
  NOR21 U27 ( .A(B[23]), .B(n143), .Q(n142) );
  AOI211 U28 ( .A(n28), .B(n29), .C(n30), .Q(n18) );
  NOR21 U29 ( .A(n38), .B(n39), .Q(n29) );
  NAND31 U30 ( .A(n31), .B(n32), .C(n33), .Q(n30) );
  OAI2111 U31 ( .A(n56), .B(n57), .C(n58), .D(n59), .Q(n28) );
  NAND31 U32 ( .A(n13), .B(n14), .C(n15), .Q(n1) );
  NAND22 U33 ( .A(A[28]), .B(n16), .Q(n15) );
  NAND22 U34 ( .A(A[29]), .B(n10), .Q(n14) );
  OAI2111 U35 ( .A(n17), .B(n18), .C(n19), .D(n20), .Q(n13) );
  AOI211 U36 ( .A(n1), .B(n2), .C(n3), .Q(LT_LE) );
  AOI2111 U37 ( .A(B[30]), .B(n8), .C(n11), .D(n9), .Q(n2) );
  NAND22 U38 ( .A(n144), .B(n145), .Q(n36) );
  NAND22 U39 ( .A(B[24]), .B(n146), .Q(n144) );
  NAND22 U40 ( .A(B[23]), .B(n143), .Q(n145) );
  INV3 U41 ( .A(A[24]), .Q(n146) );
  NAND22 U42 ( .A(n131), .B(n132), .Q(n63) );
  NAND22 U43 ( .A(A[15]), .B(n134), .Q(n131) );
  NAND22 U44 ( .A(A[14]), .B(n133), .Q(n132) );
  INV3 U45 ( .A(B[15]), .Q(n134) );
  INV3 U46 ( .A(A[11]), .Q(n127) );
  NOR21 U47 ( .A(A[8]), .B(n81), .Q(n71) );
  AOI2111 U48 ( .A(n21), .B(B[26]), .C(n22), .D(n23), .Q(n20) );
  NOR21 U49 ( .A(A[27]), .B(n150), .Q(n23) );
  NOR21 U50 ( .A(A[28]), .B(n16), .Q(n22) );
  NOR21 U51 ( .A(A[26]), .B(n24), .Q(n21) );
  NOR21 U52 ( .A(n49), .B(n50), .Q(n35) );
  NOR21 U53 ( .A(B[21]), .B(n51), .Q(n50) );
  NOR21 U54 ( .A(B[20]), .B(n52), .Q(n49) );
  INV3 U55 ( .A(A[21]), .Q(n51) );
  NAND31 U56 ( .A(n35), .B(n52), .C(B[20]), .Q(n31) );
  NAND31 U57 ( .A(A[30]), .B(n6), .C(n7), .Q(n5) );
  INV3 U58 ( .A(B[30]), .Q(n6) );
  XNR21 U59 ( .A(B[31]), .B(A[31]), .Q(n4) );
  NAND22 U60 ( .A(n48), .B(n35), .Q(n38) );
  NOR21 U61 ( .A(n53), .B(n54), .Q(n48) );
  NOR21 U62 ( .A(B[19]), .B(n34), .Q(n54) );
  NOR21 U63 ( .A(B[18]), .B(n55), .Q(n53) );
  NAND22 U64 ( .A(n40), .B(n41), .Q(n39) );
  NAND22 U65 ( .A(n45), .B(n43), .Q(n40) );
  NAND22 U66 ( .A(n42), .B(n43), .Q(n41) );
  NAND22 U67 ( .A(n61), .B(n62), .Q(n46) );
  NAND22 U68 ( .A(B[18]), .B(n55), .Q(n61) );
  NAND22 U69 ( .A(B[17]), .B(n44), .Q(n62) );
  NAND22 U70 ( .A(n147), .B(n148), .Q(n24) );
  NAND22 U71 ( .A(A[27]), .B(n150), .Q(n147) );
  NAND22 U72 ( .A(A[26]), .B(n149), .Q(n148) );
  INV3 U73 ( .A(B[27]), .Q(n150) );
  INV3 U74 ( .A(A[17]), .Q(n44) );
  INV3 U75 ( .A(A[18]), .Q(n55) );
  INV3 U76 ( .A(A[10]), .Q(n76) );
  INV3 U77 ( .A(B[25]), .Q(n27) );
  INV3 U78 ( .A(B[29]), .Q(n10) );
  INV3 U79 ( .A(A[22]), .Q(n37) );
  INV3 U80 ( .A(n11), .Q(n7) );
  NOR21 U81 ( .A(A[31]), .B(n12), .Q(n11) );
  INV3 U82 ( .A(B[31]), .Q(n12) );
  NAND22 U83 ( .A(n25), .B(n26), .Q(n19) );
  NOR21 U84 ( .A(A[25]), .B(n27), .Q(n25) );
  NOR21 U85 ( .A(A[29]), .B(n10), .Q(n9) );
  NOR21 U86 ( .A(B[17]), .B(n44), .Q(n42) );
  INV3 U87 ( .A(A[16]), .Q(n47) );
  INV3 U88 ( .A(A[20]), .Q(n52) );
  INV3 U89 ( .A(B[24]), .Q(n151) );
  INV3 U90 ( .A(B[28]), .Q(n16) );
  INV3 U91 ( .A(B[26]), .Q(n149) );
  INV3 U92 ( .A(A[30]), .Q(n8) );
  AOI2111 U93 ( .A(A[7]), .B(n91), .C(n81), .D(n92), .Q(n84) );
  INV3 U94 ( .A(B[7]), .Q(n91) );
  NOR21 U95 ( .A(B[6]), .B(n116), .Q(n92) );
  NAND22 U96 ( .A(A[3]), .B(n104), .Q(n102) );
  OAI2111 U97 ( .A(n97), .B(n98), .C(n99), .D(n100), .Q(n83) );
  NAND22 U98 ( .A(n110), .B(n111), .Q(n97) );
  AOI211 U99 ( .A(B[4]), .B(n90), .C(n103), .Q(n99) );
  NAND31 U100 ( .A(n105), .B(n106), .C(n102), .Q(n98) );
  NOR21 U101 ( .A(A[3]), .B(n104), .Q(n103) );
  INV3 U102 ( .A(n68), .Q(n57) );
  NAND22 U103 ( .A(n69), .B(n70), .Q(n68) );
  OAI2111 U104 ( .A(n82), .B(n83), .C(n84), .D(n85), .Q(n69) );
  NAND31 U105 ( .A(B[2]), .B(n101), .C(n102), .Q(n100) );
  AOI2111 U106 ( .A(n64), .B(B[14]), .C(n65), .D(n66), .Q(n58) );
  NOR21 U107 ( .A(A[16]), .B(n67), .Q(n65) );
  NOR21 U108 ( .A(A[15]), .B(n134), .Q(n66) );
  NOR21 U109 ( .A(A[14]), .B(n63), .Q(n64) );
  AOI211 U110 ( .A(n60), .B(B[13]), .C(n46), .Q(n59) );
  NOR21 U111 ( .A(A[13]), .B(n63), .Q(n60) );
  AOI221 U112 ( .A(n124), .B(n125), .C(n126), .D(n125), .Q(n123) );
  NOR21 U113 ( .A(B[10]), .B(n76), .Q(n124) );
  NOR21 U114 ( .A(B[11]), .B(n127), .Q(n126) );
  NAND22 U115 ( .A(n128), .B(n129), .Q(n79) );
  NAND22 U116 ( .A(B[12]), .B(n130), .Q(n128) );
  NAND22 U117 ( .A(B[11]), .B(n127), .Q(n129) );
  INV3 U118 ( .A(A[12]), .Q(n130) );
  INV3 U119 ( .A(B[3]), .Q(n104) );
  NAND22 U120 ( .A(n114), .B(n115), .Q(n88) );
  NAND22 U121 ( .A(B[6]), .B(n116), .Q(n114) );
  NAND22 U122 ( .A(B[5]), .B(n89), .Q(n115) );
  INV3 U123 ( .A(A[6]), .Q(n116) );
  NAND22 U124 ( .A(n93), .B(n94), .Q(n81) );
  NAND22 U125 ( .A(A[9]), .B(n96), .Q(n93) );
  NAND22 U126 ( .A(A[8]), .B(n95), .Q(n94) );
  NAND22 U127 ( .A(n78), .B(n125), .Q(n72) );
  NAND22 U128 ( .A(n80), .B(B[7]), .Q(n78) );
  NOR21 U129 ( .A(A[7]), .B(n81), .Q(n80) );
  INV3 U130 ( .A(B[14]), .Q(n133) );
  NOR21 U131 ( .A(n86), .B(n87), .Q(n85) );
  NOR31 U132 ( .A(n88), .B(B[5]), .C(n89), .Q(n87) );
  NOR31 U133 ( .A(n88), .B(B[4]), .C(n90), .Q(n86) );
  INV3 U134 ( .A(A[4]), .Q(n90) );
  NAND22 U135 ( .A(n112), .B(n113), .Q(n82) );
  INV3 U136 ( .A(n88), .Q(n113) );
  NOR21 U137 ( .A(A[1]), .B(n118), .Q(n117) );
  INV3 U138 ( .A(B[2]), .Q(n119) );
  NOR21 U139 ( .A(n108), .B(n109), .Q(n105) );
  INV3 U140 ( .A(A[0]), .Q(n110) );
  INV3 U141 ( .A(B[12]), .Q(n135) );
  INV3 U142 ( .A(B[13]), .Q(n136) );
  NAND22 U143 ( .A(n74), .B(n75), .Q(n73) );
  NAND22 U144 ( .A(B[10]), .B(n76), .Q(n75) );
  INV3 U145 ( .A(A[9]), .Q(n77) );
  NAND22 U146 ( .A(A[1]), .B(n107), .Q(n106) );
  OAI212 U147 ( .A(n4), .B(n11), .C(n5), .Q(n3) );
  CLKIN3 U148 ( .A(n24), .Q(n26) );
  CLKIN3 U149 ( .A(n46), .Q(n43) );
  CLKIN3 U150 ( .A(n111), .Q(n118) );
  CLKIN3 U151 ( .A(n79), .Q(n125) );
  CLKIN3 U152 ( .A(n36), .Q(n141) );
endmodule


module E_alu_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [16:0] A;
  input [16:0] B;
  output [16:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154;

  CLKIN3 U3 ( .A(A[2]), .Q(n136) );
  NAND20 U4 ( .A(A[2]), .B(n129), .Q(n39) );
  NAND22 U5 ( .A(n93), .B(n101), .Q(n110) );
  NAND22 U6 ( .A(n63), .B(n66), .Q(n75) );
  NAND20 U7 ( .A(B[1]), .B(n137), .Q(n45) );
  NAND20 U8 ( .A(B[9]), .B(n113), .Q(n3) );
  INV0 U9 ( .A(B[8]), .Q(n10) );
  INV0 U10 ( .A(B[1]), .Q(n132) );
  INV0 U11 ( .A(B[0]), .Q(n50) );
  INV0 U12 ( .A(B[9]), .Q(n112) );
  XOR20 U13 ( .A(B[8]), .B(A[8]), .Q(n5) );
  XOR21 U14 ( .A(n46), .B(n47), .Q(DIFF[1]) );
  NAND22 U15 ( .A(n45), .B(n42), .Q(n46) );
  IMUX21 U16 ( .A(n29), .B(n30), .S(n25), .Q(DIFF[4]) );
  NOR21 U17 ( .A(n32), .B(n33), .Q(n29) );
  XOR21 U18 ( .A(n23), .B(n24), .Q(DIFF[5]) );
  NAND22 U19 ( .A(n22), .B(n19), .Q(n23) );
  AOI2111 U20 ( .A(n51), .B(n52), .C(n53), .D(n54), .Q(DIFF[16]) );
  NOR21 U21 ( .A(B[15]), .B(n55), .Q(n54) );
  INV3 U22 ( .A(n70), .Q(n51) );
  XOR21 U23 ( .A(n40), .B(n41), .Q(DIFF[2]) );
  NAND22 U24 ( .A(n37), .B(n39), .Q(n40) );
  XOR21 U25 ( .A(n17), .B(n18), .Q(DIFF[6]) );
  NAND22 U26 ( .A(n14), .B(n16), .Q(n17) );
  XNR21 U27 ( .A(n71), .B(n72), .Q(DIFF[15]) );
  XNR21 U28 ( .A(B[15]), .B(A[15]), .Q(n71) );
  AOI211 U29 ( .A(n73), .B(n63), .C(n74), .Q(n72) );
  AOI211 U30 ( .A(n33), .B(n22), .C(n147), .Q(n145) );
  AOI211 U31 ( .A(n9), .B(n3), .C(n102), .Q(n100) );
  NOR21 U32 ( .A(A[12]), .B(n60), .Q(n82) );
  XNR21 U33 ( .A(n110), .B(n108), .Q(DIFF[10]) );
  XOR21 U34 ( .A(n1), .B(n2), .Q(DIFF[9]) );
  NAND22 U35 ( .A(n3), .B(n4), .Q(n1) );
  XOR21 U36 ( .A(n80), .B(n77), .Q(DIFF[13]) );
  NAND22 U37 ( .A(n62), .B(n69), .Q(n80) );
  XNR21 U38 ( .A(n75), .B(n73), .Q(DIFF[14]) );
  AOI211 U39 ( .A(n130), .B(n45), .C(n131), .Q(n128) );
  NAND22 U40 ( .A(A[8]), .B(n10), .Q(n103) );
  NOR31 U41 ( .A(n56), .B(n57), .C(n58), .Q(n53) );
  NAND22 U42 ( .A(n62), .B(n63), .Q(n56) );
  INV3 U43 ( .A(n61), .Q(n57) );
  NAND22 U44 ( .A(n19), .B(n20), .Q(n13) );
  NAND22 U45 ( .A(n21), .B(n22), .Q(n20) );
  NOR21 U46 ( .A(n135), .B(n127), .Q(n134) );
  NAND22 U47 ( .A(n103), .B(n115), .Q(n114) );
  NAND22 U48 ( .A(n116), .B(n7), .Q(n115) );
  INV3 U49 ( .A(n152), .Q(n116) );
  AOI211 U50 ( .A(n36), .B(n37), .C(n38), .Q(n35) );
  AOI211 U51 ( .A(n67), .B(n62), .C(n68), .Q(n65) );
  INV3 U52 ( .A(n69), .Q(n68) );
  NAND22 U53 ( .A(A[12]), .B(n60), .Q(n83) );
  NAND22 U54 ( .A(n42), .B(n43), .Q(n36) );
  NAND22 U55 ( .A(n44), .B(n45), .Q(n43) );
  NOR21 U56 ( .A(A[8]), .B(n10), .Q(n152) );
  NOR21 U57 ( .A(n91), .B(n92), .Q(n90) );
  NAND22 U58 ( .A(n3), .B(n93), .Q(n92) );
  NOR21 U59 ( .A(A[15]), .B(n59), .Q(n70) );
  INV3 U60 ( .A(B[15]), .Q(n59) );
  INV3 U61 ( .A(A[11]), .Q(n98) );
  INV3 U62 ( .A(n104), .Q(n95) );
  NOR21 U63 ( .A(A[11]), .B(n94), .Q(n104) );
  INV3 U64 ( .A(A[15]), .Q(n55) );
  NAND22 U65 ( .A(n123), .B(n124), .Q(n31) );
  AOI221 U66 ( .A(A[3]), .B(n125), .C(n133), .D(n134), .Q(n123) );
  NOR21 U67 ( .A(n138), .B(n139), .Q(n133) );
  NOR21 U68 ( .A(A[0]), .B(n50), .Q(n138) );
  NOR21 U69 ( .A(A[4]), .B(n28), .Q(n26) );
  NOR21 U70 ( .A(A[3]), .B(n125), .Q(n139) );
  NAND22 U71 ( .A(A[1]), .B(n132), .Q(n42) );
  NAND22 U72 ( .A(B[6]), .B(n150), .Q(n14) );
  INV3 U73 ( .A(A[6]), .Q(n150) );
  NAND22 U74 ( .A(A[6]), .B(n146), .Q(n16) );
  INV3 U75 ( .A(B[6]), .Q(n146) );
  INV3 U76 ( .A(B[2]), .Q(n129) );
  NAND22 U77 ( .A(A[4]), .B(n28), .Q(n27) );
  XNR21 U78 ( .A(n34), .B(n35), .Q(DIFF[3]) );
  XNR21 U79 ( .A(B[3]), .B(A[3]), .Q(n34) );
  NAND22 U80 ( .A(A[5]), .B(n148), .Q(n19) );
  INV3 U81 ( .A(B[5]), .Q(n148) );
  NAND22 U82 ( .A(A[0]), .B(n50), .Q(n48) );
  INV3 U83 ( .A(A[7]), .Q(n143) );
  INV3 U84 ( .A(B[4]), .Q(n28) );
  INV3 U85 ( .A(A[1]), .Q(n137) );
  NAND22 U86 ( .A(B[2]), .B(n136), .Q(n37) );
  NAND22 U87 ( .A(B[5]), .B(n149), .Q(n22) );
  INV3 U88 ( .A(A[5]), .Q(n149) );
  NAND22 U89 ( .A(n88), .B(n89), .Q(n61) );
  AOI211 U90 ( .A(n95), .B(n96), .C(n97), .Q(n88) );
  NAND22 U91 ( .A(n7), .B(n90), .Q(n89) );
  NOR21 U92 ( .A(B[11]), .B(n98), .Q(n97) );
  INV3 U93 ( .A(B[3]), .Q(n125) );
  IMUX21 U94 ( .A(n86), .B(n87), .S(n57), .Q(DIFF[12]) );
  XOR21 U95 ( .A(B[12]), .B(A[12]), .Q(n87) );
  NOR21 U96 ( .A(n105), .B(n67), .Q(n86) );
  NOR21 U97 ( .A(A[12]), .B(n60), .Q(n105) );
  INV3 U98 ( .A(B[7]), .Q(n122) );
  XNR21 U99 ( .A(n11), .B(n12), .Q(DIFF[7]) );
  XNR21 U100 ( .A(B[7]), .B(A[7]), .Q(n11) );
  AOI211 U101 ( .A(n13), .B(n14), .C(n15), .Q(n12) );
  XNR21 U102 ( .A(n106), .B(n107), .Q(DIFF[11]) );
  XNR21 U103 ( .A(B[11]), .B(A[11]), .Q(n106) );
  AOI211 U104 ( .A(n108), .B(n93), .C(n109), .Q(n107) );
  NOR21 U105 ( .A(n120), .B(n121), .Q(n119) );
  NAND22 U106 ( .A(n22), .B(n14), .Q(n121) );
  NAND22 U107 ( .A(n117), .B(n118), .Q(n7) );
  AOI211 U108 ( .A(n140), .B(n141), .C(n142), .Q(n117) );
  NAND22 U109 ( .A(n31), .B(n119), .Q(n118) );
  NOR21 U110 ( .A(B[7]), .B(n143), .Q(n142) );
  INV3 U111 ( .A(n151), .Q(n140) );
  NOR21 U112 ( .A(A[7]), .B(n122), .Q(n151) );
  NAND22 U113 ( .A(B[10]), .B(n154), .Q(n93) );
  INV3 U114 ( .A(A[10]), .Q(n154) );
  INV3 U115 ( .A(A[9]), .Q(n113) );
  INV3 U116 ( .A(B[12]), .Q(n60) );
  NAND22 U117 ( .A(A[14]), .B(n78), .Q(n66) );
  INV3 U118 ( .A(B[14]), .Q(n78) );
  NAND22 U119 ( .A(A[9]), .B(n112), .Q(n4) );
  NAND22 U120 ( .A(n48), .B(n49), .Q(n44) );
  NOR21 U121 ( .A(A[0]), .B(n50), .Q(n49) );
  INV3 U122 ( .A(B[11]), .Q(n94) );
  IMUX21 U123 ( .A(n5), .B(n6), .S(n7), .Q(DIFF[8]) );
  NOR21 U124 ( .A(n8), .B(n9), .Q(n6) );
  NOR21 U125 ( .A(A[8]), .B(n10), .Q(n8) );
  NAND22 U126 ( .A(A[10]), .B(n153), .Q(n101) );
  INV3 U127 ( .A(B[10]), .Q(n153) );
  NAND22 U128 ( .A(A[13]), .B(n84), .Q(n69) );
  INV3 U129 ( .A(B[13]), .Q(n84) );
  NAND22 U130 ( .A(B[13]), .B(n85), .Q(n62) );
  INV3 U131 ( .A(A[13]), .Q(n85) );
  NAND22 U132 ( .A(B[14]), .B(n79), .Q(n63) );
  INV3 U133 ( .A(A[14]), .Q(n79) );
  NOR21 U134 ( .A(A[4]), .B(n28), .Q(n32) );
  XOR21 U135 ( .A(B[4]), .B(A[4]), .Q(n30) );
  CLKIN3 U136 ( .A(n16), .Q(n15) );
  CLKIN3 U137 ( .A(n13), .Q(n18) );
  CLKIN3 U138 ( .A(n21), .Q(n24) );
  OAI212 U139 ( .A(n25), .B(n26), .C(n27), .Q(n21) );
  CLKIN3 U140 ( .A(n31), .Q(n25) );
  CLKIN3 U141 ( .A(n39), .Q(n38) );
  CLKIN3 U142 ( .A(n36), .Q(n41) );
  CLKIN3 U143 ( .A(n44), .Q(n47) );
  OAI222 U144 ( .A(A[15]), .B(n59), .C(A[12]), .D(n60), .Q(n58) );
  OAI212 U145 ( .A(n64), .B(n65), .C(n66), .Q(n52) );
  CLKIN3 U146 ( .A(n63), .Q(n64) );
  CLKIN3 U147 ( .A(n66), .Q(n74) );
  OAI212 U148 ( .A(n76), .B(n77), .C(n69), .Q(n73) );
  CLKIN3 U149 ( .A(n62), .Q(n76) );
  CLKIN3 U150 ( .A(n81), .Q(n77) );
  OAI212 U151 ( .A(n57), .B(n82), .C(n83), .Q(n81) );
  OAI222 U152 ( .A(A[8]), .B(n10), .C(A[11]), .D(n94), .Q(n91) );
  OAI212 U153 ( .A(n99), .B(n100), .C(n101), .Q(n96) );
  CLKIN3 U154 ( .A(n4), .Q(n102) );
  CLKIN3 U155 ( .A(n103), .Q(n9) );
  CLKIN3 U156 ( .A(n93), .Q(n99) );
  CLKIN3 U157 ( .A(n83), .Q(n67) );
  CLKIN3 U158 ( .A(n101), .Q(n109) );
  OAI212 U159 ( .A(n2), .B(n111), .C(n4), .Q(n108) );
  CLKIN3 U160 ( .A(n3), .Q(n111) );
  CLKIN3 U161 ( .A(n114), .Q(n2) );
  OAI222 U162 ( .A(A[7]), .B(n122), .C(A[4]), .D(n28), .Q(n120) );
  OAI212 U163 ( .A(A[3]), .B(n125), .C(n126), .Q(n124) );
  OAI212 U164 ( .A(n127), .B(n128), .C(n39), .Q(n126) );
  CLKIN3 U165 ( .A(n42), .Q(n131) );
  CLKIN3 U166 ( .A(n37), .Q(n127) );
  CLKIN3 U167 ( .A(n45), .Q(n135) );
  OAI212 U168 ( .A(n144), .B(n145), .C(n16), .Q(n141) );
  CLKIN3 U169 ( .A(n19), .Q(n147) );
  CLKIN3 U170 ( .A(n27), .Q(n33) );
  CLKIN3 U171 ( .A(n14), .Q(n144) );
  OAI212 U172 ( .A(A[0]), .B(n50), .C(n48), .Q(DIFF[0]) );
  CLKIN3 U173 ( .A(n48), .Q(n130) );
endmodule


module E_alu ( o_data_AluRes, i_data_A, i_data_B, i_con_AluCtrl, i_data_shamt
 );
  output [31:0] o_data_AluRes;
  input [31:0] i_data_A;
  input [31:0] i_data_B;
  input [3:0] i_con_AluCtrl;
  input [4:0] i_data_shamt;
  wire   N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N306, n41, n42,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n426, n428, n429, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n144, n145, n146, n147, n162, n204, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n427;
  wire   [8:0] sum_1;
  wire   [8:0] pre_sum_2a;
  wire   [8:0] pre_sum_2b;
  wire   [8:0] pre_sum_3a;
  wire   [8:0] pre_sum_3b;
  wire   [7:0] pre_sum_4a;
  wire   [7:0] pre_sum_4b;
  wire   [16:0] half_sub;
  wire   [15:0] pre_suba;
  wire   [15:0] pre_subb;

  OAI222 U28 ( .A(n425), .B(n129), .C(n33), .D(n66), .Q(n137) );
  OAI222 U36 ( .A(n64), .B(n131), .C(n32), .D(n66), .Q(n152) );
  OAI222 U46 ( .A(n64), .B(n144), .C(i_data_A[7]), .D(n139), .Q(n159) );
  OAI222 U54 ( .A(n64), .B(n146), .C(i_data_A[6]), .D(n139), .Q(n167) );
  OAI222 U62 ( .A(n425), .B(n162), .C(i_data_A[5]), .D(n139), .Q(n174) );
  OAI222 U70 ( .A(n64), .B(n416), .C(i_data_A[4]), .D(n139), .Q(n181) );
  OAI222 U78 ( .A(n64), .B(n418), .C(i_data_A[3]), .D(n139), .Q(n188) );
  OAI212 U85 ( .A(n101), .B(n63), .C(i_data_B[31]), .Q(n197) );
  OAI212 U87 ( .A(n199), .B(n100), .C(n200), .Q(n195) );
  OAI212 U95 ( .A(n427), .B(n118), .C(n211), .Q(n209) );
  OAI222 U102 ( .A(n425), .B(n102), .C(i_data_A[30]), .D(n139), .Q(n214) );
  OAI222 U107 ( .A(n425), .B(n420), .C(i_data_A[2]), .D(n139), .Q(n219) );
  OAI212 U114 ( .A(n427), .B(n120), .C(n228), .Q(n226) );
  OAI222 U121 ( .A(n64), .B(n103), .C(i_data_A[29]), .D(n139), .Q(n231) );
  OAI212 U125 ( .A(n427), .B(n122), .C(n238), .Q(n236) );
  OAI222 U132 ( .A(n64), .B(n104), .C(n54), .D(n139), .Q(n241) );
  OAI212 U136 ( .A(n427), .B(n124), .C(n248), .Q(n246) );
  OAI222 U143 ( .A(n64), .B(n105), .C(i_data_A[27]), .D(n139), .Q(n251) );
  OAI212 U147 ( .A(n427), .B(n126), .C(n258), .Q(n256) );
  OAI222 U154 ( .A(n425), .B(n106), .C(n52), .D(n139), .Q(n261) );
  OAI212 U158 ( .A(n128), .B(n427), .C(n268), .Q(n266) );
  OAI222 U165 ( .A(n64), .B(n107), .C(n51), .D(n139), .Q(n271) );
  OAI212 U169 ( .A(n130), .B(n427), .C(n278), .Q(n276) );
  OAI222 U179 ( .A(n64), .B(n108), .C(n50), .D(n66), .Q(n282) );
  OAI212 U183 ( .A(n132), .B(n427), .C(n291), .Q(n289) );
  OAI222 U190 ( .A(n64), .B(n109), .C(n49), .D(n66), .Q(n295) );
  OAI212 U194 ( .A(n145), .B(n427), .C(n303), .Q(n301) );
  OAI222 U201 ( .A(n64), .B(n110), .C(n48), .D(n66), .Q(n306) );
  OAI212 U205 ( .A(n147), .B(n427), .C(n313), .Q(n311) );
  OAI222 U212 ( .A(n64), .B(n111), .C(n47), .D(n66), .Q(n316) );
  OAI212 U216 ( .A(n204), .B(n427), .C(n323), .Q(n321) );
  OAI222 U223 ( .A(n64), .B(n112), .C(n46), .D(n66), .Q(n326) );
  OAI222 U228 ( .A(n64), .B(n422), .C(i_data_A[1]), .D(n66), .Q(n331) );
  OAI212 U235 ( .A(n417), .B(n427), .C(n340), .Q(n338) );
  OAI222 U242 ( .A(n425), .B(n113), .C(n45), .D(n66), .Q(n343) );
  OAI212 U246 ( .A(n427), .B(n419), .C(n350), .Q(n348) );
  OAI212 U257 ( .A(n427), .B(n421), .C(n360), .Q(n358) );
  OAI222 U264 ( .A(n64), .B(n115), .C(n43), .D(n66), .Q(n363) );
  OAI212 U268 ( .A(n427), .B(n423), .C(n370), .Q(n368) );
  OAI222 U281 ( .A(n64), .B(n116), .C(n40), .D(n66), .Q(n373) );
  OAI222 U284 ( .A(n64), .B(n117), .C(n39), .D(n66), .Q(n378) );
  OAI222 U292 ( .A(n425), .B(n119), .C(n38), .D(n66), .Q(n385) );
  OAI222 U300 ( .A(n64), .B(n121), .C(i_data_A[13]), .D(n66), .Q(n392) );
  OAI222 U308 ( .A(n425), .B(n123), .C(i_data_A[12]), .D(n66), .Q(n399) );
  OAI222 U316 ( .A(n64), .B(n125), .C(n35), .D(n66), .Q(n406) );
  OAI222 U325 ( .A(n64), .B(n127), .C(n34), .D(n139), .Q(n413) );
  E_alu_DW01_ash_0 sll_56 ( .A({i_data_B[31:25], n25, n23, n21, n19, n17, n15, 
        n13, n11, n4, i_data_B[15:0]}), .DATA_TC(n42), .SH(i_data_shamt), 
        .SH_TC(n42), .B({N224, N223, N222, N221, N220, N219, N218, N217, N216, 
        N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, 
        N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193}) );
  E_alu_DW01_sub_0 sub_1_root_sub_35_2 ( .A({n58, n56, i_data_A[29], n54, 
        i_data_A[27], n52, n51, n50, n49, n48, n47, n46, n45, n44, n43, 
        i_data_A[16]}), .B({i_data_B[31:24], n23, n21, n19, n17, 
        i_data_B[19:16]}), .CI(n41), .DIFF(pre_subb) );
  E_alu_DW01_sub_1 sub_34 ( .A({n58, n56, n55, n54, n53, n52, n51, n50, n49, 
        n48, n47, n46, n45, n44, n43, i_data_A[16]}), .B({i_data_B[31:25], n25, 
        n23, n21, n19, n17, i_data_B[19:16]}), .CI(n42), .DIFF(pre_suba) );
  E_alu_DW01_add_0 add_1_root_add_31_2 ( .A({n57, n56, n55, n54, n53, n52, n51, 
        n50}), .B({i_data_B[31:25], n25}), .CI(n41), .SUM(pre_sum_4b) );
  E_alu_DW01_add_1 add_30 ( .A({n57, n56, n55, i_data_A[28], n53, 
        i_data_A[26:25], n50}), .B({i_data_B[31:25], n25}), .CI(n42), .SUM(
        pre_sum_4a) );
  E_alu_DW01_add_2 add_1_root_add_29_2 ( .A({n42, n49, n48, i_data_A[21], n46, 
        n45, n44, n43, n40}), .B({n42, n23, n21, i_data_B[21], n17, 
        i_data_B[19:18], n11, n4}), .CI(n41), .SUM(pre_sum_3b) );
  E_alu_DW01_add_3 add_28 ( .A({n42, n49, n48, n47, i_data_A[20], n45, n44, 
        n43, n40}), .B({n42, n23, n21, n19, n17, i_data_B[19:18], n11, n4}), 
        .CI(n42), .SUM(pre_sum_3a) );
  E_alu_DW01_add_4 add_1_root_add_27_2 ( .A({n42, n39, n38, n37, i_data_A[12], 
        n35, n34, n33, n32}), .B({n42, n8, i_data_B[14:8]}), .CI(n41), .SUM(
        pre_sum_2b) );
  E_alu_DW01_add_5 add_26 ( .A({n42, n39, i_data_A[14], n37, i_data_A[12], n35, 
        n34, n33, n32}), .B({n42, n8, i_data_B[14:8]}), .CI(n42), .SUM(
        pre_sum_2a) );
  E_alu_DW01_add_6 add_25 ( .A({n42, i_data_A[7:0]}), .B({n42, i_data_B[7:0]}), 
        .CI(n42), .SUM(sum_1) );
  E_alu_DW_rash_0 r130 ( .A({i_data_B[31:25], n25, n23, n21, n19, n17, n15, 
        n13, n11, n4, n8, i_data_B[14:0]}), .DATA_TC(n42), .SH(i_data_shamt), 
        .SH_TC(n42), .B({N256, N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, 
        N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225}) );
  E_alu_DW01_cmp2_1 r131 ( .A({n57, n56, n55, n54, n53, i_data_A[26:25], n50, 
        n49, n48, n47, n46, n45, n44, n43, n40, i_data_A[15], n38, n37, n36, 
        n35, n34, n33, i_data_A[8:0]}), .B({i_data_B[31:24], n23, n21, 
        i_data_B[21:20], n15, n13, n11, n4, i_data_B[15:0]}), .LEQ(n42), .TC(
        n42), .LT_LE(N306) );
  E_alu_DW01_sub_3 sub_33 ( .A({n42, n39, i_data_A[14], n37, n36, n35, n34, 
        i_data_A[9], n32, i_data_A[7:0]}), .B({n42, n8, i_data_B[14:0]}), .CI(
        n42), .DIFF(half_sub) );
  NAND20 U3 ( .A(i_data_A[5]), .B(n59), .Q(n176) );
  AOI2111 U4 ( .A(N222), .B(n91), .C(n226), .D(n227), .Q(n225) );
  NAND20 U5 ( .A(i_data_A[6]), .B(n59), .Q(n169) );
  INV1 U6 ( .A(i_data_B[25]), .Q(n26) );
  NAND31 U7 ( .A(i_con_AluCtrl[0]), .B(n75), .C(n82), .Q(n424) );
  XOR21 U8 ( .A(i_data_B[31]), .B(n58), .Q(n1) );
  NAND42 U9 ( .A(n205), .B(n206), .C(n207), .D(n208), .Q(o_data_AluRes[30]) );
  AOI2111 U10 ( .A(N223), .B(n91), .C(n209), .D(n210), .Q(n208) );
  OAI221 U11 ( .A(n425), .B(n114), .C(n44), .D(n66), .Q(n353) );
  CLKIN3 U12 ( .A(n44), .Q(n114) );
  OAI2110 U13 ( .A(n44), .B(n425), .C(n424), .D(n352), .Q(n351) );
  NAND21 U14 ( .A(n44), .B(n143), .Q(n352) );
  AOI2111 U15 ( .A(pre_sum_4a[7]), .B(n96), .C(n195), .D(n196), .Q(n194) );
  NAND31 U16 ( .A(n193), .B(n191), .C(n192), .Q(n2) );
  NAND22 U17 ( .A(n194), .B(n3), .Q(o_data_AluRes[31]) );
  INV0 U18 ( .A(i_data_B[16]), .Q(n9) );
  INV3 U19 ( .A(n2), .Q(n3) );
  INV1 U20 ( .A(n9), .Q(n4) );
  NAND20 U21 ( .A(pre_sum_4b[6]), .B(n201), .Q(n206) );
  NAND20 U22 ( .A(pre_sum_4b[5]), .B(n201), .Q(n223) );
  AOI220 U23 ( .A(n261), .B(n27), .C(pre_sum_4a[2]), .D(n96), .Q(n252) );
  NAND41 U24 ( .A(n222), .B(n223), .C(n224), .D(n225), .Q(o_data_AluRes[29])
         );
  BUF2 U25 ( .A(i_data_A[18]), .Q(n44) );
  CLKIN1 U26 ( .A(n10), .Q(n11) );
  NAND20 U27 ( .A(n281), .B(n92), .Q(n283) );
  CLKIN3 U29 ( .A(n284), .Q(n97) );
  NAND20 U30 ( .A(pre_sum_4b[4]), .B(n201), .Q(n233) );
  AOI220 U31 ( .A(n4), .B(n371), .C(pre_suba[0]), .D(n61), .Q(n366) );
  NAND20 U32 ( .A(pre_sum_4b[0]), .B(n201), .Q(n273) );
  NAND20 U33 ( .A(pre_sum_4b[1]), .B(n201), .Q(n263) );
  NAND20 U34 ( .A(pre_sum_4b[2]), .B(n201), .Q(n253) );
  NAND20 U35 ( .A(pre_sum_4b[3]), .B(n201), .Q(n243) );
  CLKIN3 U37 ( .A(sum_1[8]), .Q(n98) );
  OAI2110 U38 ( .A(n40), .B(n425), .C(n424), .D(n372), .Q(n371) );
  NAND20 U39 ( .A(n40), .B(n143), .Q(n372) );
  OAI2110 U40 ( .A(n45), .B(n425), .C(n424), .D(n342), .Q(n341) );
  NAND20 U41 ( .A(n45), .B(n143), .Q(n342) );
  INV0 U42 ( .A(n45), .Q(n113) );
  INV0 U43 ( .A(n40), .Q(n116) );
  BUF6 U44 ( .A(i_data_A[17]), .Q(n43) );
  AOI220 U45 ( .A(pre_sum_2b[0]), .B(n140), .C(i_data_B[8]), .D(n153), .Q(n150) );
  AOI220 U47 ( .A(pre_sum_2b[1]), .B(n140), .C(i_data_B[9]), .D(n141), .Q(n135) );
  INV0 U48 ( .A(n14), .Q(n15) );
  INV0 U49 ( .A(n12), .Q(n13) );
  INV0 U50 ( .A(i_data_B[8]), .Q(n130) );
  INV0 U51 ( .A(i_data_B[9]), .Q(n128) );
  INV0 U52 ( .A(i_data_B[1]), .Q(n421) );
  NOR21 U53 ( .A(n70), .B(n281), .Q(n201) );
  NOR21 U55 ( .A(n97), .B(n70), .Q(n296) );
  INV3 U56 ( .A(n199), .Q(n99) );
  INV3 U57 ( .A(n60), .Q(n61) );
  BUF2 U58 ( .A(n90), .Q(n6) );
  BUF2 U59 ( .A(n90), .Q(n5) );
  AOI221 U60 ( .A(pre_subb[14]), .B(n99), .C(N255), .D(n5), .Q(n211) );
  AOI221 U61 ( .A(pre_sum_3a[8]), .B(n284), .C(pre_sum_3b[8]), .D(n97), .Q(
        n281) );
  INV3 U63 ( .A(n283), .Q(n96) );
  AOI221 U64 ( .A(pre_subb[12]), .B(n99), .C(N253), .D(n5), .Q(n238) );
  NOR21 U65 ( .A(n70), .B(n284), .Q(n294) );
  NOR21 U66 ( .A(n98), .B(n70), .Q(n140) );
  INV3 U67 ( .A(n63), .Q(n62) );
  NAND22 U68 ( .A(half_sub[16]), .B(n93), .Q(n199) );
  NAND22 U69 ( .A(n94), .B(n95), .Q(n429) );
  NOR21 U71 ( .A(n62), .B(n109), .Q(n290) );
  NOR21 U72 ( .A(n62), .B(n116), .Q(n369) );
  NOR21 U73 ( .A(n62), .B(n115), .Q(n359) );
  NOR21 U74 ( .A(n62), .B(n114), .Q(n349) );
  NOR21 U75 ( .A(n62), .B(n111), .Q(n312) );
  NOR21 U76 ( .A(n62), .B(n110), .Q(n302) );
  NOR21 U77 ( .A(n62), .B(n108), .Q(n277) );
  NOR21 U79 ( .A(n62), .B(n107), .Q(n267) );
  NOR21 U80 ( .A(n62), .B(n106), .Q(n257) );
  NOR21 U81 ( .A(n62), .B(n113), .Q(n339) );
  NOR21 U82 ( .A(n62), .B(n112), .Q(n322) );
  INV3 U83 ( .A(n202), .Q(n60) );
  NOR21 U84 ( .A(n69), .B(half_sub[16]), .Q(n202) );
  BUF2 U86 ( .A(n143), .Q(n59) );
  INV3 U88 ( .A(n67), .Q(n66) );
  INV3 U89 ( .A(n65), .Q(n64) );
  INV3 U90 ( .A(n84), .Q(n90) );
  AOI221 U91 ( .A(pre_subb[13]), .B(n99), .C(N254), .D(n5), .Q(n228) );
  NAND22 U92 ( .A(n8), .B(n203), .Q(n192) );
  AOI221 U93 ( .A(N256), .B(n6), .C(n65), .D(n1), .Q(n191) );
  AOI221 U94 ( .A(N224), .B(n91), .C(n58), .D(n63), .Q(n193) );
  AOI221 U96 ( .A(n231), .B(n30), .C(pre_sum_4a[5]), .D(n96), .Q(n222) );
  AOI221 U97 ( .A(i_data_B[29]), .B(n229), .C(pre_suba[13]), .D(n61), .Q(n224)
         );
  AOI221 U98 ( .A(n214), .B(n31), .C(pre_sum_4a[6]), .D(n96), .Q(n205) );
  AOI221 U99 ( .A(i_data_B[30]), .B(n212), .C(pre_suba[14]), .D(n202), .Q(n207) );
  OAI311 U100 ( .A(n139), .B(i_data_B[31]), .C(n58), .D(n197), .Q(n196) );
  INV3 U101 ( .A(pre_subb[15]), .Q(n100) );
  AOI221 U103 ( .A(pre_sum_2a[8]), .B(n98), .C(pre_sum_2b[8]), .D(sum_1[8]), 
        .Q(n284) );
  NAND41 U104 ( .A(n272), .B(n273), .C(n274), .D(n275), .Q(o_data_AluRes[24])
         );
  AOI221 U105 ( .A(n25), .B(n279), .C(pre_suba[8]), .D(n202), .Q(n274) );
  AOI2111 U106 ( .A(N217), .B(n91), .C(n276), .D(n277), .Q(n275) );
  NAND41 U108 ( .A(n262), .B(n263), .C(n264), .D(n265), .Q(o_data_AluRes[25])
         );
  AOI221 U109 ( .A(i_data_B[25]), .B(n269), .C(pre_suba[9]), .D(n61), .Q(n264)
         );
  AOI2111 U110 ( .A(N218), .B(n91), .C(n266), .D(n267), .Q(n265) );
  NAND41 U111 ( .A(n252), .B(n253), .C(n254), .D(n255), .Q(o_data_AluRes[26])
         );
  AOI221 U112 ( .A(i_data_B[26]), .B(n259), .C(pre_suba[10]), .D(n202), .Q(
        n254) );
  AOI2111 U113 ( .A(N219), .B(n91), .C(n256), .D(n257), .Q(n255) );
  NAND41 U115 ( .A(n242), .B(n243), .C(n244), .D(n245), .Q(o_data_AluRes[27])
         );
  AOI221 U116 ( .A(i_data_B[27]), .B(n249), .C(pre_suba[11]), .D(n61), .Q(n244) );
  AOI221 U117 ( .A(n251), .B(n28), .C(pre_sum_4a[3]), .D(n96), .Q(n242) );
  NAND41 U118 ( .A(n232), .B(n233), .C(n234), .D(n235), .Q(o_data_AluRes[28])
         );
  AOI221 U119 ( .A(n241), .B(n29), .C(pre_sum_4a[4]), .D(n96), .Q(n232) );
  AOI221 U120 ( .A(i_data_B[28]), .B(n239), .C(pre_suba[12]), .D(n202), .Q(
        n234) );
  AOI221 U122 ( .A(n282), .B(n24), .C(pre_sum_4a[0]), .D(n96), .Q(n272) );
  AOI221 U123 ( .A(n271), .B(n26), .C(pre_sum_4a[1]), .D(n96), .Q(n262) );
  AOI221 U124 ( .A(pre_subb[11]), .B(n99), .C(N252), .D(n5), .Q(n248) );
  NOR21 U126 ( .A(n70), .B(sum_1[8]), .Q(n138) );
  NAND41 U127 ( .A(n148), .B(n149), .C(n150), .D(n151), .Q(o_data_AluRes[8])
         );
  AOI221 U128 ( .A(N201), .B(n91), .C(n32), .D(n63), .Q(n148) );
  AOI221 U129 ( .A(N233), .B(n6), .C(half_sub[8]), .D(n93), .Q(n149) );
  AOI221 U130 ( .A(n152), .B(n130), .C(pre_sum_2a[0]), .D(n138), .Q(n151) );
  NAND41 U131 ( .A(n133), .B(n134), .C(n135), .D(n136), .Q(o_data_AluRes[9])
         );
  AOI221 U133 ( .A(N202), .B(n91), .C(n63), .D(i_data_A[9]), .Q(n133) );
  AOI221 U134 ( .A(N234), .B(n90), .C(half_sub[9]), .D(n93), .Q(n134) );
  AOI221 U135 ( .A(n137), .B(n128), .C(pre_sum_2a[1]), .D(n138), .Q(n136) );
  NAND41 U137 ( .A(n409), .B(n410), .C(n411), .D(n412), .Q(o_data_AluRes[10])
         );
  AOI221 U138 ( .A(N203), .B(n91), .C(n34), .D(n63), .Q(n409) );
  AOI221 U139 ( .A(N235), .B(n6), .C(half_sub[10]), .D(n93), .Q(n410) );
  AOI221 U140 ( .A(n413), .B(n126), .C(pre_sum_2a[2]), .D(n138), .Q(n412) );
  NAND41 U141 ( .A(n402), .B(n403), .C(n404), .D(n405), .Q(o_data_AluRes[11])
         );
  AOI221 U142 ( .A(N204), .B(n91), .C(n35), .D(n63), .Q(n402) );
  AOI221 U144 ( .A(N236), .B(n90), .C(half_sub[11]), .D(n93), .Q(n403) );
  AOI221 U145 ( .A(n406), .B(n124), .C(pre_sum_2a[3]), .D(n138), .Q(n405) );
  NAND41 U146 ( .A(n395), .B(n396), .C(n397), .D(n398), .Q(o_data_AluRes[12])
         );
  AOI221 U148 ( .A(N205), .B(n91), .C(i_data_A[12]), .D(n63), .Q(n395) );
  AOI221 U149 ( .A(N237), .B(n6), .C(half_sub[12]), .D(n93), .Q(n396) );
  AOI221 U150 ( .A(n399), .B(n122), .C(pre_sum_2a[4]), .D(n138), .Q(n398) );
  NAND41 U151 ( .A(n388), .B(n389), .C(n390), .D(n391), .Q(o_data_AluRes[13])
         );
  AOI221 U152 ( .A(N206), .B(n91), .C(i_data_A[13]), .D(n63), .Q(n388) );
  AOI221 U153 ( .A(N238), .B(n90), .C(half_sub[13]), .D(n93), .Q(n389) );
  AOI221 U155 ( .A(n392), .B(n120), .C(pre_sum_2a[5]), .D(n138), .Q(n391) );
  NAND41 U156 ( .A(n381), .B(n382), .C(n383), .D(n384), .Q(o_data_AluRes[14])
         );
  AOI221 U157 ( .A(N207), .B(n91), .C(n38), .D(n63), .Q(n381) );
  AOI221 U159 ( .A(N239), .B(n6), .C(half_sub[14]), .D(n93), .Q(n382) );
  AOI221 U160 ( .A(n385), .B(n118), .C(pre_sum_2a[6]), .D(n138), .Q(n384) );
  NAND41 U161 ( .A(n374), .B(n375), .C(n376), .D(n377), .Q(o_data_AluRes[15])
         );
  AOI221 U162 ( .A(N208), .B(n91), .C(n39), .D(n63), .Q(n374) );
  AOI221 U163 ( .A(N240), .B(n90), .C(half_sub[15]), .D(n93), .Q(n375) );
  AOI221 U164 ( .A(n378), .B(n7), .C(pre_sum_2a[7]), .D(n138), .Q(n377) );
  NAND41 U166 ( .A(n285), .B(n286), .C(n287), .D(n288), .Q(o_data_AluRes[23])
         );
  AOI221 U167 ( .A(i_data_B[23]), .B(n292), .C(pre_suba[7]), .D(n61), .Q(n287)
         );
  AOI2111 U168 ( .A(N216), .B(n91), .C(n289), .D(n290), .Q(n288) );
  NAND22 U170 ( .A(pre_sum_3b[7]), .B(n294), .Q(n286) );
  NAND41 U171 ( .A(n364), .B(n365), .C(n366), .D(n367), .Q(o_data_AluRes[16])
         );
  AOI2111 U172 ( .A(N209), .B(n91), .C(n368), .D(n369), .Q(n367) );
  NAND22 U173 ( .A(pre_sum_3b[0]), .B(n294), .Q(n365) );
  NAND41 U174 ( .A(n354), .B(n355), .C(n356), .D(n357), .Q(o_data_AluRes[17])
         );
  AOI221 U175 ( .A(n11), .B(n361), .C(pre_suba[1]), .D(n61), .Q(n356) );
  AOI2111 U176 ( .A(N210), .B(n91), .C(n358), .D(n359), .Q(n357) );
  NAND22 U177 ( .A(pre_sum_3b[1]), .B(n294), .Q(n355) );
  NAND41 U178 ( .A(n344), .B(n345), .C(n346), .D(n347), .Q(o_data_AluRes[18])
         );
  AOI221 U180 ( .A(i_data_B[18]), .B(n351), .C(pre_suba[2]), .D(n61), .Q(n346)
         );
  AOI2111 U181 ( .A(N211), .B(n91), .C(n348), .D(n349), .Q(n347) );
  NAND22 U182 ( .A(pre_sum_3b[2]), .B(n294), .Q(n345) );
  NAND41 U184 ( .A(n334), .B(n335), .C(n336), .D(n337), .Q(o_data_AluRes[19])
         );
  AOI221 U185 ( .A(i_data_B[19]), .B(n341), .C(pre_suba[3]), .D(n61), .Q(n336)
         );
  AOI2111 U186 ( .A(N212), .B(n91), .C(n338), .D(n339), .Q(n337) );
  NAND22 U187 ( .A(pre_sum_3b[3]), .B(n294), .Q(n335) );
  NAND41 U188 ( .A(n317), .B(n318), .C(n319), .D(n320), .Q(o_data_AluRes[20])
         );
  AOI221 U189 ( .A(i_data_B[20]), .B(n324), .C(pre_suba[4]), .D(n61), .Q(n319)
         );
  AOI2111 U191 ( .A(N213), .B(n91), .C(n321), .D(n322), .Q(n320) );
  NAND22 U192 ( .A(pre_sum_3b[4]), .B(n294), .Q(n318) );
  NAND41 U193 ( .A(n307), .B(n308), .C(n309), .D(n310), .Q(o_data_AluRes[21])
         );
  AOI221 U195 ( .A(n19), .B(n314), .C(pre_suba[5]), .D(n61), .Q(n309) );
  AOI2111 U196 ( .A(N214), .B(n91), .C(n311), .D(n312), .Q(n310) );
  NAND22 U197 ( .A(pre_sum_3b[5]), .B(n294), .Q(n308) );
  NAND41 U198 ( .A(n297), .B(n298), .C(n299), .D(n300), .Q(o_data_AluRes[22])
         );
  AOI221 U199 ( .A(i_data_B[22]), .B(n304), .C(pre_suba[6]), .D(n202), .Q(n299) );
  AOI2111 U200 ( .A(N215), .B(n91), .C(n301), .D(n302), .Q(n300) );
  NAND22 U202 ( .A(pre_sum_3b[6]), .B(n294), .Q(n298) );
  AOI221 U203 ( .A(n373), .B(n9), .C(pre_sum_3a[0]), .D(n296), .Q(n364) );
  AOI221 U204 ( .A(n363), .B(n10), .C(pre_sum_3a[1]), .D(n296), .Q(n354) );
  AOI221 U206 ( .A(n353), .B(n12), .C(pre_sum_3a[2]), .D(n296), .Q(n344) );
  AOI221 U207 ( .A(n343), .B(n14), .C(pre_sum_3a[3]), .D(n296), .Q(n334) );
  AOI221 U208 ( .A(n326), .B(n16), .C(pre_sum_3a[4]), .D(n296), .Q(n317) );
  AOI221 U209 ( .A(n316), .B(n18), .C(pre_sum_3a[5]), .D(n296), .Q(n307) );
  AOI221 U210 ( .A(n306), .B(n20), .C(pre_sum_3a[6]), .D(n296), .Q(n297) );
  AOI221 U211 ( .A(n295), .B(n22), .C(pre_sum_3a[7]), .D(n296), .Q(n285) );
  AOI221 U213 ( .A(pre_subb[7]), .B(n99), .C(N248), .D(n5), .Q(n291) );
  AOI221 U214 ( .A(pre_subb[8]), .B(n99), .C(N249), .D(n5), .Q(n278) );
  AOI221 U215 ( .A(pre_subb[9]), .B(n99), .C(N250), .D(n5), .Q(n268) );
  AOI221 U217 ( .A(pre_subb[10]), .B(n99), .C(N251), .D(n5), .Q(n258) );
  AOI221 U218 ( .A(pre_sum_2b[7]), .B(n140), .C(n8), .D(n379), .Q(n376) );
  OAI2111 U219 ( .A(n39), .B(n425), .C(n424), .D(n380), .Q(n379) );
  NAND22 U220 ( .A(n39), .B(n143), .Q(n380) );
  AOI221 U221 ( .A(N226), .B(n6), .C(half_sub[1]), .D(n93), .Q(n329) );
  AOI221 U222 ( .A(N229), .B(n6), .C(half_sub[4]), .D(n93), .Q(n179) );
  AOI221 U224 ( .A(N230), .B(n90), .C(half_sub[5]), .D(n93), .Q(n172) );
  OAI2111 U225 ( .A(n49), .B(n64), .C(n62), .D(n293), .Q(n292) );
  NAND22 U226 ( .A(n49), .B(n59), .Q(n293) );
  OAI2111 U227 ( .A(i_data_A[29]), .B(n64), .C(n424), .D(n230), .Q(n229) );
  NAND22 U229 ( .A(i_data_A[29]), .B(n59), .Q(n230) );
  OAI2111 U230 ( .A(n43), .B(n64), .C(n424), .D(n362), .Q(n361) );
  NAND22 U231 ( .A(n43), .B(n143), .Q(n362) );
  OAI2111 U232 ( .A(n46), .B(n425), .C(n424), .D(n325), .Q(n324) );
  NAND22 U233 ( .A(n46), .B(n143), .Q(n325) );
  OAI2111 U234 ( .A(n47), .B(n425), .C(n62), .D(n315), .Q(n314) );
  NAND22 U236 ( .A(n47), .B(n59), .Q(n315) );
  OAI2111 U237 ( .A(n48), .B(n425), .C(n424), .D(n305), .Q(n304) );
  NAND22 U238 ( .A(n48), .B(n59), .Q(n305) );
  OAI2111 U239 ( .A(n50), .B(n64), .C(n424), .D(n280), .Q(n279) );
  NAND22 U240 ( .A(n50), .B(n59), .Q(n280) );
  OAI2111 U241 ( .A(n51), .B(n425), .C(n62), .D(n270), .Q(n269) );
  NAND22 U243 ( .A(n51), .B(n59), .Q(n270) );
  OAI2111 U244 ( .A(n52), .B(n64), .C(n424), .D(n260), .Q(n259) );
  NAND22 U245 ( .A(n52), .B(n59), .Q(n260) );
  OAI2111 U247 ( .A(i_data_A[27]), .B(n64), .C(n424), .D(n250), .Q(n249) );
  NAND22 U248 ( .A(i_data_A[27]), .B(n59), .Q(n250) );
  OAI2111 U249 ( .A(n54), .B(n64), .C(n424), .D(n240), .Q(n239) );
  NAND22 U250 ( .A(n54), .B(n59), .Q(n240) );
  OAI2111 U251 ( .A(i_data_A[30]), .B(n425), .C(n62), .D(n213), .Q(n212) );
  NAND22 U252 ( .A(i_data_A[30]), .B(n59), .Q(n213) );
  AOI221 U253 ( .A(N227), .B(n90), .C(half_sub[2]), .D(n93), .Q(n217) );
  AOI221 U254 ( .A(N231), .B(n6), .C(half_sub[6]), .D(n93), .Q(n165) );
  INV3 U255 ( .A(n424), .Q(n63) );
  AOI221 U256 ( .A(pre_subb[3]), .B(n99), .C(N244), .D(n6), .Q(n340) );
  AOI221 U258 ( .A(pre_subb[4]), .B(n99), .C(N245), .D(n90), .Q(n323) );
  AOI221 U259 ( .A(pre_subb[5]), .B(n99), .C(N246), .D(n5), .Q(n313) );
  AOI221 U260 ( .A(pre_subb[6]), .B(n99), .C(N247), .D(n5), .Q(n303) );
  AOI221 U261 ( .A(pre_subb[1]), .B(n99), .C(N242), .D(n6), .Q(n360) );
  AOI221 U262 ( .A(pre_subb[2]), .B(n99), .C(N243), .D(n5), .Q(n350) );
  INV3 U263 ( .A(n70), .Q(n92) );
  NAND31 U265 ( .A(i_con_AluCtrl[1]), .B(n72), .C(n82), .Q(n70) );
  IMUX21 U266 ( .A(n79), .B(n74), .S(n1), .Q(n76) );
  INV3 U267 ( .A(n69), .Q(n93) );
  INV3 U269 ( .A(n49), .Q(n109) );
  INV3 U270 ( .A(n203), .Q(n427) );
  NAND31 U271 ( .A(i_con_AluCtrl[1]), .B(i_con_AluCtrl[2]), .C(n94), .Q(n80)
         );
  INV3 U272 ( .A(n33), .Q(n129) );
  INV3 U273 ( .A(n35), .Q(n125) );
  INV3 U274 ( .A(n36), .Q(n123) );
  INV3 U275 ( .A(i_data_A[13]), .Q(n121) );
  INV3 U276 ( .A(n38), .Q(n119) );
  INV3 U277 ( .A(n39), .Q(n117) );
  INV3 U278 ( .A(n32), .Q(n131) );
  INV3 U279 ( .A(n34), .Q(n127) );
  NOR21 U280 ( .A(n429), .B(i_con_AluCtrl[1]), .Q(n143) );
  INV3 U282 ( .A(n198), .Q(n101) );
  NAND22 U283 ( .A(n59), .B(n58), .Q(n198) );
  INV3 U285 ( .A(n425), .Q(n65) );
  NOR21 U286 ( .A(n95), .B(i_con_AluCtrl[1]), .Q(n426) );
  INV3 U287 ( .A(n139), .Q(n67) );
  INV3 U288 ( .A(i_data_A[29]), .Q(n103) );
  INV3 U289 ( .A(n50), .Q(n108) );
  INV3 U290 ( .A(n43), .Q(n115) );
  INV3 U291 ( .A(n48), .Q(n110) );
  INV3 U293 ( .A(n46), .Q(n112) );
  INV3 U294 ( .A(n47), .Q(n111) );
  INV3 U295 ( .A(n51), .Q(n107) );
  INV3 U296 ( .A(n52), .Q(n106) );
  INV3 U297 ( .A(i_data_A[27]), .Q(n105) );
  INV3 U298 ( .A(n54), .Q(n104) );
  INV3 U299 ( .A(i_data_A[30]), .Q(n102) );
  NOR21 U301 ( .A(n62), .B(n103), .Q(n227) );
  NOR21 U302 ( .A(n62), .B(n102), .Q(n210) );
  AOI2111 U303 ( .A(N220), .B(n91), .C(n246), .D(n247), .Q(n245) );
  NOR21 U304 ( .A(n62), .B(n105), .Q(n247) );
  AOI2111 U305 ( .A(N221), .B(n91), .C(n236), .D(n237), .Q(n235) );
  NOR21 U306 ( .A(n62), .B(n104), .Q(n237) );
  BUF2 U307 ( .A(i_data_A[19]), .Q(n45) );
  BUF2 U309 ( .A(i_data_A[20]), .Q(n46) );
  INV3 U310 ( .A(n16), .Q(n17) );
  INV3 U311 ( .A(n18), .Q(n19) );
  OAI2111 U312 ( .A(n32), .B(n425), .C(n62), .D(n154), .Q(n153) );
  NAND22 U313 ( .A(n32), .B(n59), .Q(n154) );
  OAI2111 U314 ( .A(i_data_A[9]), .B(n425), .C(n62), .D(n142), .Q(n141) );
  NAND22 U315 ( .A(n59), .B(i_data_A[9]), .Q(n142) );
  AOI221 U317 ( .A(pre_sum_2b[2]), .B(n140), .C(i_data_B[10]), .D(n414), .Q(
        n411) );
  OAI2111 U318 ( .A(n34), .B(n425), .C(n62), .D(n415), .Q(n414) );
  NAND22 U319 ( .A(n34), .B(n143), .Q(n415) );
  AOI221 U320 ( .A(pre_sum_2b[3]), .B(n140), .C(i_data_B[11]), .D(n407), .Q(
        n404) );
  OAI2111 U321 ( .A(n35), .B(n425), .C(n62), .D(n408), .Q(n407) );
  NAND22 U322 ( .A(n35), .B(n143), .Q(n408) );
  AOI221 U323 ( .A(pre_sum_2b[4]), .B(n140), .C(i_data_B[12]), .D(n400), .Q(
        n397) );
  OAI2111 U324 ( .A(i_data_A[12]), .B(n425), .C(n424), .D(n401), .Q(n400) );
  NAND22 U326 ( .A(i_data_A[12]), .B(n143), .Q(n401) );
  AOI221 U327 ( .A(pre_sum_2b[5]), .B(n140), .C(i_data_B[13]), .D(n393), .Q(
        n390) );
  OAI2111 U328 ( .A(i_data_A[13]), .B(n425), .C(n424), .D(n394), .Q(n393) );
  NAND22 U329 ( .A(i_data_A[13]), .B(n143), .Q(n394) );
  AOI221 U330 ( .A(pre_sum_2b[6]), .B(n140), .C(i_data_B[14]), .D(n386), .Q(
        n383) );
  OAI2111 U331 ( .A(n38), .B(n425), .C(n424), .D(n387), .Q(n386) );
  NAND22 U332 ( .A(n38), .B(n143), .Q(n387) );
  BUF2 U333 ( .A(i_data_A[22]), .Q(n48) );
  BUF2 U334 ( .A(i_data_A[10]), .Q(n34) );
  BUF2 U335 ( .A(i_data_A[8]), .Q(n32) );
  INV3 U336 ( .A(n24), .Q(n25) );
  BUF2 U337 ( .A(i_data_A[21]), .Q(n47) );
  BUF2 U338 ( .A(i_data_A[16]), .Q(n40) );
  INV3 U339 ( .A(n20), .Q(n21) );
  INV3 U340 ( .A(n22), .Q(n23) );
  BUF2 U341 ( .A(i_data_A[9]), .Q(n33) );
  AOI221 U342 ( .A(N225), .B(n6), .C(half_sub[0]), .D(n93), .Q(n87) );
  OAI2111 U343 ( .A(i_data_A[4]), .B(n64), .C(n62), .D(n183), .Q(n182) );
  NAND22 U344 ( .A(i_data_A[4]), .B(n59), .Q(n183) );
  OAI2111 U345 ( .A(i_data_A[7]), .B(n425), .C(n62), .D(n161), .Q(n160) );
  NAND22 U346 ( .A(i_data_A[7]), .B(n59), .Q(n161) );
  OAI2111 U347 ( .A(i_data_A[3]), .B(n425), .C(n62), .D(n190), .Q(n189) );
  NAND22 U348 ( .A(i_data_A[3]), .B(n59), .Q(n190) );
  OAI2111 U349 ( .A(i_data_A[0]), .B(n425), .C(n428), .D(n424), .Q(n85) );
  NAND22 U350 ( .A(i_data_A[0]), .B(n143), .Q(n428) );
  OAI2111 U351 ( .A(i_data_A[1]), .B(n64), .C(n424), .D(n333), .Q(n332) );
  NAND22 U352 ( .A(i_data_A[1]), .B(n143), .Q(n333) );
  OAI2111 U353 ( .A(i_data_A[6]), .B(n425), .C(n62), .D(n169), .Q(n168) );
  OAI2111 U354 ( .A(i_data_A[2]), .B(n64), .C(n62), .D(n221), .Q(n220) );
  NAND22 U355 ( .A(i_data_A[2]), .B(n59), .Q(n221) );
  OAI2111 U356 ( .A(i_data_A[5]), .B(n425), .C(n62), .D(n176), .Q(n175) );
  NAND41 U357 ( .A(n89), .B(n88), .C(n87), .D(n86), .Q(o_data_AluRes[0]) );
  IMUX30 U358 ( .A(n67), .B(n65), .C(n85), .S0(i_data_A[0]), .S1(i_data_B[0]), 
        .Q(n86) );
  AOI221 U359 ( .A(i_con_AluCtrl[0]), .B(n81), .C(sum_1[0]), .D(n92), .Q(n89)
         );
  AOI221 U360 ( .A(N193), .B(n91), .C(i_data_A[0]), .D(n63), .Q(n88) );
  NAND41 U361 ( .A(n327), .B(n328), .C(n329), .D(n330), .Q(o_data_AluRes[1])
         );
  NAND22 U362 ( .A(i_data_A[1]), .B(n63), .Q(n328) );
  AOI221 U363 ( .A(n331), .B(n421), .C(i_data_B[1]), .D(n332), .Q(n330) );
  AOI221 U364 ( .A(N194), .B(n91), .C(sum_1[1]), .D(n92), .Q(n327) );
  NAND41 U365 ( .A(n215), .B(n216), .C(n217), .D(n218), .Q(o_data_AluRes[2])
         );
  NAND22 U366 ( .A(i_data_A[2]), .B(n63), .Q(n216) );
  AOI221 U367 ( .A(n219), .B(n419), .C(i_data_B[2]), .D(n220), .Q(n218) );
  AOI221 U368 ( .A(N195), .B(n91), .C(sum_1[2]), .D(n92), .Q(n215) );
  NAND41 U369 ( .A(n184), .B(n185), .C(n186), .D(n187), .Q(o_data_AluRes[3])
         );
  NAND22 U370 ( .A(i_data_A[3]), .B(n63), .Q(n185) );
  AOI221 U371 ( .A(N196), .B(n91), .C(sum_1[3]), .D(n92), .Q(n184) );
  AOI221 U372 ( .A(n188), .B(n417), .C(i_data_B[3]), .D(n189), .Q(n187) );
  NAND41 U373 ( .A(n177), .B(n178), .C(n179), .D(n180), .Q(o_data_AluRes[4])
         );
  NAND22 U374 ( .A(i_data_A[4]), .B(n63), .Q(n178) );
  AOI221 U375 ( .A(n181), .B(n204), .C(i_data_B[4]), .D(n182), .Q(n180) );
  AOI221 U376 ( .A(N197), .B(n91), .C(sum_1[4]), .D(n92), .Q(n177) );
  NAND41 U377 ( .A(n170), .B(n171), .C(n172), .D(n173), .Q(o_data_AluRes[5])
         );
  NAND22 U378 ( .A(i_data_A[5]), .B(n63), .Q(n171) );
  AOI221 U379 ( .A(n174), .B(n147), .C(i_data_B[5]), .D(n175), .Q(n173) );
  AOI221 U380 ( .A(N198), .B(n91), .C(sum_1[5]), .D(n92), .Q(n170) );
  NAND41 U381 ( .A(n163), .B(n164), .C(n165), .D(n166), .Q(o_data_AluRes[6])
         );
  NAND22 U382 ( .A(i_data_A[6]), .B(n63), .Q(n164) );
  AOI221 U383 ( .A(n167), .B(n145), .C(i_data_B[6]), .D(n168), .Q(n166) );
  AOI221 U384 ( .A(N199), .B(n91), .C(sum_1[6]), .D(n92), .Q(n163) );
  NAND41 U385 ( .A(n155), .B(n156), .C(n157), .D(n158), .Q(o_data_AluRes[7])
         );
  NAND22 U386 ( .A(i_data_A[7]), .B(n63), .Q(n156) );
  AOI221 U387 ( .A(n159), .B(n132), .C(i_data_B[7]), .D(n160), .Q(n158) );
  AOI221 U388 ( .A(N232), .B(n90), .C(half_sub[7]), .D(n93), .Q(n157) );
  AOI221 U389 ( .A(N228), .B(n90), .C(half_sub[3]), .D(n93), .Q(n186) );
  AOI221 U390 ( .A(N200), .B(n91), .C(sum_1[7]), .D(n92), .Q(n155) );
  BUF2 U391 ( .A(i_data_A[24]), .Q(n50) );
  AOI221 U392 ( .A(pre_subb[0]), .B(n99), .C(N241), .D(n90), .Q(n370) );
  BUF2 U393 ( .A(i_data_A[12]), .Q(n36) );
  BUF2 U394 ( .A(i_data_A[11]), .Q(n35) );
  INV3 U395 ( .A(n7), .Q(n8) );
  BUF2 U396 ( .A(i_data_A[25]), .Q(n51) );
  BUF2 U397 ( .A(i_data_A[26]), .Q(n52) );
  BUF2 U398 ( .A(i_data_A[13]), .Q(n37) );
  BUF2 U399 ( .A(i_data_A[27]), .Q(n53) );
  NOR40 U400 ( .A(n94), .B(i_con_AluCtrl[0]), .C(i_con_AluCtrl[1]), .D(
        i_con_AluCtrl[2]), .Q(n203) );
  INV3 U401 ( .A(i_data_A[4]), .Q(n416) );
  INV3 U402 ( .A(i_data_A[7]), .Q(n144) );
  INV3 U403 ( .A(i_data_A[3]), .Q(n418) );
  INV3 U404 ( .A(i_data_A[1]), .Q(n422) );
  INV3 U405 ( .A(i_data_A[6]), .Q(n146) );
  INV3 U406 ( .A(i_data_A[2]), .Q(n420) );
  INV3 U407 ( .A(i_data_A[5]), .Q(n162) );
  NAND31 U408 ( .A(i_con_AluCtrl[0]), .B(i_con_AluCtrl[1]), .C(n82), .Q(n83)
         );
  BUF2 U409 ( .A(i_data_A[15]), .Q(n39) );
  BUF2 U410 ( .A(i_data_A[28]), .Q(n54) );
  BUF2 U411 ( .A(i_data_A[31]), .Q(n58) );
  BUF2 U412 ( .A(i_data_A[30]), .Q(n56) );
  BUF2 U413 ( .A(i_data_A[14]), .Q(n38) );
  BUF2 U414 ( .A(i_data_A[31]), .Q(n57) );
  BUF2 U415 ( .A(i_data_A[29]), .Q(n55) );
  INV3 U416 ( .A(i_data_B[11]), .Q(n124) );
  INV3 U417 ( .A(i_data_B[7]), .Q(n132) );
  INV3 U418 ( .A(i_data_B[12]), .Q(n122) );
  INV3 U419 ( .A(i_data_B[10]), .Q(n126) );
  INV3 U420 ( .A(i_data_B[14]), .Q(n118) );
  INV3 U421 ( .A(i_data_B[13]), .Q(n120) );
  INV3 U422 ( .A(i_data_B[4]), .Q(n204) );
  INV3 U423 ( .A(i_data_B[6]), .Q(n145) );
  INV3 U424 ( .A(i_data_B[5]), .Q(n147) );
  INV3 U425 ( .A(i_data_B[3]), .Q(n417) );
  INV3 U426 ( .A(i_data_B[2]), .Q(n419) );
  INV3 U427 ( .A(i_data_B[18]), .Q(n12) );
  INV3 U428 ( .A(i_data_B[17]), .Q(n10) );
  INV3 U429 ( .A(i_data_B[21]), .Q(n18) );
  INV3 U430 ( .A(i_data_B[20]), .Q(n16) );
  INV3 U431 ( .A(i_data_B[19]), .Q(n14) );
  INV3 U432 ( .A(i_data_B[24]), .Q(n24) );
  INV3 U433 ( .A(i_data_B[22]), .Q(n20) );
  INV3 U434 ( .A(i_data_B[23]), .Q(n22) );
  INV3 U435 ( .A(i_data_B[28]), .Q(n29) );
  INV3 U436 ( .A(i_data_B[26]), .Q(n27) );
  INV3 U437 ( .A(i_data_B[27]), .Q(n28) );
  INV3 U438 ( .A(i_data_B[30]), .Q(n31) );
  INV3 U439 ( .A(i_data_B[29]), .Q(n30) );
  INV3 U440 ( .A(i_data_B[15]), .Q(n7) );
  LOGIC0 U441 ( .Q(n42) );
  LOGIC1 U442 ( .Q(n41) );
  BUF2 U443 ( .A(i_data_A[23]), .Q(n49) );
  AOI221 U444 ( .A(pre_sum_4b[7]), .B(n201), .C(pre_suba[15]), .D(n61), .Q(
        n200) );
  CLKIN3 U445 ( .A(i_con_AluCtrl[3]), .Q(n94) );
  CLKIN3 U446 ( .A(n80), .Q(n68) );
  CLKIN3 U447 ( .A(i_con_AluCtrl[0]), .Q(n72) );
  NAND22 U448 ( .A(n68), .B(n72), .Q(n69) );
  CLKIN3 U449 ( .A(n429), .Q(n82) );
  CLKIN3 U450 ( .A(i_con_AluCtrl[1]), .Q(n75) );
  NAND22 U451 ( .A(n426), .B(i_con_AluCtrl[3]), .Q(n71) );
  CLKIN3 U452 ( .A(n71), .Q(n73) );
  NAND22 U453 ( .A(n73), .B(n72), .Q(n139) );
  NAND22 U454 ( .A(n73), .B(i_con_AluCtrl[0]), .Q(n425) );
  CLKIN3 U455 ( .A(N306), .Q(n79) );
  CLKIN3 U456 ( .A(n58), .Q(n74) );
  NAND22 U457 ( .A(n76), .B(n75), .Q(n78) );
  CLKIN3 U458 ( .A(i_con_AluCtrl[2]), .Q(n95) );
  NAND22 U459 ( .A(i_con_AluCtrl[3]), .B(n95), .Q(n77) );
  OAI222 U460 ( .A(n80), .B(n79), .C(n78), .D(n77), .Q(n81) );
  CLKIN3 U461 ( .A(n83), .Q(n91) );
  NAND22 U462 ( .A(n426), .B(n94), .Q(n84) );
  CLKIN3 U463 ( .A(i_data_B[0]), .Q(n423) );
endmodule


module E_alu_control ( o_con_AluCtrl, i_con_AluOp, i_con_FuncCode );
  output [3:0] o_con_AluCtrl;
  input [5:0] i_con_AluOp;
  input [5:0] i_con_FuncCode;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21;

  OAI212 U4 ( .A(n25), .B(n26), .C(n9), .Q(n23) );
  OAI212 U12 ( .A(n35), .B(n40), .C(n9), .Q(n36) );
  OAI2111 U3 ( .A(n27), .B(n28), .C(n29), .D(n2), .Q(o_con_AluCtrl[2]) );
  INV3 U5 ( .A(n30), .Q(n2) );
  NOR40 U6 ( .A(n12), .B(n31), .C(n16), .D(n26), .Q(n27) );
  INV3 U7 ( .A(n33), .Q(n16) );
  OAI2111 U8 ( .A(n20), .B(n32), .C(n11), .D(n18), .Q(n26) );
  OAI2111 U9 ( .A(n10), .B(n22), .C(n23), .D(n24), .Q(o_con_AluCtrl[3]) );
  NAND31 U10 ( .A(n21), .B(n20), .C(n47), .Q(n49) );
  NOR21 U11 ( .A(n21), .B(n14), .Q(n31) );
  INV3 U13 ( .A(n50), .Q(n11) );
  NOR40 U14 ( .A(n25), .B(n35), .C(n31), .D(n51), .Q(n50) );
  NAND31 U15 ( .A(n49), .B(n32), .C(n33), .Q(n51) );
  NAND41 U16 ( .A(n49), .B(n13), .C(n11), .D(n18), .Q(n40) );
  INV3 U17 ( .A(n31), .Q(n13) );
  NAND41 U18 ( .A(n36), .B(n29), .C(n6), .D(n37), .Q(o_con_AluCtrl[1]) );
  INV3 U19 ( .A(n39), .Q(n6) );
  NOR21 U20 ( .A(n8), .B(n1), .Q(n37) );
  INV3 U21 ( .A(n22), .Q(n4) );
  INV3 U22 ( .A(n38), .Q(n1) );
  INV3 U23 ( .A(n28), .Q(n9) );
  NOR31 U24 ( .A(i_con_FuncCode[3]), .B(i_con_FuncCode[5]), .C(
        i_con_FuncCode[2]), .Q(n47) );
  NOR21 U25 ( .A(n14), .B(i_con_FuncCode[0]), .Q(n25) );
  INV3 U26 ( .A(i_con_FuncCode[1]), .Q(n20) );
  INV3 U27 ( .A(n53), .Q(n14) );
  NOR40 U28 ( .A(n15), .B(n19), .C(n20), .D(i_con_FuncCode[2]), .Q(n53) );
  INV3 U29 ( .A(i_con_FuncCode[5]), .Q(n15) );
  INV3 U30 ( .A(i_con_FuncCode[3]), .Q(n19) );
  OAI2111 U31 ( .A(n41), .B(n28), .C(n24), .D(n42), .Q(o_con_AluCtrl[0]) );
  AOI311 U32 ( .A(i_con_AluOp[3]), .B(i_con_AluOp[0]), .C(n43), .D(n3), .Q(n42) );
  AOI2111 U33 ( .A(n47), .B(i_con_FuncCode[0]), .C(n48), .D(n40), .Q(n41) );
  INV3 U34 ( .A(n29), .Q(n3) );
  NAND31 U35 ( .A(i_con_FuncCode[5]), .B(n19), .C(i_con_FuncCode[2]), .Q(n32)
         );
  NOR40 U36 ( .A(n5), .B(n7), .C(i_con_AluOp[3]), .D(i_con_AluOp[4]), .Q(n44)
         );
  NOR31 U37 ( .A(i_con_FuncCode[2]), .B(i_con_FuncCode[3]), .C(n15), .Q(n35)
         );
  AOI211 U38 ( .A(n8), .B(i_con_AluOp[0]), .C(n46), .Q(n38) );
  NOR40 U39 ( .A(n10), .B(n43), .C(n44), .D(n4), .Q(n46) );
  AOI311 U40 ( .A(n4), .B(n7), .C(i_con_AluOp[0]), .D(n30), .Q(n24) );
  NAND31 U41 ( .A(i_con_AluOp[3]), .B(n5), .C(i_con_AluOp[4]), .Q(n22) );
  OAI311 U42 ( .A(n32), .B(i_con_FuncCode[1]), .C(n21), .D(n52), .Q(n48) );
  AOI311 U43 ( .A(i_con_FuncCode[1]), .B(n21), .C(n17), .D(n25), .Q(n52) );
  INV3 U44 ( .A(n32), .Q(n17) );
  NOR21 U45 ( .A(i_con_AluOp[5]), .B(i_con_AluOp[4]), .Q(n43) );
  NAND22 U46 ( .A(n44), .B(i_con_AluOp[0]), .Q(n29) );
  NAND22 U47 ( .A(i_con_AluOp[1]), .B(n10), .Q(n28) );
  INV3 U48 ( .A(i_con_AluOp[0]), .Q(n10) );
  NAND22 U49 ( .A(n47), .B(i_con_FuncCode[1]), .Q(n33) );
  INV3 U50 ( .A(i_con_FuncCode[0]), .Q(n21) );
  NAND22 U51 ( .A(n38), .B(n45), .Q(n30) );
  NAND41 U52 ( .A(n43), .B(i_con_AluOp[2]), .C(i_con_AluOp[3]), .D(
        i_con_AluOp[0]), .Q(n45) );
  INV3 U53 ( .A(i_con_AluOp[2]), .Q(n7) );
  INV3 U54 ( .A(i_con_AluOp[5]), .Q(n5) );
  INV3 U55 ( .A(i_con_AluOp[1]), .Q(n8) );
  INV3 U56 ( .A(i_con_FuncCode[4]), .Q(n18) );
  INV3 U57 ( .A(n34), .Q(n12) );
  NAND22 U58 ( .A(i_con_FuncCode[1]), .B(n35), .Q(n34) );
  NOR31 U59 ( .A(i_con_AluOp[2]), .B(i_con_AluOp[3]), .C(n10), .Q(n39) );
endmodule


module E_famux5 ( i_data_rs, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fa, o_data_alusra );
  input [31:0] i_data_rs;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fa;
  output [31:0] o_data_alusra;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  CLKBU4 U1 ( .A(n3), .Q(n5) );
  BUF2 U2 ( .A(n114), .Q(n10) );
  AOI221 U3 ( .A(i_data_lwM[16]), .B(n1), .C(i_data_lwW[16]), .D(n10), .Q(n67)
         );
  NAND31 U4 ( .A(n24), .B(n23), .C(n22), .Q(o_data_alusra[1]) );
  NAND31 U5 ( .A(n27), .B(n26), .C(n25), .Q(o_data_alusra[2]) );
  NAND31 U6 ( .A(n36), .B(n35), .C(n34), .Q(o_data_alusra[5]) );
  NAND31 U7 ( .A(i_con_fa[2]), .B(n15), .C(n17), .Q(n16) );
  NAND31 U8 ( .A(n39), .B(n38), .C(n37), .Q(o_data_alusra[6]) );
  NAND31 U9 ( .A(n21), .B(n20), .C(n19), .Q(o_data_alusra[0]) );
  INV3 U10 ( .A(n16), .Q(n1) );
  CLKIN3 U11 ( .A(i_con_fa[0]), .Q(n15) );
  AOI221 U12 ( .A(i_data_lwM[18]), .B(n1), .C(i_data_lwW[18]), .D(n10), .Q(n73) );
  BUF6 U13 ( .A(n113), .Q(n2) );
  NAND30 U14 ( .A(i_con_fa[1]), .B(n13), .C(n15), .Q(n14) );
  INV2 U15 ( .A(n18), .Q(n114) );
  AOI220 U16 ( .A(i_data_lwM[4]), .B(n1), .C(i_data_lwW[4]), .D(n8), .Q(n31)
         );
  AOI220 U17 ( .A(i_data_lwM[7]), .B(n1), .C(i_data_lwW[7]), .D(n8), .Q(n40)
         );
  AOI220 U18 ( .A(i_data_lwM[3]), .B(n1), .C(i_data_lwW[3]), .D(n8), .Q(n28)
         );
  AOI220 U19 ( .A(i_data_lwM[0]), .B(n1), .C(i_data_lwW[0]), .D(n8), .Q(n19)
         );
  AOI220 U20 ( .A(i_data_lwM[9]), .B(n1), .C(i_data_lwW[9]), .D(n8), .Q(n46)
         );
  AOI220 U21 ( .A(i_data_lwM[10]), .B(n1), .C(i_data_lwW[10]), .D(n8), .Q(n49)
         );
  AOI220 U22 ( .A(i_data_lwM[1]), .B(n1), .C(i_data_lwW[1]), .D(n8), .Q(n22)
         );
  NAND30 U23 ( .A(i_con_fa[0]), .B(n13), .C(n17), .Q(n12) );
  AOI220 U24 ( .A(i_data_rs[18]), .B(n5), .C(i_data_writeres[18]), .D(n112), 
        .Q(n75) );
  AOI220 U25 ( .A(i_data_rs[19]), .B(n5), .C(i_data_writeres[19]), .D(n7), .Q(
        n78) );
  AOI220 U26 ( .A(i_data_lwM[19]), .B(n1), .C(i_data_lwW[19]), .D(n9), .Q(n76)
         );
  AOI220 U27 ( .A(i_data_lwM[8]), .B(n1), .C(i_data_lwW[8]), .D(n8), .Q(n43)
         );
  AOI220 U28 ( .A(i_data_rs[20]), .B(n5), .C(i_data_writeres[20]), .D(n6), .Q(
        n81) );
  AOI220 U29 ( .A(i_data_lwM[20]), .B(n1), .C(i_data_lwW[20]), .D(n10), .Q(n79) );
  AOI220 U30 ( .A(i_data_rs[21]), .B(n5), .C(i_data_writeres[21]), .D(n7), .Q(
        n84) );
  AOI220 U31 ( .A(i_data_lwM[21]), .B(n1), .C(i_data_lwW[21]), .D(n9), .Q(n82)
         );
  AOI220 U32 ( .A(i_data_rs[22]), .B(n5), .C(i_data_writeres[22]), .D(n6), .Q(
        n87) );
  AOI220 U33 ( .A(i_data_lwM[22]), .B(n1), .C(i_data_lwW[22]), .D(n10), .Q(n85) );
  AOI220 U34 ( .A(i_data_rs[23]), .B(n5), .C(i_data_writeres[23]), .D(n7), .Q(
        n90) );
  AOI220 U35 ( .A(i_data_lwM[23]), .B(n1), .C(i_data_lwW[23]), .D(n9), .Q(n88)
         );
  AOI220 U36 ( .A(i_data_rs[31]), .B(n5), .C(i_data_writeres[31]), .D(n7), .Q(
        n117) );
  AOI220 U37 ( .A(i_data_lwM[31]), .B(n1), .C(i_data_lwW[31]), .D(n9), .Q(n115) );
  NAND30 U38 ( .A(i_con_fa[2]), .B(i_con_fa[0]), .C(n17), .Q(n18) );
  AOI220 U39 ( .A(i_data_lwM[6]), .B(n1), .C(i_data_lwW[6]), .D(n8), .Q(n37)
         );
  AOI220 U40 ( .A(i_data_lwM[2]), .B(n1), .C(i_data_lwW[2]), .D(n8), .Q(n25)
         );
  AOI220 U41 ( .A(i_data_lwM[5]), .B(n1), .C(i_data_lwW[5]), .D(n8), .Q(n34)
         );
  AOI220 U42 ( .A(i_data_rs[11]), .B(n4), .C(i_data_writeres[11]), .D(n7), .Q(
        n54) );
  AOI220 U43 ( .A(i_data_lwM[11]), .B(n1), .C(i_data_lwW[11]), .D(n9), .Q(n52)
         );
  AOI220 U44 ( .A(i_data_rs[12]), .B(n4), .C(i_data_writeres[12]), .D(n6), .Q(
        n57) );
  AOI220 U45 ( .A(i_data_lwM[12]), .B(n1), .C(i_data_lwW[12]), .D(n10), .Q(n55) );
  AOI220 U46 ( .A(i_data_rs[13]), .B(n4), .C(i_data_writeres[13]), .D(n7), .Q(
        n60) );
  AOI220 U47 ( .A(i_data_lwM[13]), .B(n1), .C(i_data_lwW[13]), .D(n9), .Q(n58)
         );
  AOI220 U48 ( .A(i_data_rs[14]), .B(n4), .C(i_data_writeres[14]), .D(n6), .Q(
        n63) );
  AOI220 U49 ( .A(i_data_lwM[14]), .B(n1), .C(i_data_lwW[14]), .D(n10), .Q(n61) );
  AOI220 U50 ( .A(i_data_rs[15]), .B(n4), .C(i_data_writeres[15]), .D(n7), .Q(
        n66) );
  AOI220 U51 ( .A(i_data_lwM[15]), .B(n1), .C(i_data_lwW[15]), .D(n9), .Q(n64)
         );
  AOI220 U52 ( .A(i_data_rs[27]), .B(n5), .C(i_data_writeres[27]), .D(n7), .Q(
        n102) );
  AOI220 U53 ( .A(i_data_lwM[27]), .B(n1), .C(i_data_lwW[27]), .D(n9), .Q(n100) );
  AOI220 U54 ( .A(i_data_rs[28]), .B(n5), .C(i_data_writeres[28]), .D(n112), 
        .Q(n105) );
  AOI220 U55 ( .A(i_data_lwM[28]), .B(n1), .C(i_data_lwW[28]), .D(n10), .Q(
        n103) );
  AOI220 U56 ( .A(i_data_rs[29]), .B(n5), .C(i_data_writeres[29]), .D(n7), .Q(
        n108) );
  AOI220 U57 ( .A(i_data_lwM[29]), .B(n1), .C(i_data_lwW[29]), .D(n9), .Q(n106) );
  AOI220 U58 ( .A(i_data_rs[30]), .B(n5), .C(i_data_writeres[30]), .D(n112), 
        .Q(n111) );
  AOI220 U59 ( .A(i_data_lwM[30]), .B(n1), .C(i_data_lwW[30]), .D(n10), .Q(
        n109) );
  AOI220 U60 ( .A(i_data_rs[25]), .B(n5), .C(i_data_writeres[25]), .D(n7), .Q(
        n96) );
  AOI220 U61 ( .A(i_data_lwM[25]), .B(n1), .C(i_data_lwW[25]), .D(n9), .Q(n94)
         );
  AOI220 U62 ( .A(i_data_rs[24]), .B(n5), .C(i_data_writeres[24]), .D(n112), 
        .Q(n93) );
  AOI220 U63 ( .A(i_data_lwM[24]), .B(n1), .C(i_data_lwW[24]), .D(n10), .Q(n91) );
  AOI220 U64 ( .A(i_data_rs[26]), .B(n5), .C(i_data_writeres[26]), .D(n112), 
        .Q(n99) );
  AOI220 U65 ( .A(i_data_lwM[26]), .B(n1), .C(i_data_lwW[26]), .D(n10), .Q(n97) );
  BUF2 U66 ( .A(n3), .Q(n4) );
  XOR21 U67 ( .A(n17), .B(n11), .Q(n3) );
  BUF2 U68 ( .A(n112), .Q(n7) );
  BUF2 U69 ( .A(n114), .Q(n9) );
  BUF2 U70 ( .A(n114), .Q(n8) );
  BUF2 U71 ( .A(n112), .Q(n6) );
  INV3 U72 ( .A(n14), .Q(n113) );
  NAND31 U73 ( .A(n69), .B(n68), .C(n67), .Q(o_data_alusra[16]) );
  AOI221 U74 ( .A(i_data_rs[16]), .B(n5), .C(i_data_writeres[16]), .D(n112), 
        .Q(n69) );
  NAND31 U75 ( .A(n72), .B(n71), .C(n70), .Q(o_data_alusra[17]) );
  AOI221 U76 ( .A(i_data_lwM[17]), .B(n1), .C(i_data_lwW[17]), .D(n9), .Q(n70)
         );
  AOI221 U77 ( .A(i_data_rs[17]), .B(n5), .C(i_data_writeres[17]), .D(n7), .Q(
        n72) );
  NAND31 U78 ( .A(n75), .B(n74), .C(n73), .Q(o_data_alusra[18]) );
  INV3 U79 ( .A(n12), .Q(n112) );
  AOI221 U80 ( .A(i_data_rs[4]), .B(n4), .C(i_data_writeres[4]), .D(n6), .Q(
        n33) );
  AOI221 U81 ( .A(i_data_rs[7]), .B(n4), .C(i_data_writeres[7]), .D(n6), .Q(
        n42) );
  AOI221 U82 ( .A(i_data_rs[0]), .B(n4), .C(i_data_writeres[0]), .D(n6), .Q(
        n21) );
  AOI221 U83 ( .A(i_data_rs[3]), .B(n4), .C(i_data_writeres[3]), .D(n6), .Q(
        n30) );
  AOI221 U84 ( .A(i_data_rs[1]), .B(n4), .C(i_data_writeres[1]), .D(n6), .Q(
        n24) );
  NAND31 U85 ( .A(n81), .B(n80), .C(n79), .Q(o_data_alusra[20]) );
  NAND31 U86 ( .A(n78), .B(n77), .C(n76), .Q(o_data_alusra[19]) );
  NAND31 U87 ( .A(n90), .B(n89), .C(n88), .Q(o_data_alusra[23]) );
  AOI221 U88 ( .A(i_data_rs[6]), .B(n4), .C(i_data_writeres[6]), .D(n6), .Q(
        n39) );
  AOI221 U89 ( .A(i_data_rs[2]), .B(n4), .C(i_data_writeres[2]), .D(n6), .Q(
        n27) );
  AOI221 U90 ( .A(i_data_rs[5]), .B(n4), .C(i_data_writeres[5]), .D(n6), .Q(
        n36) );
  NAND31 U91 ( .A(n54), .B(n53), .C(n52), .Q(o_data_alusra[11]) );
  NAND31 U92 ( .A(n57), .B(n56), .C(n55), .Q(o_data_alusra[12]) );
  NAND31 U93 ( .A(n60), .B(n59), .C(n58), .Q(o_data_alusra[13]) );
  NAND31 U94 ( .A(n63), .B(n62), .C(n61), .Q(o_data_alusra[14]) );
  NAND31 U95 ( .A(n66), .B(n65), .C(n64), .Q(o_data_alusra[15]) );
  NAND31 U96 ( .A(n102), .B(n101), .C(n100), .Q(o_data_alusra[27]) );
  NAND31 U97 ( .A(n105), .B(n104), .C(n103), .Q(o_data_alusra[28]) );
  NAND31 U98 ( .A(n111), .B(n110), .C(n109), .Q(o_data_alusra[30]) );
  NAND31 U99 ( .A(n96), .B(n95), .C(n94), .Q(o_data_alusra[25]) );
  NAND31 U100 ( .A(n99), .B(n98), .C(n97), .Q(o_data_alusra[26]) );
  NAND31 U101 ( .A(n51), .B(n50), .C(n49), .Q(o_data_alusra[10]) );
  AOI221 U102 ( .A(i_data_rs[10]), .B(n4), .C(i_data_writeres[10]), .D(n6), 
        .Q(n51) );
  NAND31 U103 ( .A(n87), .B(n86), .C(n85), .Q(o_data_alusra[22]) );
  NAND31 U104 ( .A(n93), .B(n92), .C(n91), .Q(o_data_alusra[24]) );
  NAND31 U105 ( .A(n45), .B(n44), .C(n43), .Q(o_data_alusra[8]) );
  AOI221 U106 ( .A(i_data_rs[8]), .B(n4), .C(i_data_writeres[8]), .D(n6), .Q(
        n45) );
  NAND31 U107 ( .A(n48), .B(n47), .C(n46), .Q(o_data_alusra[9]) );
  AOI221 U108 ( .A(i_data_rs[9]), .B(n4), .C(i_data_writeres[9]), .D(n6), .Q(
        n48) );
  NAND31 U109 ( .A(n84), .B(n83), .C(n82), .Q(o_data_alusra[21]) );
  NAND31 U110 ( .A(n108), .B(n107), .C(n106), .Q(o_data_alusra[29]) );
  NAND31 U111 ( .A(n117), .B(n116), .C(n115), .Q(o_data_alusra[31]) );
  CLKIN3 U112 ( .A(i_con_fa[1]), .Q(n17) );
  CLKIN3 U113 ( .A(i_con_fa[2]), .Q(n13) );
  NAND22 U114 ( .A(n13), .B(n15), .Q(n11) );
  NAND22 U115 ( .A(i_data_alures[0]), .B(n2), .Q(n20) );
  NAND22 U116 ( .A(i_data_alures[1]), .B(n2), .Q(n23) );
  NAND22 U117 ( .A(i_data_alures[2]), .B(n2), .Q(n26) );
  NAND22 U118 ( .A(i_data_alures[3]), .B(n2), .Q(n29) );
  NAND33 U119 ( .A(n30), .B(n29), .C(n28), .Q(o_data_alusra[3]) );
  NAND22 U120 ( .A(i_data_alures[4]), .B(n2), .Q(n32) );
  NAND33 U121 ( .A(n33), .B(n32), .C(n31), .Q(o_data_alusra[4]) );
  NAND22 U122 ( .A(i_data_alures[5]), .B(n2), .Q(n35) );
  NAND22 U123 ( .A(i_data_alures[6]), .B(n2), .Q(n38) );
  NAND22 U124 ( .A(i_data_alures[7]), .B(n2), .Q(n41) );
  NAND33 U125 ( .A(n42), .B(n41), .C(n40), .Q(o_data_alusra[7]) );
  NAND22 U126 ( .A(i_data_alures[8]), .B(n2), .Q(n44) );
  NAND22 U127 ( .A(i_data_alures[9]), .B(n2), .Q(n47) );
  NAND22 U128 ( .A(i_data_alures[10]), .B(n2), .Q(n50) );
  NAND22 U129 ( .A(i_data_alures[11]), .B(n2), .Q(n53) );
  NAND22 U130 ( .A(i_data_alures[12]), .B(n2), .Q(n56) );
  NAND22 U131 ( .A(i_data_alures[13]), .B(n2), .Q(n59) );
  NAND22 U132 ( .A(i_data_alures[14]), .B(n2), .Q(n62) );
  NAND22 U133 ( .A(i_data_alures[15]), .B(n2), .Q(n65) );
  NAND22 U134 ( .A(i_data_alures[16]), .B(n113), .Q(n68) );
  NAND22 U135 ( .A(i_data_alures[17]), .B(n113), .Q(n71) );
  NAND22 U136 ( .A(i_data_alures[18]), .B(n113), .Q(n74) );
  NAND22 U137 ( .A(i_data_alures[19]), .B(n2), .Q(n77) );
  NAND22 U138 ( .A(i_data_alures[20]), .B(n2), .Q(n80) );
  NAND22 U139 ( .A(i_data_alures[21]), .B(n2), .Q(n83) );
  NAND22 U140 ( .A(i_data_alures[22]), .B(n2), .Q(n86) );
  NAND22 U141 ( .A(i_data_alures[23]), .B(n2), .Q(n89) );
  NAND22 U142 ( .A(i_data_alures[24]), .B(n2), .Q(n92) );
  NAND22 U143 ( .A(i_data_alures[25]), .B(n2), .Q(n95) );
  NAND22 U144 ( .A(i_data_alures[26]), .B(n2), .Q(n98) );
  NAND22 U145 ( .A(i_data_alures[27]), .B(n2), .Q(n101) );
  NAND22 U146 ( .A(i_data_alures[28]), .B(n2), .Q(n104) );
  NAND22 U147 ( .A(i_data_alures[29]), .B(n2), .Q(n107) );
  NAND22 U148 ( .A(i_data_alures[30]), .B(n2), .Q(n110) );
  NAND22 U149 ( .A(i_data_alures[31]), .B(n2), .Q(n116) );
endmodule


module E_fbmux5 ( i_data_rt, i_data_alures, i_data_writeres, i_data_lwM, 
        i_data_lwW, i_con_fb, o_data_alusrb );
  input [31:0] i_data_rt;
  input [31:0] i_data_alures;
  input [31:0] i_data_writeres;
  input [31:0] i_data_lwM;
  input [31:0] i_data_lwW;
  input [2:0] i_con_fb;
  output [31:0] o_data_alusrb;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118;

  NAND22 U1 ( .A(n15), .B(n5), .Q(n14) );
  CLKIN3 U2 ( .A(n14), .Q(n113) );
  CLKIN2 U3 ( .A(n14), .Q(n2) );
  XOR21 U4 ( .A(n17), .B(n11), .Q(n8) );
  BUF6 U5 ( .A(n8), .Q(n9) );
  BUF6 U6 ( .A(n114), .Q(n10) );
  NAND22 U7 ( .A(n71), .B(n7), .Q(o_data_alusrb[17]) );
  INV6 U8 ( .A(i_con_fb[0]), .Q(n15) );
  AOI221 U9 ( .A(i_data_rt[17]), .B(n9), .C(i_data_writeres[17]), .D(n112), 
        .Q(n72) );
  INV3 U10 ( .A(n12), .Q(n1) );
  INV3 U11 ( .A(n12), .Q(n112) );
  CLKIN6 U12 ( .A(i_con_fb[2]), .Q(n13) );
  NAND30 U13 ( .A(i_con_fb[0]), .B(n13), .C(n17), .Q(n12) );
  NAND31 U14 ( .A(n69), .B(n68), .C(n67), .Q(o_data_alusrb[16]) );
  AOI220 U15 ( .A(i_data_writeres[16]), .B(n112), .C(i_data_alures[16]), .D(
        n113), .Q(n69) );
  NAND31 U16 ( .A(n48), .B(n47), .C(n46), .Q(o_data_alusrb[9]) );
  NAND20 U17 ( .A(i_data_alures[17]), .B(n113), .Q(n71) );
  CLKIN3 U18 ( .A(n16), .Q(n115) );
  INV6 U19 ( .A(n16), .Q(n3) );
  NAND30 U20 ( .A(i_con_fb[2]), .B(n15), .C(n17), .Q(n16) );
  NAND20 U21 ( .A(n13), .B(i_con_fb[1]), .Q(n4) );
  INV2 U22 ( .A(n4), .Q(n5) );
  NAND22 U23 ( .A(n72), .B(n70), .Q(n6) );
  INV3 U24 ( .A(n6), .Q(n7) );
  AOI220 U25 ( .A(i_data_lwM[17]), .B(n115), .C(i_data_lwW[17]), .D(n10), .Q(
        n70) );
  CLKIN6 U26 ( .A(i_con_fb[1]), .Q(n17) );
  AOI220 U27 ( .A(i_data_rt[8]), .B(n9), .C(i_data_writeres[8]), .D(n1), .Q(
        n45) );
  AOI220 U28 ( .A(i_data_lwM[8]), .B(n3), .C(i_data_lwW[8]), .D(n10), .Q(n43)
         );
  AOI220 U29 ( .A(i_data_rt[18]), .B(n9), .C(i_data_writeres[18]), .D(n112), 
        .Q(n75) );
  AOI220 U30 ( .A(i_data_lwM[18]), .B(n115), .C(i_data_lwW[18]), .D(n10), .Q(
        n73) );
  AOI220 U31 ( .A(i_data_rt[19]), .B(n9), .C(i_data_writeres[19]), .D(n1), .Q(
        n78) );
  AOI220 U32 ( .A(i_data_lwM[19]), .B(n115), .C(i_data_lwW[19]), .D(n10), .Q(
        n76) );
  AOI220 U33 ( .A(i_data_rt[20]), .B(n9), .C(i_data_writeres[20]), .D(n1), .Q(
        n81) );
  AOI220 U34 ( .A(i_data_lwM[20]), .B(n3), .C(i_data_lwW[20]), .D(n10), .Q(n79) );
  AOI220 U35 ( .A(i_data_rt[3]), .B(n9), .C(i_data_writeres[3]), .D(n1), .Q(
        n30) );
  AOI220 U36 ( .A(i_data_lwM[3]), .B(n3), .C(i_data_lwW[3]), .D(n10), .Q(n28)
         );
  AOI220 U37 ( .A(i_data_rt[4]), .B(n9), .C(i_data_writeres[4]), .D(n1), .Q(
        n33) );
  AOI220 U38 ( .A(i_data_lwM[4]), .B(n3), .C(i_data_lwW[4]), .D(n10), .Q(n31)
         );
  AOI220 U39 ( .A(i_data_rt[21]), .B(n9), .C(i_data_writeres[21]), .D(n1), .Q(
        n84) );
  AOI220 U40 ( .A(i_data_lwM[21]), .B(n3), .C(i_data_lwW[21]), .D(n10), .Q(n82) );
  AOI220 U41 ( .A(i_data_rt[22]), .B(n9), .C(i_data_writeres[22]), .D(n1), .Q(
        n87) );
  AOI220 U42 ( .A(i_data_lwM[22]), .B(n3), .C(i_data_lwW[22]), .D(n10), .Q(n85) );
  AOI220 U43 ( .A(i_data_rt[0]), .B(n9), .C(i_data_writeres[0]), .D(n1), .Q(
        n21) );
  AOI220 U44 ( .A(i_data_lwM[0]), .B(n3), .C(i_data_lwW[0]), .D(n10), .Q(n19)
         );
  AOI220 U45 ( .A(i_data_rt[1]), .B(n9), .C(i_data_writeres[1]), .D(n1), .Q(
        n24) );
  AOI220 U46 ( .A(i_data_lwM[1]), .B(n3), .C(i_data_lwW[1]), .D(n10), .Q(n22)
         );
  AOI220 U47 ( .A(i_data_rt[9]), .B(n9), .C(i_data_writeres[9]), .D(n1), .Q(
        n48) );
  AOI220 U48 ( .A(i_data_lwM[9]), .B(n3), .C(i_data_lwW[9]), .D(n10), .Q(n46)
         );
  AOI220 U49 ( .A(i_data_rt[2]), .B(n9), .C(i_data_writeres[2]), .D(n1), .Q(
        n27) );
  AOI220 U50 ( .A(i_data_lwM[2]), .B(n3), .C(i_data_lwW[2]), .D(n10), .Q(n25)
         );
  AOI220 U51 ( .A(i_data_rt[10]), .B(n9), .C(i_data_writeres[10]), .D(n1), .Q(
        n51) );
  AOI220 U52 ( .A(i_data_lwM[10]), .B(n3), .C(i_data_lwW[10]), .D(n10), .Q(n49) );
  AOI220 U53 ( .A(i_data_rt[11]), .B(n9), .C(i_data_writeres[11]), .D(n1), .Q(
        n54) );
  AOI220 U54 ( .A(i_data_lwM[11]), .B(n3), .C(i_data_lwW[11]), .D(n10), .Q(n52) );
  CLKIN3 U55 ( .A(n18), .Q(n114) );
  NAND30 U56 ( .A(i_con_fb[2]), .B(i_con_fb[0]), .C(n17), .Q(n18) );
  AOI220 U57 ( .A(i_data_rt[5]), .B(n9), .C(i_data_writeres[5]), .D(n1), .Q(
        n36) );
  AOI220 U58 ( .A(i_data_lwM[5]), .B(n3), .C(i_data_lwW[5]), .D(n10), .Q(n34)
         );
  AOI220 U59 ( .A(i_data_rt[6]), .B(n9), .C(i_data_writeres[6]), .D(n1), .Q(
        n39) );
  AOI220 U60 ( .A(i_data_lwM[6]), .B(n3), .C(i_data_lwW[6]), .D(n10), .Q(n37)
         );
  AOI220 U61 ( .A(i_data_rt[7]), .B(n9), .C(i_data_writeres[7]), .D(n1), .Q(
        n42) );
  AOI220 U62 ( .A(i_data_lwM[7]), .B(n3), .C(i_data_lwW[7]), .D(n10), .Q(n40)
         );
  AOI220 U63 ( .A(i_data_rt[12]), .B(n9), .C(i_data_writeres[12]), .D(n1), .Q(
        n57) );
  AOI220 U64 ( .A(i_data_lwM[12]), .B(n3), .C(i_data_lwW[12]), .D(n10), .Q(n55) );
  AOI220 U65 ( .A(i_data_rt[13]), .B(n9), .C(i_data_writeres[13]), .D(n1), .Q(
        n60) );
  AOI220 U66 ( .A(i_data_lwM[13]), .B(n3), .C(i_data_lwW[13]), .D(n10), .Q(n58) );
  AOI220 U67 ( .A(i_data_rt[14]), .B(n9), .C(i_data_writeres[14]), .D(n1), .Q(
        n63) );
  AOI220 U68 ( .A(i_data_lwM[14]), .B(n3), .C(i_data_lwW[14]), .D(n10), .Q(n61) );
  AOI220 U69 ( .A(i_data_rt[15]), .B(n9), .C(i_data_writeres[15]), .D(n1), .Q(
        n66) );
  AOI220 U70 ( .A(i_data_lwM[15]), .B(n3), .C(i_data_lwW[15]), .D(n10), .Q(n64) );
  AOI220 U71 ( .A(i_data_rt[23]), .B(n9), .C(i_data_writeres[23]), .D(n1), .Q(
        n90) );
  AOI220 U72 ( .A(i_data_lwM[23]), .B(n3), .C(i_data_lwW[23]), .D(n10), .Q(n88) );
  AOI220 U73 ( .A(i_data_rt[24]), .B(n9), .C(i_data_writeres[24]), .D(n1), .Q(
        n93) );
  AOI220 U74 ( .A(i_data_lwM[24]), .B(n3), .C(i_data_lwW[24]), .D(n10), .Q(n91) );
  AOI220 U75 ( .A(i_data_rt[25]), .B(n9), .C(i_data_writeres[25]), .D(n1), .Q(
        n96) );
  AOI220 U76 ( .A(i_data_lwM[25]), .B(n3), .C(i_data_lwW[25]), .D(n10), .Q(n94) );
  AOI220 U77 ( .A(i_data_rt[26]), .B(n9), .C(i_data_writeres[26]), .D(n1), .Q(
        n99) );
  AOI220 U78 ( .A(i_data_lwM[26]), .B(n3), .C(i_data_lwW[26]), .D(n10), .Q(n97) );
  AOI220 U79 ( .A(i_data_rt[27]), .B(n9), .C(i_data_writeres[27]), .D(n1), .Q(
        n102) );
  AOI220 U80 ( .A(i_data_lwM[27]), .B(n3), .C(i_data_lwW[27]), .D(n10), .Q(
        n100) );
  AOI220 U81 ( .A(i_data_rt[28]), .B(n9), .C(i_data_writeres[28]), .D(n1), .Q(
        n105) );
  AOI220 U82 ( .A(i_data_lwM[28]), .B(n3), .C(i_data_lwW[28]), .D(n10), .Q(
        n103) );
  AOI220 U83 ( .A(i_data_rt[29]), .B(n9), .C(i_data_writeres[29]), .D(n1), .Q(
        n108) );
  AOI220 U84 ( .A(i_data_lwM[29]), .B(n3), .C(i_data_lwW[29]), .D(n10), .Q(
        n106) );
  AOI220 U85 ( .A(i_data_rt[30]), .B(n9), .C(i_data_writeres[30]), .D(n1), .Q(
        n111) );
  AOI220 U86 ( .A(i_data_lwM[30]), .B(n3), .C(i_data_lwW[30]), .D(n10), .Q(
        n109) );
  AOI220 U87 ( .A(i_data_rt[31]), .B(n9), .C(i_data_writeres[31]), .D(n1), .Q(
        n118) );
  AOI220 U88 ( .A(i_data_lwM[31]), .B(n3), .C(i_data_lwW[31]), .D(n10), .Q(
        n116) );
  NAND22 U89 ( .A(n13), .B(n15), .Q(n11) );
  NAND31 U90 ( .A(n75), .B(n74), .C(n73), .Q(o_data_alusrb[18]) );
  AOI221 U91 ( .A(i_data_lwM[16]), .B(n115), .C(i_data_lwW[16]), .D(n10), .Q(
        n68) );
  NAND22 U92 ( .A(i_data_rt[16]), .B(n9), .Q(n67) );
  NAND31 U93 ( .A(n21), .B(n20), .C(n19), .Q(o_data_alusrb[0]) );
  NAND31 U94 ( .A(n24), .B(n23), .C(n22), .Q(o_data_alusrb[1]) );
  NAND31 U95 ( .A(n78), .B(n77), .C(n76), .Q(o_data_alusrb[19]) );
  NAND31 U96 ( .A(n81), .B(n80), .C(n79), .Q(o_data_alusrb[20]) );
  NAND31 U97 ( .A(n84), .B(n83), .C(n82), .Q(o_data_alusrb[21]) );
  NAND31 U98 ( .A(n27), .B(n26), .C(n25), .Q(o_data_alusrb[2]) );
  NAND31 U99 ( .A(n30), .B(n29), .C(n28), .Q(o_data_alusrb[3]) );
  NAND31 U100 ( .A(n45), .B(n44), .C(n43), .Q(o_data_alusrb[8]) );
  NAND31 U101 ( .A(n51), .B(n50), .C(n49), .Q(o_data_alusrb[10]) );
  NAND31 U102 ( .A(n54), .B(n53), .C(n52), .Q(o_data_alusrb[11]) );
  NAND31 U103 ( .A(n87), .B(n86), .C(n85), .Q(o_data_alusrb[22]) );
  NAND31 U104 ( .A(n90), .B(n89), .C(n88), .Q(o_data_alusrb[23]) );
  NAND31 U105 ( .A(n93), .B(n92), .C(n91), .Q(o_data_alusrb[24]) );
  NAND31 U106 ( .A(n102), .B(n101), .C(n100), .Q(o_data_alusrb[27]) );
  NAND31 U107 ( .A(n118), .B(n117), .C(n116), .Q(o_data_alusrb[31]) );
  NAND31 U108 ( .A(n33), .B(n32), .C(n31), .Q(o_data_alusrb[4]) );
  NAND31 U109 ( .A(n36), .B(n35), .C(n34), .Q(o_data_alusrb[5]) );
  NAND31 U110 ( .A(n42), .B(n41), .C(n40), .Q(o_data_alusrb[7]) );
  NAND31 U111 ( .A(n66), .B(n65), .C(n64), .Q(o_data_alusrb[15]) );
  NAND31 U112 ( .A(n96), .B(n95), .C(n94), .Q(o_data_alusrb[25]) );
  NAND31 U113 ( .A(n99), .B(n98), .C(n97), .Q(o_data_alusrb[26]) );
  NAND31 U114 ( .A(n105), .B(n104), .C(n103), .Q(o_data_alusrb[28]) );
  NAND31 U115 ( .A(n108), .B(n107), .C(n106), .Q(o_data_alusrb[29]) );
  NAND31 U116 ( .A(n111), .B(n110), .C(n109), .Q(o_data_alusrb[30]) );
  NAND31 U117 ( .A(n39), .B(n38), .C(n37), .Q(o_data_alusrb[6]) );
  NAND31 U118 ( .A(n57), .B(n56), .C(n55), .Q(o_data_alusrb[12]) );
  NAND31 U119 ( .A(n60), .B(n59), .C(n58), .Q(o_data_alusrb[13]) );
  NAND31 U120 ( .A(n63), .B(n62), .C(n61), .Q(o_data_alusrb[14]) );
  NAND22 U121 ( .A(i_data_alures[0]), .B(n2), .Q(n20) );
  NAND22 U122 ( .A(i_data_alures[1]), .B(n2), .Q(n23) );
  NAND22 U123 ( .A(i_data_alures[2]), .B(n113), .Q(n26) );
  NAND22 U124 ( .A(i_data_alures[3]), .B(n2), .Q(n29) );
  NAND22 U125 ( .A(i_data_alures[4]), .B(n113), .Q(n32) );
  NAND22 U126 ( .A(i_data_alures[5]), .B(n2), .Q(n35) );
  NAND22 U127 ( .A(i_data_alures[6]), .B(n2), .Q(n38) );
  NAND22 U128 ( .A(i_data_alures[7]), .B(n113), .Q(n41) );
  NAND22 U129 ( .A(i_data_alures[8]), .B(n113), .Q(n44) );
  NAND22 U130 ( .A(i_data_alures[9]), .B(n2), .Q(n47) );
  NAND22 U131 ( .A(i_data_alures[10]), .B(n113), .Q(n50) );
  NAND22 U132 ( .A(i_data_alures[11]), .B(n113), .Q(n53) );
  NAND22 U133 ( .A(i_data_alures[12]), .B(n2), .Q(n56) );
  NAND22 U134 ( .A(i_data_alures[13]), .B(n2), .Q(n59) );
  NAND22 U135 ( .A(i_data_alures[14]), .B(n2), .Q(n62) );
  NAND22 U136 ( .A(i_data_alures[15]), .B(n2), .Q(n65) );
  NAND22 U137 ( .A(i_data_alures[18]), .B(n113), .Q(n74) );
  NAND22 U138 ( .A(i_data_alures[19]), .B(n2), .Q(n77) );
  NAND22 U139 ( .A(i_data_alures[20]), .B(n113), .Q(n80) );
  NAND22 U140 ( .A(i_data_alures[21]), .B(n2), .Q(n83) );
  NAND22 U141 ( .A(i_data_alures[22]), .B(n2), .Q(n86) );
  NAND22 U142 ( .A(i_data_alures[23]), .B(n113), .Q(n89) );
  NAND22 U143 ( .A(i_data_alures[24]), .B(n2), .Q(n92) );
  NAND22 U144 ( .A(i_data_alures[25]), .B(n113), .Q(n95) );
  NAND22 U145 ( .A(i_data_alures[26]), .B(n2), .Q(n98) );
  NAND22 U146 ( .A(i_data_alures[27]), .B(n113), .Q(n101) );
  NAND22 U147 ( .A(i_data_alures[28]), .B(n2), .Q(n104) );
  NAND22 U148 ( .A(i_data_alures[29]), .B(n113), .Q(n107) );
  NAND22 U149 ( .A(i_data_alures[30]), .B(n2), .Q(n110) );
  NAND22 U150 ( .A(i_data_alures[31]), .B(n2), .Q(n117) );
endmodule


module E_alubmux ( i_data_fb, i_data_imm, i_con_imm, o_data_alub );
  input [31:0] i_data_fb;
  input [31:0] i_data_imm;
  output [31:0] o_data_alub;
  input i_con_imm;
  wire   n1, n2, n3;

  NAND22 U1 ( .A(n2), .B(n3), .Q(o_data_alub[9]) );
  NAND22 U2 ( .A(i_data_fb[9]), .B(n1), .Q(n2) );
  MUX24 U3 ( .A(i_data_fb[16]), .B(i_data_imm[16]), .S(i_con_imm), .Q(
        o_data_alub[16]) );
  NAND22 U4 ( .A(i_data_imm[9]), .B(i_con_imm), .Q(n3) );
  INV2 U5 ( .A(i_con_imm), .Q(n1) );
  MUX21 U6 ( .A(i_data_fb[20]), .B(i_data_imm[20]), .S(i_con_imm), .Q(
        o_data_alub[20]) );
  MUX22 U7 ( .A(i_data_fb[17]), .B(i_data_imm[17]), .S(i_con_imm), .Q(
        o_data_alub[17]) );
  MUX21 U8 ( .A(i_data_fb[21]), .B(i_data_imm[21]), .S(i_con_imm), .Q(
        o_data_alub[21]) );
  MUX21 U9 ( .A(i_data_fb[22]), .B(i_data_imm[22]), .S(i_con_imm), .Q(
        o_data_alub[22]) );
  MUX21 U10 ( .A(i_data_fb[24]), .B(i_data_imm[24]), .S(i_con_imm), .Q(
        o_data_alub[24]) );
  MUX21 U11 ( .A(i_data_fb[25]), .B(i_data_imm[25]), .S(i_con_imm), .Q(
        o_data_alub[25]) );
  MUX21 U12 ( .A(i_data_fb[23]), .B(i_data_imm[23]), .S(i_con_imm), .Q(
        o_data_alub[23]) );
  MUX21 U13 ( .A(i_data_fb[15]), .B(i_data_imm[15]), .S(i_con_imm), .Q(
        o_data_alub[15]) );
  MUX22 U14 ( .A(i_data_fb[18]), .B(i_data_imm[18]), .S(i_con_imm), .Q(
        o_data_alub[18]) );
  MUX22 U15 ( .A(i_data_fb[0]), .B(i_data_imm[0]), .S(i_con_imm), .Q(
        o_data_alub[0]) );
  MUX22 U16 ( .A(i_data_fb[1]), .B(i_data_imm[1]), .S(i_con_imm), .Q(
        o_data_alub[1]) );
  MUX22 U17 ( .A(i_data_fb[19]), .B(i_data_imm[19]), .S(i_con_imm), .Q(
        o_data_alub[19]) );
  MUX22 U18 ( .A(i_data_fb[8]), .B(i_data_imm[8]), .S(i_con_imm), .Q(
        o_data_alub[8]) );
  MUX22 U19 ( .A(i_data_fb[11]), .B(i_data_imm[11]), .S(i_con_imm), .Q(
        o_data_alub[11]) );
  MUX22 U20 ( .A(i_data_fb[10]), .B(i_data_imm[10]), .S(i_con_imm), .Q(
        o_data_alub[10]) );
  MUX22 U21 ( .A(i_data_fb[3]), .B(i_data_imm[3]), .S(i_con_imm), .Q(
        o_data_alub[3]) );
  MUX22 U22 ( .A(i_data_fb[2]), .B(i_data_imm[2]), .S(i_con_imm), .Q(
        o_data_alub[2]) );
  MUX22 U23 ( .A(i_data_fb[7]), .B(i_data_imm[7]), .S(i_con_imm), .Q(
        o_data_alub[7]) );
  MUX22 U24 ( .A(i_data_fb[12]), .B(i_data_imm[12]), .S(i_con_imm), .Q(
        o_data_alub[12]) );
  MUX22 U25 ( .A(i_data_fb[14]), .B(i_data_imm[14]), .S(i_con_imm), .Q(
        o_data_alub[14]) );
  MUX22 U26 ( .A(i_data_fb[13]), .B(i_data_imm[13]), .S(i_con_imm), .Q(
        o_data_alub[13]) );
  MUX22 U27 ( .A(i_data_fb[4]), .B(i_data_imm[4]), .S(i_con_imm), .Q(
        o_data_alub[4]) );
  MUX22 U28 ( .A(i_data_fb[6]), .B(i_data_imm[6]), .S(i_con_imm), .Q(
        o_data_alub[6]) );
  MUX22 U29 ( .A(i_data_fb[5]), .B(i_data_imm[5]), .S(i_con_imm), .Q(
        o_data_alub[5]) );
  MUX22 U30 ( .A(i_data_fb[28]), .B(i_data_imm[28]), .S(i_con_imm), .Q(
        o_data_alub[28]) );
  MUX22 U31 ( .A(i_data_fb[26]), .B(i_data_imm[26]), .S(i_con_imm), .Q(
        o_data_alub[26]) );
  MUX22 U32 ( .A(i_data_fb[27]), .B(i_data_imm[27]), .S(i_con_imm), .Q(
        o_data_alub[27]) );
  MUX22 U33 ( .A(i_data_fb[30]), .B(i_data_imm[30]), .S(i_con_imm), .Q(
        o_data_alub[30]) );
  MUX22 U34 ( .A(i_data_fb[29]), .B(i_data_imm[29]), .S(i_con_imm), .Q(
        o_data_alub[29]) );
  MUX22 U35 ( .A(i_data_fb[31]), .B(i_data_imm[31]), .S(i_con_imm), .Q(
        o_data_alub[31]) );
endmodule


module E_rdmux ( i_data_rtE, i_data_rdE, i_con_regdst, i_con_aluPC4, 
        o_data_writeE );
  input [4:0] i_data_rtE;
  input [4:0] i_data_rdE;
  output [4:0] o_data_writeE;
  input i_con_regdst, i_con_aluPC4;
  wire   n7, n8, n9, n10, n11, n1, n2, n3, n4, n5, n6;

  OAI2111 U2 ( .A(i_con_regdst), .B(n5), .C(n6), .D(n11), .Q(o_data_writeE[0])
         );
  INV3 U3 ( .A(i_data_rtE[0]), .Q(n5) );
  NAND22 U4 ( .A(i_data_rdE[0]), .B(i_con_regdst), .Q(n11) );
  OAI2111 U5 ( .A(i_con_regdst), .B(n4), .C(n6), .D(n10), .Q(o_data_writeE[1])
         );
  INV3 U6 ( .A(i_data_rtE[1]), .Q(n4) );
  NAND22 U7 ( .A(i_data_rdE[1]), .B(i_con_regdst), .Q(n10) );
  OAI2111 U8 ( .A(i_con_regdst), .B(n3), .C(n6), .D(n9), .Q(o_data_writeE[2])
         );
  INV3 U9 ( .A(i_data_rtE[2]), .Q(n3) );
  NAND22 U10 ( .A(i_data_rdE[2]), .B(i_con_regdst), .Q(n9) );
  OAI2111 U11 ( .A(i_con_regdst), .B(n2), .C(n6), .D(n8), .Q(o_data_writeE[3])
         );
  INV3 U12 ( .A(i_data_rtE[3]), .Q(n2) );
  NAND22 U13 ( .A(i_data_rdE[3]), .B(i_con_regdst), .Q(n8) );
  OAI2111 U14 ( .A(i_con_regdst), .B(n1), .C(n6), .D(n7), .Q(o_data_writeE[4])
         );
  INV3 U15 ( .A(i_data_rtE[4]), .Q(n1) );
  NAND22 U16 ( .A(i_data_rdE[4]), .B(i_con_regdst), .Q(n7) );
  INV3 U17 ( .A(i_con_aluPC4), .Q(n6) );
endmodule


module D_compare_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49;

  INV0 U1 ( .A(B[0]), .Q(n4) );
  INV3 U2 ( .A(n5), .Q(EQ) );
  INV3 U3 ( .A(n28), .Q(n2) );
  INV3 U4 ( .A(A[1]), .Q(n3) );
  NAND20 U5 ( .A(n6), .B(n7), .Q(n5) );
  NOR40 U6 ( .A(n8), .B(n9), .C(n10), .D(n11), .Q(n7) );
  NAND40 U7 ( .A(n12), .B(n13), .C(n14), .D(n15), .Q(n11) );
  XNR20 U8 ( .A(B[11]), .B(A[11]), .Q(n15) );
  XNR20 U9 ( .A(B[12]), .B(A[12]), .Q(n14) );
  XNR20 U10 ( .A(B[13]), .B(A[13]), .Q(n13) );
  XNR20 U11 ( .A(B[14]), .B(A[14]), .Q(n12) );
  NAND40 U12 ( .A(n16), .B(n17), .C(n18), .D(n19), .Q(n10) );
  XNR20 U13 ( .A(B[7]), .B(A[7]), .Q(n19) );
  XNR20 U14 ( .A(B[8]), .B(A[8]), .Q(n18) );
  XNR20 U15 ( .A(B[9]), .B(A[9]), .Q(n17) );
  XNR20 U16 ( .A(B[10]), .B(A[10]), .Q(n16) );
  NAND40 U17 ( .A(n20), .B(n21), .C(n22), .D(n23), .Q(n9) );
  XNR20 U18 ( .A(B[3]), .B(A[3]), .Q(n23) );
  XNR20 U19 ( .A(B[4]), .B(A[4]), .Q(n22) );
  XNR20 U20 ( .A(B[5]), .B(A[5]), .Q(n21) );
  XNR20 U21 ( .A(B[6]), .B(A[6]), .Q(n20) );
  NAND40 U22 ( .A(n24), .B(n25), .C(n2), .D(n26), .Q(n8) );
  OAI220 U23 ( .A(n27), .B(n3), .C(B[1]), .D(n27), .Q(n26) );
  NOR20 U24 ( .A(n4), .B(A[0]), .Q(n27) );
  AOI220 U25 ( .A(n3), .B(n29), .C(n29), .D(B[1]), .Q(n28) );
  NAND20 U26 ( .A(A[0]), .B(n4), .Q(n29) );
  XNR20 U27 ( .A(B[31]), .B(A[31]), .Q(n25) );
  XNR20 U28 ( .A(B[2]), .B(A[2]), .Q(n24) );
  NOR40 U29 ( .A(n30), .B(n31), .C(n32), .D(n33), .Q(n6) );
  NAND40 U30 ( .A(n34), .B(n35), .C(n36), .D(n37), .Q(n33) );
  XNR20 U31 ( .A(B[27]), .B(A[27]), .Q(n37) );
  XNR20 U32 ( .A(B[28]), .B(A[28]), .Q(n36) );
  XNR20 U33 ( .A(B[29]), .B(A[29]), .Q(n35) );
  XNR20 U34 ( .A(B[30]), .B(A[30]), .Q(n34) );
  NAND40 U35 ( .A(n38), .B(n39), .C(n40), .D(n41), .Q(n32) );
  XNR20 U36 ( .A(B[23]), .B(A[23]), .Q(n41) );
  XNR20 U37 ( .A(B[24]), .B(A[24]), .Q(n40) );
  XNR20 U38 ( .A(B[25]), .B(A[25]), .Q(n39) );
  XNR20 U39 ( .A(B[26]), .B(A[26]), .Q(n38) );
  NAND40 U40 ( .A(n42), .B(n43), .C(n44), .D(n45), .Q(n31) );
  XNR20 U41 ( .A(B[19]), .B(A[19]), .Q(n45) );
  XNR20 U42 ( .A(B[20]), .B(A[20]), .Q(n44) );
  XNR20 U43 ( .A(B[21]), .B(A[21]), .Q(n43) );
  XNR20 U44 ( .A(B[22]), .B(A[22]), .Q(n42) );
  NAND40 U45 ( .A(n46), .B(n47), .C(n48), .D(n49), .Q(n30) );
  XNR20 U46 ( .A(B[15]), .B(A[15]), .Q(n49) );
  XNR20 U47 ( .A(B[16]), .B(A[16]), .Q(n48) );
  XNR20 U48 ( .A(B[17]), .B(A[17]), .Q(n47) );
  XNR20 U49 ( .A(B[18]), .B(A[18]), .Q(n46) );
endmodule


module D_compare ( o_con_ifbranch, i_data_rs, i_data_rt, i_con_bop );
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [2:0] i_con_bop;
  output o_con_ifbranch;
  wire   equal, n3, n7, n8, n9, n10, n1, n2, n4;

  OAI222 U3 ( .A(n7), .B(n2), .C(i_con_bop[2]), .D(n8), .Q(o_con_ifbranch) );
  D_compare_DW01_cmp6_0 eq_34 ( .A(i_data_rs), .B(i_data_rt), .TC(n3), .EQ(
        equal) );
  INV3 U2 ( .A(i_con_bop[2]), .Q(n2) );
  AOI311 U4 ( .A(i_con_bop[0]), .B(n4), .C(i_data_rs[31]), .D(n10), .Q(n7) );
  AOI221 U5 ( .A(n9), .B(i_con_bop[1]), .C(equal), .D(i_con_bop[0]), .Q(n8) );
  AOI2111 U6 ( .A(equal), .B(n4), .C(i_data_rs[31]), .D(i_con_bop[0]), .Q(n10)
         );
  AOI211 U7 ( .A(i_con_bop[0]), .B(n1), .C(equal), .Q(n9) );
  INV3 U8 ( .A(i_data_rs[31]), .Q(n1) );
  INV3 U9 ( .A(i_con_bop[1]), .Q(n4) );
  LOGIC0 U10 ( .Q(n3) );
endmodule


module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Efamux, i_con_Efbmux, 
        i_con_Ealuop, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread, 
        i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_bop, o_data_pc4, o_data_alures, o_data_rt, o_addr_regdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_addr_Erd, o_addr_Mrt, o_con_ifbranch );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [5:0] i_con_Ealuop;
  input [2:0] i_con_bop;
  output [31:0] o_data_pc4;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch;
  wire   n1;
  wire   [31:0] alu_o_data_AluRes;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;

  DFC3 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC3 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC3 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC3 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC3 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC3 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[31]) );
  DFC3 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[30]) );
  DFC3 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[29]) );
  DFC3 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[28]) );
  DFC3 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[27]) );
  DFC3 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[26]) );
  DFC3 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[25]) );
  DFC3 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[24]) );
  DFC3 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[23]) );
  DFC3 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[22]) );
  DFC3 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[21]) );
  DFC3 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[20]) );
  DFC3 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[19]) );
  DFC3 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[18]) );
  DFC3 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[17]) );
  DFC3 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[16]) );
  DFC3 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[15]) );
  DFC3 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[14]) );
  DFC3 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[13]) );
  DFC3 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[12]) );
  DFC3 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[11]) );
  DFC3 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[10]) );
  DFC3 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[9]) );
  DFC3 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[8]) );
  DFC3 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[7]) );
  DFC3 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[6]) );
  DFC3 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[5]) );
  DFC3 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[4]) );
  DFC3 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[3]) );
  DFC3 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[2]) );
  DFC3 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[1]) );
  DFC3 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[0]) );
  DFC3 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC3 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC3 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC3 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC3 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC3 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC3 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC3 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC3 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC3 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC3 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC3 pipe_alures_reg_15_ ( .D(alu_o_data_AluRes[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[15]) );
  DFC3 pipe_alures_reg_14_ ( .D(alu_o_data_AluRes[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[14]) );
  DFC3 pipe_alures_reg_13_ ( .D(alu_o_data_AluRes[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[13]) );
  DFC3 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC3 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC3 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC3 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC3 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC3 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC3 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC3 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC3 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC3 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC3 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC3 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC3 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC3 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC3 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC3 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC3 pipe_rt_reg_28_ ( .D(compare_i_data_rt[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[28]) );
  DFC3 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  DFC3 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC3 pipe_rt_reg_25_ ( .D(compare_i_data_rt[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[25]) );
  DFC3 pipe_rt_reg_24_ ( .D(compare_i_data_rt[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[24]) );
  DFC3 pipe_rt_reg_23_ ( .D(compare_i_data_rt[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[23]) );
  DFC3 pipe_rt_reg_22_ ( .D(compare_i_data_rt[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[22]) );
  DFC3 pipe_rt_reg_21_ ( .D(compare_i_data_rt[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[21]) );
  DFC3 pipe_rt_reg_20_ ( .D(compare_i_data_rt[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[20]) );
  DFC3 pipe_rt_reg_16_ ( .D(n1), .C(i_clk), .RN(i_nrst), .Q(o_data_rt[16]) );
  DFC3 pipe_rt_reg_15_ ( .D(compare_i_data_rt[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[15]) );
  DFC3 pipe_rt_reg_14_ ( .D(compare_i_data_rt[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[14]) );
  DFC3 pipe_rt_reg_13_ ( .D(compare_i_data_rt[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[13]) );
  DFC3 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC3 pipe_rt_reg_11_ ( .D(compare_i_data_rt[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[11]) );
  DFC3 pipe_rt_reg_10_ ( .D(compare_i_data_rt[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[10]) );
  DFC3 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC3 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC3 pipe_rt_reg_5_ ( .D(compare_i_data_rt[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[5]) );
  DFC3 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(compare_i_data_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[2]) );
  DFC3 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC3 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC3 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC3 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC3 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC3 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC3 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC3 pipe_con_Malupc8_reg ( .D(i_con_Malupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Malupc8) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  E_alu u_alu ( .o_data_AluRes(alu_o_data_AluRes), .i_data_A(compare_i_data_rs), .i_data_B(alu_i_data_B), .i_con_AluCtrl(alu_i_con_AluCtrl), .i_data_shamt(
        i_data_immext[10:6]) );
  E_alu_control u_alu_control ( .o_con_AluCtrl(alu_i_con_AluCtrl), 
        .i_con_AluOp(i_con_Ealuop), .i_con_FuncCode(i_data_immext[5:0]) );
  E_famux5 u_famux5 ( .i_data_rs(i_data_rs), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fa(i_con_Efamux), .o_data_alusra(
        compare_i_data_rs) );
  E_fbmux5 u_fbmux ( .i_data_rt(i_data_rt), .i_data_alures(i_data_FEalures), 
        .i_data_writeres(i_data_FMalures), .i_data_lwM(i_data_FMmemout), 
        .i_data_lwW(i_data_FWmemout), .i_con_fb(i_con_Efbmux), .o_data_alusrb(
        compare_i_data_rt) );
  E_alubmux u_alubmux ( .i_data_fb(compare_i_data_rt), .i_data_imm(
        i_data_immext), .i_con_imm(i_con_Ealusrc), .o_data_alub(alu_i_data_B)
         );
  E_rdmux u_rdmux ( .i_data_rtE(i_addr_rt), .i_data_rdE(i_addr_rd), 
        .i_con_regdst(i_con_Eregdst), .i_con_aluPC4(i_con_Malupc8), 
        .o_data_writeE(o_addr_Erd) );
  D_compare u_compare ( .o_con_ifbranch(o_con_ifbranch), .i_data_rs(
        compare_i_data_rs), .i_data_rt({compare_i_data_rt[31:17], n1, 
        compare_i_data_rt[15:0]}), .i_con_bop(i_con_bop) );
  DFC1 pipe_rt_reg_19_ ( .D(compare_i_data_rt[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[19]) );
  DFC1 pipe_rt_reg_18_ ( .D(compare_i_data_rt[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[18]) );
  DFC1 pipe_rt_reg_17_ ( .D(compare_i_data_rt[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[17]) );
  DFC1 pipe_rt_reg_9_ ( .D(compare_i_data_rt[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[9]) );
  DFC1 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC1 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC1 pipe_rt_reg_0_ ( .D(compare_i_data_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[0]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  BUF2 U3 ( .A(compare_i_data_rt[16]), .Q(n1) );
endmodule


module M_resmux ( i_data_alures, i_data_pc8, i_con_pc8, o_data_alu );
  input [31:0] i_data_alures;
  input [31:0] i_data_pc8;
  output [31:0] o_data_alu;
  input i_con_pc8;
  wire   n34, n35, n36, n37, n38, n39, n40, n43, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n1;

  INV3 U1 ( .A(n40), .Q(o_data_alu[3]) );
  INV3 U2 ( .A(n39), .Q(o_data_alu[4]) );
  INV3 U3 ( .A(n36), .Q(o_data_alu[7]) );
  INV3 U4 ( .A(n35), .Q(o_data_alu[8]) );
  INV3 U5 ( .A(n34), .Q(o_data_alu[9]) );
  INV3 U6 ( .A(n63), .Q(o_data_alu[11]) );
  INV3 U7 ( .A(n62), .Q(o_data_alu[12]) );
  INV3 U8 ( .A(n61), .Q(o_data_alu[13]) );
  INV3 U9 ( .A(n59), .Q(o_data_alu[15]) );
  INV3 U10 ( .A(n58), .Q(o_data_alu[16]) );
  INV3 U11 ( .A(n57), .Q(o_data_alu[17]) );
  INV3 U12 ( .A(n55), .Q(o_data_alu[19]) );
  INV3 U13 ( .A(n53), .Q(o_data_alu[20]) );
  INV3 U14 ( .A(n52), .Q(o_data_alu[21]) );
  INV3 U15 ( .A(n50), .Q(o_data_alu[23]) );
  INV3 U16 ( .A(n49), .Q(o_data_alu[24]) );
  INV3 U17 ( .A(n48), .Q(o_data_alu[25]) );
  MUX22 U18 ( .A(i_data_alures[30]), .B(i_data_pc8[30]), .S(i_con_pc8), .Q(
        o_data_alu[30]) );
  AOI221 U19 ( .A(i_data_alures[23]), .B(n1), .C(i_data_pc8[23]), .D(i_con_pc8), .Q(n50) );
  AOI221 U20 ( .A(i_data_alures[20]), .B(n1), .C(i_data_pc8[20]), .D(i_con_pc8), .Q(n53) );
  AOI221 U21 ( .A(i_data_alures[21]), .B(n1), .C(i_data_pc8[21]), .D(i_con_pc8), .Q(n52) );
  AOI221 U22 ( .A(i_data_alures[24]), .B(n1), .C(i_data_pc8[24]), .D(i_con_pc8), .Q(n49) );
  AOI221 U23 ( .A(i_data_alures[11]), .B(n1), .C(i_data_pc8[11]), .D(i_con_pc8), .Q(n63) );
  AOI221 U24 ( .A(i_data_alures[15]), .B(n1), .C(i_data_pc8[15]), .D(i_con_pc8), .Q(n59) );
  AOI221 U25 ( .A(i_data_alures[16]), .B(n1), .C(i_data_pc8[16]), .D(i_con_pc8), .Q(n58) );
  AOI221 U26 ( .A(i_data_alures[17]), .B(n1), .C(i_data_pc8[17]), .D(i_con_pc8), .Q(n57) );
  AOI221 U27 ( .A(i_data_alures[19]), .B(n1), .C(i_data_pc8[19]), .D(i_con_pc8), .Q(n55) );
  AOI221 U28 ( .A(i_data_alures[25]), .B(n1), .C(i_data_pc8[25]), .D(i_con_pc8), .Q(n48) );
  AOI221 U29 ( .A(i_data_alures[9]), .B(n1), .C(i_data_pc8[9]), .D(i_con_pc8), 
        .Q(n34) );
  AOI221 U30 ( .A(i_data_alures[12]), .B(n1), .C(i_data_pc8[12]), .D(i_con_pc8), .Q(n62) );
  AOI221 U31 ( .A(i_data_alures[13]), .B(n1), .C(i_data_pc8[13]), .D(i_con_pc8), .Q(n61) );
  AOI221 U32 ( .A(i_data_alures[3]), .B(n1), .C(i_data_pc8[3]), .D(i_con_pc8), 
        .Q(n40) );
  AOI221 U33 ( .A(i_data_alures[4]), .B(n1), .C(i_data_pc8[4]), .D(i_con_pc8), 
        .Q(n39) );
  AOI221 U34 ( .A(i_data_alures[7]), .B(n1), .C(i_data_pc8[7]), .D(i_con_pc8), 
        .Q(n36) );
  AOI221 U35 ( .A(i_data_alures[8]), .B(n1), .C(i_data_pc8[8]), .D(i_con_pc8), 
        .Q(n35) );
  MUX22 U36 ( .A(i_data_alures[31]), .B(i_data_pc8[31]), .S(i_con_pc8), .Q(
        o_data_alu[31]) );
  INV3 U37 ( .A(n60), .Q(o_data_alu[14]) );
  AOI221 U38 ( .A(i_data_alures[14]), .B(n1), .C(i_data_pc8[14]), .D(i_con_pc8), .Q(n60) );
  INV3 U39 ( .A(n56), .Q(o_data_alu[18]) );
  AOI221 U40 ( .A(i_data_alures[18]), .B(n1), .C(i_data_pc8[18]), .D(i_con_pc8), .Q(n56) );
  INV3 U41 ( .A(n51), .Q(o_data_alu[22]) );
  AOI221 U42 ( .A(i_data_alures[22]), .B(n1), .C(i_data_pc8[22]), .D(i_con_pc8), .Q(n51) );
  INV3 U43 ( .A(n47), .Q(o_data_alu[26]) );
  AOI221 U44 ( .A(i_data_alures[26]), .B(n1), .C(i_data_pc8[26]), .D(i_con_pc8), .Q(n47) );
  MUX22 U45 ( .A(i_data_alures[27]), .B(i_data_pc8[27]), .S(i_con_pc8), .Q(
        o_data_alu[27]) );
  MUX22 U46 ( .A(i_data_alures[28]), .B(i_data_pc8[28]), .S(i_con_pc8), .Q(
        o_data_alu[28]) );
  MUX22 U47 ( .A(i_data_alures[29]), .B(i_data_pc8[29]), .S(i_con_pc8), .Q(
        o_data_alu[29]) );
  INV3 U48 ( .A(n38), .Q(o_data_alu[5]) );
  AOI221 U49 ( .A(i_data_alures[5]), .B(n1), .C(i_data_pc8[5]), .D(i_con_pc8), 
        .Q(n38) );
  INV3 U50 ( .A(n37), .Q(o_data_alu[6]) );
  AOI221 U51 ( .A(i_data_alures[6]), .B(n1), .C(i_data_pc8[6]), .D(i_con_pc8), 
        .Q(n37) );
  INV3 U52 ( .A(n64), .Q(o_data_alu[10]) );
  AOI221 U53 ( .A(i_data_alures[10]), .B(n1), .C(i_data_pc8[10]), .D(i_con_pc8), .Q(n64) );
  INV3 U54 ( .A(i_con_pc8), .Q(n1) );
  INV3 U55 ( .A(n65), .Q(o_data_alu[0]) );
  AOI221 U56 ( .A(i_data_alures[0]), .B(n1), .C(i_data_pc8[0]), .D(i_con_pc8), 
        .Q(n65) );
  INV3 U57 ( .A(n54), .Q(o_data_alu[1]) );
  AOI221 U58 ( .A(i_data_alures[1]), .B(n1), .C(i_data_pc8[1]), .D(i_con_pc8), 
        .Q(n54) );
  INV3 U59 ( .A(n43), .Q(o_data_alu[2]) );
  AOI221 U60 ( .A(i_data_alures[2]), .B(n1), .C(i_data_pc8[2]), .D(i_con_pc8), 
        .Q(n43) );
endmodule


module mem_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INV3 U2 ( .A(n53), .Q(n54) );
  INV3 U3 ( .A(n41), .Q(n42) );
  INV3 U4 ( .A(n29), .Q(n30) );
  INV3 U5 ( .A(n66), .Q(n67) );
  INV3 U6 ( .A(n77), .Q(n78) );
  NOR21 U7 ( .A(n82), .B(n83), .Q(n81) );
  INV3 U8 ( .A(n84), .Q(n82) );
  NOR31 U9 ( .A(n9), .B(n85), .C(n6), .Q(n84) );
  NAND22 U10 ( .A(n35), .B(n36), .Q(n34) );
  NOR31 U11 ( .A(n39), .B(n37), .C(n38), .Q(n36) );
  NOR21 U12 ( .A(n22), .B(n34), .Q(n21) );
  INV3 U13 ( .A(n23), .Q(n22) );
  NOR31 U14 ( .A(n26), .B(n24), .C(n25), .Q(n23) );
  INV3 U15 ( .A(n58), .Q(n47) );
  NAND31 U16 ( .A(n59), .B(n60), .C(n61), .Q(n58) );
  NOR21 U17 ( .A(n63), .B(n64), .Q(n59) );
  INV3 U18 ( .A(n62), .Q(n60) );
  NOR21 U19 ( .A(n51), .B(n55), .Q(n53) );
  NOR21 U20 ( .A(n39), .B(n43), .Q(n41) );
  NOR21 U21 ( .A(n26), .B(n31), .Q(n29) );
  NOR21 U22 ( .A(n64), .B(n68), .Q(n66) );
  NAND22 U23 ( .A(n66), .B(A[14]), .Q(n65) );
  NAND22 U24 ( .A(n53), .B(A[18]), .Q(n52) );
  NAND22 U25 ( .A(n41), .B(A[22]), .Q(n40) );
  NOR21 U26 ( .A(n79), .B(n2), .Q(n77) );
  NAND22 U27 ( .A(n5), .B(A[6]), .Q(n4) );
  NAND22 U28 ( .A(n77), .B(A[10]), .Q(n76) );
  INV3 U29 ( .A(n7), .Q(n5) );
  NAND22 U30 ( .A(n8), .B(A[5]), .Q(n7) );
  INV3 U31 ( .A(n8), .Q(n10) );
  NAND22 U32 ( .A(A[3]), .B(A[2]), .Q(n83) );
  NOR21 U33 ( .A(n19), .B(n20), .Q(n18) );
  INV3 U34 ( .A(A[28]), .Q(n20) );
  NOR21 U35 ( .A(n72), .B(n3), .Q(n61) );
  INV3 U36 ( .A(n73), .Q(n72) );
  NOR31 U37 ( .A(n2), .B(n74), .C(n75), .Q(n73) );
  NAND22 U38 ( .A(A[11]), .B(A[8]), .Q(n74) );
  NOR21 U39 ( .A(n15), .B(n17), .Q(n14) );
  INV3 U40 ( .A(A[2]), .Q(SUM[2]) );
  INV3 U41 ( .A(n46), .Q(n35) );
  NAND22 U42 ( .A(n47), .B(n48), .Q(n46) );
  NOR31 U43 ( .A(n51), .B(n49), .C(n50), .Q(n48) );
  NAND22 U44 ( .A(A[19]), .B(A[16]), .Q(n49) );
  XOR21 U45 ( .A(A[30]), .B(n14), .Q(SUM[30]) );
  XOR21 U46 ( .A(n12), .B(n13), .Q(SUM[31]) );
  INV3 U47 ( .A(A[31]), .Q(n12) );
  NAND22 U48 ( .A(A[30]), .B(n14), .Q(n13) );
  INV3 U49 ( .A(A[17]), .Q(n51) );
  NOR21 U50 ( .A(n34), .B(n33), .Q(n32) );
  INV3 U51 ( .A(A[24]), .Q(n33) );
  INV3 U52 ( .A(A[9]), .Q(n2) );
  INV3 U53 ( .A(A[13]), .Q(n64) );
  NOR21 U54 ( .A(n70), .B(n71), .Q(n69) );
  INV3 U55 ( .A(A[12]), .Q(n71) );
  INV3 U56 ( .A(A[5]), .Q(n9) );
  INV3 U57 ( .A(A[14]), .Q(n63) );
  NOR21 U58 ( .A(n58), .B(n57), .Q(n56) );
  INV3 U59 ( .A(A[16]), .Q(n57) );
  NOR21 U60 ( .A(n46), .B(n45), .Q(n44) );
  INV3 U61 ( .A(A[20]), .Q(n45) );
  INV3 U62 ( .A(A[6]), .Q(n6) );
  INV3 U63 ( .A(A[10]), .Q(n75) );
  NAND22 U64 ( .A(A[7]), .B(A[4]), .Q(n85) );
  NAND22 U65 ( .A(A[15]), .B(A[12]), .Q(n62) );
  XNR21 U66 ( .A(n67), .B(A[14]), .Q(SUM[14]) );
  XNR21 U67 ( .A(A[15]), .B(n65), .Q(SUM[15]) );
  XNR21 U68 ( .A(n56), .B(n51), .Q(SUM[17]) );
  XNR21 U69 ( .A(n54), .B(A[18]), .Q(SUM[18]) );
  XNR21 U70 ( .A(A[19]), .B(n52), .Q(SUM[19]) );
  XNR21 U71 ( .A(A[20]), .B(n46), .Q(SUM[20]) );
  XNR21 U72 ( .A(n44), .B(n39), .Q(SUM[21]) );
  XNR21 U73 ( .A(n42), .B(A[22]), .Q(SUM[22]) );
  XNR21 U74 ( .A(A[23]), .B(n40), .Q(SUM[23]) );
  XNR21 U75 ( .A(A[24]), .B(n34), .Q(SUM[24]) );
  XNR21 U76 ( .A(n32), .B(n26), .Q(SUM[25]) );
  XNR21 U77 ( .A(n30), .B(A[26]), .Q(SUM[26]) );
  XOR21 U78 ( .A(n27), .B(n28), .Q(SUM[27]) );
  INV3 U79 ( .A(A[27]), .Q(n27) );
  NAND22 U80 ( .A(n29), .B(A[26]), .Q(n28) );
  XOR21 U81 ( .A(n20), .B(n19), .Q(SUM[28]) );
  XOR21 U82 ( .A(n17), .B(n15), .Q(SUM[29]) );
  INV3 U83 ( .A(A[29]), .Q(n17) );
  NOR21 U84 ( .A(n83), .B(n11), .Q(n8) );
  INV3 U85 ( .A(A[4]), .Q(n11) );
  NOR21 U86 ( .A(n3), .B(n80), .Q(n1) );
  INV3 U87 ( .A(A[8]), .Q(n80) );
  INV3 U88 ( .A(A[21]), .Q(n39) );
  INV3 U89 ( .A(A[25]), .Q(n26) );
  INV3 U90 ( .A(A[18]), .Q(n50) );
  INV3 U91 ( .A(A[22]), .Q(n38) );
  INV3 U92 ( .A(A[26]), .Q(n25) );
  NAND22 U93 ( .A(A[27]), .B(A[24]), .Q(n24) );
  NAND22 U94 ( .A(A[23]), .B(A[20]), .Q(n37) );
  XNR21 U95 ( .A(A[16]), .B(n58), .Q(SUM[16]) );
  XNR21 U96 ( .A(n10), .B(A[5]), .Q(SUM[5]) );
  XNR21 U97 ( .A(n7), .B(A[6]), .Q(SUM[6]) );
  XNR21 U98 ( .A(A[7]), .B(n4), .Q(SUM[7]) );
  XNR21 U99 ( .A(A[8]), .B(n3), .Q(SUM[8]) );
  XNR21 U100 ( .A(n1), .B(n2), .Q(SUM[9]) );
  XNR21 U101 ( .A(n78), .B(A[10]), .Q(SUM[10]) );
  XNR21 U102 ( .A(A[11]), .B(n76), .Q(SUM[11]) );
  XNR21 U103 ( .A(A[12]), .B(n70), .Q(SUM[12]) );
  XNR21 U104 ( .A(n69), .B(n64), .Q(SUM[13]) );
  XNR21 U105 ( .A(A[3]), .B(SUM[2]), .Q(SUM[3]) );
  XNR21 U106 ( .A(A[4]), .B(n83), .Q(SUM[4]) );
  CLKIN3 U107 ( .A(n18), .Q(n15) );
  CLKIN3 U108 ( .A(n21), .Q(n19) );
  CLKIN3 U109 ( .A(n32), .Q(n31) );
  CLKIN3 U110 ( .A(n44), .Q(n43) );
  CLKIN3 U111 ( .A(n56), .Q(n55) );
  CLKIN3 U112 ( .A(n69), .Q(n68) );
  CLKIN3 U113 ( .A(n61), .Q(n70) );
  CLKIN3 U114 ( .A(n1), .Q(n79) );
  CLKIN3 U115 ( .A(n81), .Q(n3) );
endmodule


module mem ( i_clk, i_nrst, i_data_pc4, i_data_alures, i_data_memout, 
        i_addr_regdst, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_FWmemread, i_addr_Mrt, o_data_alures, o_data_memout, 
        o_addr_regdst, o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread, 
        o_addr_Wrt );
  input [31:0] i_data_pc4;
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  input [4:0] i_addr_regdst;
  input [4:0] i_addr_Mrt;
  output [31:0] o_data_alures;
  output [31:0] o_data_memout;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Wrt;
  input i_clk, i_nrst, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite,
         i_con_FWmemread;
  output o_con_Wmemtoreg, o_con_Wregwrite, o_con_FWmemread;
  wire   n_Logic1_, n_Logic0_;
  wire   [31:0] pc8;
  wire   [31:0] resmux_o_data_alu;

  DFC3 pipe_rt_reg_4_ ( .D(i_addr_Mrt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[4]) );
  DFC3 pipe_rt_reg_3_ ( .D(i_addr_Mrt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[3]) );
  DFC3 pipe_rt_reg_2_ ( .D(i_addr_Mrt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[2]) );
  DFC3 pipe_rt_reg_1_ ( .D(i_addr_Mrt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[1]) );
  DFC3 pipe_rt_reg_0_ ( .D(i_addr_Mrt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Wrt[0]) );
  DFC3 pipe_data_alures_reg_31_ ( .D(resmux_o_data_alu[31]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[31]) );
  DFC3 pipe_data_alures_reg_30_ ( .D(resmux_o_data_alu[30]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[30]) );
  DFC3 pipe_data_alures_reg_29_ ( .D(resmux_o_data_alu[29]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[29]) );
  DFC3 pipe_data_alures_reg_28_ ( .D(resmux_o_data_alu[28]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[28]) );
  DFC3 pipe_data_alures_reg_27_ ( .D(resmux_o_data_alu[27]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[27]) );
  DFC3 pipe_data_alures_reg_26_ ( .D(resmux_o_data_alu[26]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[26]) );
  DFC3 pipe_data_alures_reg_25_ ( .D(resmux_o_data_alu[25]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[25]) );
  DFC3 pipe_data_alures_reg_24_ ( .D(resmux_o_data_alu[24]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[24]) );
  DFC3 pipe_data_alures_reg_23_ ( .D(resmux_o_data_alu[23]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[23]) );
  DFC3 pipe_data_alures_reg_22_ ( .D(resmux_o_data_alu[22]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[22]) );
  DFC3 pipe_data_alures_reg_21_ ( .D(resmux_o_data_alu[21]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[21]) );
  DFC3 pipe_data_alures_reg_20_ ( .D(resmux_o_data_alu[20]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[20]) );
  DFC3 pipe_data_alures_reg_19_ ( .D(resmux_o_data_alu[19]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[19]) );
  DFC3 pipe_data_alures_reg_18_ ( .D(resmux_o_data_alu[18]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[18]) );
  DFC3 pipe_data_alures_reg_17_ ( .D(resmux_o_data_alu[17]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[17]) );
  DFC3 pipe_data_alures_reg_16_ ( .D(resmux_o_data_alu[16]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[16]) );
  DFC3 pipe_data_alures_reg_15_ ( .D(resmux_o_data_alu[15]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[15]) );
  DFC3 pipe_data_alures_reg_14_ ( .D(resmux_o_data_alu[14]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[14]) );
  DFC3 pipe_data_alures_reg_13_ ( .D(resmux_o_data_alu[13]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[13]) );
  DFC3 pipe_data_alures_reg_12_ ( .D(resmux_o_data_alu[12]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[12]) );
  DFC3 pipe_data_alures_reg_11_ ( .D(resmux_o_data_alu[11]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[11]) );
  DFC3 pipe_data_alures_reg_10_ ( .D(resmux_o_data_alu[10]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[10]) );
  DFC3 pipe_data_alures_reg_9_ ( .D(resmux_o_data_alu[9]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[9]) );
  DFC3 pipe_data_alures_reg_8_ ( .D(resmux_o_data_alu[8]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[8]) );
  DFC3 pipe_data_alures_reg_7_ ( .D(resmux_o_data_alu[7]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[7]) );
  DFC3 pipe_data_alures_reg_6_ ( .D(resmux_o_data_alu[6]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[6]) );
  DFC3 pipe_data_alures_reg_5_ ( .D(resmux_o_data_alu[5]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[5]) );
  DFC3 pipe_data_alures_reg_4_ ( .D(resmux_o_data_alu[4]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[4]) );
  DFC3 pipe_data_alures_reg_3_ ( .D(resmux_o_data_alu[3]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[3]) );
  DFC3 pipe_data_alures_reg_2_ ( .D(resmux_o_data_alu[2]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[2]) );
  DFC3 pipe_data_alures_reg_1_ ( .D(resmux_o_data_alu[1]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[1]) );
  DFC3 pipe_data_alures_reg_0_ ( .D(resmux_o_data_alu[0]), .C(i_clk), .RN(
        i_nrst), .Q(o_data_alures[0]) );
  DFC3 pipe_data_memout_reg_31_ ( .D(i_data_memout[31]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[31]) );
  DFC3 pipe_data_memout_reg_30_ ( .D(i_data_memout[30]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[30]) );
  DFC3 pipe_data_memout_reg_29_ ( .D(i_data_memout[29]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[29]) );
  DFC3 pipe_data_memout_reg_28_ ( .D(i_data_memout[28]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[28]) );
  DFC3 pipe_data_memout_reg_27_ ( .D(i_data_memout[27]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[27]) );
  DFC3 pipe_data_memout_reg_26_ ( .D(i_data_memout[26]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[26]) );
  DFC3 pipe_data_memout_reg_25_ ( .D(i_data_memout[25]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[25]) );
  DFC3 pipe_data_memout_reg_24_ ( .D(i_data_memout[24]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[24]) );
  DFC3 pipe_data_memout_reg_23_ ( .D(i_data_memout[23]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[23]) );
  DFC3 pipe_data_memout_reg_22_ ( .D(i_data_memout[22]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[22]) );
  DFC3 pipe_data_memout_reg_21_ ( .D(i_data_memout[21]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[21]) );
  DFC3 pipe_data_memout_reg_20_ ( .D(i_data_memout[20]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[20]) );
  DFC3 pipe_data_memout_reg_19_ ( .D(i_data_memout[19]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[19]) );
  DFC3 pipe_data_memout_reg_18_ ( .D(i_data_memout[18]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[18]) );
  DFC3 pipe_data_memout_reg_17_ ( .D(i_data_memout[17]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[17]) );
  DFC3 pipe_data_memout_reg_16_ ( .D(i_data_memout[16]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[16]) );
  DFC3 pipe_data_memout_reg_15_ ( .D(i_data_memout[15]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[15]) );
  DFC3 pipe_data_memout_reg_14_ ( .D(i_data_memout[14]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[14]) );
  DFC3 pipe_data_memout_reg_13_ ( .D(i_data_memout[13]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[13]) );
  DFC3 pipe_data_memout_reg_12_ ( .D(i_data_memout[12]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[12]) );
  DFC3 pipe_data_memout_reg_11_ ( .D(i_data_memout[11]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[11]) );
  DFC3 pipe_data_memout_reg_10_ ( .D(i_data_memout[10]), .C(i_clk), .RN(i_nrst), .Q(o_data_memout[10]) );
  DFC3 pipe_data_memout_reg_9_ ( .D(i_data_memout[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[9]) );
  DFC3 pipe_data_memout_reg_8_ ( .D(i_data_memout[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[8]) );
  DFC3 pipe_data_memout_reg_7_ ( .D(i_data_memout[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[7]) );
  DFC3 pipe_data_memout_reg_6_ ( .D(i_data_memout[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[6]) );
  DFC3 pipe_data_memout_reg_5_ ( .D(i_data_memout[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[5]) );
  DFC3 pipe_data_memout_reg_4_ ( .D(i_data_memout[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[4]) );
  DFC3 pipe_data_memout_reg_3_ ( .D(i_data_memout[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[3]) );
  DFC3 pipe_data_memout_reg_2_ ( .D(i_data_memout[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[2]) );
  DFC3 pipe_data_memout_reg_1_ ( .D(i_data_memout[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[1]) );
  DFC3 pipe_data_memout_reg_0_ ( .D(i_data_memout[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_memout[0]) );
  DFC3 pipe_addr_regdst_reg_4_ ( .D(i_addr_regdst[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[4]) );
  DFC3 pipe_addr_regdst_reg_3_ ( .D(i_addr_regdst[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[3]) );
  DFC3 pipe_addr_regdst_reg_2_ ( .D(i_addr_regdst[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[2]) );
  DFC3 pipe_addr_regdst_reg_1_ ( .D(i_addr_regdst[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[1]) );
  DFC3 pipe_addr_regdst_reg_0_ ( .D(i_addr_regdst[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_addr_regdst[0]) );
  DFC3 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC3 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_con_FWmemread_reg ( .D(i_con_FWmemread), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_FWmemread) );
  M_resmux u_resmux ( .i_data_alures(i_data_alures), .i_data_pc8(pc8), 
        .i_con_pc8(i_con_Malupc8), .o_data_alu(resmux_o_data_alu) );
  mem_DW01_add_1 add_27 ( .A(i_data_pc4), .B({n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, n_Logic0_, 
        n_Logic0_, n_Logic0_, n_Logic1_, n_Logic0_, n_Logic0_}), .CI(n_Logic0_), .SUM(pc8) );
  LOGIC0 U3 ( .Q(n_Logic0_) );
  LOGIC1 U4 ( .Q(n_Logic1_) );
endmodule


module W_datamux ( i_data_alu, i_data_load, i_con_memtoreg, o_data_toreg );
  input [31:0] i_data_alu;
  input [31:0] i_data_load;
  output [31:0] o_data_toreg;
  input i_con_memtoreg;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n1;

  INV3 U1 ( .A(n65), .Q(o_data_toreg[0]) );
  AOI221 U2 ( .A(i_data_alu[0]), .B(n1), .C(i_data_load[0]), .D(i_con_memtoreg), .Q(n65) );
  INV3 U3 ( .A(n54), .Q(o_data_toreg[1]) );
  AOI221 U4 ( .A(i_data_alu[1]), .B(n1), .C(i_data_load[1]), .D(i_con_memtoreg), .Q(n54) );
  INV3 U5 ( .A(n43), .Q(o_data_toreg[2]) );
  AOI221 U6 ( .A(i_data_alu[2]), .B(n1), .C(i_data_load[2]), .D(i_con_memtoreg), .Q(n43) );
  INV3 U7 ( .A(n40), .Q(o_data_toreg[3]) );
  AOI221 U8 ( .A(i_data_alu[3]), .B(n1), .C(i_data_load[3]), .D(i_con_memtoreg), .Q(n40) );
  INV3 U9 ( .A(n64), .Q(o_data_toreg[10]) );
  AOI221 U10 ( .A(i_data_alu[10]), .B(n1), .C(i_data_load[10]), .D(
        i_con_memtoreg), .Q(n64) );
  INV3 U11 ( .A(n63), .Q(o_data_toreg[11]) );
  AOI221 U12 ( .A(i_data_alu[11]), .B(n1), .C(i_data_load[11]), .D(
        i_con_memtoreg), .Q(n63) );
  INV3 U13 ( .A(n62), .Q(o_data_toreg[12]) );
  AOI221 U14 ( .A(i_data_alu[12]), .B(n1), .C(i_data_load[12]), .D(
        i_con_memtoreg), .Q(n62) );
  INV3 U15 ( .A(n61), .Q(o_data_toreg[13]) );
  AOI221 U16 ( .A(i_data_alu[13]), .B(n1), .C(i_data_load[13]), .D(
        i_con_memtoreg), .Q(n61) );
  INV3 U17 ( .A(n60), .Q(o_data_toreg[14]) );
  AOI221 U18 ( .A(i_data_alu[14]), .B(n1), .C(i_data_load[14]), .D(
        i_con_memtoreg), .Q(n60) );
  INV3 U19 ( .A(n59), .Q(o_data_toreg[15]) );
  AOI221 U20 ( .A(i_data_alu[15]), .B(n1), .C(i_data_load[15]), .D(
        i_con_memtoreg), .Q(n59) );
  INV3 U21 ( .A(n58), .Q(o_data_toreg[16]) );
  AOI221 U22 ( .A(i_data_alu[16]), .B(n1), .C(i_data_load[16]), .D(
        i_con_memtoreg), .Q(n58) );
  INV3 U23 ( .A(n57), .Q(o_data_toreg[17]) );
  AOI221 U24 ( .A(i_data_alu[17]), .B(n1), .C(i_data_load[17]), .D(
        i_con_memtoreg), .Q(n57) );
  INV3 U25 ( .A(n56), .Q(o_data_toreg[18]) );
  AOI221 U26 ( .A(i_data_alu[18]), .B(n1), .C(i_data_load[18]), .D(
        i_con_memtoreg), .Q(n56) );
  INV3 U27 ( .A(n55), .Q(o_data_toreg[19]) );
  AOI221 U28 ( .A(i_data_alu[19]), .B(n1), .C(i_data_load[19]), .D(
        i_con_memtoreg), .Q(n55) );
  INV3 U29 ( .A(n53), .Q(o_data_toreg[20]) );
  AOI221 U30 ( .A(i_data_alu[20]), .B(n1), .C(i_data_load[20]), .D(
        i_con_memtoreg), .Q(n53) );
  INV3 U31 ( .A(n52), .Q(o_data_toreg[21]) );
  AOI221 U32 ( .A(i_data_alu[21]), .B(n1), .C(i_data_load[21]), .D(
        i_con_memtoreg), .Q(n52) );
  INV3 U33 ( .A(n51), .Q(o_data_toreg[22]) );
  AOI221 U34 ( .A(i_data_alu[22]), .B(n1), .C(i_data_load[22]), .D(
        i_con_memtoreg), .Q(n51) );
  INV3 U35 ( .A(n50), .Q(o_data_toreg[23]) );
  AOI221 U36 ( .A(i_data_alu[23]), .B(n1), .C(i_data_load[23]), .D(
        i_con_memtoreg), .Q(n50) );
  INV3 U37 ( .A(n49), .Q(o_data_toreg[24]) );
  AOI221 U38 ( .A(i_data_alu[24]), .B(n1), .C(i_data_load[24]), .D(
        i_con_memtoreg), .Q(n49) );
  INV3 U39 ( .A(n48), .Q(o_data_toreg[25]) );
  AOI221 U40 ( .A(i_data_alu[25]), .B(n1), .C(i_data_load[25]), .D(
        i_con_memtoreg), .Q(n48) );
  INV3 U41 ( .A(n47), .Q(o_data_toreg[26]) );
  AOI221 U42 ( .A(i_data_alu[26]), .B(n1), .C(i_data_load[26]), .D(
        i_con_memtoreg), .Q(n47) );
  INV3 U43 ( .A(n46), .Q(o_data_toreg[27]) );
  AOI221 U44 ( .A(i_data_alu[27]), .B(n1), .C(i_data_load[27]), .D(
        i_con_memtoreg), .Q(n46) );
  INV3 U45 ( .A(n45), .Q(o_data_toreg[28]) );
  AOI221 U46 ( .A(i_data_alu[28]), .B(n1), .C(i_data_load[28]), .D(
        i_con_memtoreg), .Q(n45) );
  INV3 U47 ( .A(n44), .Q(o_data_toreg[29]) );
  AOI221 U48 ( .A(i_data_alu[29]), .B(n1), .C(i_data_load[29]), .D(
        i_con_memtoreg), .Q(n44) );
  INV3 U49 ( .A(n42), .Q(o_data_toreg[30]) );
  AOI221 U50 ( .A(i_data_alu[30]), .B(n1), .C(i_data_load[30]), .D(
        i_con_memtoreg), .Q(n42) );
  INV3 U51 ( .A(n41), .Q(o_data_toreg[31]) );
  AOI221 U52 ( .A(i_data_alu[31]), .B(n1), .C(i_data_load[31]), .D(
        i_con_memtoreg), .Q(n41) );
  INV3 U53 ( .A(n39), .Q(o_data_toreg[4]) );
  AOI221 U54 ( .A(i_data_alu[4]), .B(n1), .C(i_data_load[4]), .D(
        i_con_memtoreg), .Q(n39) );
  INV3 U55 ( .A(n38), .Q(o_data_toreg[5]) );
  AOI221 U56 ( .A(i_data_alu[5]), .B(n1), .C(i_data_load[5]), .D(
        i_con_memtoreg), .Q(n38) );
  INV3 U57 ( .A(n37), .Q(o_data_toreg[6]) );
  AOI221 U58 ( .A(i_data_alu[6]), .B(n1), .C(i_data_load[6]), .D(
        i_con_memtoreg), .Q(n37) );
  INV3 U59 ( .A(n36), .Q(o_data_toreg[7]) );
  AOI221 U60 ( .A(i_data_alu[7]), .B(n1), .C(i_data_load[7]), .D(
        i_con_memtoreg), .Q(n36) );
  INV3 U61 ( .A(n35), .Q(o_data_toreg[8]) );
  AOI221 U62 ( .A(i_data_alu[8]), .B(n1), .C(i_data_load[8]), .D(
        i_con_memtoreg), .Q(n35) );
  INV3 U63 ( .A(n34), .Q(o_data_toreg[9]) );
  AOI221 U64 ( .A(i_data_alu[9]), .B(n1), .C(i_data_load[9]), .D(
        i_con_memtoreg), .Q(n34) );
  INV3 U65 ( .A(i_con_memtoreg), .Q(n1) );
endmodule


module writeback ( i_data_alures, i_data_memout, i_con_Wmemtoreg, 
        o_data_regwrite );
  input [31:0] i_data_alures;
  input [31:0] i_data_memout;
  output [31:0] o_data_regwrite;
  input i_con_Wmemtoreg;


  W_datamux u_datamux ( .i_data_alu(i_data_alures), .i_data_load(i_data_memout), .i_con_memtoreg(i_con_Wmemtoreg), .o_data_toreg(o_data_regwrite) );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Mmemread, ex_con_Mmemwrite, ex_con_Malupc8, ex_con_Wmemtoreg,
         mem_con_Malupc8, mem_con_Wmemtoreg, wb_con_Wmemtoreg, n1,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2;
  wire   [31:0] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [31:0] id_addr_pc4;
  wire   [31:0] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] wb_data_memout;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] mem_data_alures;
  wire   [31:0] mem_data_pc4;

  fetch u_fetch ( .i_clk(clk), .i_nrst(rst_n), .i_addr_b(if_addr_b), 
        .i_addr_j({if_addr_j, n1, n1}), .i_addr_jr(id_data_jr), .i_con_b(
        if_con_b), .i_con_j(if_con_j), .i_data_instr(read_instruction), 
        .i_con_ifstall(if_con_ifstall), .o_addr_pc(instruction_address), 
        .o_addr_pc4(id_addr_pc4), .o_data_instr(id_data_instr) );
  decode u_decode ( .i_clk(clk), .i_nrst(rst_n), .i_addr_pc4(id_addr_pc4), 
        .i_data_instr(id_data_instr), .i_con_Wregwrite(id_con_Wregwrite), 
        .i_data_Wregwrite(id_data_Wregwrite), .i_addr_Wregwrite(
        id_addr_Wregwrite), .i_addr_Erd(for_o_addr_Erd), .i_addr_Mrd(
        mem_addr_regdst), .i_con_Eregwrite(ex_con_Wregwrite), 
        .i_con_Mregwrite(mem_con_Wregwrite), .i_addr_rtM(for_addr_rtM), 
        .i_addr_rtW(for_addr_rtW), .i_con_memreadM(mem_read), .i_con_memreadW(
        for_FWmemread), .i_data_Wmemout(wb_data_memout), .o_data_rs(id_data_rs), .o_data_rt(ex_data_rt), .o_addr_rd(ex_addr_rd), .o_addr_rt(ex_addr_rt), 
        .o_data_jr(id_data_jr), .o_con_jump(if_con_j), .o_addr_pc4(ex_data_pc4), .o_addr_branch(if_addr_b), .o_addr_jump({if_addr_j, SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2}), .o_con_Ealuop(ex_con_Ealuop), 
        .o_con_Ealusrc(ex_con_Ealusrc), .o_con_Eregdst(ex_con_Eregdst), 
        .o_con_Mmemread(ex_con_Mmemread), .o_con_Mmemwrite(ex_con_Mmemwrite), 
        .o_con_Malupc8(ex_con_Malupc8), .o_con_Wmemtoreg(ex_con_Wmemtoreg), 
        .o_con_Wregwrite(ex_con_Wregwrite), .o_con_ifstall(if_con_ifstall), 
        .o_con_Ebop(ex_con_bop), .o_data_signext(ex_data_immext), 
        .o_con_Efamux(for_o_con_Efamux), .o_con_Efbmux(for_o_con_Efbmux), 
        .o_data_Fmemout(for_memout) );
  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext(
        ex_data_immext), .i_addr_rt(ex_addr_rt), .i_addr_rd(ex_addr_rd), 
        .i_data_FEalures(data_address), .i_data_FMalures(mem_data_alures), 
        .i_data_FMmemout(wb_data_memout), .i_data_FWmemout(for_memout), 
        .i_con_Efamux(for_o_con_Efamux), .i_con_Efbmux(for_o_con_Efbmux), 
        .i_con_Ealuop(ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), 
        .i_con_Eregdst(ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), 
        .i_con_Mmemwrite(ex_con_Mmemwrite), .i_con_Malupc8(ex_con_Malupc8), 
        .i_con_Wmemtoreg(ex_con_Wmemtoreg), .i_con_Wregwrite(ex_con_Wregwrite), 
        .i_con_bop(ex_con_bop), .o_data_pc4(mem_data_pc4), .o_data_alures(
        data_address), .o_data_rt(write_data), .o_addr_regdst(mem_addr_regdst), 
        .o_con_Mmemread(mem_read), .o_con_Mmemwrite(mem_write), 
        .o_con_Malupc8(mem_con_Malupc8), .o_con_Wmemtoreg(mem_con_Wmemtoreg), 
        .o_con_Wregwrite(mem_con_Wregwrite), .o_addr_Erd(for_o_addr_Erd), 
        .o_addr_Mrt(for_addr_rtM), .o_con_ifbranch(if_con_b) );
  mem u_mem ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(mem_data_pc4), 
        .i_data_alures(data_address), .i_data_memout(read_data), 
        .i_addr_regdst(mem_addr_regdst), .i_con_Malupc8(mem_con_Malupc8), 
        .i_con_Wmemtoreg(mem_con_Wmemtoreg), .i_con_Wregwrite(
        mem_con_Wregwrite), .i_con_FWmemread(ex_con_Mmemread), .i_addr_Mrt(
        for_addr_rtM), .o_data_alures(mem_data_alures), .o_data_memout(
        wb_data_memout), .o_addr_regdst(id_addr_Wregwrite), .o_con_Wmemtoreg(
        wb_con_Wmemtoreg), .o_con_Wregwrite(id_con_Wregwrite), 
        .o_con_FWmemread(for_FWmemread), .o_addr_Wrt(for_addr_rtW) );
  writeback u_writeback ( .i_data_alures(mem_data_alures), .i_data_memout(
        wb_data_memout), .i_con_Wmemtoreg(wb_con_Wmemtoreg), .o_data_regwrite(
        id_data_Wregwrite) );
  LOGIC0 U1 ( .Q(n1) );
endmodule

