`timescale 1ns / 1ps

module E_mula(input logic [15:0]A, input logic [31:0]B, output logic [31:0]C);

	assign C = A + B; 
endmodule 