
module execute ( i_clk, i_nrst, i_data_pc4, i_data_rs, i_data_rt, 
        i_data_immext, i_addr_rt, i_addr_rd, i_data_FEalures, i_data_FMalures, 
        i_data_FMmemout, i_data_FWmemout, i_con_Efamux, i_con_Efbmux, 
        i_con_Ealuop, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread, 
        i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite, 
        i_con_bop, o_data_pc4, o_data_alures, o_data_rt, o_addr_regdst, 
        o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg, 
        o_con_Wregwrite, o_addr_Erd, o_addr_Mrt, o_con_ifbranch );
  input [31:0] i_data_pc4;
  input [31:0] i_data_rs;
  input [31:0] i_data_rt;
  input [31:0] i_data_immext;
  input [4:0] i_addr_rt;
  input [4:0] i_addr_rd;
  input [31:0] i_data_FEalures;
  input [31:0] i_data_FMalures;
  input [31:0] i_data_FMmemout;
  input [31:0] i_data_FWmemout;
  input [2:0] i_con_Efamux;
  input [2:0] i_con_Efbmux;
  input [5:0] i_con_Ealuop;
  input [2:0] i_con_bop;
  output [31:0] o_data_pc4;
  output [31:0] o_data_alures;
  output [31:0] o_data_rt;
  output [4:0] o_addr_regdst;
  output [4:0] o_addr_Erd;
  output [4:0] o_addr_Mrt;
  input i_clk, i_nrst, i_con_Ealusrc, i_con_Eregdst, i_con_Mmemread,
         i_con_Mmemwrite, i_con_Malupc8, i_con_Wmemtoreg, i_con_Wregwrite;
  output o_con_Mmemread, o_con_Mmemwrite, o_con_Malupc8, o_con_Wmemtoreg,
         o_con_Wregwrite, o_con_ifbranch;
  wire   u_alu_N306, u_alu_N256, u_alu_N253, u_alu_N252, u_alu_N250,
         u_alu_N249, u_alu_N248, u_alu_N247, u_alu_N246, u_alu_N245,
         u_alu_N241, u_alu_N240, u_alu_N235, u_alu_N234, u_alu_N233,
         u_alu_N232, u_alu_N231, u_alu_N230, u_alu_N229, u_alu_N228,
         u_alu_N227, u_alu_N226, u_alu_N225, u_alu_N224, u_alu_N222,
         u_alu_N221, u_alu_N220, u_alu_N219, u_alu_N218, u_alu_N217,
         u_alu_N216, u_alu_N215, u_alu_N214, u_alu_N213, u_alu_N209,
         u_alu_N203, u_alu_N202, u_alu_N201, u_alu_N200, u_alu_N199,
         u_alu_N198, u_alu_N197, u_alu_N196, u_alu_N195, u_alu_N194,
         u_alu_N193, u_alu_N173, u_alu_N172, u_alu_N171, u_alu_N170,
         u_alu_N169, u_alu_N168, u_alu_N167, u_alu_N166, u_alu_N165,
         u_alu_half_sub_0_, u_alu_half_sub_1_, u_alu_half_sub_2_,
         u_alu_half_sub_3_, u_alu_half_sub_4_, u_alu_half_sub_5_,
         u_alu_half_sub_6_, u_alu_half_sub_7_, u_alu_half_sub_8_,
         u_alu_half_sub_9_, u_alu_half_sub_10_, u_alu_half_sub_11_,
         u_alu_half_sub_12_, u_alu_half_sub_13_, u_alu_half_sub_14_,
         u_alu_half_sub_15_, u_alu_half_sub_16_, u_alu_sum_1_0_,
         u_alu_sum_1_1_, u_alu_sum_1_2_, u_alu_sum_1_3_, u_alu_sum_1_4_,
         u_alu_sum_1_5_, u_alu_sum_1_6_, u_alu_sum_1_7_, u_alu_sum_1_8_,
         u_alu_ashr_4_SH_3_, u_alu_ashr_4_SH_1_, u_alu_add_x_1_n50,
         u_alu_add_x_1_n49, u_alu_add_x_1_n48, u_alu_add_x_1_n47,
         u_alu_add_x_1_n46, u_alu_add_x_1_n45, u_alu_add_x_1_n44,
         u_alu_add_x_1_n43, u_alu_add_x_1_n41, u_alu_add_x_1_n40,
         u_alu_add_x_1_n39, u_alu_add_x_1_n38, u_alu_add_x_1_n37,
         u_alu_add_x_1_n36, u_alu_add_x_1_n35, u_alu_add_x_1_n34,
         u_alu_add_x_1_n33, u_alu_add_x_1_n32, u_alu_add_x_1_n31,
         u_alu_add_x_1_n30, u_alu_add_x_1_n29, u_alu_add_x_1_n28,
         u_alu_add_x_1_n27, u_alu_add_x_1_n26, u_alu_add_x_1_n24,
         u_alu_add_x_1_n23, u_alu_add_x_1_n22, u_alu_add_x_1_n21,
         u_alu_add_x_1_n20, u_alu_add_x_1_n19, u_alu_add_x_1_n18,
         u_alu_add_x_1_n17, u_alu_add_x_1_n16, u_alu_add_x_1_n15,
         u_alu_add_x_1_n14, u_alu_add_x_1_n13, u_alu_add_x_1_n12,
         u_alu_add_x_1_n11, u_alu_add_x_1_n10, u_alu_add_x_1_n8,
         u_alu_add_x_1_n7, u_alu_add_x_1_n6, u_alu_add_x_1_n5,
         u_alu_add_x_1_n4, u_alu_add_x_1_n3, u_alu_add_x_1_n2,
         u_alu_add_x_1_n1, u_alu_DP_OP_85J3_126_1427_n46,
         u_alu_DP_OP_85J3_126_1427_n45, u_alu_DP_OP_85J3_126_1427_n44,
         u_alu_DP_OP_85J3_126_1427_n43, u_alu_DP_OP_85J3_126_1427_n42,
         u_alu_DP_OP_85J3_126_1427_n41, u_alu_DP_OP_85J3_126_1427_n40,
         u_alu_DP_OP_85J3_126_1427_n39, u_alu_DP_OP_85J3_126_1427_n38,
         u_alu_DP_OP_85J3_126_1427_n37, u_alu_DP_OP_85J3_126_1427_n36,
         u_alu_DP_OP_85J3_126_1427_n35, u_alu_DP_OP_85J3_126_1427_n34,
         u_alu_DP_OP_85J3_126_1427_n33, u_alu_DP_OP_85J3_126_1427_n32,
         u_alu_DP_OP_84J3_125_2615_n15, u_alu_DP_OP_84J3_125_2615_n14,
         u_alu_DP_OP_84J3_125_2615_n13, u_alu_DP_OP_84J3_125_2615_n12,
         u_alu_DP_OP_84J3_125_2615_n11, u_alu_DP_OP_84J3_125_2615_n10,
         u_alu_DP_OP_84J3_125_2615_n9, u_alu_DP_OP_84J3_125_2615_n6,
         u_alu_DP_OP_84J3_125_2615_n5, u_alu_DP_OP_84J3_125_2615_n4,
         u_alu_DP_OP_84J3_125_2615_n3, u_alu_DP_OP_84J3_125_2615_n2,
         u_alu_DP_OP_84J3_125_2615_n1, u_alu_DP_OP_83J3_124_3384_n15,
         u_alu_DP_OP_83J3_124_3384_n14, u_alu_DP_OP_83J3_124_3384_n13,
         u_alu_DP_OP_83J3_124_3384_n12, u_alu_DP_OP_83J3_124_3384_n11,
         u_alu_DP_OP_83J3_124_3384_n10, u_alu_DP_OP_83J3_124_3384_n9,
         u_alu_DP_OP_83J3_124_3384_n7, u_alu_DP_OP_83J3_124_3384_n6,
         u_alu_DP_OP_83J3_124_3384_n5, u_alu_DP_OP_83J3_124_3384_n4,
         u_alu_DP_OP_83J3_124_3384_n3, u_alu_DP_OP_83J3_124_3384_n2,
         u_alu_DP_OP_83J3_124_3384_n1, u_alu_lt_x_11_B_10_, u_alu_lt_x_11_B_7_,
         u_alu_lt_x_11_B_1_, u_alu_sub_x_2_n17, u_alu_sub_x_2_n16,
         u_alu_sub_x_2_n15, u_alu_sub_x_2_n14, u_alu_sub_x_2_n13,
         u_alu_sub_x_2_n12, u_alu_sub_x_2_n11, u_alu_sub_x_2_n10,
         u_alu_sub_x_2_n9, u_alu_sub_x_2_n8, u_alu_sub_x_2_n7,
         u_alu_sub_x_2_n6, u_alu_sub_x_2_n5, u_alu_sub_x_2_n4,
         u_alu_sub_x_2_n3, u_alu_sub_x_2_n2, DP_OP_77_130_260_I3,
         DP_OP_77_130_260_n46, DP_OP_77_130_260_n45, DP_OP_77_130_260_n44,
         DP_OP_77_130_260_n43, DP_OP_77_130_260_n42, DP_OP_77_130_260_n41,
         DP_OP_77_130_260_n40, DP_OP_77_130_260_n39, DP_OP_77_130_260_n37,
         DP_OP_77_130_260_n36, DP_OP_77_130_260_n35, DP_OP_77_130_260_n34,
         DP_OP_77_130_260_n33, DP_OP_77_130_260_n32, DP_OP_77_130_260_n31,
         DP_OP_77_130_260_n30, DP_OP_77_130_260_n29, DP_OP_77_130_260_n23,
         DP_OP_77_130_260_n22, DP_OP_77_130_260_n21, DP_OP_77_130_260_n20,
         DP_OP_77_130_260_n19, DP_OP_77_130_260_n18, DP_OP_77_130_260_n17,
         DP_OP_77_130_260_n16, DP_OP_77_130_260_n15, DP_OP_77_130_260_n14,
         DP_OP_77_130_260_n13, DP_OP_77_130_260_n12, DP_OP_77_130_260_n11,
         DP_OP_77_130_260_n10, DP_OP_77_130_260_n9, DP_OP_77_130_260_n8,
         DP_OP_77_130_260_n7, DP_OP_77_130_260_n6, DP_OP_77_130_260_n5,
         DP_OP_77_130_260_n4, DP_OP_77_130_260_n3, DP_OP_77_130_260_n2,
         DP_OP_77_130_260_n1, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306;
  wire   [31:0] alu_o_data_AluRes;
  wire   [31:0] compare_i_data_rs;
  wire   [31:0] compare_i_data_rt;
  wire   [31:0] alu_i_data_B;
  wire   [3:0] alu_i_con_AluCtrl;
  wire   [15:0] u_alu_pre_subb;
  wire   [15:1] u_alu_pre_suba;
  wire   [7:1] u_alu_pre_sum_4b;
  wire   [7:0] u_alu_pre_sum_4a;
  wire   [8:1] u_alu_pre_sum_3b;
  wire   [8:0] u_alu_pre_sum_3a;

  DFC1 pipe_addr_rt_reg_4_ ( .D(i_addr_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[4]) );
  DFC1 pipe_addr_rt_reg_3_ ( .D(i_addr_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[3]) );
  DFC1 pipe_addr_rt_reg_2_ ( .D(i_addr_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[2]) );
  DFC1 pipe_addr_rt_reg_1_ ( .D(i_addr_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[1]) );
  DFC1 pipe_addr_rt_reg_0_ ( .D(i_addr_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_Mrt[0]) );
  DFC1 pipe_pc4_reg_31_ ( .D(i_data_pc4[31]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[31]) );
  DFC1 pipe_pc4_reg_30_ ( .D(i_data_pc4[30]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[30]) );
  DFC1 pipe_pc4_reg_29_ ( .D(i_data_pc4[29]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[29]) );
  DFC1 pipe_pc4_reg_28_ ( .D(i_data_pc4[28]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[28]) );
  DFC1 pipe_pc4_reg_27_ ( .D(i_data_pc4[27]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[27]) );
  DFC1 pipe_pc4_reg_26_ ( .D(i_data_pc4[26]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[26]) );
  DFC1 pipe_pc4_reg_25_ ( .D(i_data_pc4[25]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[25]) );
  DFC1 pipe_pc4_reg_24_ ( .D(i_data_pc4[24]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[24]) );
  DFC1 pipe_pc4_reg_23_ ( .D(i_data_pc4[23]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[23]) );
  DFC1 pipe_pc4_reg_22_ ( .D(i_data_pc4[22]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[22]) );
  DFC1 pipe_pc4_reg_21_ ( .D(i_data_pc4[21]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[21]) );
  DFC1 pipe_pc4_reg_20_ ( .D(i_data_pc4[20]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[20]) );
  DFC1 pipe_pc4_reg_19_ ( .D(i_data_pc4[19]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[19]) );
  DFC1 pipe_pc4_reg_18_ ( .D(i_data_pc4[18]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[18]) );
  DFC1 pipe_pc4_reg_17_ ( .D(i_data_pc4[17]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[17]) );
  DFC1 pipe_pc4_reg_16_ ( .D(i_data_pc4[16]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[16]) );
  DFC1 pipe_pc4_reg_15_ ( .D(i_data_pc4[15]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[15]) );
  DFC1 pipe_pc4_reg_14_ ( .D(i_data_pc4[14]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[14]) );
  DFC1 pipe_pc4_reg_13_ ( .D(i_data_pc4[13]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[13]) );
  DFC1 pipe_pc4_reg_12_ ( .D(i_data_pc4[12]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[12]) );
  DFC1 pipe_pc4_reg_11_ ( .D(i_data_pc4[11]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[11]) );
  DFC1 pipe_pc4_reg_10_ ( .D(i_data_pc4[10]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[10]) );
  DFC1 pipe_pc4_reg_9_ ( .D(i_data_pc4[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[9]) );
  DFC1 pipe_pc4_reg_8_ ( .D(i_data_pc4[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[8]) );
  DFC1 pipe_pc4_reg_7_ ( .D(i_data_pc4[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[7]) );
  DFC1 pipe_pc4_reg_6_ ( .D(i_data_pc4[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[6]) );
  DFC1 pipe_pc4_reg_5_ ( .D(i_data_pc4[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[5]) );
  DFC1 pipe_pc4_reg_4_ ( .D(i_data_pc4[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[4]) );
  DFC1 pipe_pc4_reg_1_ ( .D(i_data_pc4[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[1]) );
  DFC1 pipe_pc4_reg_0_ ( .D(i_data_pc4[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[0]) );
  DFC1 pipe_alures_reg_31_ ( .D(alu_o_data_AluRes[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[31]) );
  DFC1 pipe_alures_reg_30_ ( .D(alu_o_data_AluRes[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[30]) );
  DFC1 pipe_alures_reg_29_ ( .D(alu_o_data_AluRes[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[29]) );
  DFC1 pipe_alures_reg_28_ ( .D(alu_o_data_AluRes[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[28]) );
  DFC1 pipe_alures_reg_27_ ( .D(alu_o_data_AluRes[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[27]) );
  DFC1 pipe_alures_reg_26_ ( .D(alu_o_data_AluRes[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[26]) );
  DFC1 pipe_alures_reg_25_ ( .D(alu_o_data_AluRes[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[25]) );
  DFC1 pipe_alures_reg_24_ ( .D(alu_o_data_AluRes[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[24]) );
  DFC1 pipe_alures_reg_23_ ( .D(alu_o_data_AluRes[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[23]) );
  DFC1 pipe_alures_reg_22_ ( .D(alu_o_data_AluRes[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[22]) );
  DFC1 pipe_alures_reg_21_ ( .D(alu_o_data_AluRes[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[21]) );
  DFC1 pipe_alures_reg_20_ ( .D(alu_o_data_AluRes[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[20]) );
  DFC1 pipe_alures_reg_19_ ( .D(alu_o_data_AluRes[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[19]) );
  DFC1 pipe_alures_reg_18_ ( .D(alu_o_data_AluRes[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[18]) );
  DFC1 pipe_alures_reg_17_ ( .D(alu_o_data_AluRes[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[17]) );
  DFC1 pipe_alures_reg_16_ ( .D(alu_o_data_AluRes[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[16]) );
  DFC1 pipe_alures_reg_15_ ( .D(alu_o_data_AluRes[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[15]) );
  DFC1 pipe_alures_reg_14_ ( .D(alu_o_data_AluRes[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[14]) );
  DFC1 pipe_alures_reg_13_ ( .D(alu_o_data_AluRes[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[13]) );
  DFC1 pipe_alures_reg_12_ ( .D(alu_o_data_AluRes[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[12]) );
  DFC1 pipe_alures_reg_11_ ( .D(alu_o_data_AluRes[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[11]) );
  DFC1 pipe_alures_reg_10_ ( .D(alu_o_data_AluRes[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[10]) );
  DFC1 pipe_alures_reg_9_ ( .D(alu_o_data_AluRes[9]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[9]) );
  DFC1 pipe_alures_reg_8_ ( .D(alu_o_data_AluRes[8]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[8]) );
  DFC1 pipe_alures_reg_7_ ( .D(alu_o_data_AluRes[7]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[7]) );
  DFC1 pipe_alures_reg_6_ ( .D(alu_o_data_AluRes[6]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[6]) );
  DFC1 pipe_alures_reg_5_ ( .D(alu_o_data_AluRes[5]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[5]) );
  DFC1 pipe_alures_reg_4_ ( .D(alu_o_data_AluRes[4]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[4]) );
  DFC1 pipe_alures_reg_3_ ( .D(alu_o_data_AluRes[3]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[3]) );
  DFC1 pipe_alures_reg_2_ ( .D(alu_o_data_AluRes[2]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[2]) );
  DFC1 pipe_alures_reg_1_ ( .D(alu_o_data_AluRes[1]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[1]) );
  DFC1 pipe_alures_reg_0_ ( .D(alu_o_data_AluRes[0]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_alures[0]) );
  DFC1 pipe_rt_reg_31_ ( .D(compare_i_data_rt[31]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[31]) );
  DFC1 pipe_rt_reg_30_ ( .D(compare_i_data_rt[30]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[30]) );
  DFC1 pipe_rt_reg_29_ ( .D(compare_i_data_rt[29]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[29]) );
  DFC1 pipe_rt_reg_28_ ( .D(compare_i_data_rt[28]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[28]) );
  DFC1 pipe_rt_reg_27_ ( .D(compare_i_data_rt[27]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[27]) );
  DFC1 pipe_rt_reg_26_ ( .D(compare_i_data_rt[26]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[26]) );
  DFC1 pipe_rt_reg_25_ ( .D(compare_i_data_rt[25]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[25]) );
  DFC1 pipe_rt_reg_24_ ( .D(compare_i_data_rt[24]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[24]) );
  DFC1 pipe_rt_reg_23_ ( .D(compare_i_data_rt[23]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[23]) );
  DFC1 pipe_rt_reg_22_ ( .D(compare_i_data_rt[22]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[22]) );
  DFC1 pipe_rt_reg_21_ ( .D(compare_i_data_rt[21]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[21]) );
  DFC1 pipe_rt_reg_20_ ( .D(compare_i_data_rt[20]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[20]) );
  DFC1 pipe_rt_reg_19_ ( .D(compare_i_data_rt[19]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[19]) );
  DFC1 pipe_rt_reg_18_ ( .D(compare_i_data_rt[18]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[18]) );
  DFC1 pipe_rt_reg_17_ ( .D(compare_i_data_rt[17]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[17]) );
  DFC1 pipe_rt_reg_16_ ( .D(compare_i_data_rt[16]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[16]) );
  DFC1 pipe_rt_reg_15_ ( .D(compare_i_data_rt[15]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[15]) );
  DFC1 pipe_rt_reg_14_ ( .D(compare_i_data_rt[14]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[14]) );
  DFC1 pipe_rt_reg_13_ ( .D(compare_i_data_rt[13]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[13]) );
  DFC1 pipe_rt_reg_12_ ( .D(compare_i_data_rt[12]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[12]) );
  DFC1 pipe_rt_reg_11_ ( .D(compare_i_data_rt[11]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[11]) );
  DFC1 pipe_rt_reg_10_ ( .D(compare_i_data_rt[10]), .C(i_clk), .RN(i_nrst), 
        .Q(o_data_rt[10]) );
  DFC1 pipe_rt_reg_9_ ( .D(compare_i_data_rt[9]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[9]) );
  DFC1 pipe_rt_reg_8_ ( .D(compare_i_data_rt[8]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[8]) );
  DFC1 pipe_rt_reg_7_ ( .D(compare_i_data_rt[7]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[7]) );
  DFC1 pipe_rt_reg_6_ ( .D(compare_i_data_rt[6]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[6]) );
  DFC1 pipe_rt_reg_5_ ( .D(compare_i_data_rt[5]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[5]) );
  DFC1 pipe_rt_reg_4_ ( .D(compare_i_data_rt[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[4]) );
  DFC1 pipe_rt_reg_3_ ( .D(compare_i_data_rt[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[3]) );
  DFC1 pipe_rt_reg_2_ ( .D(compare_i_data_rt[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[2]) );
  DFC1 pipe_rt_reg_1_ ( .D(compare_i_data_rt[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[1]) );
  DFC1 pipe_rt_reg_0_ ( .D(compare_i_data_rt[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_rt[0]) );
  DFC1 pipe_regdst_reg_4_ ( .D(o_addr_Erd[4]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[4]) );
  DFC1 pipe_regdst_reg_3_ ( .D(o_addr_Erd[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[3]) );
  DFC1 pipe_regdst_reg_2_ ( .D(o_addr_Erd[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[2]) );
  DFC1 pipe_regdst_reg_1_ ( .D(o_addr_Erd[1]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[1]) );
  DFC1 pipe_regdst_reg_0_ ( .D(o_addr_Erd[0]), .C(i_clk), .RN(i_nrst), .Q(
        o_addr_regdst[0]) );
  DFC1 pipe_con_Mmemread_reg ( .D(i_con_Mmemread), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Mmemread) );
  DFC1 pipe_con_Mmemwrite_reg ( .D(i_con_Mmemwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Mmemwrite) );
  DFC1 pipe_con_Wmemtoreg_reg ( .D(i_con_Wmemtoreg), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wmemtoreg) );
  DFC1 pipe_con_Wregwrite_reg ( .D(i_con_Wregwrite), .C(i_clk), .RN(i_nrst), 
        .Q(o_con_Wregwrite) );
  DFC3 pipe_pc4_reg_2_ ( .D(i_data_pc4[2]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[2]) );
  DFC3 pipe_pc4_reg_3_ ( .D(i_data_pc4[3]), .C(i_clk), .RN(i_nrst), .Q(
        o_data_pc4[3]) );
  DFC3 pipe_con_Malupc8_reg ( .D(i_con_Malupc8), .C(i_clk), .RN(i_nrst), .Q(
        o_con_Malupc8) );
  AOI210 u_alu_add_x_1_U19 ( .A(u_alu_add_x_1_n29), .B(u_alu_add_x_1_n20), .C(
        u_alu_add_x_1_n21), .Q(u_alu_add_x_1_n19) );
  XNR21 u_alu_add_x_1_U34 ( .A(u_alu_add_x_1_n5), .B(u_alu_add_x_1_n35), .Q(
        u_alu_sum_1_3_) );
  XNR21 u_alu_add_x_1_U26 ( .A(u_alu_add_x_1_n4), .B(u_alu_add_x_1_n29), .Q(
        u_alu_sum_1_4_) );
  NAND20 u_alu_add_x_1_U8 ( .A(u_alu_add_x_1_n44), .B(u_alu_add_x_1_n15), .Q(
        u_alu_add_x_1_n1) );
  OAI210 u_alu_add_x_1_U13 ( .A(u_alu_add_x_1_n17), .B(u_alu_add_x_1_n19), .C(
        u_alu_add_x_1_n18), .Q(u_alu_add_x_1_n16) );
  XNR21 u_alu_add_x_1_U2 ( .A(u_alu_add_x_1_n1), .B(u_alu_add_x_1_n16), .Q(
        u_alu_sum_1_7_) );
  NAND22 u_alu_add_x_1_U4 ( .A(u_alu_add_x_1_n20), .B(u_alu_add_x_1_n12), .Q(
        u_alu_add_x_1_n10) );
  NAND22 u_alu_add_x_1_U60 ( .A(alu_i_data_B[0]), .B(compare_i_data_rs[0]), 
        .Q(u_alu_add_x_1_n43) );
  OAI212 u_alu_add_x_1_U51 ( .A(u_alu_add_x_1_n43), .B(u_alu_add_x_1_n40), .C(
        u_alu_add_x_1_n41), .Q(u_alu_add_x_1_n39) );
  OAI212 u_alu_add_x_1_U21 ( .A(u_alu_add_x_1_n28), .B(u_alu_add_x_1_n22), .C(
        u_alu_add_x_1_n23), .Q(u_alu_add_x_1_n21) );
  OAI212 u_alu_add_x_1_U3 ( .A(u_alu_add_x_1_n10), .B(u_alu_add_x_1_n30), .C(
        u_alu_add_x_1_n11), .Q(u_alu_sum_1_8_) );
  AOI211 u_alu_add_x_1_U27 ( .A(u_alu_add_x_1_n29), .B(u_alu_add_x_1_n47), .C(
        u_alu_add_x_1_n26), .Q(u_alu_add_x_1_n24) );
  XOR21 u_alu_add_x_1_U18 ( .A(u_alu_add_x_1_n3), .B(u_alu_add_x_1_n24), .Q(
        u_alu_sum_1_5_) );
  XOR21 u_alu_add_x_1_U12 ( .A(u_alu_add_x_1_n2), .B(u_alu_add_x_1_n19), .Q(
        u_alu_sum_1_6_) );
  XOR21 u_alu_add_x_1_U43 ( .A(u_alu_add_x_1_n6), .B(u_alu_add_x_1_n38), .Q(
        u_alu_sum_1_2_) );
  NOR21 u_alu_add_x_1_U54 ( .A(compare_i_data_rs[1]), .B(u_alu_lt_x_11_B_1_), 
        .Q(u_alu_add_x_1_n40) );
  NAND22 u_alu_add_x_1_U55 ( .A(u_alu_lt_x_11_B_1_), .B(compare_i_data_rs[1]), 
        .Q(u_alu_add_x_1_n41) );
  NAND22 u_alu_add_x_1_U42 ( .A(alu_i_data_B[3]), .B(compare_i_data_rs[3]), 
        .Q(u_alu_add_x_1_n34) );
  OAI212 u_alu_add_x_1_U38 ( .A(u_alu_add_x_1_n37), .B(u_alu_add_x_1_n33), .C(
        u_alu_add_x_1_n34), .Q(u_alu_add_x_1_n32) );
  NAND22 u_alu_add_x_1_U33 ( .A(alu_i_data_B[4]), .B(compare_i_data_rs[4]), 
        .Q(u_alu_add_x_1_n28) );
  NAND22 u_alu_add_x_1_U17 ( .A(alu_i_data_B[6]), .B(compare_i_data_rs[6]), 
        .Q(u_alu_add_x_1_n18) );
  AOI212 u_alu_add_x_1_U36 ( .A(u_alu_add_x_1_n39), .B(u_alu_add_x_1_n31), .C(
        u_alu_add_x_1_n32), .Q(u_alu_add_x_1_n30) );
  NAND20 u_alu_add_x_1_U22 ( .A(u_alu_add_x_1_n46), .B(u_alu_add_x_1_n23), .Q(
        u_alu_add_x_1_n3) );
  XOR20 u_alu_add_x_1_U49 ( .A(u_alu_add_x_1_n43), .B(u_alu_add_x_1_n7), .Q(
        u_alu_sum_1_1_) );
  NAND20 u_alu_add_x_1_U14 ( .A(u_alu_add_x_1_n45), .B(u_alu_add_x_1_n18), .Q(
        u_alu_add_x_1_n2) );
  NAND22 u_alu_add_x_1_U11 ( .A(u_alu_lt_x_11_B_7_), .B(compare_i_data_rs[7]), 
        .Q(u_alu_add_x_1_n15) );
  OAI212 u_alu_add_x_1_U7 ( .A(u_alu_add_x_1_n18), .B(u_alu_add_x_1_n14), .C(
        u_alu_add_x_1_n15), .Q(u_alu_add_x_1_n13) );
  NOR22 u_alu_add_x_1_U41 ( .A(compare_i_data_rs[3]), .B(alu_i_data_B[3]), .Q(
        u_alu_add_x_1_n33) );
  NAND22 u_alu_add_x_1_U25 ( .A(n294), .B(compare_i_data_rs[5]), .Q(
        u_alu_add_x_1_n23) );
  NOR22 u_alu_add_x_1_U24 ( .A(compare_i_data_rs[5]), .B(n294), .Q(
        u_alu_add_x_1_n22) );
  NOR22 u_alu_add_x_1_U6 ( .A(u_alu_add_x_1_n17), .B(u_alu_add_x_1_n14), .Q(
        u_alu_add_x_1_n12) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U49 ( .A(n143), .B(compare_i_data_rs[28]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n35), .CO(u_alu_DP_OP_85J3_126_1427_n34), 
        .S(u_alu_pre_suba[12]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U2 ( .A(u_alu_pre_sum_4a[6]), .B(
        u_alu_DP_OP_84J3_125_2615_n2), .CO(u_alu_DP_OP_84J3_125_2615_n1), .S(
        u_alu_pre_sum_4b[6]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U4 ( .A(u_alu_pre_sum_4a[4]), .B(
        u_alu_DP_OP_84J3_125_2615_n4), .CO(u_alu_DP_OP_84J3_125_2615_n3), .S(
        u_alu_pre_sum_4b[4]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U5 ( .A(u_alu_pre_sum_4a[3]), .B(
        u_alu_DP_OP_84J3_125_2615_n5), .CO(u_alu_DP_OP_84J3_125_2615_n4), .S(
        u_alu_pre_sum_4b[3]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U6 ( .A(u_alu_pre_sum_4a[2]), .B(
        u_alu_DP_OP_84J3_125_2615_n6), .CO(u_alu_DP_OP_84J3_125_2615_n5), .S(
        u_alu_pre_sum_4b[2]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U7 ( .A(u_alu_pre_sum_4a[1]), .B(
        u_alu_pre_sum_4a[0]), .CO(u_alu_DP_OP_84J3_125_2615_n6), .S(
        u_alu_pre_sum_4b[1]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U3 ( .A(u_alu_pre_sum_4a[5]), .B(
        u_alu_DP_OP_84J3_125_2615_n3), .CO(u_alu_DP_OP_84J3_125_2615_n2), .S(
        u_alu_pre_sum_4b[5]) );
  ADD31 u_alu_DP_OP_83J3_124_3384_U15 ( .A(compare_i_data_rs[18]), .B(
        alu_i_data_B[18]), .CI(u_alu_DP_OP_83J3_124_3384_n14), .CO(
        u_alu_DP_OP_83J3_124_3384_n13), .S(u_alu_pre_sum_3a[2]) );
  ADD31 u_alu_DP_OP_83J3_124_3384_U14 ( .A(compare_i_data_rs[19]), .B(
        alu_i_data_B[19]), .CI(u_alu_DP_OP_83J3_124_3384_n13), .CO(
        u_alu_DP_OP_83J3_124_3384_n12), .S(u_alu_pre_sum_3a[3]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U10 ( .A(compare_i_data_rs[23]), .B(
        alu_i_data_B[23]), .CI(u_alu_DP_OP_83J3_124_3384_n9), .CO(
        u_alu_pre_sum_3a[8]), .S(u_alu_pre_sum_3a[7]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U5 ( .A(u_alu_pre_sum_3a[4]), .B(
        u_alu_DP_OP_83J3_124_3384_n5), .CO(u_alu_DP_OP_83J3_124_3384_n4), .S(
        u_alu_pre_sum_3b[4]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U6 ( .A(u_alu_pre_sum_3a[3]), .B(
        u_alu_DP_OP_83J3_124_3384_n6), .CO(u_alu_DP_OP_83J3_124_3384_n5), .S(
        u_alu_pre_sum_3b[3]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U7 ( .A(u_alu_pre_sum_3a[2]), .B(
        u_alu_DP_OP_83J3_124_3384_n7), .CO(u_alu_DP_OP_83J3_124_3384_n6), .S(
        u_alu_pre_sum_3b[2]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U8 ( .A(u_alu_pre_sum_3a[1]), .B(
        u_alu_pre_sum_3a[0]), .CO(u_alu_DP_OP_83J3_124_3384_n7), .S(
        u_alu_pre_sum_3b[1]) );
  ADD31 u_alu_sub_x_2_U11 ( .A(n173), .B(compare_i_data_rs[6]), .CI(
        u_alu_sub_x_2_n12), .CO(u_alu_sub_x_2_n11), .S(u_alu_half_sub_6_) );
  AOI221 DP_OP_77_130_260_U25 ( .A(compare_i_data_rs[9]), .B(
        DP_OP_77_130_260_I3), .C(n170), .D(DP_OP_77_130_260_n39), .Q(
        DP_OP_77_130_260_n16) );
  ADD21 DP_OP_77_130_260_U34 ( .A(compare_i_data_rs[9]), .B(
        compare_i_data_rs[8]), .CO(DP_OP_77_130_260_n23), .S(
        DP_OP_77_130_260_n39) );
  ADD22 DP_OP_77_130_260_U30 ( .A(DP_OP_77_130_260_n20), .B(
        compare_i_data_rs[13]), .CO(DP_OP_77_130_260_n19), .S(
        DP_OP_77_130_260_n43) );
  ADD22 DP_OP_77_130_260_U29 ( .A(DP_OP_77_130_260_n19), .B(
        compare_i_data_rs[14]), .CO(DP_OP_77_130_260_n18), .S(
        DP_OP_77_130_260_n44) );
  AOI221 DP_OP_77_130_260_U23 ( .A(compare_i_data_rs[10]), .B(
        DP_OP_77_130_260_I3), .C(n170), .D(DP_OP_77_130_260_n40), .Q(
        DP_OP_77_130_260_n15) );
  ADD22 DP_OP_77_130_260_U28 ( .A(DP_OP_77_130_260_n18), .B(
        compare_i_data_rs[15]), .CO(DP_OP_77_130_260_n46), .S(
        DP_OP_77_130_260_n45) );
  AOI221 DP_OP_77_130_260_U21 ( .A(compare_i_data_rs[11]), .B(
        DP_OP_77_130_260_I3), .C(DP_OP_77_130_260_n41), .D(n170), .Q(
        DP_OP_77_130_260_n14) );
  AOI221 DP_OP_77_130_260_U19 ( .A(compare_i_data_rs[12]), .B(
        DP_OP_77_130_260_I3), .C(DP_OP_77_130_260_n42), .D(n170), .Q(
        DP_OP_77_130_260_n13) );
  AOI221 DP_OP_77_130_260_U17 ( .A(compare_i_data_rs[13]), .B(
        DP_OP_77_130_260_I3), .C(DP_OP_77_130_260_n43), .D(n170), .Q(
        DP_OP_77_130_260_n12) );
  INV3 DP_OP_77_130_260_U10 ( .A(DP_OP_77_130_260_n9), .Q(DP_OP_77_130_260_n37) );
  NAND22 DP_OP_77_130_260_U11 ( .A(DP_OP_77_130_260_n46), .B(n170), .Q(
        DP_OP_77_130_260_n9) );
  INV3 DP_OP_77_130_260_U26 ( .A(DP_OP_77_130_260_n17), .Q(
        DP_OP_77_130_260_n29) );
  INV3 DP_OP_77_130_260_U24 ( .A(DP_OP_77_130_260_n16), .Q(
        DP_OP_77_130_260_n30) );
  INV3 DP_OP_77_130_260_U22 ( .A(DP_OP_77_130_260_n15), .Q(
        DP_OP_77_130_260_n31) );
  INV3 DP_OP_77_130_260_U20 ( .A(DP_OP_77_130_260_n14), .Q(
        DP_OP_77_130_260_n32) );
  INV3 DP_OP_77_130_260_U18 ( .A(DP_OP_77_130_260_n13), .Q(
        DP_OP_77_130_260_n33) );
  INV3 DP_OP_77_130_260_U16 ( .A(DP_OP_77_130_260_n12), .Q(
        DP_OP_77_130_260_n34) );
  INV3 DP_OP_77_130_260_U14 ( .A(DP_OP_77_130_260_n11), .Q(
        DP_OP_77_130_260_n35) );
  AOI221 DP_OP_77_130_260_U15 ( .A(compare_i_data_rs[14]), .B(
        DP_OP_77_130_260_I3), .C(DP_OP_77_130_260_n44), .D(n170), .Q(
        DP_OP_77_130_260_n11) );
  INV3 DP_OP_77_130_260_U12 ( .A(DP_OP_77_130_260_n10), .Q(
        DP_OP_77_130_260_n36) );
  AOI221 DP_OP_77_130_260_U13 ( .A(compare_i_data_rs[15]), .B(
        DP_OP_77_130_260_I3), .C(DP_OP_77_130_260_n45), .D(n170), .Q(
        DP_OP_77_130_260_n10) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U17 ( .A(compare_i_data_rs[16]), .B(
        alu_i_data_B[16]), .CO(u_alu_DP_OP_83J3_124_3384_n15), .S(
        u_alu_pre_sum_3a[0]) );
  ADD22 u_alu_DP_OP_84J3_125_2615_U17 ( .A(compare_i_data_rs[24]), .B(
        alu_i_data_B[24]), .CO(u_alu_DP_OP_84J3_125_2615_n15), .S(
        u_alu_pre_sum_4a[0]) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U16 ( .A(compare_i_data_rs[25]), .B(
        alu_i_data_B[25]), .CI(u_alu_DP_OP_84J3_125_2615_n15), .CO(
        u_alu_DP_OP_84J3_125_2615_n14), .S(u_alu_pre_sum_4a[1]) );
  NAND21 u_alu_add_x_1_U30 ( .A(u_alu_add_x_1_n47), .B(u_alu_add_x_1_n28), .Q(
        u_alu_add_x_1_n4) );
  ADD22 DP_OP_77_130_260_U32 ( .A(DP_OP_77_130_260_n22), .B(
        compare_i_data_rs[11]), .CO(DP_OP_77_130_260_n21), .S(
        DP_OP_77_130_260_n41) );
  NAND21 u_alu_add_x_1_U39 ( .A(u_alu_add_x_1_n48), .B(u_alu_add_x_1_n34), .Q(
        u_alu_add_x_1_n5) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U15 ( .A(compare_i_data_rs[26]), .B(
        alu_i_data_B[26]), .CI(u_alu_DP_OP_84J3_125_2615_n14), .CO(
        u_alu_DP_OP_84J3_125_2615_n13), .S(u_alu_pre_sum_4a[2]) );
  ADD22 DP_OP_77_130_260_U31 ( .A(DP_OP_77_130_260_n21), .B(
        compare_i_data_rs[12]), .CO(DP_OP_77_130_260_n20), .S(
        DP_OP_77_130_260_n42) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U14 ( .A(compare_i_data_rs[27]), .B(
        alu_i_data_B[27]), .CI(u_alu_DP_OP_84J3_125_2615_n13), .CO(
        u_alu_DP_OP_84J3_125_2615_n12), .S(u_alu_pre_sum_4a[3]) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U13 ( .A(compare_i_data_rs[28]), .B(
        alu_i_data_B[28]), .CI(u_alu_DP_OP_84J3_125_2615_n12), .CO(
        u_alu_DP_OP_84J3_125_2615_n11), .S(u_alu_pre_sum_4a[4]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U13 ( .A(compare_i_data_rs[20]), .B(
        alu_i_data_B[20]), .CI(u_alu_DP_OP_83J3_124_3384_n12), .CO(
        u_alu_DP_OP_83J3_124_3384_n11), .S(u_alu_pre_sum_3a[4]) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U12 ( .A(compare_i_data_rs[29]), .B(
        alu_i_data_B[29]), .CI(u_alu_DP_OP_84J3_125_2615_n11), .CO(
        u_alu_DP_OP_84J3_125_2615_n10), .S(u_alu_pre_sum_4a[5]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U12 ( .A(compare_i_data_rs[21]), .B(
        alu_i_data_B[21]), .CI(u_alu_DP_OP_83J3_124_3384_n11), .CO(
        u_alu_DP_OP_83J3_124_3384_n10), .S(u_alu_pre_sum_3a[5]) );
  ADD32 u_alu_DP_OP_84J3_125_2615_U11 ( .A(compare_i_data_rs[30]), .B(
        alu_i_data_B[30]), .CI(u_alu_DP_OP_84J3_125_2615_n10), .CO(
        u_alu_DP_OP_84J3_125_2615_n9), .S(u_alu_pre_sum_4a[6]) );
  ADD32 u_alu_DP_OP_83J3_124_3384_U11 ( .A(compare_i_data_rs[22]), .B(
        alu_i_data_B[22]), .CI(u_alu_DP_OP_83J3_124_3384_n10), .CO(
        u_alu_DP_OP_83J3_124_3384_n9), .S(u_alu_pre_sum_3a[6]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U4 ( .A(u_alu_pre_sum_3a[5]), .B(
        u_alu_DP_OP_83J3_124_3384_n4), .CO(u_alu_DP_OP_83J3_124_3384_n3), .S(
        u_alu_pre_sum_3b[5]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U3 ( .A(u_alu_pre_sum_3a[6]), .B(
        u_alu_DP_OP_83J3_124_3384_n3), .CO(u_alu_DP_OP_83J3_124_3384_n2), .S(
        u_alu_pre_sum_3b[6]) );
  ADD32 u_alu_DP_OP_85J3_126_1427_U56 ( .A(n127), .B(compare_i_data_rs[21]), 
        .CI(u_alu_DP_OP_85J3_126_1427_n42), .CO(u_alu_DP_OP_85J3_126_1427_n41), 
        .S(u_alu_pre_suba[5]) );
  ADD22 u_alu_DP_OP_83J3_124_3384_U2 ( .A(u_alu_pre_sum_3a[7]), .B(
        u_alu_DP_OP_83J3_124_3384_n2), .CO(u_alu_DP_OP_83J3_124_3384_n1), .S(
        u_alu_pre_sum_3b[7]) );
  NAND20 u_alu_add_x_1_U45 ( .A(u_alu_add_x_1_n49), .B(u_alu_add_x_1_n37), .Q(
        u_alu_add_x_1_n6) );
  NAND20 u_alu_add_x_1_U52 ( .A(u_alu_add_x_1_n50), .B(u_alu_add_x_1_n41), .Q(
        u_alu_add_x_1_n7) );
  ADD22 DP_OP_77_130_260_U33 ( .A(DP_OP_77_130_260_n23), .B(
        compare_i_data_rs[10]), .CO(DP_OP_77_130_260_n22), .S(
        DP_OP_77_130_260_n40) );
  NAND24 U3 ( .A(n808), .B(n807), .Q(alu_i_data_B[16]) );
  BUF6 U4 ( .A(n861), .Q(n168) );
  AOI211 U5 ( .A(n1168), .B(u_alu_pre_sum_4a[2]), .C(n1117), .Q(n1119) );
  INV6 U6 ( .A(n839), .Q(n300) );
  INV3 U7 ( .A(compare_i_data_rs[16]), .Q(n138) );
  NOR22 U8 ( .A(u_alu_add_x_1_n27), .B(u_alu_add_x_1_n22), .Q(
        u_alu_add_x_1_n20) );
  INV3 U9 ( .A(alu_i_data_B[2]), .Q(n133) );
  BUF2 U10 ( .A(n839), .Q(n299) );
  BUF2 U11 ( .A(n842), .Q(n298) );
  NAND33 U12 ( .A(n725), .B(n724), .C(n723), .Q(compare_i_data_rs[0]) );
  MUX22 U13 ( .A(compare_i_data_rt[4]), .B(i_data_immext[4]), .S(n305), .Q(
        alu_i_data_B[4]) );
  NOR21 U14 ( .A(n880), .B(n881), .Q(n1179) );
  INV3 U15 ( .A(n576), .Q(n141) );
  BUF2 U16 ( .A(n1181), .Q(n575) );
  NAND41 U17 ( .A(n1102), .B(n1101), .C(n1100), .D(n1099), .Q(n1103) );
  NAND41 U18 ( .A(n1130), .B(n1129), .C(n1128), .D(n1127), .Q(n1131) );
  INV8 U19 ( .A(n574), .Q(n140) );
  BUF6 U20 ( .A(n722), .Q(n169) );
  NAND31 U21 ( .A(n851), .B(n850), .C(n849), .Q(compare_i_data_rt[5]) );
  NAND31 U22 ( .A(n797), .B(n796), .C(n795), .Q(compare_i_data_rt[18]) );
  OAI2111 U23 ( .A(u_alu_pre_subb[0]), .B(n304), .C(n1012), .D(n1011), .Q(
        alu_o_data_AluRes[16]) );
  AOI211 U24 ( .A(n1158), .B(u_alu_pre_subb[8]), .C(n1091), .Q(n1093) );
  NAND31 U25 ( .A(n1120), .B(n1119), .C(n1118), .Q(alu_o_data_AluRes[26]) );
  CLKIN0 U26 ( .A(alu_i_con_AluCtrl[0]), .Q(n1) );
  CLKIN0 U27 ( .A(compare_i_data_rs[29]), .Q(n2) );
  AOI2110 U28 ( .A(n1), .B(n2), .C(n129), .D(n1184), .Q(n3) );
  IMUX20 U29 ( .A(n2), .B(compare_i_data_rs[29]), .S(alu_i_data_B[29]), .Q(n4)
         );
  AOI220 U30 ( .A(compare_i_data_rs[29]), .B(n141), .C(n1179), .D(n4), .Q(n5)
         );
  OAI310 U31 ( .A(alu_i_data_B[29]), .B(compare_i_data_rs[29]), .C(n1144), .D(
        n5), .Q(n6) );
  AOI2110 U32 ( .A(alu_i_data_B[13]), .B(n1161), .C(n3), .D(n6), .Q(n1148) );
  MUX22 U33 ( .A(compare_i_data_rt[7]), .B(u_alu_ashr_4_SH_1_), .S(n305), .Q(
        u_alu_lt_x_11_B_7_) );
  CLKIN0 U34 ( .A(u_alu_half_sub_11_), .Q(n7) );
  NOR20 U35 ( .A(n303), .B(compare_i_data_rs[11]), .Q(n8) );
  AOI2110 U36 ( .A(compare_i_data_rs[11]), .B(n577), .C(n141), .D(n8), .Q(n9)
         );
  NOR20 U37 ( .A(alu_i_data_B[11]), .B(n1144), .Q(n10) );
  OAI210 U38 ( .A(alu_i_data_B[11]), .B(n303), .C(n576), .Q(n11) );
  IMUX20 U39 ( .A(n10), .B(n11), .S(compare_i_data_rs[11]), .Q(n12) );
  IMUX20 U40 ( .A(n530), .B(n489), .S(u_alu_ashr_4_SH_3_), .Q(n13) );
  MUX21 U41 ( .A(n13), .B(n511), .S(i_data_immext[10]), .Q(n14) );
  NAND20 U42 ( .A(n1180), .B(n14), .Q(n15) );
  OAI2110 U43 ( .A(n134), .B(n9), .C(n12), .D(n15), .Q(n16) );
  AOI210 U44 ( .A(u_alu_N168), .B(n998), .C(n16), .Q(n17) );
  CLKIN0 U45 ( .A(n437), .Q(n18) );
  NAND30 U46 ( .A(n575), .B(n390), .C(n18), .Q(n19) );
  OAI2110 U47 ( .A(n999), .B(n7), .C(n17), .D(n19), .Q(alu_o_data_AluRes[11])
         );
  IMUX20 U48 ( .A(n375), .B(n378), .S(u_alu_ashr_4_SH_3_), .Q(n20) );
  IMUX20 U49 ( .A(n20), .B(n345), .S(n437), .Q(n21) );
  CLKIN0 U50 ( .A(n575), .Q(n22) );
  CLKIN0 U51 ( .A(compare_i_data_rs[17]), .Q(n23) );
  IMUX20 U52 ( .A(compare_i_data_rs[17]), .B(n23), .S(alu_i_data_B[17]), .Q(
        n24) );
  OAI220 U53 ( .A(n303), .B(n24), .C(n171), .D(n1023), .Q(n25) );
  AOI210 U54 ( .A(compare_i_data_rs[17]), .B(n141), .C(n25), .Q(n26) );
  CLKIN0 U55 ( .A(i_data_immext[10]), .Q(n27) );
  CLKIN0 U56 ( .A(n1184), .Q(n28) );
  OAI2110 U57 ( .A(compare_i_data_rs[17]), .B(alu_i_con_AluCtrl[0]), .C(
        alu_i_data_B[17]), .D(n28), .Q(n29) );
  OAI310 U58 ( .A(alu_i_data_B[17]), .B(compare_i_data_rs[17]), .C(n1144), .D(
        n29), .Q(n30) );
  AOI310 U59 ( .A(n1180), .B(n495), .C(n27), .D(n30), .Q(n31) );
  OAI2110 U60 ( .A(n21), .B(n22), .C(n26), .D(n31), .Q(n1013) );
  CLKIN0 U61 ( .A(u_alu_half_sub_12_), .Q(n32) );
  NOR30 U62 ( .A(alu_i_data_B[12]), .B(compare_i_data_rs[12]), .C(n1144), .Q(
        n33) );
  NOR20 U63 ( .A(n303), .B(compare_i_data_rs[12]), .Q(n34) );
  AOI2110 U64 ( .A(compare_i_data_rs[12]), .B(n577), .C(n141), .D(n34), .Q(n35) );
  OAI210 U65 ( .A(alu_i_data_B[12]), .B(n303), .C(n576), .Q(n36) );
  IMUX20 U66 ( .A(n534), .B(n499), .S(u_alu_ashr_4_SH_3_), .Q(n37) );
  IMUX20 U67 ( .A(n37), .B(n512), .S(i_data_immext[10]), .Q(n38) );
  AOI220 U68 ( .A(compare_i_data_rs[12]), .B(n36), .C(n1180), .D(n38), .Q(n39)
         );
  OAI210 U69 ( .A(n137), .B(n35), .C(n39), .Q(n40) );
  AOI2110 U70 ( .A(n998), .B(u_alu_N169), .C(n33), .D(n40), .Q(n41) );
  CLKIN0 U71 ( .A(i_data_immext[10]), .Q(n42) );
  NAND30 U72 ( .A(n575), .B(n397), .C(n42), .Q(n43) );
  OAI2110 U73 ( .A(n999), .B(n32), .C(n41), .D(n43), .Q(alu_o_data_AluRes[12])
         );
  IMUX20 U74 ( .A(n382), .B(n339), .S(u_alu_ashr_4_SH_3_), .Q(n44) );
  IMUX20 U75 ( .A(n44), .B(n406), .S(n437), .Q(n45) );
  CLKIN0 U76 ( .A(n575), .Q(n46) );
  CLKIN0 U77 ( .A(compare_i_data_rs[18]), .Q(n47) );
  IMUX20 U78 ( .A(compare_i_data_rs[18]), .B(n47), .S(alu_i_data_B[18]), .Q(
        n48) );
  OAI220 U79 ( .A(n303), .B(n48), .C(n133), .D(n1023), .Q(n49) );
  AOI210 U80 ( .A(compare_i_data_rs[18]), .B(n141), .C(n49), .Q(n50) );
  CLKIN0 U81 ( .A(i_data_immext[10]), .Q(n51) );
  CLKIN0 U82 ( .A(n1184), .Q(n52) );
  OAI2110 U83 ( .A(compare_i_data_rs[18]), .B(alu_i_con_AluCtrl[0]), .C(
        alu_i_data_B[18]), .D(n52), .Q(n53) );
  OAI310 U84 ( .A(alu_i_data_B[18]), .B(compare_i_data_rs[18]), .C(n1144), .D(
        n53), .Q(n54) );
  AOI310 U85 ( .A(n1180), .B(n521), .C(n51), .D(n54), .Q(n55) );
  OAI2110 U86 ( .A(n45), .B(n46), .C(n50), .D(n55), .Q(n1018) );
  AOI2110 U87 ( .A(compare_i_data_rs[21]), .B(n141), .C(n1046), .D(n1047), .Q(
        n56) );
  AOI220 U88 ( .A(n1180), .B(u_alu_N246), .C(n575), .D(u_alu_N214), .Q(n57) );
  NAND30 U89 ( .A(n56), .B(n1048), .C(n57), .Q(n1049) );
  CLKIN0 U90 ( .A(u_alu_half_sub_13_), .Q(n58) );
  NOR20 U91 ( .A(n303), .B(compare_i_data_rs[13]), .Q(n59) );
  AOI2110 U92 ( .A(compare_i_data_rs[13]), .B(n577), .C(n141), .D(n59), .Q(n60) );
  OAI210 U93 ( .A(alu_i_data_B[13]), .B(n303), .C(n576), .Q(n61) );
  NOR20 U94 ( .A(alu_i_data_B[13]), .B(n1144), .Q(n62) );
  IMUX20 U95 ( .A(n62), .B(n61), .S(compare_i_data_rs[13]), .Q(n63) );
  IMUX20 U96 ( .A(n541), .B(n501), .S(u_alu_ashr_4_SH_3_), .Q(n64) );
  MUX21 U97 ( .A(n64), .B(n513), .S(i_data_immext[10]), .Q(n65) );
  NAND20 U98 ( .A(n1180), .B(n65), .Q(n66) );
  OAI2110 U99 ( .A(n162), .B(n60), .C(n63), .D(n66), .Q(n67) );
  AOI210 U100 ( .A(n998), .B(u_alu_N170), .C(n67), .Q(n68) );
  CLKIN0 U101 ( .A(n437), .Q(n69) );
  NAND30 U102 ( .A(n575), .B(n404), .C(n69), .Q(n70) );
  OAI2110 U103 ( .A(n999), .B(n58), .C(n68), .D(n70), .Q(alu_o_data_AluRes[13]) );
  NOR20 U104 ( .A(n914), .B(n921), .Q(n71) );
  AOI310 U105 ( .A(n1247), .B(n913), .C(n71), .D(i_data_immext[4]), .Q(n1177)
         );
  OAI210 U106 ( .A(alu_i_data_B[0]), .B(compare_i_data_rs[0]), .C(
        u_alu_add_x_1_n43), .Q(u_alu_add_x_1_n8) );
  IMUX20 U107 ( .A(n388), .B(n343), .S(u_alu_ashr_4_SH_3_), .Q(n72) );
  IMUX20 U108 ( .A(n72), .B(n419), .S(n437), .Q(n73) );
  CLKIN0 U109 ( .A(n575), .Q(n74) );
  CLKIN0 U110 ( .A(compare_i_data_rs[19]), .Q(n75) );
  IMUX20 U111 ( .A(compare_i_data_rs[19]), .B(n75), .S(alu_i_data_B[19]), .Q(
        n76) );
  OAI220 U112 ( .A(n303), .B(n76), .C(n153), .D(n1023), .Q(n77) );
  AOI210 U113 ( .A(compare_i_data_rs[19]), .B(n141), .C(n77), .Q(n78) );
  CLKIN0 U114 ( .A(i_data_immext[10]), .Q(n79) );
  CLKIN0 U115 ( .A(n1184), .Q(n80) );
  OAI2110 U116 ( .A(compare_i_data_rs[19]), .B(alu_i_con_AluCtrl[0]), .C(
        alu_i_data_B[19]), .D(n80), .Q(n81) );
  OAI310 U117 ( .A(alu_i_data_B[19]), .B(compare_i_data_rs[19]), .C(n1144), 
        .D(n81), .Q(n82) );
  AOI310 U118 ( .A(n1180), .B(n532), .C(n79), .D(n82), .Q(n83) );
  OAI2110 U119 ( .A(n73), .B(n74), .C(n78), .D(n83), .Q(n1024) );
  AOI2110 U120 ( .A(compare_i_data_rs[22]), .B(n141), .C(n1056), .D(n1057), 
        .Q(n84) );
  AOI220 U121 ( .A(n1180), .B(u_alu_N247), .C(n575), .D(u_alu_N215), .Q(n85)
         );
  NAND30 U122 ( .A(n84), .B(n1058), .C(n85), .Q(n1059) );
  NAND22 U123 ( .A(u_alu_pre_sum_4b[4]), .B(n1167), .Q(n86) );
  AOI220 U124 ( .A(n575), .B(u_alu_N221), .C(n1180), .D(u_alu_N253), .Q(n87)
         );
  AOI2110 U125 ( .A(compare_i_data_rs[28]), .B(n141), .C(n1138), .D(n1139), 
        .Q(n88) );
  NAND30 U126 ( .A(n86), .B(n87), .C(n88), .Q(n1140) );
  NAND20 U127 ( .A(i_data_FWmemout[2]), .B(n863), .Q(n89) );
  AOI221 U128 ( .A(n301), .B(i_data_FMmemout[2]), .C(n139), .D(i_data_rt[2]), 
        .Q(n90) );
  AOI220 U129 ( .A(n302), .B(i_data_FMalures[2]), .C(n300), .D(
        i_data_FEalures[2]), .Q(n91) );
  NAND31 U130 ( .A(n89), .B(n90), .C(n91), .Q(compare_i_data_rt[2]) );
  CLKIN0 U131 ( .A(u_alu_half_sub_14_), .Q(n92) );
  AOI2110 U132 ( .A(compare_i_data_rs[14]), .B(n577), .C(n141), .D(n990), .Q(
        n93) );
  IMUX20 U133 ( .A(n475), .B(n523), .S(i_data_immext[10]), .Q(n94) );
  AOI220 U134 ( .A(compare_i_data_rs[14]), .B(n992), .C(n1180), .D(n94), .Q(
        n95) );
  OAI210 U135 ( .A(n156), .B(n93), .C(n95), .Q(n96) );
  AOI2110 U136 ( .A(n998), .B(u_alu_N171), .C(n991), .D(n96), .Q(n97) );
  CLKIN0 U137 ( .A(i_data_immext[10]), .Q(n98) );
  NAND30 U138 ( .A(n575), .B(n410), .C(n98), .Q(n99) );
  OAI2110 U139 ( .A(n999), .B(n92), .C(n97), .D(n99), .Q(alu_o_data_AluRes[14]) );
  OAI210 U140 ( .A(n440), .B(n311), .C(i_data_immext[8]), .Q(n100) );
  OAI210 U141 ( .A(n328), .B(i_data_immext[8]), .C(n100), .Q(n349) );
  CLKIN0 U142 ( .A(i_data_immext[10]), .Q(n101) );
  NAND30 U143 ( .A(n1180), .B(n510), .C(n101), .Q(n1115) );
  CLKIN0 U144 ( .A(i_data_immext[10]), .Q(n102) );
  NAND30 U145 ( .A(n1180), .B(n513), .C(n102), .Q(n1146) );
  AOI2110 U146 ( .A(compare_i_data_rs[23]), .B(n141), .C(n1066), .D(n1067), 
        .Q(n103) );
  AOI220 U147 ( .A(n1180), .B(u_alu_N248), .C(n575), .D(u_alu_N216), .Q(n104)
         );
  NAND30 U148 ( .A(n103), .B(n1068), .C(n104), .Q(n1069) );
  CLKIN0 U149 ( .A(n575), .Q(n105) );
  IMUX20 U150 ( .A(alu_i_data_B[30]), .B(alu_i_data_B[29]), .S(
        i_data_immext[6]), .Q(n106) );
  IMUX20 U151 ( .A(n106), .B(n407), .S(n440), .Q(n107) );
  IMUX20 U152 ( .A(n107), .B(n408), .S(i_data_immext[8]), .Q(n108) );
  IMUX20 U153 ( .A(n108), .B(n409), .S(u_alu_ashr_4_SH_3_), .Q(n109) );
  IMUX20 U154 ( .A(n109), .B(n410), .S(n437), .Q(n110) );
  NOR20 U155 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[30]), .Q(n111)
         );
  NAND20 U156 ( .A(alu_i_data_B[14]), .B(n1161), .Q(n112) );
  OAI310 U157 ( .A(n1184), .B(n111), .C(n130), .D(n112), .Q(n113) );
  CLKIN0 U158 ( .A(n1180), .Q(n114) );
  CLKIN0 U159 ( .A(n1179), .Q(n115) );
  IMAJ30 U160 ( .A(n115), .B(alu_i_data_B[30]), .C(compare_i_data_rs[30]), .Q(
        n116) );
  OAI310 U161 ( .A(alu_i_data_B[30]), .B(compare_i_data_rs[30]), .C(n1178), 
        .D(n116), .Q(n117) );
  OAI310 U162 ( .A(i_data_immext[10]), .B(n523), .C(n114), .D(n117), .Q(n118)
         );
  AOI2110 U163 ( .A(compare_i_data_rs[30]), .B(n141), .C(n113), .D(n118), .Q(
        n119) );
  OAI210 U164 ( .A(n105), .B(n110), .C(n119), .Q(n1153) );
  CLKIN0 U165 ( .A(u_alu_half_sub_15_), .Q(n120) );
  NAND20 U166 ( .A(n1180), .B(u_alu_N240), .Q(n121) );
  OAI2110 U167 ( .A(n135), .B(n997), .C(n996), .D(n121), .Q(n122) );
  AOI210 U168 ( .A(u_alu_N172), .B(n998), .C(n122), .Q(n123) );
  CLKIN0 U169 ( .A(i_data_immext[10]), .Q(n124) );
  NAND30 U170 ( .A(n575), .B(n417), .C(n124), .Q(n125) );
  OAI2110 U171 ( .A(n999), .B(n120), .C(n123), .D(n125), .Q(
        alu_o_data_AluRes[15]) );
  NOR24 U172 ( .A(i_con_Efamux[2]), .B(i_con_Efamux[0]), .Q(n581) );
  NAND33 U173 ( .A(n648), .B(n647), .C(n646), .Q(compare_i_data_rs[16]) );
  NOR23 U174 ( .A(compare_i_data_rs[6]), .B(alu_i_data_B[6]), .Q(
        u_alu_add_x_1_n17) );
  NOR24 U175 ( .A(n582), .B(n573), .Q(n720) );
  NAND33 U176 ( .A(n285), .B(n284), .C(n176), .Q(u_alu_DP_OP_85J3_126_1427_n33) );
  NOR22 U177 ( .A(compare_i_data_rs[4]), .B(alu_i_data_B[4]), .Q(
        u_alu_add_x_1_n27) );
  MUX21 U178 ( .A(n905), .B(n904), .S(compare_i_data_rs[0]), .Q(n908) );
  AOI210 U179 ( .A(n297), .B(i_data_rs[15]), .C(n650), .Q(n651) );
  AOI210 U180 ( .A(n297), .B(i_data_rs[13]), .C(n656), .Q(n657) );
  AOI210 U181 ( .A(n297), .B(i_data_rs[11]), .C(n662), .Q(n663) );
  AOI210 U182 ( .A(n297), .B(i_data_rs[28]), .C(n595), .Q(n596) );
  AOI210 U183 ( .A(n297), .B(i_data_rs[22]), .C(n613), .Q(n614) );
  AOI210 U184 ( .A(n297), .B(i_data_rs[10]), .C(n665), .Q(n666) );
  AOI210 U185 ( .A(n297), .B(i_data_rs[21]), .C(n616), .Q(n617) );
  AOI210 U186 ( .A(n297), .B(i_data_rs[31]), .C(n586), .Q(n587) );
  AOI210 U187 ( .A(n297), .B(i_data_rs[30]), .C(n589), .Q(n590) );
  AOI210 U188 ( .A(n297), .B(i_data_rs[8]), .C(n671), .Q(n672) );
  AOI210 U189 ( .A(n297), .B(i_data_rs[9]), .C(n668), .Q(n669) );
  AOI210 U190 ( .A(n297), .B(i_data_rs[24]), .C(n607), .Q(n608) );
  AOI210 U191 ( .A(n297), .B(i_data_rs[27]), .C(n598), .Q(n599) );
  AOI210 U192 ( .A(n297), .B(i_data_rs[26]), .C(n601), .Q(n602) );
  AOI210 U193 ( .A(n297), .B(i_data_rs[25]), .C(n604), .Q(n605) );
  INV6 U194 ( .A(compare_i_data_rs[0]), .Q(n152) );
  NAND26 U195 ( .A(n693), .B(n692), .Q(compare_i_data_rs[5]) );
  NAND28 U196 ( .A(n1076), .B(n1075), .Q(n1167) );
  NAND24 U197 ( .A(u_alu_pre_sum_3a[8]), .B(n1074), .Q(n1075) );
  NAND28 U198 ( .A(n719), .B(n718), .Q(compare_i_data_rs[1]) );
  NAND23 U199 ( .A(n296), .B(i_data_rs[1]), .Q(n719) );
  ADD32 U200 ( .A(n150), .B(compare_i_data_rs[4]), .CI(u_alu_sub_x_2_n14), 
        .CO(u_alu_sub_x_2_n13), .S(u_alu_half_sub_4_) );
  NOR24 U201 ( .A(n999), .B(u_alu_half_sub_16_), .Q(n1174) );
  NAND42 U202 ( .A(n1172), .B(n1171), .C(n1170), .D(n1169), .Q(n1173) );
  CLKIN4 U203 ( .A(u_alu_sub_x_2_n2), .Q(u_alu_half_sub_16_) );
  OAI2110 U204 ( .A(compare_i_data_rs[4]), .B(n1205), .C(n1206), .D(n1207), 
        .Q(alu_o_data_AluRes[4]) );
  AOI210 U205 ( .A(u_alu_pre_sum_3b[4]), .B(n1073), .C(n1038), .Q(n1040) );
  AOI210 U206 ( .A(u_alu_pre_sum_3b[6]), .B(n1073), .C(n1059), .Q(n1061) );
  AOI210 U207 ( .A(u_alu_pre_sum_3b[5]), .B(n1073), .C(n1049), .Q(n1051) );
  AOI210 U208 ( .A(u_alu_pre_sum_3b[7]), .B(n1073), .C(n1069), .Q(n1071) );
  OAI210 U209 ( .A(n141), .B(n1208), .C(compare_i_data_rs[4]), .Q(n1207) );
  AOI210 U210 ( .A(n1073), .B(u_alu_pre_sum_3b[1]), .C(n1013), .Q(n1017) );
  AOI210 U211 ( .A(n1073), .B(u_alu_pre_sum_3b[2]), .C(n1018), .Q(n1022) );
  AOI210 U212 ( .A(n1073), .B(u_alu_pre_sum_3b[3]), .C(n1024), .Q(n1028) );
  NAND24 U213 ( .A(u_alu_pre_sum_3b[8]), .B(n1073), .Q(n1076) );
  AOI210 U214 ( .A(n296), .B(i_data_rs[29]), .C(n592), .Q(n593) );
  NOR24 U215 ( .A(n999), .B(u_alu_sub_x_2_n2), .Q(n1158) );
  ADD31 U216 ( .A(n172), .B(compare_i_data_rs[5]), .CI(u_alu_sub_x_2_n13), 
        .CO(u_alu_sub_x_2_n12), .S(u_alu_half_sub_5_) );
  NAND23 U217 ( .A(n297), .B(i_data_rs[0]), .Q(n725) );
  NAND28 U218 ( .A(n707), .B(n706), .Q(compare_i_data_rs[3]) );
  NAND28 U219 ( .A(n581), .B(i_con_Efamux[1]), .Q(n711) );
  NOR33 U220 ( .A(n584), .B(i_con_Efamux[1]), .C(i_con_Efamux[2]), .Q(n721) );
  INV3 U221 ( .A(n711), .Q(n573) );
  INV3 U222 ( .A(n1174), .Q(n304) );
  INV3 U223 ( .A(n720), .Q(n295) );
  BUF6 U224 ( .A(alu_i_data_B[1]), .Q(u_alu_lt_x_11_B_1_) );
  NOR21 U225 ( .A(n1240), .B(n141), .Q(n904) );
  MUX22 U226 ( .A(n533), .B(n532), .S(n437), .Q(u_alu_N228) );
  MUX22 U227 ( .A(n360), .B(n422), .S(n437), .Q(u_alu_N215) );
  MUX22 U228 ( .A(n522), .B(n521), .S(n437), .Q(u_alu_N227) );
  MUX22 U229 ( .A(n350), .B(n420), .S(n437), .Q(u_alu_N213) );
  MUX22 U230 ( .A(n355), .B(n421), .S(n437), .Q(u_alu_N214) );
  INV3 U231 ( .A(alu_i_data_B[26]), .Q(n132) );
  INV3 U232 ( .A(alu_i_data_B[29]), .Q(n129) );
  NAND20 U233 ( .A(alu_i_data_B[14]), .B(n164), .Q(n209) );
  NAND20 U234 ( .A(n157), .B(alu_i_data_B[28]), .Q(n175) );
  INV3 U235 ( .A(alu_i_data_B[27]), .Q(n128) );
  INV3 U236 ( .A(alu_i_data_B[24]), .Q(n131) );
  INV3 U237 ( .A(alu_i_data_B[30]), .Q(n130) );
  INV3 U238 ( .A(alu_i_data_B[21]), .Q(n127) );
  INV3 U239 ( .A(alu_i_data_B[11]), .Q(n134) );
  INV3 U240 ( .A(alu_i_data_B[12]), .Q(n137) );
  INV3 U241 ( .A(alu_i_data_B[8]), .Q(n136) );
  INV3 U242 ( .A(alu_i_data_B[15]), .Q(n135) );
  NAND22 U243 ( .A(compare_i_data_rt[21]), .B(n806), .Q(n787) );
  OAI211 U244 ( .A(n842), .B(n1283), .C(n746), .Q(compare_i_data_rt[29]) );
  AOI211 U245 ( .A(n139), .B(i_data_rt[14]), .C(n815), .Q(n816) );
  AOI211 U246 ( .A(n139), .B(i_data_rt[15]), .C(n811), .Q(n812) );
  AOI211 U247 ( .A(n139), .B(i_data_rt[30]), .C(n740), .Q(n741) );
  NAND22 U248 ( .A(n139), .B(i_data_rt[17]), .Q(n801) );
  OAI210 U249 ( .A(n299), .B(n734), .C(n733), .Q(n735) );
  BUF12 U250 ( .A(n861), .Q(n139) );
  OAI211 U251 ( .A(n711), .B(n810), .C(n649), .Q(n650) );
  NOR21 U252 ( .A(i_con_Ealuop[2]), .B(n1251), .Q(n1252) );
  INV1 U253 ( .A(i_data_immext[6]), .Q(n572) );
  INV3 U254 ( .A(i_data_FEalures[22]), .Q(n779) );
  INV2 U255 ( .A(i_data_FEalures[19]), .Q(n625) );
  NOR22 U256 ( .A(i_con_Efbmux[2]), .B(i_con_Efbmux[0]), .Q(n729) );
  INV3 U257 ( .A(i_data_FEalures[21]), .Q(n784) );
  INV3 U258 ( .A(i_data_FEalures[23]), .Q(n774) );
  INV2 U259 ( .A(i_data_FEalures[3]), .Q(n701) );
  INV2 U260 ( .A(i_data_FEalures[20]), .Q(n618) );
  INV2 U261 ( .A(i_data_FEalures[1]), .Q(n712) );
  INV2 U262 ( .A(i_con_Efamux[2]), .Q(n583) );
  NAND31 U263 ( .A(n1134), .B(n1133), .C(n1132), .Q(alu_o_data_AluRes[27]) );
  NAND41 U264 ( .A(n1116), .B(n1115), .C(n1114), .D(n1113), .Q(n1117) );
  AOI211 U265 ( .A(u_alu_lt_x_11_B_7_), .B(n141), .C(n1194), .Q(n1191) );
  OAI211 U266 ( .A(n141), .B(n1198), .C(compare_i_data_rs[6]), .Q(n1197) );
  OAI211 U267 ( .A(n141), .B(n1219), .C(compare_i_data_rs[2]), .Q(n1218) );
  AOI211 U268 ( .A(alu_i_data_B[4]), .B(n141), .C(n1209), .Q(n1206) );
  OAI211 U269 ( .A(n141), .B(n1213), .C(compare_i_data_rs[3]), .Q(n1212) );
  AOI211 U270 ( .A(alu_i_data_B[3]), .B(n141), .C(n1214), .Q(n1211) );
  AOI211 U271 ( .A(u_alu_lt_x_11_B_1_), .B(n141), .C(n1233), .Q(n1230) );
  AOI211 U272 ( .A(n294), .B(n141), .C(n1204), .Q(n1201) );
  AOI211 U273 ( .A(alu_i_data_B[2]), .B(n141), .C(n1220), .Q(n1217) );
  OAI211 U274 ( .A(n141), .B(n1232), .C(compare_i_data_rs[1]), .Q(n1231) );
  OAI211 U275 ( .A(n141), .B(n1193), .C(compare_i_data_rs[7]), .Q(n1192) );
  OAI211 U276 ( .A(n141), .B(n1203), .C(compare_i_data_rs[5]), .Q(n1202) );
  NAND21 U277 ( .A(i_con_bop[1]), .B(n1303), .Q(n1304) );
  NAND20 U278 ( .A(u_alu_N250), .B(n1180), .Q(n1100) );
  NAND20 U279 ( .A(u_alu_N252), .B(n1180), .Q(n1128) );
  NAND21 U280 ( .A(u_alu_N197), .B(n575), .Q(n894) );
  NAND21 U281 ( .A(u_alu_N195), .B(n575), .Q(n900) );
  INV3 U282 ( .A(n1179), .Q(n303) );
  INV2 U283 ( .A(n999), .Q(n906) );
  INV3 U284 ( .A(n384), .Q(n436) );
  IMUX21 U285 ( .A(n443), .B(n556), .S(u_alu_ashr_4_SH_3_), .Q(n444) );
  IMUX21 U286 ( .A(n276), .B(u_alu_pre_subb[0]), .S(u_alu_pre_suba[1]), .Q(
        u_alu_pre_subb[1]) );
  AOI211 U287 ( .A(u_alu_add_x_1_n21), .B(u_alu_add_x_1_n12), .C(
        u_alu_add_x_1_n13), .Q(u_alu_add_x_1_n11) );
  INV3 U288 ( .A(alu_i_data_B[18]), .Q(n144) );
  NOR20 U289 ( .A(alu_i_data_B[13]), .B(n154), .Q(n190) );
  INV3 U290 ( .A(u_alu_lt_x_11_B_7_), .Q(n147) );
  NOR20 U291 ( .A(alu_i_data_B[31]), .B(n158), .Q(n174) );
  INV6 U292 ( .A(alu_i_data_B[17]), .Q(n126) );
  NOR20 U293 ( .A(alu_i_data_B[25]), .B(n166), .Q(n241) );
  NOR20 U294 ( .A(alu_i_data_B[24]), .B(n161), .Q(n242) );
  INV0 U295 ( .A(u_alu_add_x_1_n28), .Q(u_alu_add_x_1_n26) );
  IMUX21 U296 ( .A(u_alu_lt_x_11_B_1_), .B(alu_i_data_B[0]), .S(
        i_data_immext[6]), .Q(n317) );
  INV3 U297 ( .A(alu_i_data_B[0]), .Q(n1235) );
  XNR21 U298 ( .A(compare_i_data_rt[29]), .B(compare_i_data_rs[29]), .Q(n948)
         );
  INV2 U299 ( .A(compare_i_data_rs[25]), .Q(n166) );
  INV3 U300 ( .A(compare_i_data_rs[31]), .Q(n158) );
  IMUX21 U301 ( .A(alu_i_data_B[3]), .B(alu_i_data_B[2]), .S(i_data_immext[6]), 
        .Q(n315) );
  INV3 U302 ( .A(compare_i_data_rs[21]), .Q(n1043) );
  INV3 U303 ( .A(compare_i_data_rs[9]), .Q(n167) );
  INV3 U304 ( .A(compare_i_data_rs[8]), .Q(n151) );
  INV3 U305 ( .A(compare_i_data_rs[2]), .Q(n936) );
  INV3 U306 ( .A(compare_i_data_rs[11]), .Q(n155) );
  INV3 U307 ( .A(compare_i_data_rs[14]), .Q(n164) );
  INV2 U308 ( .A(compare_i_data_rs[15]), .Q(n925) );
  INV3 U309 ( .A(compare_i_data_rs[13]), .Q(n154) );
  NAND23 U310 ( .A(n679), .B(n678), .Q(compare_i_data_rs[7]) );
  NAND22 U311 ( .A(n700), .B(n699), .Q(compare_i_data_rs[4]) );
  NAND22 U312 ( .A(compare_i_data_rt[26]), .B(n806), .Q(n762) );
  NAND22 U313 ( .A(compare_i_data_rt[25]), .B(n806), .Q(n767) );
  NAND22 U314 ( .A(compare_i_data_rt[24]), .B(n806), .Q(n772) );
  NAND22 U315 ( .A(compare_i_data_rt[16]), .B(n806), .Q(n808) );
  NAND31 U316 ( .A(n805), .B(n804), .C(n803), .Q(compare_i_data_rt[16]) );
  AOI2111 U317 ( .A(i_data_FMalures[7]), .B(n721), .C(n677), .D(n676), .Q(n678) );
  OAI211 U318 ( .A(n842), .B(n1282), .C(n751), .Q(compare_i_data_rt[28]) );
  AOI2111 U319 ( .A(i_data_FMalures[1]), .B(n721), .C(n717), .D(n716), .Q(n718) );
  NAND22 U320 ( .A(n168), .B(i_data_rt[16]), .Q(n805) );
  OAI211 U321 ( .A(n711), .B(n834), .C(n667), .Q(n668) );
  OAI211 U322 ( .A(n711), .B(n838), .C(n670), .Q(n671) );
  AOI221 U323 ( .A(n169), .B(i_data_FMmemout[2]), .C(n574), .D(
        i_data_FWmemout[2]), .Q(n708) );
  OAI211 U324 ( .A(n711), .B(n754), .C(n597), .Q(n598) );
  OAI211 U325 ( .A(n711), .B(n779), .C(n612), .Q(n613) );
  OAI211 U326 ( .A(n711), .B(n784), .C(n615), .Q(n616) );
  OAI211 U327 ( .A(n711), .B(n759), .C(n600), .Q(n601) );
  OAI211 U328 ( .A(n711), .B(n774), .C(n609), .Q(n610) );
  OAI211 U329 ( .A(n711), .B(n749), .C(n594), .Q(n595) );
  OAI211 U330 ( .A(n711), .B(n764), .C(n603), .Q(n604) );
  OAI212 U331 ( .A(n734), .B(n711), .C(n585), .Q(n586) );
  OAI211 U332 ( .A(n711), .B(n769), .C(n606), .Q(n607) );
  OAI211 U333 ( .A(n711), .B(n814), .C(n652), .Q(n653) );
  OAI211 U334 ( .A(n711), .B(n818), .C(n655), .Q(n656) );
  OAI211 U335 ( .A(n711), .B(n830), .C(n664), .Q(n665) );
  AOI221 U336 ( .A(n169), .B(i_data_FMmemout[0]), .C(n574), .D(
        i_data_FWmemout[0]), .Q(n723) );
  OAI211 U337 ( .A(n711), .B(n822), .C(n658), .Q(n659) );
  OAI211 U338 ( .A(n711), .B(n826), .C(n661), .Q(n662) );
  NOR21 U339 ( .A(n618), .B(n711), .Q(n622) );
  OAI211 U340 ( .A(n711), .B(n744), .C(n591), .Q(n592) );
  OAI211 U341 ( .A(n711), .B(n739), .C(n588), .Q(n589) );
  NAND22 U342 ( .A(n728), .B(n727), .Q(n842) );
  BUF12 U343 ( .A(n864), .Q(n301) );
  OAI211 U344 ( .A(i_con_Ealuop[5]), .B(n1252), .C(i_con_Ealuop[0]), .Q(n1253)
         );
  AOI221 U345 ( .A(i_con_Ealuop[4]), .B(n1251), .C(i_con_Ealuop[5]), .D(n1248), 
        .Q(n1249) );
  NOR31 U346 ( .A(n583), .B(i_con_Efamux[1]), .C(i_con_Efamux[0]), .Q(n722) );
  BUF8 U347 ( .A(i_con_Ealusrc), .Q(n305) );
  INV2 U348 ( .A(i_data_FWmemout[4]), .Q(n696) );
  INV2 U349 ( .A(i_data_FEalures[4]), .Q(n694) );
  INV1 U350 ( .A(i_con_bop[2]), .Q(n967) );
  INV2 U351 ( .A(i_data_FWmemout[5]), .Q(n689) );
  INV2 U352 ( .A(i_data_FEalures[5]), .Q(n687) );
  INV2 U353 ( .A(i_con_Efamux[0]), .Q(n584) );
  INV2 U354 ( .A(i_data_FWmemout[3]), .Q(n703) );
  INV2 U355 ( .A(i_data_FWmemout[6]), .Q(n682) );
  INV2 U356 ( .A(i_data_FEalures[6]), .Q(n680) );
  NAND42 U357 ( .A(n1017), .B(n1016), .C(n1015), .D(n1014), .Q(
        alu_o_data_AluRes[17]) );
  NAND42 U358 ( .A(n1022), .B(n1021), .C(n1020), .D(n1019), .Q(
        alu_o_data_AluRes[18]) );
  NAND42 U359 ( .A(n1157), .B(n1156), .C(n1155), .D(n1154), .Q(
        alu_o_data_AluRes[30]) );
  NAND42 U360 ( .A(n1028), .B(n1027), .C(n1026), .D(n1025), .Q(
        alu_o_data_AluRes[19]) );
  INV2 U361 ( .A(n1167), .Q(n1090) );
  INV2 U362 ( .A(u_alu_pre_suba[14]), .Q(n291) );
  INV2 U363 ( .A(n1073), .Q(n1009) );
  INV2 U364 ( .A(n274), .Q(n292) );
  NAND21 U365 ( .A(u_alu_pre_sum_3a[7]), .B(n1074), .Q(n1068) );
  NAND21 U366 ( .A(u_alu_pre_sum_3a[5]), .B(n1074), .Q(n1048) );
  NAND21 U367 ( .A(u_alu_pre_sum_3a[6]), .B(n1074), .Q(n1058) );
  IMUX21 U368 ( .A(n283), .B(u_alu_pre_suba[13]), .S(n272), .Q(
        u_alu_pre_subb[13]) );
  INV2 U369 ( .A(u_alu_pre_suba[13]), .Q(n283) );
  IMUX21 U370 ( .A(n282), .B(u_alu_pre_suba[11]), .S(n270), .Q(
        u_alu_pre_subb[11]) );
  IMUX21 U371 ( .A(n281), .B(u_alu_pre_suba[9]), .S(n268), .Q(
        u_alu_pre_subb[9]) );
  OAI211 U372 ( .A(n1185), .B(compare_i_data_rs[8]), .C(n1186), .Q(
        alu_o_data_AluRes[8]) );
  OAI221 U373 ( .A(n1234), .B(n1241), .C(n1242), .D(n1243), .Q(n1238) );
  IMUX21 U374 ( .A(n280), .B(u_alu_pre_suba[7]), .S(n266), .Q(
        u_alu_pre_subb[7]) );
  OAI2111 U375 ( .A(compare_i_data_rs[5]), .B(n1200), .C(n1201), .D(n1202), 
        .Q(alu_o_data_AluRes[5]) );
  AOI311 U376 ( .A(n1302), .B(i_con_bop[2]), .C(i_con_bop[0]), .D(n1305), .Q(
        n969) );
  IMUX21 U377 ( .A(n279), .B(u_alu_pre_suba[5]), .S(n264), .Q(
        u_alu_pre_subb[5]) );
  OAI2111 U378 ( .A(compare_i_data_rs[1]), .B(n1229), .C(n1230), .D(n1231), 
        .Q(alu_o_data_AluRes[1]) );
  OAI2111 U379 ( .A(compare_i_data_rs[3]), .B(n1210), .C(n1211), .D(n1212), 
        .Q(alu_o_data_AluRes[3]) );
  NAND21 U380 ( .A(u_alu_N166), .B(n998), .Q(n973) );
  OAI2111 U381 ( .A(compare_i_data_rs[2]), .B(n1216), .C(n1217), .D(n1218), 
        .Q(alu_o_data_AluRes[2]) );
  INV2 U382 ( .A(u_alu_pre_sum_3a[8]), .Q(n1077) );
  NOR21 U383 ( .A(i_con_bop[2]), .B(n1304), .Q(n1305) );
  NAND21 U384 ( .A(u_alu_half_sub_7_), .B(n906), .Q(n885) );
  INV1 U385 ( .A(u_alu_pre_sum_4a[7]), .Q(n260) );
  OAI211 U386 ( .A(n245), .B(n244), .C(n243), .Q(n246) );
  AOI210 U387 ( .A(n1180), .B(u_alu_N256), .C(n1166), .Q(n1172) );
  NAND21 U388 ( .A(u_alu_half_sub_6_), .B(n906), .Q(n888) );
  AOI220 U389 ( .A(n998), .B(u_alu_sum_1_7_), .C(u_alu_N232), .D(n1180), .Q(
        n884) );
  IMAJ30 U390 ( .A(i_con_bop[2]), .B(i_con_bop[1]), .C(n1303), .Q(n1306) );
  INV2 U391 ( .A(n1303), .Q(n966) );
  AOI220 U392 ( .A(n998), .B(u_alu_sum_1_6_), .C(u_alu_N231), .D(n1180), .Q(
        n887) );
  NAND21 U393 ( .A(u_alu_N201), .B(n575), .Q(n878) );
  NAND21 U394 ( .A(u_alu_N220), .B(n575), .Q(n1129) );
  NAND21 U395 ( .A(u_alu_N199), .B(n575), .Q(n886) );
  NAND21 U396 ( .A(u_alu_N200), .B(n575), .Q(n883) );
  AOI220 U397 ( .A(n998), .B(u_alu_sum_1_5_), .C(u_alu_N230), .D(n1180), .Q(
        n890) );
  NAND21 U398 ( .A(u_alu_N219), .B(n575), .Q(n1114) );
  NAND21 U399 ( .A(u_alu_half_sub_5_), .B(n906), .Q(n891) );
  NAND31 U400 ( .A(n1301), .B(n1300), .C(n1299), .Q(n1303) );
  NAND21 U401 ( .A(u_alu_N233), .B(n1180), .Q(n877) );
  NAND21 U402 ( .A(u_alu_N198), .B(n575), .Q(n889) );
  NAND20 U403 ( .A(u_alu_N217), .B(n575), .Q(n1085) );
  NAND21 U404 ( .A(u_alu_N218), .B(n575), .Q(n1101) );
  NAND21 U405 ( .A(u_alu_N222), .B(n575), .Q(n1147) );
  NAND21 U406 ( .A(u_alu_N224), .B(n575), .Q(n1170) );
  NAND21 U407 ( .A(u_alu_N213), .B(n575), .Q(n1036) );
  NAND21 U408 ( .A(u_alu_N194), .B(n575), .Q(n903) );
  NAND21 U409 ( .A(u_alu_N196), .B(n575), .Q(n897) );
  AOI220 U410 ( .A(n998), .B(u_alu_sum_1_3_), .C(u_alu_half_sub_3_), .D(n906), 
        .Q(n896) );
  MUX22 U411 ( .A(n444), .B(n481), .S(i_data_immext[10]), .Q(u_alu_N225) );
  INV3 U412 ( .A(n964), .Q(n1299) );
  INV2 U413 ( .A(n481), .Q(n566) );
  MUX22 U414 ( .A(n562), .B(n561), .S(i_data_immext[10]), .Q(u_alu_N234) );
  NAND21 U415 ( .A(u_alu_half_sub_4_), .B(n906), .Q(n893) );
  AOI220 U416 ( .A(n998), .B(u_alu_sum_1_2_), .C(n906), .D(u_alu_half_sub_2_), 
        .Q(n899) );
  MUX22 U417 ( .A(n496), .B(n495), .S(n437), .Q(u_alu_N226) );
  NOR21 U418 ( .A(i_data_immext[10]), .B(n436), .Q(u_alu_N203) );
  AOI220 U419 ( .A(n906), .B(u_alu_half_sub_1_), .C(n998), .D(u_alu_sum_1_1_), 
        .Q(n902) );
  INV2 U420 ( .A(n557), .Q(n565) );
  INV2 U421 ( .A(n345), .Q(n427) );
  INV1 U422 ( .A(u_alu_pre_suba[2]), .Q(n277) );
  INV2 U423 ( .A(n543), .Q(n568) );
  INV2 U424 ( .A(n511), .Q(n570) );
  INV2 U425 ( .A(n561), .Q(n567) );
  INV2 U426 ( .A(n420), .Q(n430) );
  IMUX21 U427 ( .A(n560), .B(n559), .S(u_alu_ashr_4_SH_3_), .Q(n562) );
  INV2 U428 ( .A(n422), .Q(n432) );
  INV2 U429 ( .A(n419), .Q(n429) );
  INV2 U430 ( .A(n423), .Q(n433) );
  INV2 U431 ( .A(n421), .Q(n431) );
  INV2 U432 ( .A(n406), .Q(n428) );
  NAND31 U433 ( .A(n963), .B(n962), .C(n961), .Q(n964) );
  NOR20 U434 ( .A(i_data_immext[8]), .B(n564), .Q(n498) );
  NOR20 U435 ( .A(i_data_immext[8]), .B(n563), .Q(n503) );
  OAI211 U436 ( .A(n215), .B(n214), .C(n223), .Q(n216) );
  NOR40 U437 ( .A(n960), .B(n959), .C(n958), .D(n957), .Q(n961) );
  NOR20 U438 ( .A(i_data_immext[8]), .B(n569), .Q(n506) );
  INV1 U439 ( .A(n232), .Q(n257) );
  INV1 U440 ( .A(u_alu_add_x_1_n30), .Q(u_alu_add_x_1_n29) );
  IMUX20 U441 ( .A(n471), .B(n474), .S(i_data_immext[8]), .Q(n487) );
  MUX21 U442 ( .A(n479), .B(n478), .S(i_data_immext[8]), .Q(n507) );
  IMUX21 U443 ( .A(n539), .B(n493), .S(i_data_immext[8]), .Q(n560) );
  INV1 U444 ( .A(n505), .Q(n569) );
  INV1 U445 ( .A(n230), .Q(n254) );
  INV2 U446 ( .A(u_alu_add_x_1_n8), .Q(u_alu_sum_1_0_) );
  INV1 U447 ( .A(u_alu_add_x_1_n39), .Q(u_alu_add_x_1_n38) );
  IMUX21 U448 ( .A(n535), .B(n458), .S(i_data_immext[8]), .Q(n556) );
  NAND21 U449 ( .A(alu_i_con_AluCtrl[3]), .B(n1245), .Q(n1234) );
  INV2 U450 ( .A(n239), .Q(n259) );
  IMUX20 U451 ( .A(n476), .B(n479), .S(i_data_immext[8]), .Q(n489) );
  INV2 U452 ( .A(n178), .Q(n258) );
  INV1 U453 ( .A(n502), .Q(n563) );
  MUX21 U454 ( .A(n460), .B(n459), .S(i_data_immext[8]), .Q(n499) );
  INV1 U455 ( .A(n497), .Q(n564) );
  MUX21 U456 ( .A(n474), .B(n473), .S(i_data_immext[8]), .Q(n504) );
  IMUX21 U457 ( .A(n470), .B(n469), .S(n440), .Q(n484) );
  XOR21 U458 ( .A(compare_i_data_rs[29]), .B(n129), .Q(n286) );
  IMUX20 U459 ( .A(n527), .B(n492), .S(u_alu_ashr_4_SH_1_), .Q(n539) );
  INV2 U460 ( .A(u_alu_pre_subb[0]), .Q(n276) );
  IMUX20 U461 ( .A(n399), .B(n386), .S(u_alu_ashr_4_SH_1_), .Q(n413) );
  NOR40 U462 ( .A(n944), .B(n943), .C(n942), .D(n941), .Q(n962) );
  IMUX20 U463 ( .A(n392), .B(n380), .S(u_alu_ashr_4_SH_1_), .Q(n408) );
  NOR40 U464 ( .A(n929), .B(n928), .C(n927), .D(n926), .Q(n1301) );
  IMUX21 U465 ( .A(n309), .B(n311), .S(n440), .Q(n320) );
  IMUX20 U466 ( .A(n380), .B(n366), .S(u_alu_ashr_4_SH_1_), .Q(n393) );
  INV2 U467 ( .A(n228), .Q(n255) );
  IMUX21 U468 ( .A(n315), .B(n317), .S(n440), .Q(n324) );
  IMUX20 U469 ( .A(n525), .B(n528), .S(u_alu_ashr_4_SH_1_), .Q(n540) );
  INV2 U470 ( .A(n330), .Q(n426) );
  INV1 U471 ( .A(n237), .Q(n256) );
  IMUX20 U472 ( .A(n528), .B(n527), .S(u_alu_ashr_4_SH_1_), .Q(n552) );
  IMUX20 U473 ( .A(n386), .B(n373), .S(u_alu_ashr_4_SH_1_), .Q(n400) );
  NOR40 U474 ( .A(n940), .B(n939), .C(n938), .D(n937), .Q(n963) );
  INV2 U475 ( .A(alu_i_data_B[31]), .Q(n1159) );
  NAND21 U476 ( .A(alu_i_con_AluCtrl[3]), .B(alu_i_con_AluCtrl[0]), .Q(n880)
         );
  IMUX20 U477 ( .A(n492), .B(n462), .S(u_alu_ashr_4_SH_1_), .Q(n551) );
  IMUX20 U478 ( .A(n332), .B(n322), .S(u_alu_ashr_4_SH_1_), .Q(n342) );
  IMUX21 U479 ( .A(alu_i_data_B[2]), .B(u_alu_lt_x_11_B_1_), .S(
        i_data_immext[6]), .Q(n309) );
  INV3 U480 ( .A(alu_i_data_B[25]), .Q(n142) );
  INV3 U481 ( .A(alu_i_data_B[28]), .Q(n143) );
  INV2 U482 ( .A(compare_i_data_rs[12]), .Q(n930) );
  INV3 U483 ( .A(alu_i_data_B[20]), .Q(n145) );
  INV3 U484 ( .A(alu_i_data_B[22]), .Q(n146) );
  INV2 U485 ( .A(compare_i_data_rs[27]), .Q(n1122) );
  INV3 U486 ( .A(alu_i_data_B[23]), .Q(n148) );
  INV2 U487 ( .A(compare_i_data_rs[26]), .Q(n1108) );
  INV1 U488 ( .A(alu_i_con_AluCtrl[3]), .Q(n882) );
  NAND22 U489 ( .A(alu_i_data_B[0]), .B(n572), .Q(n311) );
  INV3 U490 ( .A(compare_i_data_rs[10]), .Q(n149) );
  INV3 U491 ( .A(alu_i_data_B[4]), .Q(n150) );
  NAND21 U492 ( .A(compare_i_data_rt[20]), .B(n806), .Q(n791) );
  INV1 U493 ( .A(n1263), .Q(n1256) );
  OAI2112 U494 ( .A(n1254), .B(n1261), .C(n1266), .D(n1253), .Q(
        alu_i_con_AluCtrl[0]) );
  INV3 U495 ( .A(alu_i_data_B[3]), .Q(n153) );
  NAND21 U496 ( .A(compare_i_data_rt[30]), .B(n806), .Q(n742) );
  NAND21 U497 ( .A(compare_i_data_rt[28]), .B(n806), .Q(n752) );
  NAND21 U498 ( .A(compare_i_data_rt[31]), .B(n806), .Q(n737) );
  INV3 U499 ( .A(alu_i_data_B[14]), .Q(n156) );
  INV3 U500 ( .A(compare_i_data_rs[28]), .Q(n157) );
  NAND21 U501 ( .A(compare_i_data_rt[29]), .B(n806), .Q(n747) );
  INV3 U502 ( .A(compare_i_data_rs[23]), .Q(n159) );
  INV3 U503 ( .A(alu_i_data_B[9]), .Q(n160) );
  INV2 U504 ( .A(compare_i_data_rs[24]), .Q(n161) );
  INV3 U505 ( .A(alu_i_data_B[13]), .Q(n162) );
  INV3 U506 ( .A(compare_i_data_rs[22]), .Q(n163) );
  INV1 U507 ( .A(compare_i_data_rs[20]), .Q(n165) );
  MUX26 U508 ( .A(compare_i_data_rt[5]), .B(i_data_immext[5]), .S(n305), .Q(
        n294) );
  OAI211 U509 ( .A(n298), .B(n1285), .C(n736), .Q(compare_i_data_rt[31]) );
  NAND31 U510 ( .A(n854), .B(n853), .C(n852), .Q(compare_i_data_rt[4]) );
  NAND31 U511 ( .A(n857), .B(n856), .C(n855), .Q(compare_i_data_rt[3]) );
  OAI211 U512 ( .A(n924), .B(n923), .C(n1264), .Q(n1265) );
  NAND33 U513 ( .A(n860), .B(n859), .C(n858), .Q(compare_i_data_rt[1]) );
  OAI211 U514 ( .A(n922), .B(n921), .C(n1264), .Q(n1262) );
  OAI211 U515 ( .A(n140), .B(n627), .C(n626), .Q(n628) );
  INV2 U516 ( .A(n1177), .Q(n1255) );
  AOI211 U517 ( .A(n917), .B(n909), .C(n919), .Q(n871) );
  OAI211 U518 ( .A(n620), .B(n140), .C(n619), .Q(n621) );
  INV3 U519 ( .A(n295), .Q(n296) );
  OAI211 U520 ( .A(n140), .B(n634), .C(n633), .Q(n635) );
  NAND22 U521 ( .A(n920), .B(n913), .Q(n919) );
  INV2 U522 ( .A(n920), .Q(n922) );
  OAI211 U523 ( .A(n299), .B(n826), .C(n825), .Q(n827) );
  OAI211 U524 ( .A(n299), .B(n838), .C(n837), .Q(n840) );
  OAI211 U525 ( .A(n299), .B(n834), .C(n833), .Q(n835) );
  OAI211 U526 ( .A(n299), .B(n779), .C(n778), .Q(n780) );
  OAI211 U527 ( .A(n299), .B(n784), .C(n783), .Q(n785) );
  OAI211 U528 ( .A(n299), .B(n774), .C(n773), .Q(n775) );
  OAI211 U529 ( .A(n299), .B(n749), .C(n748), .Q(n750) );
  OAI211 U530 ( .A(n299), .B(n769), .C(n768), .Q(n770) );
  OAI211 U531 ( .A(n299), .B(n764), .C(n763), .Q(n765) );
  OAI211 U532 ( .A(n299), .B(n759), .C(n758), .Q(n760) );
  OAI211 U533 ( .A(n299), .B(n754), .C(n753), .Q(n755) );
  OAI211 U534 ( .A(n299), .B(n744), .C(n743), .Q(n745) );
  OAI211 U535 ( .A(n299), .B(n739), .C(n738), .Q(n740) );
  OAI211 U536 ( .A(n299), .B(n818), .C(n817), .Q(n819) );
  OAI211 U537 ( .A(n299), .B(n810), .C(n809), .Q(n811) );
  OAI211 U538 ( .A(n299), .B(n830), .C(n829), .Q(n831) );
  OAI211 U539 ( .A(n299), .B(n814), .C(n813), .Q(n815) );
  OAI211 U540 ( .A(n299), .B(n822), .C(n821), .Q(n823) );
  AOI2111 U541 ( .A(n1247), .B(i_data_immext[2]), .C(n917), .D(n916), .Q(n918)
         );
  AOI311 U542 ( .A(i_con_Ealuop[3]), .B(i_con_Ealuop[2]), .C(n1250), .D(n1259), 
        .Q(n1266) );
  NAND22 U543 ( .A(n914), .B(i_data_immext[0]), .Q(n920) );
  INV6 U544 ( .A(n714), .Q(n574) );
  INV6 U545 ( .A(n842), .Q(n863) );
  BUF12 U546 ( .A(n862), .Q(n302) );
  AOI211 U547 ( .A(i_con_Ealuop[1]), .B(n1249), .C(n1267), .Q(n1259) );
  INV3 U548 ( .A(n868), .Q(n917) );
  NOR21 U549 ( .A(i_con_Ealuop[4]), .B(n1267), .Q(n1250) );
  INV2 U550 ( .A(u_alu_ashr_4_SH_3_), .Q(n571) );
  NOR21 U551 ( .A(n1257), .B(i_con_Ealuop[0]), .Q(n1264) );
  INV3 U552 ( .A(i_data_FWmemout[14]), .Q(n1273) );
  INV3 U553 ( .A(i_data_FWmemout[15]), .Q(n1274) );
  INV2 U554 ( .A(i_con_Ealuop[3]), .Q(n1251) );
  INV3 U555 ( .A(i_data_FEalures[14]), .Q(n814) );
  INV2 U556 ( .A(i_con_Ealuop[4]), .Q(n1268) );
  INV1 U557 ( .A(i_data_FEalures[17]), .Q(n639) );
  INV3 U558 ( .A(i_data_FEalures[11]), .Q(n826) );
  INV2 U559 ( .A(i_data_FEalures[24]), .Q(n769) );
  INV2 U560 ( .A(i_data_FWmemout[17]), .Q(n641) );
  INV3 U561 ( .A(i_data_FWmemout[22]), .Q(n1276) );
  INV3 U562 ( .A(i_data_FWmemout[11]), .Q(n1270) );
  INV2 U563 ( .A(i_data_FWmemout[7]), .Q(n675) );
  INV3 U564 ( .A(i_con_Malupc8), .Q(n1293) );
  INV3 U565 ( .A(i_data_FEalures[9]), .Q(n834) );
  INV3 U566 ( .A(i_data_FWmemout[13]), .Q(n1272) );
  INV3 U567 ( .A(i_data_FWmemout[26]), .Q(n1280) );
  INV3 U568 ( .A(i_data_FWmemout[12]), .Q(n1271) );
  INV3 U569 ( .A(i_data_FEalures[13]), .Q(n818) );
  INV2 U570 ( .A(i_data_FEalures[26]), .Q(n759) );
  INV2 U571 ( .A(i_data_FWmemout[20]), .Q(n620) );
  INV2 U572 ( .A(i_data_FEalures[25]), .Q(n764) );
  INV3 U573 ( .A(i_data_FEalures[12]), .Q(n822) );
  INV3 U574 ( .A(i_data_FWmemout[21]), .Q(n1275) );
  INV3 U575 ( .A(i_data_FWmemout[27]), .Q(n1281) );
  INV3 U576 ( .A(i_data_FWmemout[23]), .Q(n1277) );
  INV3 U577 ( .A(i_con_Efamux[1]), .Q(n580) );
  INV3 U578 ( .A(i_data_FWmemout[25]), .Q(n1279) );
  INV2 U579 ( .A(i_data_FEalures[27]), .Q(n754) );
  INV3 U580 ( .A(i_data_FEalures[10]), .Q(n830) );
  INV2 U581 ( .A(i_data_FWmemout[1]), .Q(n715) );
  INV3 U582 ( .A(i_data_FWmemout[29]), .Q(n1283) );
  INV2 U583 ( .A(i_data_FWmemout[18]), .Q(n634) );
  INV3 U584 ( .A(i_con_Ealuop[1]), .Q(n1257) );
  INV3 U585 ( .A(i_data_FWmemout[10]), .Q(n1269) );
  INV3 U586 ( .A(i_data_FWmemout[31]), .Q(n1285) );
  INV1 U587 ( .A(i_data_FEalures[18]), .Q(n632) );
  INV2 U588 ( .A(i_data_FEalures[28]), .Q(n749) );
  INV3 U589 ( .A(i_data_FWmemout[8]), .Q(n1286) );
  INV3 U590 ( .A(i_data_FEalures[31]), .Q(n734) );
  NAND21 U591 ( .A(i_data_immext[1]), .B(i_data_immext[3]), .Q(n869) );
  INV2 U592 ( .A(i_con_bop[1]), .Q(n1302) );
  INV2 U593 ( .A(i_data_FEalures[30]), .Q(n739) );
  INV3 U594 ( .A(i_data_FEalures[8]), .Q(n838) );
  INV2 U595 ( .A(i_data_FWmemout[19]), .Q(n627) );
  INV3 U596 ( .A(i_data_FWmemout[30]), .Q(n1284) );
  INV1 U597 ( .A(i_data_immext[0]), .Q(n916) );
  INV1 U598 ( .A(i_con_Ealuop[2]), .Q(n1248) );
  INV3 U599 ( .A(i_data_FWmemout[24]), .Q(n1278) );
  INV3 U600 ( .A(i_data_FEalures[15]), .Q(n810) );
  INV2 U601 ( .A(i_data_FEalures[29]), .Q(n744) );
  INV3 U602 ( .A(i_data_FWmemout[9]), .Q(n1287) );
  INV2 U603 ( .A(i_data_FEalures[7]), .Q(n673) );
  INV3 U604 ( .A(i_con_Ealuop[0]), .Q(n1267) );
  INV3 U605 ( .A(i_data_FWmemout[28]), .Q(n1282) );
  BUF6 U606 ( .A(i_data_immext[10]), .Q(n437) );
  XOR22 U607 ( .A(DP_OP_77_130_260_n1), .B(DP_OP_77_130_260_n37), .Q(
        u_alu_N173) );
  AOI222 U608 ( .A(compare_i_data_rs[8]), .B(DP_OP_77_130_260_I3), .C(n170), 
        .D(n151), .Q(DP_OP_77_130_260_n17) );
  BUF6 U609 ( .A(u_alu_sum_1_8_), .Q(n170) );
  ADD32 U610 ( .A(DP_OP_77_130_260_n35), .B(alu_i_data_B[14]), .CI(
        DP_OP_77_130_260_n3), .CO(DP_OP_77_130_260_n2), .S(u_alu_N171) );
  ADD32 U611 ( .A(DP_OP_77_130_260_n36), .B(alu_i_data_B[15]), .CI(
        DP_OP_77_130_260_n2), .CO(DP_OP_77_130_260_n1), .S(u_alu_N172) );
  ADD32 U612 ( .A(DP_OP_77_130_260_n33), .B(alu_i_data_B[12]), .CI(
        DP_OP_77_130_260_n5), .CO(DP_OP_77_130_260_n4), .S(u_alu_N169) );
  ADD32 U613 ( .A(DP_OP_77_130_260_n34), .B(alu_i_data_B[13]), .CI(
        DP_OP_77_130_260_n4), .CO(DP_OP_77_130_260_n3), .S(u_alu_N170) );
  ADD32 U614 ( .A(DP_OP_77_130_260_n31), .B(u_alu_lt_x_11_B_10_), .CI(
        DP_OP_77_130_260_n7), .CO(DP_OP_77_130_260_n6), .S(u_alu_N167) );
  ADD32 U615 ( .A(DP_OP_77_130_260_n32), .B(alu_i_data_B[11]), .CI(
        DP_OP_77_130_260_n6), .CO(DP_OP_77_130_260_n5), .S(u_alu_N168) );
  ADD22 U616 ( .A(DP_OP_77_130_260_n29), .B(alu_i_data_B[8]), .CO(
        DP_OP_77_130_260_n8), .S(u_alu_N165) );
  ADD32 U617 ( .A(DP_OP_77_130_260_n30), .B(alu_i_data_B[9]), .CI(
        DP_OP_77_130_260_n8), .CO(DP_OP_77_130_260_n7), .S(u_alu_N166) );
  IMUX20 U618 ( .A(n152), .B(compare_i_data_rs[0]), .S(alu_i_data_B[0]), .Q(
        u_alu_half_sub_0_) );
  INV3 U619 ( .A(alu_i_data_B[6]), .Q(n173) );
  INV3 U620 ( .A(n294), .Q(n172) );
  NAND22 U621 ( .A(alu_i_data_B[0]), .B(n152), .Q(u_alu_sub_x_2_n17) );
  INV3 U622 ( .A(alu_i_data_B[1]), .Q(n171) );
  ADD32 U623 ( .A(n293), .B(compare_i_data_rs[10]), .CI(u_alu_sub_x_2_n8), 
        .CO(u_alu_sub_x_2_n7), .S(u_alu_half_sub_10_) );
  ADD32 U624 ( .A(n134), .B(compare_i_data_rs[11]), .CI(u_alu_sub_x_2_n7), 
        .CO(u_alu_sub_x_2_n6), .S(u_alu_half_sub_11_) );
  ADD32 U625 ( .A(n137), .B(compare_i_data_rs[12]), .CI(u_alu_sub_x_2_n6), 
        .CO(u_alu_sub_x_2_n5), .S(u_alu_half_sub_12_) );
  ADD32 U626 ( .A(n160), .B(compare_i_data_rs[9]), .CI(u_alu_sub_x_2_n9), .CO(
        u_alu_sub_x_2_n8), .S(u_alu_half_sub_9_) );
  ADD32 U627 ( .A(n162), .B(compare_i_data_rs[13]), .CI(u_alu_sub_x_2_n5), 
        .CO(u_alu_sub_x_2_n4), .S(u_alu_half_sub_13_) );
  ADD32 U628 ( .A(n156), .B(compare_i_data_rs[14]), .CI(u_alu_sub_x_2_n4), 
        .CO(u_alu_sub_x_2_n3), .S(u_alu_half_sub_14_) );
  ADD32 U629 ( .A(n133), .B(compare_i_data_rs[2]), .CI(u_alu_sub_x_2_n16), 
        .CO(u_alu_sub_x_2_n15), .S(u_alu_half_sub_2_) );
  ADD32 U630 ( .A(n153), .B(compare_i_data_rs[3]), .CI(u_alu_sub_x_2_n15), 
        .CO(u_alu_sub_x_2_n14), .S(u_alu_half_sub_3_) );
  ADD32 U631 ( .A(n147), .B(compare_i_data_rs[7]), .CI(u_alu_sub_x_2_n11), 
        .CO(u_alu_sub_x_2_n10), .S(u_alu_half_sub_7_) );
  ADD32 U632 ( .A(n136), .B(compare_i_data_rs[8]), .CI(u_alu_sub_x_2_n10), 
        .CO(u_alu_sub_x_2_n9), .S(u_alu_half_sub_8_) );
  ADD32 U633 ( .A(n135), .B(compare_i_data_rs[15]), .CI(u_alu_sub_x_2_n3), 
        .CO(u_alu_sub_x_2_n2), .S(u_alu_half_sub_15_) );
  ADD32 U634 ( .A(n171), .B(compare_i_data_rs[1]), .CI(u_alu_sub_x_2_n17), 
        .CO(u_alu_sub_x_2_n16), .S(u_alu_half_sub_1_) );
  IMAJ30 U635 ( .A(n129), .B(compare_i_data_rs[29]), .C(n175), .Q(n185) );
  NAND20 U636 ( .A(compare_i_data_rs[29]), .B(n129), .Q(n176) );
  AOI220 U637 ( .A(n128), .B(compare_i_data_rs[27]), .C(n132), .D(
        compare_i_data_rs[26]), .Q(n239) );
  NOR20 U638 ( .A(compare_i_data_rs[24]), .B(n131), .Q(n177) );
  MAJ31 U639 ( .A(alu_i_data_B[25]), .B(n166), .C(n177), .Q(n180) );
  NOR20 U640 ( .A(compare_i_data_rs[26]), .B(n132), .Q(n178) );
  IMAJ30 U641 ( .A(n128), .B(compare_i_data_rs[27]), .C(n258), .Q(n179) );
  NOR20 U642 ( .A(compare_i_data_rs[30]), .B(n130), .Q(n182) );
  MAJ31 U643 ( .A(alu_i_data_B[31]), .B(n158), .C(n182), .Q(n183) );
  NOR20 U644 ( .A(alu_i_data_B[17]), .B(n252), .Q(n226) );
  OAI220 U645 ( .A(n159), .B(alu_i_data_B[23]), .C(n163), .D(alu_i_data_B[22]), 
        .Q(n237) );
  NAND20 U646 ( .A(compare_i_data_rs[21]), .B(n127), .Q(n187) );
  NOR20 U647 ( .A(alu_i_data_B[19]), .B(n253), .Q(n188) );
  AOI210 U648 ( .A(compare_i_data_rs[18]), .B(n144), .C(n188), .Q(n230) );
  OAI210 U649 ( .A(alu_i_data_B[16]), .B(n138), .C(n230), .Q(n225) );
  NAND20 U650 ( .A(compare_i_data_rs[15]), .B(n135), .Q(n189) );
  AOI2110 U651 ( .A(compare_i_data_rs[12]), .B(n137), .C(n190), .D(n218), .Q(
        n223) );
  NOR20 U652 ( .A(alu_i_data_B[9]), .B(n167), .Q(n191) );
  OAI220 U653 ( .A(alu_i_data_B[11]), .B(n155), .C(u_alu_lt_x_11_B_10_), .D(
        n149), .Q(n212) );
  AOI2110 U654 ( .A(compare_i_data_rs[8]), .B(n136), .C(n191), .D(n212), .Q(
        n222) );
  NAND20 U655 ( .A(compare_i_data_rs[7]), .B(n147), .Q(n192) );
  OAI210 U656 ( .A(alu_i_data_B[6]), .B(n251), .C(n192), .Q(n207) );
  NOR20 U657 ( .A(n294), .B(n250), .Q(n200) );
  NOR20 U658 ( .A(alu_i_data_B[3]), .B(n249), .Q(n193) );
  AOI210 U659 ( .A(compare_i_data_rs[2]), .B(n133), .C(n193), .Q(n198) );
  OAI210 U660 ( .A(u_alu_lt_x_11_B_1_), .B(n248), .C(alu_i_data_B[0]), .Q(n194) );
  OAI220 U661 ( .A(compare_i_data_rs[0]), .B(n194), .C(compare_i_data_rs[1]), 
        .D(n171), .Q(n197) );
  NOR20 U662 ( .A(compare_i_data_rs[2]), .B(n133), .Q(n195) );
  MAJ31 U663 ( .A(alu_i_data_B[3]), .B(n249), .C(n195), .Q(n196) );
  AOI2110 U664 ( .A(compare_i_data_rs[4]), .B(n150), .C(n200), .D(n199), .Q(
        n203) );
  NOR20 U665 ( .A(compare_i_data_rs[4]), .B(n150), .Q(n201) );
  MAJ31 U666 ( .A(n294), .B(n250), .C(n201), .Q(n202) );
  NAND20 U667 ( .A(alu_i_data_B[6]), .B(n251), .Q(n204) );
  MAJ31 U668 ( .A(compare_i_data_rs[7]), .B(n147), .C(n204), .Q(n205) );
  NOR20 U669 ( .A(n137), .B(compare_i_data_rs[12]), .Q(n208) );
  MAJ31 U670 ( .A(compare_i_data_rs[15]), .B(n135), .C(n209), .Q(n217) );
  NAND20 U671 ( .A(n149), .B(u_alu_lt_x_11_B_10_), .Q(n210) );
  IMAJ30 U672 ( .A(n134), .B(compare_i_data_rs[11]), .C(n210), .Q(n215) );
  NOR20 U673 ( .A(n136), .B(compare_i_data_rs[8]), .Q(n211) );
  IMAJ30 U674 ( .A(n167), .B(alu_i_data_B[9]), .C(n211), .Q(n213) );
  NOR40 U675 ( .A(n226), .B(n232), .C(n225), .D(n224), .Q(n245) );
  NAND20 U676 ( .A(alu_i_data_B[20]), .B(n165), .Q(n227) );
  MAJ31 U677 ( .A(compare_i_data_rs[21]), .B(n127), .C(n227), .Q(n238) );
  NOR20 U678 ( .A(compare_i_data_rs[18]), .B(n144), .Q(n229) );
  MAJ31 U679 ( .A(alu_i_data_B[19]), .B(n253), .C(n229), .Q(n234) );
  MAJ31 U680 ( .A(compare_i_data_rs[17]), .B(n126), .C(
        u_alu_DP_OP_85J3_126_1427_n46), .Q(n231) );
  NOR40 U681 ( .A(n242), .B(n241), .C(n240), .D(n259), .Q(n243) );
  INV0 U682 ( .A(compare_i_data_rs[17]), .Q(n252) );
  INV0 U683 ( .A(compare_i_data_rs[19]), .Q(n253) );
  INV0 U684 ( .A(compare_i_data_rs[6]), .Q(n251) );
  INV0 U685 ( .A(compare_i_data_rs[5]), .Q(n250) );
  INV0 U686 ( .A(compare_i_data_rs[3]), .Q(n249) );
  INV0 U687 ( .A(compare_i_data_rs[1]), .Q(n248) );
  AOI211 U688 ( .A(n239), .B(n180), .C(n179), .Q(n181) );
  NOR21 U689 ( .A(n240), .B(n181), .Q(n184) );
  AOI2111 U690 ( .A(n186), .B(n185), .C(n184), .D(n183), .Q(n247) );
  AOI211 U691 ( .A(n198), .B(n197), .C(n196), .Q(n199) );
  NOR21 U692 ( .A(n203), .B(n202), .Q(n206) );
  OAI212 U693 ( .A(n207), .B(n206), .C(n205), .Q(n221) );
  NOR21 U694 ( .A(n213), .B(n212), .Q(n214) );
  OAI2111 U695 ( .A(n219), .B(n218), .C(n217), .D(n216), .Q(n220) );
  AOI311 U696 ( .A(n223), .B(n222), .C(n221), .D(n220), .Q(n224) );
  NOR21 U697 ( .A(n231), .B(n254), .Q(n233) );
  OAI212 U698 ( .A(n234), .B(n233), .C(n257), .Q(n235) );
  OAI2111 U699 ( .A(n238), .B(n237), .C(n236), .D(n235), .Q(n244) );
  NAND22 U700 ( .A(n247), .B(n246), .Q(u_alu_N306) );
  OAI2111 U701 ( .A(alu_i_data_B[28]), .B(n157), .C(n186), .D(n176), .Q(n240)
         );
  AOI210 U702 ( .A(compare_i_data_rs[30]), .B(n130), .C(n174), .Q(n186) );
  OAI2111 U703 ( .A(alu_i_data_B[20]), .B(n165), .C(n256), .D(n187), .Q(n232)
         );
  OAI210 U704 ( .A(alu_i_data_B[14]), .B(n164), .C(n189), .Q(n218) );
  IMAJ30 U705 ( .A(n154), .B(alu_i_data_B[13]), .C(n208), .Q(n219) );
  NAND20 U706 ( .A(alu_i_data_B[22]), .B(n163), .Q(n228) );
  IMAJ30 U707 ( .A(n159), .B(alu_i_data_B[23]), .C(n255), .Q(n236) );
  XOR21 U708 ( .A(u_alu_pre_sum_3a[8]), .B(u_alu_DP_OP_83J3_124_3384_n1), .Q(
        u_alu_pre_sum_3b[8]) );
  ADD31 U709 ( .A(compare_i_data_rs[17]), .B(alu_i_data_B[17]), .CI(
        u_alu_DP_OP_83J3_124_3384_n15), .CO(u_alu_DP_OP_83J3_124_3384_n14), 
        .S(u_alu_pre_sum_3a[1]) );
  XOR31 U710 ( .A(alu_i_data_B[31]), .B(u_alu_DP_OP_84J3_125_2615_n9), .C(
        compare_i_data_rs[31]), .Q(u_alu_pre_sum_4a[7]) );
  IMUX21 U711 ( .A(n260), .B(u_alu_pre_sum_4a[7]), .S(
        u_alu_DP_OP_84J3_125_2615_n1), .Q(u_alu_pre_sum_4b[7]) );
  XNR31 U712 ( .A(alu_i_data_B[31]), .B(u_alu_DP_OP_85J3_126_1427_n32), .C(
        compare_i_data_rs[31]), .Q(u_alu_pre_suba[15]) );
  XNR21 U713 ( .A(alu_i_data_B[16]), .B(compare_i_data_rs[16]), .Q(
        u_alu_pre_subb[0]) );
  XOR31 U714 ( .A(u_alu_DP_OP_85J3_126_1427_n43), .B(compare_i_data_rs[20]), 
        .C(n145), .Q(u_alu_pre_suba[4]) );
  XNR21 U715 ( .A(u_alu_pre_suba[14]), .B(n274), .Q(u_alu_pre_subb[14]) );
  XNR21 U716 ( .A(u_alu_pre_suba[4]), .B(n263), .Q(u_alu_pre_subb[4]) );
  XNR21 U717 ( .A(u_alu_pre_suba[10]), .B(n269), .Q(u_alu_pre_subb[10]) );
  XNR21 U718 ( .A(u_alu_pre_suba[12]), .B(n271), .Q(u_alu_pre_subb[12]) );
  XNR21 U719 ( .A(u_alu_pre_suba[6]), .B(n265), .Q(u_alu_pre_subb[6]) );
  XNR21 U720 ( .A(u_alu_pre_suba[8]), .B(n267), .Q(u_alu_pre_subb[8]) );
  INV3 U721 ( .A(alu_i_data_B[19]), .Q(n275) );
  NAND22 U722 ( .A(alu_i_data_B[16]), .B(n138), .Q(
        u_alu_DP_OP_85J3_126_1427_n46) );
  NAND22 U723 ( .A(u_alu_DP_OP_85J3_126_1427_n43), .B(compare_i_data_rs[20]), 
        .Q(n289) );
  NAND22 U724 ( .A(u_alu_DP_OP_85J3_126_1427_n43), .B(n145), .Q(n288) );
  NAND22 U725 ( .A(compare_i_data_rs[20]), .B(n145), .Q(n287) );
  NOR31 U726 ( .A(u_alu_pre_suba[2]), .B(u_alu_pre_suba[1]), .C(n276), .Q(n262) );
  INV3 U727 ( .A(u_alu_pre_suba[3]), .Q(n278) );
  NAND22 U728 ( .A(n262), .B(n278), .Q(n263) );
  NOR21 U729 ( .A(u_alu_pre_suba[4]), .B(n263), .Q(n264) );
  INV3 U730 ( .A(u_alu_pre_suba[5]), .Q(n279) );
  NAND22 U731 ( .A(n264), .B(n279), .Q(n265) );
  NOR21 U732 ( .A(u_alu_pre_suba[6]), .B(n265), .Q(n266) );
  INV3 U733 ( .A(u_alu_pre_suba[7]), .Q(n280) );
  NAND22 U734 ( .A(n266), .B(n280), .Q(n267) );
  NOR21 U735 ( .A(u_alu_pre_suba[8]), .B(n267), .Q(n268) );
  INV3 U736 ( .A(u_alu_pre_suba[9]), .Q(n281) );
  NAND22 U737 ( .A(n268), .B(n281), .Q(n269) );
  NOR21 U738 ( .A(u_alu_pre_suba[10]), .B(n269), .Q(n270) );
  INV3 U739 ( .A(u_alu_pre_suba[11]), .Q(n282) );
  NAND22 U740 ( .A(n270), .B(n282), .Q(n271) );
  NOR21 U741 ( .A(u_alu_pre_suba[12]), .B(n271), .Q(n272) );
  XOR21 U742 ( .A(u_alu_DP_OP_85J3_126_1427_n34), .B(n286), .Q(
        u_alu_pre_suba[13]) );
  NAND22 U743 ( .A(n272), .B(n283), .Q(n274) );
  NAND22 U744 ( .A(n292), .B(n291), .Q(n290) );
  OAI311 U745 ( .A(n274), .B(u_alu_pre_suba[14]), .C(u_alu_pre_suba[15]), .D(
        n273), .Q(u_alu_pre_subb[15]) );
  NOR21 U746 ( .A(u_alu_pre_suba[1]), .B(n276), .Q(n261) );
  NAND22 U747 ( .A(u_alu_DP_OP_85J3_126_1427_n34), .B(compare_i_data_rs[29]), 
        .Q(n285) );
  NAND22 U748 ( .A(u_alu_DP_OP_85J3_126_1427_n34), .B(n129), .Q(n284) );
  IMUX21 U749 ( .A(n277), .B(u_alu_pre_suba[2]), .S(n261), .Q(
        u_alu_pre_subb[2]) );
  NAND22 U750 ( .A(n290), .B(u_alu_pre_suba[15]), .Q(n273) );
  NAND33 U751 ( .A(n289), .B(n288), .C(n287), .Q(u_alu_DP_OP_85J3_126_1427_n42) );
  IMUX21 U752 ( .A(n278), .B(u_alu_pre_suba[3]), .S(n262), .Q(
        u_alu_pre_subb[3]) );
  ADD32 U753 ( .A(n130), .B(compare_i_data_rs[30]), .CI(
        u_alu_DP_OP_85J3_126_1427_n33), .CO(u_alu_DP_OP_85J3_126_1427_n32), 
        .S(u_alu_pre_suba[14]) );
  ADD32 U754 ( .A(n132), .B(compare_i_data_rs[26]), .CI(
        u_alu_DP_OP_85J3_126_1427_n37), .CO(u_alu_DP_OP_85J3_126_1427_n36), 
        .S(u_alu_pre_suba[10]) );
  ADD32 U755 ( .A(n128), .B(compare_i_data_rs[27]), .CI(
        u_alu_DP_OP_85J3_126_1427_n36), .CO(u_alu_DP_OP_85J3_126_1427_n35), 
        .S(u_alu_pre_suba[11]) );
  ADD32 U756 ( .A(n144), .B(compare_i_data_rs[18]), .CI(
        u_alu_DP_OP_85J3_126_1427_n45), .CO(u_alu_DP_OP_85J3_126_1427_n44), 
        .S(u_alu_pre_suba[2]) );
  ADD32 U757 ( .A(n275), .B(compare_i_data_rs[19]), .CI(
        u_alu_DP_OP_85J3_126_1427_n44), .CO(u_alu_DP_OP_85J3_126_1427_n43), 
        .S(u_alu_pre_suba[3]) );
  ADD32 U758 ( .A(n131), .B(compare_i_data_rs[24]), .CI(
        u_alu_DP_OP_85J3_126_1427_n39), .CO(u_alu_DP_OP_85J3_126_1427_n38), 
        .S(u_alu_pre_suba[8]) );
  ADD32 U759 ( .A(n142), .B(compare_i_data_rs[25]), .CI(
        u_alu_DP_OP_85J3_126_1427_n38), .CO(u_alu_DP_OP_85J3_126_1427_n37), 
        .S(u_alu_pre_suba[9]) );
  ADD32 U760 ( .A(n126), .B(compare_i_data_rs[17]), .CI(
        u_alu_DP_OP_85J3_126_1427_n46), .CO(u_alu_DP_OP_85J3_126_1427_n45), 
        .S(u_alu_pre_suba[1]) );
  ADD32 U761 ( .A(n148), .B(compare_i_data_rs[23]), .CI(
        u_alu_DP_OP_85J3_126_1427_n40), .CO(u_alu_DP_OP_85J3_126_1427_n39), 
        .S(u_alu_pre_suba[7]) );
  ADD32 U762 ( .A(n146), .B(compare_i_data_rs[22]), .CI(
        u_alu_DP_OP_85J3_126_1427_n41), .CO(u_alu_DP_OP_85J3_126_1427_n40), 
        .S(u_alu_pre_suba[6]) );
  NAND23 U763 ( .A(n729), .B(i_con_Efbmux[1]), .Q(n839) );
  NOR24 U764 ( .A(n730), .B(n300), .Q(n861) );
  NOR23 U765 ( .A(compare_i_data_rs[7]), .B(u_alu_lt_x_11_B_7_), .Q(
        u_alu_add_x_1_n14) );
  AOI221 U766 ( .A(n302), .B(i_data_FMalures[17]), .C(n300), .D(
        i_data_FEalures[17]), .Q(n800) );
  NAND33 U767 ( .A(n801), .B(n800), .C(n799), .Q(compare_i_data_rt[17]) );
  AOI220 U768 ( .A(n998), .B(u_alu_sum_1_4_), .C(u_alu_N229), .D(n1180), .Q(
        n892) );
  OAI2111 U769 ( .A(compare_i_data_rs[6]), .B(n1195), .C(n1196), .D(n1197), 
        .Q(alu_o_data_AluRes[6]) );
  AOI211 U770 ( .A(alu_i_data_B[6]), .B(n141), .C(n1199), .Q(n1196) );
  NAND20 U771 ( .A(u_alu_N226), .B(n1180), .Q(n901) );
  AOI210 U772 ( .A(n995), .B(compare_i_data_rs[15]), .C(n994), .Q(n996) );
  IMUX20 U773 ( .A(alu_i_data_B[13]), .B(alu_i_data_B[14]), .S(
        i_data_immext[6]), .Q(n462) );
  AOI211 U774 ( .A(compare_i_data_rs[8]), .B(n1187), .C(n1188), .Q(n1186) );
  IMUX20 U775 ( .A(alu_i_data_B[14]), .B(alu_i_data_B[15]), .S(
        i_data_immext[6]), .Q(n448) );
  IMUX20 U776 ( .A(alu_i_data_B[12]), .B(alu_i_data_B[13]), .S(
        i_data_immext[6]), .Q(n445) );
  IMUX21 U777 ( .A(n507), .B(n506), .S(u_alu_ashr_4_SH_3_), .Q(n553) );
  IMUX21 U778 ( .A(n501), .B(n500), .S(u_alu_ashr_4_SH_3_), .Q(n543) );
  IMUX21 U779 ( .A(n489), .B(n488), .S(u_alu_ashr_4_SH_3_), .Q(n532) );
  IMUX21 U780 ( .A(n378), .B(n377), .S(u_alu_ashr_4_SH_3_), .Q(n425) );
  IMUX21 U781 ( .A(n343), .B(n344), .S(u_alu_ashr_4_SH_3_), .Q(n390) );
  IMUX21 U782 ( .A(n353), .B(n354), .S(u_alu_ashr_4_SH_3_), .Q(n404) );
  IMUX21 U783 ( .A(n555), .B(n508), .S(u_alu_ashr_4_SH_3_), .Q(n481) );
  IMUX21 U784 ( .A(n371), .B(n370), .S(u_alu_ashr_4_SH_3_), .Q(n424) );
  IMUX21 U785 ( .A(n487), .B(n486), .S(u_alu_ashr_4_SH_3_), .Q(n521) );
  IMUX21 U786 ( .A(n504), .B(n503), .S(u_alu_ashr_4_SH_3_), .Q(n548) );
  IMUX21 U787 ( .A(n348), .B(n349), .S(u_alu_ashr_4_SH_3_), .Q(n397) );
  IMUX21 U788 ( .A(n339), .B(n340), .S(u_alu_ashr_4_SH_3_), .Q(n384) );
  IMUX21 U789 ( .A(n499), .B(n498), .S(u_alu_ashr_4_SH_3_), .Q(n537) );
  IMUX20 U790 ( .A(alu_i_data_B[28]), .B(alu_i_data_B[29]), .S(
        i_data_immext[6]), .Q(n453) );
  IMUX20 U791 ( .A(alu_i_data_B[26]), .B(alu_i_data_B[27]), .S(
        i_data_immext[6]), .Q(n454) );
  IMUX21 U792 ( .A(n358), .B(n359), .S(u_alu_ashr_4_SH_3_), .Q(n410) );
  IMUX20 U793 ( .A(alu_i_data_B[14]), .B(alu_i_data_B[13]), .S(
        i_data_immext[6]), .Q(n326) );
  IMUX20 U794 ( .A(alu_i_data_B[28]), .B(alu_i_data_B[27]), .S(
        i_data_immext[6]), .Q(n407) );
  IMUX21 U795 ( .A(n559), .B(n509), .S(u_alu_ashr_4_SH_3_), .Q(n495) );
  IMUX20 U796 ( .A(alu_i_data_B[29]), .B(alu_i_data_B[30]), .S(
        i_data_immext[6]), .Q(n470) );
  IMUX20 U797 ( .A(alu_i_data_B[27]), .B(alu_i_data_B[28]), .S(
        i_data_immext[6]), .Q(n467) );
  IMUX21 U798 ( .A(n363), .B(n364), .S(u_alu_ashr_4_SH_3_), .Q(n417) );
  IMUX20 U799 ( .A(alu_i_data_B[13]), .B(alu_i_data_B[12]), .S(
        i_data_immext[6]), .Q(n322) );
  IMUX20 U800 ( .A(alu_i_data_B[15]), .B(alu_i_data_B[14]), .S(
        i_data_immext[6]), .Q(n332) );
  IMUX20 U801 ( .A(alu_i_data_B[27]), .B(alu_i_data_B[26]), .S(
        i_data_immext[6]), .Q(n399) );
  IMUX20 U802 ( .A(alu_i_data_B[29]), .B(alu_i_data_B[28]), .S(
        i_data_immext[6]), .Q(n411) );
  NOR23 U803 ( .A(n1078), .B(u_alu_N173), .Q(n1074) );
  AOI221 U804 ( .A(n721), .B(i_data_FMalures[0]), .C(n573), .D(
        i_data_FEalures[0]), .Q(n724) );
  AOI221 U805 ( .A(n301), .B(i_data_FMmemout[0]), .C(n863), .D(
        i_data_FWmemout[0]), .Q(n865) );
  NOR21 U806 ( .A(n712), .B(n711), .Q(n717) );
  MUX22 U807 ( .A(compare_i_data_rt[1]), .B(i_data_immext[1]), .S(n305), .Q(
        alu_i_data_B[1]) );
  AOI221 U808 ( .A(n301), .B(i_data_FMmemout[1]), .C(n863), .D(
        i_data_FWmemout[1]), .Q(n858) );
  NAND33 U809 ( .A(n710), .B(n709), .C(n708), .Q(compare_i_data_rs[2]) );
  AOI2111 U810 ( .A(i_data_FMalures[3]), .B(n721), .C(n705), .D(n704), .Q(n706) );
  AOI221 U811 ( .A(n302), .B(i_data_FMalures[4]), .C(n300), .D(
        i_data_FEalures[4]), .Q(n853) );
  NAND20 U812 ( .A(n169), .B(i_data_FMmemout[5]), .Q(n688) );
  NAND22 U813 ( .A(n296), .B(i_data_rs[5]), .Q(n693) );
  AOI220 U814 ( .A(n302), .B(i_data_FMalures[5]), .C(n300), .D(
        i_data_FEalures[5]), .Q(n850) );
  NAND20 U815 ( .A(n169), .B(i_data_FMmemout[6]), .Q(n681) );
  NAND20 U816 ( .A(n169), .B(i_data_FMmemout[7]), .Q(n674) );
  AOI220 U817 ( .A(n302), .B(i_data_FMalures[7]), .C(n300), .D(
        i_data_FEalures[7]), .Q(n844) );
  BUF6 U818 ( .A(i_data_immext[9]), .Q(u_alu_ashr_4_SH_3_) );
  AOI211 U819 ( .A(n139), .B(i_data_rt[11]), .C(n827), .Q(n828) );
  AOI211 U820 ( .A(n168), .B(i_data_rt[12]), .C(n823), .Q(n824) );
  AOI211 U821 ( .A(n139), .B(i_data_rt[13]), .C(n819), .Q(n820) );
  AOI211 U822 ( .A(n720), .B(i_data_rs[14]), .C(n653), .Q(n654) );
  MUX22 U823 ( .A(compare_i_data_rt[15]), .B(i_data_immext[15]), .S(n305), .Q(
        alu_i_data_B[15]) );
  NOR21 U824 ( .A(i_data_immext[3]), .B(i_data_immext[1]), .Q(n1246) );
  NAND22 U825 ( .A(n168), .B(i_data_rt[20]), .Q(n790) );
  NAND22 U826 ( .A(n296), .B(i_data_rs[20]), .Q(n624) );
  AOI220 U827 ( .A(n169), .B(i_data_FMmemout[16]), .C(n574), .D(
        i_data_FWmemout[16]), .Q(n646) );
  AOI220 U828 ( .A(n301), .B(i_data_FMmemout[16]), .C(n863), .D(
        i_data_FWmemout[16]), .Q(n803) );
  AOI220 U829 ( .A(n301), .B(i_data_FMmemout[18]), .C(n863), .D(
        i_data_FWmemout[18]), .Q(n795) );
  NOR21 U830 ( .A(n625), .B(n711), .Q(n629) );
  NAND22 U831 ( .A(n296), .B(i_data_rs[19]), .Q(n631) );
  NAND22 U832 ( .A(n168), .B(i_data_rt[19]), .Q(n794) );
  AOI211 U833 ( .A(n139), .B(i_data_rt[23]), .C(n775), .Q(n776) );
  AOI211 U834 ( .A(n139), .B(i_data_rt[25]), .C(n765), .Q(n766) );
  AOI211 U835 ( .A(n168), .B(i_data_rt[27]), .C(n755), .Q(n756) );
  NAND22 U836 ( .A(n580), .B(n579), .Q(n714) );
  AOI211 U837 ( .A(n168), .B(i_data_rt[28]), .C(n750), .Q(n751) );
  NOR31 U838 ( .A(n732), .B(i_con_Efbmux[1]), .C(i_con_Efbmux[2]), .Q(n862) );
  AOI221 U839 ( .A(n169), .B(i_data_FMmemout[9]), .C(n721), .D(
        i_data_FMalures[9]), .Q(n667) );
  IMUX20 U840 ( .A(n493), .B(n483), .S(i_data_immext[8]), .Q(n541) );
  IMUX20 U841 ( .A(n551), .B(n477), .S(i_data_immext[8]), .Q(n530) );
  IMUX20 U842 ( .A(n546), .B(n472), .S(i_data_immext[8]), .Q(n519) );
  IMUX20 U843 ( .A(n362), .B(n342), .S(i_data_immext[8]), .Q(n388) );
  IMUX21 U844 ( .A(n334), .B(n336), .S(i_data_immext[8]), .Q(n354) );
  IMUX20 U845 ( .A(n374), .B(n352), .S(i_data_immext[8]), .Q(n402) );
  AOI311 U846 ( .A(i_con_bop[0]), .B(n967), .C(n966), .D(n965), .Q(n968) );
  NOR40 U847 ( .A(n934), .B(n933), .C(n932), .D(n931), .Q(n1300) );
  IMUX21 U848 ( .A(n329), .B(n328), .S(i_data_immext[8]), .Q(n371) );
  IMUX20 U849 ( .A(n347), .B(n327), .S(i_data_immext[8]), .Q(n368) );
  IMUX20 U850 ( .A(n357), .B(n338), .S(i_data_immext[8]), .Q(n382) );
  IMUX20 U851 ( .A(n367), .B(n347), .S(i_data_immext[8]), .Q(n395) );
  IMUX21 U852 ( .A(n321), .B(n320), .S(i_data_immext[8]), .Q(n359) );
  IMUX20 U853 ( .A(n381), .B(n357), .S(i_data_immext[8]), .Q(n409) );
  IMUX21 U854 ( .A(n485), .B(n484), .S(i_data_immext[8]), .Q(n509) );
  IMUX21 U855 ( .A(n335), .B(n334), .S(i_data_immext[8]), .Q(n378) );
  IMUX20 U856 ( .A(n352), .B(n333), .S(i_data_immext[8]), .Q(n375) );
  IMUX21 U857 ( .A(n325), .B(n324), .S(i_data_immext[8]), .Q(n364) );
  IMUX20 U858 ( .A(n387), .B(n362), .S(i_data_immext[8]), .Q(n415) );
  MUX26 U859 ( .A(compare_i_data_rt[0]), .B(i_data_immext[0]), .S(n305), .Q(
        alu_i_data_B[0]) );
  NAND33 U860 ( .A(n867), .B(n866), .C(n865), .Q(compare_i_data_rt[0]) );
  AOI221 U861 ( .A(n302), .B(i_data_FMalures[0]), .C(n300), .D(
        i_data_FEalures[0]), .Q(n866) );
  OAI212 U862 ( .A(n715), .B(n714), .C(n713), .Q(n716) );
  AOI220 U863 ( .A(n169), .B(i_data_FMmemout[10]), .C(n721), .D(
        i_data_FMalures[10]), .Q(n664) );
  NOR32 U864 ( .A(n731), .B(i_con_Efbmux[1]), .C(i_con_Efbmux[0]), .Q(n864) );
  IMUX21 U865 ( .A(n482), .B(n485), .S(i_data_immext[8]), .Q(n501) );
  IMUX21 U866 ( .A(n478), .B(n505), .S(i_data_immext[8]), .Q(n488) );
  IMUX21 U867 ( .A(n323), .B(n325), .S(i_data_immext[8]), .Q(n343) );
  IMUX21 U868 ( .A(n333), .B(n335), .S(i_data_immext[8]), .Q(n353) );
  IMUX21 U869 ( .A(n319), .B(n321), .S(i_data_immext[8]), .Q(n339) );
  IMUX21 U870 ( .A(n473), .B(n502), .S(i_data_immext[8]), .Q(n486) );
  IMUX21 U871 ( .A(n338), .B(n319), .S(i_data_immext[8]), .Q(n358) );
  IMUX21 U872 ( .A(n322), .B(n312), .S(u_alu_ashr_4_SH_1_), .Q(n333) );
  AOI221 U873 ( .A(n302), .B(i_data_FMalures[1]), .C(n300), .D(
        i_data_FEalures[1]), .Q(n859) );
  NAND22 U874 ( .A(n169), .B(i_data_FMmemout[3]), .Q(n702) );
  AOI221 U875 ( .A(n302), .B(i_data_FMalures[3]), .C(n300), .D(
        i_data_FEalures[3]), .Q(n856) );
  AOI220 U876 ( .A(n169), .B(i_data_FMmemout[11]), .C(n721), .D(
        i_data_FMalures[11]), .Q(n661) );
  OAI212 U877 ( .A(n140), .B(n641), .C(n640), .Q(n642) );
  NOR21 U878 ( .A(n639), .B(n711), .Q(n643) );
  AOI221 U879 ( .A(n301), .B(i_data_FMmemout[17]), .C(n863), .D(
        i_data_FWmemout[17]), .Q(n799) );
  IMUX20 U880 ( .A(n526), .B(n525), .S(u_alu_ashr_4_SH_1_), .Q(n529) );
  IMUX20 U881 ( .A(n517), .B(n516), .S(n440), .Q(n547) );
  IMUX20 U882 ( .A(n461), .B(n464), .S(n440), .Q(n477) );
  IMUX20 U883 ( .A(n462), .B(n461), .S(n440), .Q(n493) );
  IMUX20 U884 ( .A(n448), .B(n447), .S(n440), .Q(n472) );
  IMUX20 U885 ( .A(n446), .B(n445), .S(n440), .Q(n546) );
  IMUX20 U886 ( .A(n514), .B(n517), .S(n440), .Q(n536) );
  IMUX20 U887 ( .A(n441), .B(n515), .S(u_alu_ashr_4_SH_1_), .Q(n442) );
  IMUX20 U888 ( .A(n445), .B(n448), .S(n440), .Q(n458) );
  IMUX20 U889 ( .A(n516), .B(n446), .S(n440), .Q(n535) );
  IMUX20 U890 ( .A(n465), .B(n468), .S(n440), .Q(n479) );
  IMUX20 U891 ( .A(n463), .B(n466), .S(n440), .Q(n476) );
  IMUX20 U892 ( .A(n361), .B(n351), .S(n440), .Q(n374) );
  IMUX20 U893 ( .A(n411), .B(n399), .S(u_alu_ashr_4_SH_1_), .Q(n401) );
  IMUX20 U894 ( .A(n447), .B(n450), .S(n440), .Q(n457) );
  IMUX21 U895 ( .A(n459), .B(n497), .S(i_data_immext[8]), .Q(n508) );
  IMUX20 U896 ( .A(n450), .B(n449), .S(n440), .Q(n471) );
  IMUX20 U897 ( .A(n452), .B(n451), .S(n440), .Q(n474) );
  IMUX20 U898 ( .A(n407), .B(n392), .S(u_alu_ashr_4_SH_1_), .Q(n394) );
  IMUX20 U899 ( .A(n449), .B(n452), .S(n440), .Q(n460) );
  IMUX20 U900 ( .A(n318), .B(n306), .S(n440), .Q(n327) );
  IMUX20 U901 ( .A(n337), .B(n326), .S(n440), .Q(n347) );
  IMUX20 U902 ( .A(n356), .B(n346), .S(n440), .Q(n367) );
  IMUX20 U903 ( .A(n326), .B(n318), .S(n440), .Q(n338) );
  IMUX20 U904 ( .A(n346), .B(n337), .S(n440), .Q(n357) );
  IMUX20 U905 ( .A(n366), .B(n356), .S(n440), .Q(n381) );
  IMUX21 U906 ( .A(alu_i_data_B[30]), .B(alu_i_data_B[31]), .S(
        i_data_immext[6]), .Q(n455) );
  IMUX20 U907 ( .A(n466), .B(n465), .S(n440), .Q(n482) );
  IMUX20 U908 ( .A(n464), .B(n463), .S(n440), .Q(n483) );
  IMUX20 U909 ( .A(n341), .B(n332), .S(n440), .Q(n352) );
  IMUX21 U910 ( .A(n342), .B(n323), .S(i_data_immext[8]), .Q(n363) );
  IMUX20 U911 ( .A(n351), .B(n341), .S(n440), .Q(n362) );
  IMUX20 U912 ( .A(n373), .B(n361), .S(n440), .Q(n387) );
  NOR31 U913 ( .A(n882), .B(alu_i_con_AluCtrl[0]), .C(n881), .Q(n1178) );
  INV3 U914 ( .A(n1182), .Q(n576) );
  NAND22 U915 ( .A(n139), .B(i_data_rt[0]), .Q(n867) );
  NAND22 U916 ( .A(n169), .B(i_data_FMmemout[1]), .Q(n713) );
  NAND22 U917 ( .A(n168), .B(i_data_rt[1]), .Q(n860) );
  AOI221 U918 ( .A(n721), .B(i_data_FMalures[2]), .C(n573), .D(
        i_data_FEalures[2]), .Q(n709) );
  NAND22 U919 ( .A(n169), .B(i_data_FMmemout[4]), .Q(n695) );
  AOI220 U920 ( .A(n169), .B(i_data_FMmemout[12]), .C(n721), .D(
        i_data_FMalures[12]), .Q(n658) );
  NOR31 U921 ( .A(n1183), .B(alu_i_con_AluCtrl[0]), .C(alu_i_con_AluCtrl[3]), 
        .Q(n875) );
  OAI2111 U922 ( .A(n1268), .B(n1267), .C(n1266), .D(n1265), .Q(
        alu_i_con_AluCtrl[3]) );
  NOR21 U923 ( .A(n869), .B(n868), .Q(n914) );
  AOI2111 U924 ( .A(n721), .B(i_data_FMalures[17]), .C(n643), .D(n642), .Q(
        n644) );
  IMUX21 U925 ( .A(n327), .B(n329), .S(i_data_immext[8]), .Q(n348) );
  INV6 U926 ( .A(u_alu_sum_1_8_), .Q(DP_OP_77_130_260_I3) );
  INV3 U927 ( .A(n439), .Q(n440) );
  NOR22 U928 ( .A(n881), .B(alu_i_con_AluCtrl[3]), .Q(n1180) );
  MUX26 U929 ( .A(compare_i_data_rt[2]), .B(i_data_immext[2]), .S(n305), .Q(
        alu_i_data_B[2]) );
  OAI212 U930 ( .A(n703), .B(n140), .C(n702), .Q(n704) );
  MUX26 U931 ( .A(compare_i_data_rt[3]), .B(i_data_immext[3]), .S(n305), .Q(
        alu_i_data_B[3]) );
  AOI221 U932 ( .A(n301), .B(i_data_FMmemout[3]), .C(n863), .D(
        i_data_FWmemout[3]), .Q(n855) );
  OAI212 U933 ( .A(n696), .B(n140), .C(n695), .Q(n697) );
  AOI221 U934 ( .A(n301), .B(i_data_FMmemout[4]), .C(n863), .D(
        i_data_FWmemout[4]), .Q(n852) );
  MUX26 U935 ( .A(compare_i_data_rt[6]), .B(i_data_immext[6]), .S(n305), .Q(
        alu_i_data_B[6]) );
  BUF2 U936 ( .A(i_data_immext[7]), .Q(u_alu_ashr_4_SH_1_) );
  AOI221 U937 ( .A(n169), .B(i_data_FMmemout[8]), .C(n721), .D(
        i_data_FMalures[8]), .Q(n670) );
  NAND31 U938 ( .A(n1263), .B(n1266), .C(n1262), .Q(alu_i_con_AluCtrl[2]) );
  AOI220 U939 ( .A(n169), .B(i_data_FMmemout[31]), .C(i_data_FMalures[31]), 
        .D(n721), .Q(n585) );
  NAND22 U940 ( .A(n296), .B(i_data_rs[17]), .Q(n645) );
  OAI212 U941 ( .A(n305), .B(n802), .C(n807), .Q(alu_i_data_B[17]) );
  AOI2111 U942 ( .A(n721), .B(i_data_FMalures[18]), .C(n636), .D(n635), .Q(
        n637) );
  IMUX20 U943 ( .A(n1179), .B(n1178), .S(n136), .Q(n1185) );
  NAND22 U944 ( .A(n1074), .B(u_alu_pre_sum_3a[4]), .Q(n1034) );
  NOR24 U945 ( .A(n1078), .B(n1000), .Q(n1073) );
  NOR21 U946 ( .A(n874), .B(n1184), .Q(n1182) );
  NAND22 U947 ( .A(n296), .B(i_data_rs[3]), .Q(n707) );
  NAND22 U948 ( .A(n139), .B(i_data_rt[3]), .Q(n857) );
  NOR21 U949 ( .A(n694), .B(n711), .Q(n698) );
  OAI212 U950 ( .A(n689), .B(n140), .C(n688), .Q(n690) );
  AOI221 U951 ( .A(n301), .B(i_data_FMmemout[5]), .C(n863), .D(
        i_data_FWmemout[5]), .Q(n849) );
  OAI212 U952 ( .A(n682), .B(n140), .C(n681), .Q(n683) );
  AOI221 U953 ( .A(n301), .B(i_data_FMmemout[6]), .C(n863), .D(
        i_data_FWmemout[6]), .Q(n846) );
  AOI221 U954 ( .A(n301), .B(i_data_FMmemout[7]), .C(n863), .D(
        i_data_FWmemout[7]), .Q(n843) );
  NAND22 U955 ( .A(n875), .B(alu_i_con_AluCtrl[2]), .Q(n999) );
  INV3 U956 ( .A(compare_i_data_rt[17]), .Q(n802) );
  NOR21 U957 ( .A(n632), .B(n711), .Q(n636) );
  NAND22 U958 ( .A(n305), .B(i_data_immext[16]), .Q(n807) );
  INV3 U959 ( .A(n305), .Q(n806) );
  IMUX21 U960 ( .A(n457), .B(n460), .S(i_data_immext[8]), .Q(n555) );
  NAND22 U961 ( .A(n1168), .B(u_alu_pre_sum_4a[0]), .Q(n1089) );
  IMUX21 U962 ( .A(n483), .B(n482), .S(i_data_immext[8]), .Q(n559) );
  NAND22 U963 ( .A(n1168), .B(u_alu_pre_sum_4a[7]), .Q(n1169) );
  AOI2112 U964 ( .A(u_alu_pre_sum_3b[8]), .B(u_alu_N173), .C(n1079), .D(n1078), 
        .Q(n1168) );
  NOR21 U965 ( .A(u_alu_N173), .B(n1077), .Q(n1079) );
  AOI2111 U966 ( .A(i_data_FMalures[4]), .B(n721), .C(n698), .D(n697), .Q(n699) );
  OAI212 U967 ( .A(n675), .B(n140), .C(n674), .Q(n676) );
  NOR31 U968 ( .A(i_data_immext[2]), .B(i_data_immext[0]), .C(i_data_immext[1]), .Q(n870) );
  AOI2111 U969 ( .A(i_data_FMalures[20]), .B(n721), .C(n622), .D(n621), .Q(
        n623) );
  AOI220 U970 ( .A(n302), .B(i_data_FMalures[16]), .C(n300), .D(
        i_data_FEalures[16]), .Q(n804) );
  AOI2111 U971 ( .A(n721), .B(i_data_FMalures[19]), .C(n629), .D(n628), .Q(
        n630) );
  INV3 U972 ( .A(i_con_Efbmux[0]), .Q(n732) );
  INV3 U973 ( .A(i_con_Efbmux[2]), .Q(n731) );
  IMUX20 U974 ( .A(n1178), .B(n1179), .S(u_alu_lt_x_11_B_1_), .Q(n1229) );
  AOI210 U975 ( .A(n972), .B(compare_i_data_rs[9]), .C(n971), .Q(n974) );
  AOI210 U976 ( .A(n982), .B(compare_i_data_rs[10]), .C(n981), .Q(n984) );
  AOI211 U977 ( .A(alu_i_con_AluCtrl[0]), .B(n1238), .C(n1239), .Q(n1237) );
  AOI221 U978 ( .A(n906), .B(u_alu_half_sub_0_), .C(n998), .D(u_alu_sum_1_0_), 
        .Q(n907) );
  AOI211 U979 ( .A(n575), .B(u_alu_N209), .C(n1006), .Q(n1008) );
  OAI2111 U980 ( .A(n1023), .B(n1235), .C(n1005), .D(n1004), .Q(n1006) );
  NAND22 U981 ( .A(n1158), .B(u_alu_pre_subb[0]), .Q(n1012) );
  IMUX21 U982 ( .A(n453), .B(n455), .S(n440), .Q(n497) );
  NAND22 U983 ( .A(alu_i_data_B[2]), .B(compare_i_data_rs[2]), .Q(
        u_alu_add_x_1_n37) );
  NOR21 U984 ( .A(compare_i_data_rs[2]), .B(alu_i_data_B[2]), .Q(
        u_alu_add_x_1_n36) );
  AOI2111 U985 ( .A(i_data_FMalures[5]), .B(n721), .C(n691), .D(n690), .Q(n692) );
  AOI2111 U986 ( .A(i_data_FMalures[6]), .B(n721), .C(n684), .D(n683), .Q(n685) );
  NOR21 U987 ( .A(n914), .B(n924), .Q(n915) );
  INV3 U988 ( .A(compare_i_data_rt[18]), .Q(n798) );
  INV3 U989 ( .A(compare_i_data_rt[19]), .Q(n935) );
  AOI220 U990 ( .A(n301), .B(i_data_FMmemout[19]), .C(n863), .D(
        i_data_FWmemout[19]), .Q(n792) );
  INV6 U991 ( .A(n295), .Q(n297) );
  NAND22 U992 ( .A(n1293), .B(n1288), .Q(o_addr_Erd[0]) );
  NAND22 U993 ( .A(n1293), .B(n1290), .Q(o_addr_Erd[2]) );
  NAND22 U994 ( .A(n1293), .B(n1292), .Q(o_addr_Erd[4]) );
  NAND22 U995 ( .A(n1293), .B(n1291), .Q(o_addr_Erd[3]) );
  NAND22 U996 ( .A(n1293), .B(n1289), .Q(o_addr_Erd[1]) );
  OAI2111 U997 ( .A(compare_i_data_rs[7]), .B(n1190), .C(n1191), .D(n1192), 
        .Q(alu_o_data_AluRes[7]) );
  NAND31 U998 ( .A(n885), .B(n884), .C(n883), .Q(n1194) );
  IMUX20 U999 ( .A(n303), .B(n1184), .S(alu_i_data_B[2]), .Q(n1219) );
  NAND31 U1000 ( .A(n900), .B(n899), .C(n898), .Q(n1220) );
  IMUX20 U1001 ( .A(n1178), .B(n1179), .S(alu_i_data_B[2]), .Q(n1216) );
  IMUX20 U1002 ( .A(n303), .B(n1184), .S(alu_i_data_B[4]), .Q(n1208) );
  NAND31 U1003 ( .A(n894), .B(n893), .C(n892), .Q(n1209) );
  IMUX20 U1004 ( .A(n1178), .B(n1179), .S(alu_i_data_B[4]), .Q(n1205) );
  IMUX20 U1005 ( .A(n303), .B(n1184), .S(alu_i_data_B[3]), .Q(n1213) );
  NAND31 U1006 ( .A(n897), .B(n896), .C(n895), .Q(n1214) );
  IMUX20 U1007 ( .A(n1178), .B(n1179), .S(alu_i_data_B[3]), .Q(n1210) );
  IMUX20 U1008 ( .A(n303), .B(n1184), .S(alu_i_data_B[6]), .Q(n1198) );
  NAND31 U1009 ( .A(n888), .B(n887), .C(n886), .Q(n1199) );
  IMUX20 U1010 ( .A(n1178), .B(n1179), .S(alu_i_data_B[6]), .Q(n1195) );
  NAND31 U1011 ( .A(n903), .B(n902), .C(n901), .Q(n1233) );
  IMUX20 U1012 ( .A(alu_i_data_B[3]), .B(alu_i_data_B[4]), .S(i_data_immext[6]), .Q(n526) );
  IMUX20 U1013 ( .A(u_alu_lt_x_11_B_1_), .B(alu_i_data_B[2]), .S(
        i_data_immext[6]), .Q(n490) );
  IMUX20 U1014 ( .A(n303), .B(n1184), .S(n294), .Q(n1203) );
  NAND31 U1015 ( .A(n891), .B(n890), .C(n889), .Q(n1204) );
  IMUX20 U1016 ( .A(u_alu_lt_x_11_B_7_), .B(alu_i_data_B[8]), .S(
        i_data_immext[6]), .Q(n528) );
  IMUX20 U1017 ( .A(n294), .B(alu_i_data_B[6]), .S(i_data_immext[6]), .Q(n525)
         );
  IMUX20 U1018 ( .A(n1178), .B(n1179), .S(n294), .Q(n1200) );
  IMUX20 U1019 ( .A(n480), .B(n524), .S(i_data_immext[10]), .Q(u_alu_N240) );
  OAI2111 U1020 ( .A(n999), .B(n979), .C(n978), .D(n977), .Q(
        alu_o_data_AluRes[9]) );
  NAND22 U1021 ( .A(u_alu_N202), .B(n575), .Q(n977) );
  NOR21 U1022 ( .A(n437), .B(n435), .Q(u_alu_N202) );
  INV3 U1023 ( .A(n425), .Q(n435) );
  AOI211 U1024 ( .A(n1180), .B(u_alu_N234), .C(n976), .Q(n978) );
  OAI2111 U1025 ( .A(n975), .B(n160), .C(n974), .D(n973), .Q(n976) );
  IMUX20 U1026 ( .A(alu_i_data_B[15]), .B(alu_i_data_B[16]), .S(
        i_data_immext[6]), .Q(n461) );
  IMUX20 U1027 ( .A(alu_i_data_B[11]), .B(alu_i_data_B[12]), .S(
        i_data_immext[6]), .Q(n492) );
  IMUX20 U1028 ( .A(alu_i_data_B[9]), .B(u_alu_lt_x_11_B_10_), .S(
        i_data_immext[6]), .Q(n527) );
  INV3 U1029 ( .A(u_alu_half_sub_9_), .Q(n979) );
  OAI2111 U1030 ( .A(n999), .B(n989), .C(n988), .D(n987), .Q(
        alu_o_data_AluRes[10]) );
  NAND22 U1031 ( .A(u_alu_N203), .B(n575), .Q(n987) );
  AOI211 U1032 ( .A(n998), .B(u_alu_N167), .C(n986), .Q(n988) );
  OAI2111 U1033 ( .A(n985), .B(n293), .C(n984), .D(n983), .Q(n986) );
  MUX21 U1034 ( .A(n456), .B(n510), .S(i_data_immext[10]), .Q(u_alu_N235) );
  INV3 U1035 ( .A(u_alu_half_sub_10_), .Q(n989) );
  OAI2111 U1036 ( .A(n576), .B(n1235), .C(n1236), .D(n1237), .Q(
        alu_o_data_AluRes[0]) );
  NAND22 U1037 ( .A(n908), .B(n907), .Q(n1239) );
  IMUX20 U1038 ( .A(n1184), .B(n303), .S(n1235), .Q(n1240) );
  IMUX20 U1039 ( .A(n1179), .B(n1178), .S(n1235), .Q(n905) );
  INV3 U1040 ( .A(u_alu_N306), .Q(n1242) );
  AOI221 U1041 ( .A(n575), .B(u_alu_N193), .C(n1180), .D(u_alu_N225), .Q(n1236) );
  IMUX20 U1042 ( .A(alu_i_data_B[6]), .B(u_alu_lt_x_11_B_7_), .S(
        i_data_immext[6]), .Q(n517) );
  IMUX20 U1043 ( .A(alu_i_data_B[4]), .B(n294), .S(i_data_immext[6]), .Q(n514)
         );
  IMUX20 U1044 ( .A(alu_i_data_B[2]), .B(alu_i_data_B[3]), .S(i_data_immext[6]), .Q(n515) );
  IMUX20 U1045 ( .A(alu_i_data_B[0]), .B(u_alu_lt_x_11_B_1_), .S(
        i_data_immext[6]), .Q(n441) );
  NOR21 U1046 ( .A(n437), .B(n426), .Q(u_alu_N193) );
  NAND41 U1047 ( .A(n879), .B(n878), .C(n877), .D(n876), .Q(n1188) );
  NAND22 U1048 ( .A(u_alu_half_sub_8_), .B(n906), .Q(n876) );
  MUX21 U1049 ( .A(n558), .B(n557), .S(i_data_immext[10]), .Q(u_alu_N233) );
  IMUX20 U1050 ( .A(u_alu_lt_x_11_B_10_), .B(alu_i_data_B[11]), .S(
        i_data_immext[6]), .Q(n446) );
  IMUX20 U1051 ( .A(alu_i_data_B[8]), .B(alu_i_data_B[9]), .S(i_data_immext[6]), .Q(n516) );
  NOR21 U1052 ( .A(n437), .B(n434), .Q(u_alu_N201) );
  INV3 U1053 ( .A(n424), .Q(n434) );
  NAND31 U1054 ( .A(n1072), .B(n1071), .C(n1070), .Q(alu_o_data_AluRes[23]) );
  NAND22 U1055 ( .A(n1174), .B(u_alu_pre_suba[7]), .Q(n1070) );
  NOR21 U1056 ( .A(n437), .B(n553), .Q(u_alu_N248) );
  NOR21 U1057 ( .A(u_alu_ashr_4_SH_3_), .B(n364), .Q(n423) );
  NAND22 U1058 ( .A(n1158), .B(u_alu_pre_subb[7]), .Q(n1072) );
  NAND31 U1059 ( .A(n1052), .B(n1051), .C(n1050), .Q(alu_o_data_AluRes[21]) );
  NAND22 U1060 ( .A(n1174), .B(u_alu_pre_suba[5]), .Q(n1050) );
  NOR21 U1061 ( .A(n437), .B(n568), .Q(u_alu_N246) );
  NOR21 U1062 ( .A(u_alu_ashr_4_SH_3_), .B(n354), .Q(n421) );
  NAND22 U1063 ( .A(n1158), .B(u_alu_pre_subb[5]), .Q(n1052) );
  NAND22 U1064 ( .A(n1158), .B(u_alu_pre_subb[3]), .Q(n1025) );
  NAND22 U1065 ( .A(n1174), .B(u_alu_pre_suba[3]), .Q(n1026) );
  NAND22 U1066 ( .A(n1074), .B(u_alu_pre_sum_3a[3]), .Q(n1027) );
  NOR21 U1067 ( .A(u_alu_ashr_4_SH_3_), .B(n344), .Q(n419) );
  NAND31 U1068 ( .A(n1106), .B(n1105), .C(n1104), .Q(alu_o_data_AluRes[25]) );
  NAND22 U1069 ( .A(n1174), .B(u_alu_pre_suba[9]), .Q(n1104) );
  AOI211 U1070 ( .A(n1168), .B(u_alu_pre_sum_4a[1]), .C(n1103), .Q(n1105) );
  NAND22 U1071 ( .A(n1167), .B(u_alu_pre_sum_4b[1]), .Q(n1099) );
  NOR21 U1072 ( .A(n437), .B(n567), .Q(u_alu_N250) );
  NOR21 U1073 ( .A(u_alu_ashr_4_SH_3_), .B(n509), .Q(n561) );
  NAND22 U1074 ( .A(n1158), .B(u_alu_pre_subb[9]), .Q(n1106) );
  NAND22 U1075 ( .A(n1174), .B(u_alu_pre_suba[11]), .Q(n1132) );
  AOI211 U1076 ( .A(n1168), .B(u_alu_pre_sum_4a[3]), .C(n1131), .Q(n1133) );
  NAND22 U1077 ( .A(n1167), .B(u_alu_pre_sum_4b[3]), .Q(n1127) );
  NOR21 U1078 ( .A(n437), .B(n570), .Q(u_alu_N252) );
  NOR21 U1079 ( .A(u_alu_ashr_4_SH_3_), .B(n488), .Q(n511) );
  NAND22 U1080 ( .A(n438), .B(n324), .Q(n344) );
  NAND22 U1081 ( .A(n1158), .B(u_alu_pre_subb[11]), .Q(n1134) );
  NAND31 U1082 ( .A(n1152), .B(n1151), .C(n1150), .Q(alu_o_data_AluRes[29]) );
  NAND22 U1083 ( .A(n1174), .B(u_alu_pre_suba[13]), .Q(n1150) );
  AOI211 U1084 ( .A(n1168), .B(u_alu_pre_sum_4a[5]), .C(n1149), .Q(n1151) );
  NAND41 U1085 ( .A(n1148), .B(n1147), .C(n1146), .D(n1145), .Q(n1149) );
  NAND22 U1086 ( .A(n1167), .B(u_alu_pre_sum_4b[5]), .Q(n1145) );
  NOR21 U1087 ( .A(u_alu_ashr_4_SH_3_), .B(n500), .Q(n513) );
  NAND22 U1088 ( .A(n438), .B(n484), .Q(n500) );
  NAND22 U1089 ( .A(n1158), .B(u_alu_pre_subb[13]), .Q(n1152) );
  NOR31 U1090 ( .A(i_con_bop[0]), .B(compare_i_data_rs[31]), .C(n1306), .Q(
        n965) );
  NAND41 U1091 ( .A(n956), .B(n955), .C(n954), .D(n953), .Q(n957) );
  NAND41 U1092 ( .A(n952), .B(n951), .C(n950), .D(n949), .Q(n958) );
  NAND22 U1093 ( .A(n948), .B(n947), .Q(n959) );
  NAND31 U1094 ( .A(n946), .B(n1298), .C(n945), .Q(n960) );
  AOI211 U1095 ( .A(n1074), .B(u_alu_pre_sum_3a[0]), .C(n1010), .Q(n1011) );
  OAI2111 U1096 ( .A(u_alu_pre_sum_3a[0]), .B(n1009), .C(n1008), .D(n1007), 
        .Q(n1010) );
  IMUX20 U1097 ( .A(n303), .B(n1184), .S(compare_i_data_rs[16]), .Q(n1003) );
  NAND22 U1098 ( .A(n1093), .B(n1092), .Q(alu_o_data_AluRes[24]) );
  NAND22 U1099 ( .A(n1174), .B(u_alu_pre_suba[8]), .Q(n1092) );
  OAI2111 U1100 ( .A(n1090), .B(u_alu_pre_sum_4a[0]), .C(n1089), .D(n1088), 
        .Q(n1091) );
  AOI211 U1101 ( .A(n1180), .B(u_alu_N249), .C(n1087), .Q(n1088) );
  OAI2111 U1102 ( .A(n131), .B(n1086), .C(n1085), .D(n1084), .Q(n1087) );
  NOR21 U1103 ( .A(n437), .B(n565), .Q(u_alu_N249) );
  NOR21 U1104 ( .A(u_alu_ashr_4_SH_3_), .B(n508), .Q(n557) );
  NAND22 U1105 ( .A(n1158), .B(u_alu_pre_subb[2]), .Q(n1019) );
  NAND22 U1106 ( .A(n1174), .B(u_alu_pre_suba[2]), .Q(n1020) );
  NAND22 U1107 ( .A(n1074), .B(u_alu_pre_sum_3a[2]), .Q(n1021) );
  IMUX20 U1108 ( .A(alu_i_data_B[18]), .B(alu_i_data_B[19]), .S(
        i_data_immext[6]), .Q(n450) );
  NOR21 U1109 ( .A(u_alu_ashr_4_SH_3_), .B(n340), .Q(n406) );
  NAND31 U1110 ( .A(n1062), .B(n1061), .C(n1060), .Q(alu_o_data_AluRes[22]) );
  NAND22 U1111 ( .A(n1174), .B(u_alu_pre_suba[6]), .Q(n1060) );
  NOR21 U1112 ( .A(n437), .B(n548), .Q(u_alu_N247) );
  NOR21 U1113 ( .A(u_alu_ashr_4_SH_3_), .B(n359), .Q(n422) );
  NAND22 U1114 ( .A(n1158), .B(u_alu_pre_subb[6]), .Q(n1062) );
  NAND31 U1115 ( .A(n1143), .B(n1142), .C(n1141), .Q(alu_o_data_AluRes[28]) );
  NAND22 U1116 ( .A(n1174), .B(u_alu_pre_suba[12]), .Q(n1141) );
  AOI211 U1117 ( .A(n1168), .B(u_alu_pre_sum_4a[4]), .C(n1140), .Q(n1142) );
  NOR21 U1118 ( .A(n437), .B(n512), .Q(u_alu_N253) );
  NAND31 U1119 ( .A(n571), .B(n438), .C(n497), .Q(n512) );
  NAND22 U1120 ( .A(n1158), .B(u_alu_pre_subb[12]), .Q(n1143) );
  NAND22 U1121 ( .A(n1174), .B(u_alu_pre_suba[10]), .Q(n1118) );
  NAND22 U1122 ( .A(n1167), .B(u_alu_pre_sum_4b[2]), .Q(n1113) );
  NAND22 U1123 ( .A(n438), .B(n320), .Q(n340) );
  NOR21 U1124 ( .A(u_alu_ashr_4_SH_3_), .B(n486), .Q(n510) );
  NAND22 U1125 ( .A(n1158), .B(u_alu_pre_subb[10]), .Q(n1120) );
  NAND31 U1126 ( .A(n1041), .B(n1040), .C(n1039), .Q(alu_o_data_AluRes[20]) );
  NAND22 U1127 ( .A(n1174), .B(u_alu_pre_suba[4]), .Q(n1039) );
  NAND41 U1128 ( .A(n1037), .B(n1036), .C(n1035), .D(n1034), .Q(n1038) );
  IMUX20 U1129 ( .A(alu_i_data_B[24]), .B(alu_i_data_B[25]), .S(
        i_data_immext[6]), .Q(n451) );
  IMUX20 U1130 ( .A(alu_i_data_B[22]), .B(alu_i_data_B[23]), .S(
        i_data_immext[6]), .Q(n452) );
  IMUX20 U1131 ( .A(alu_i_data_B[20]), .B(alu_i_data_B[21]), .S(
        i_data_immext[6]), .Q(n449) );
  NOR21 U1132 ( .A(u_alu_ashr_4_SH_3_), .B(n349), .Q(n420) );
  NAND22 U1133 ( .A(n1158), .B(u_alu_pre_subb[4]), .Q(n1041) );
  NAND22 U1134 ( .A(u_alu_pre_subb[14]), .B(n1158), .Q(n1154) );
  NAND22 U1135 ( .A(n1168), .B(u_alu_pre_sum_4a[6]), .Q(n1155) );
  NAND22 U1136 ( .A(n1174), .B(u_alu_pre_suba[14]), .Q(n1156) );
  AOI211 U1137 ( .A(n1167), .B(u_alu_pre_sum_4b[6]), .C(n1153), .Q(n1157) );
  IMUX20 U1138 ( .A(alu_i_data_B[4]), .B(alu_i_data_B[3]), .S(i_data_immext[6]), .Q(n310) );
  IMUX20 U1139 ( .A(alu_i_data_B[6]), .B(n294), .S(i_data_immext[6]), .Q(n307)
         );
  IMUX20 U1140 ( .A(alu_i_data_B[8]), .B(u_alu_lt_x_11_B_7_), .S(
        i_data_immext[6]), .Q(n308) );
  IMUX20 U1141 ( .A(u_alu_lt_x_11_B_10_), .B(alu_i_data_B[9]), .S(
        i_data_immext[6]), .Q(n306) );
  IMUX20 U1142 ( .A(alu_i_data_B[12]), .B(alu_i_data_B[11]), .S(
        i_data_immext[6]), .Q(n318) );
  IMUX20 U1143 ( .A(alu_i_data_B[16]), .B(alu_i_data_B[15]), .S(
        i_data_immext[6]), .Q(n337) );
  IMUX20 U1144 ( .A(alu_i_data_B[20]), .B(alu_i_data_B[19]), .S(
        i_data_immext[6]), .Q(n356) );
  IMUX20 U1145 ( .A(alu_i_data_B[22]), .B(alu_i_data_B[21]), .S(
        i_data_immext[6]), .Q(n366) );
  IMUX20 U1146 ( .A(alu_i_data_B[24]), .B(alu_i_data_B[23]), .S(
        i_data_immext[6]), .Q(n380) );
  IMUX20 U1147 ( .A(alu_i_data_B[26]), .B(alu_i_data_B[25]), .S(
        i_data_immext[6]), .Q(n392) );
  NAND31 U1148 ( .A(n502), .B(n571), .C(n438), .Q(n523) );
  NOR21 U1149 ( .A(n440), .B(n455), .Q(n502) );
  NAND22 U1150 ( .A(n1158), .B(u_alu_pre_subb[1]), .Q(n1014) );
  NAND22 U1151 ( .A(n1174), .B(u_alu_pre_suba[1]), .Q(n1015) );
  NAND22 U1152 ( .A(n1074), .B(u_alu_pre_sum_3a[1]), .Q(n1016) );
  IMUX20 U1153 ( .A(alu_i_data_B[25]), .B(alu_i_data_B[26]), .S(
        i_data_immext[6]), .Q(n468) );
  IMUX20 U1154 ( .A(alu_i_data_B[23]), .B(alu_i_data_B[24]), .S(
        i_data_immext[6]), .Q(n465) );
  IMUX20 U1155 ( .A(alu_i_data_B[21]), .B(alu_i_data_B[22]), .S(
        i_data_immext[6]), .Q(n466) );
  IMUX20 U1156 ( .A(alu_i_data_B[19]), .B(alu_i_data_B[20]), .S(
        i_data_immext[6]), .Q(n463) );
  NOR21 U1157 ( .A(u_alu_ashr_4_SH_3_), .B(n377), .Q(n345) );
  NAND22 U1158 ( .A(n336), .B(n438), .Q(n377) );
  INV3 U1159 ( .A(i_data_immext[8]), .Q(n438) );
  NOR21 U1160 ( .A(n440), .B(n317), .Q(n336) );
  INV3 U1161 ( .A(n1178), .Q(n1144) );
  INV3 U1162 ( .A(n1161), .Q(n1023) );
  NAND22 U1163 ( .A(n1176), .B(n1175), .Q(alu_o_data_AluRes[31]) );
  AOI211 U1164 ( .A(u_alu_pre_suba[15]), .B(n1174), .C(n1173), .Q(n1175) );
  IMUX20 U1165 ( .A(n294), .B(alu_i_data_B[4]), .S(i_data_immext[6]), .Q(n316)
         );
  IMUX20 U1166 ( .A(u_alu_lt_x_11_B_7_), .B(alu_i_data_B[6]), .S(
        i_data_immext[6]), .Q(n313) );
  IMUX20 U1167 ( .A(alu_i_data_B[9]), .B(alu_i_data_B[8]), .S(i_data_immext[6]), .Q(n314) );
  IMUX20 U1168 ( .A(alu_i_data_B[11]), .B(u_alu_lt_x_11_B_10_), .S(
        i_data_immext[6]), .Q(n312) );
  IMUX20 U1169 ( .A(alu_i_data_B[19]), .B(alu_i_data_B[18]), .S(
        i_data_immext[6]), .Q(n351) );
  IMUX20 U1170 ( .A(alu_i_data_B[21]), .B(alu_i_data_B[20]), .S(
        i_data_immext[6]), .Q(n361) );
  IMUX20 U1171 ( .A(alu_i_data_B[23]), .B(alu_i_data_B[22]), .S(
        i_data_immext[6]), .Q(n373) );
  IMUX20 U1172 ( .A(alu_i_data_B[25]), .B(alu_i_data_B[24]), .S(
        i_data_immext[6]), .Q(n386) );
  IMUX20 U1173 ( .A(alu_i_data_B[31]), .B(alu_i_data_B[30]), .S(
        i_data_immext[6]), .Q(n412) );
  NAND22 U1174 ( .A(n1167), .B(u_alu_pre_sum_4b[7]), .Q(n1171) );
  INV3 U1175 ( .A(u_alu_N173), .Q(n1000) );
  NOR21 U1176 ( .A(u_alu_add_x_1_n36), .B(u_alu_add_x_1_n33), .Q(
        u_alu_add_x_1_n31) );
  NOR21 U1177 ( .A(alu_i_con_AluCtrl[0]), .B(n1234), .Q(n1161) );
  NOR21 U1178 ( .A(alu_i_con_AluCtrl[1]), .B(alu_i_con_AluCtrl[3]), .Q(n872)
         );
  NAND31 U1179 ( .A(n505), .B(n571), .C(n438), .Q(n524) );
  NOR21 U1180 ( .A(n440), .B(n469), .Q(n505) );
  NAND22 U1181 ( .A(alu_i_data_B[31]), .B(n572), .Q(n469) );
  INV3 U1182 ( .A(u_alu_ashr_4_SH_1_), .Q(n439) );
  NAND22 U1183 ( .A(u_alu_pre_subb[15]), .B(n1158), .Q(n1176) );
  NAND22 U1184 ( .A(n297), .B(i_data_rs[2]), .Q(n710) );
  NOR21 U1185 ( .A(n701), .B(n711), .Q(n705) );
  NAND22 U1186 ( .A(n296), .B(i_data_rs[4]), .Q(n700) );
  NAND22 U1187 ( .A(n139), .B(i_data_rt[4]), .Q(n854) );
  NOR21 U1188 ( .A(n687), .B(n711), .Q(n691) );
  NAND22 U1189 ( .A(n168), .B(i_data_rt[5]), .Q(n851) );
  NAND22 U1190 ( .A(n686), .B(n685), .Q(compare_i_data_rs[6]) );
  NOR21 U1191 ( .A(n680), .B(n711), .Q(n684) );
  NAND22 U1192 ( .A(n296), .B(i_data_rs[6]), .Q(n686) );
  NAND31 U1193 ( .A(n848), .B(n847), .C(n846), .Q(compare_i_data_rt[6]) );
  NAND22 U1194 ( .A(n168), .B(i_data_rt[6]), .Q(n848) );
  NOR21 U1195 ( .A(n673), .B(n711), .Q(n677) );
  NAND22 U1196 ( .A(n296), .B(i_data_rs[7]), .Q(n679) );
  NAND31 U1197 ( .A(n845), .B(n844), .C(n843), .Q(compare_i_data_rt[7]) );
  NAND22 U1198 ( .A(n139), .B(i_data_rt[7]), .Q(n845) );
  OAI212 U1199 ( .A(n140), .B(n1286), .C(n672), .Q(compare_i_data_rs[8]) );
  MUX22 U1200 ( .A(compare_i_data_rt[8]), .B(i_data_immext[8]), .S(n305), .Q(
        alu_i_data_B[8]) );
  OAI212 U1201 ( .A(n298), .B(n1286), .C(n841), .Q(compare_i_data_rt[8]) );
  AOI211 U1202 ( .A(n139), .B(i_data_rt[8]), .C(n840), .Q(n841) );
  OAI212 U1203 ( .A(n140), .B(n1287), .C(n669), .Q(compare_i_data_rs[9]) );
  MUX22 U1204 ( .A(compare_i_data_rt[9]), .B(u_alu_ashr_4_SH_3_), .S(n305), 
        .Q(alu_i_data_B[9]) );
  OAI212 U1205 ( .A(n298), .B(n1287), .C(n836), .Q(compare_i_data_rt[9]) );
  AOI211 U1206 ( .A(n139), .B(i_data_rt[9]), .C(n835), .Q(n836) );
  OAI212 U1207 ( .A(n140), .B(n1269), .C(n666), .Q(compare_i_data_rs[10]) );
  INV3 U1208 ( .A(n293), .Q(u_alu_lt_x_11_B_10_) );
  IMUX21 U1209 ( .A(compare_i_data_rt[10]), .B(i_data_immext[10]), .S(n305), 
        .Q(n293) );
  OAI212 U1210 ( .A(n298), .B(n1269), .C(n832), .Q(compare_i_data_rt[10]) );
  AOI211 U1211 ( .A(n168), .B(i_data_rt[10]), .C(n831), .Q(n832) );
  OAI212 U1212 ( .A(n140), .B(n1270), .C(n663), .Q(compare_i_data_rs[11]) );
  MUX22 U1213 ( .A(compare_i_data_rt[11]), .B(i_data_immext[11]), .S(n305), 
        .Q(alu_i_data_B[11]) );
  OAI212 U1214 ( .A(n298), .B(n1270), .C(n828), .Q(compare_i_data_rt[11]) );
  OAI212 U1215 ( .A(n140), .B(n1271), .C(n660), .Q(compare_i_data_rs[12]) );
  AOI211 U1216 ( .A(n720), .B(i_data_rs[12]), .C(n659), .Q(n660) );
  MUX22 U1217 ( .A(compare_i_data_rt[12]), .B(i_data_immext[12]), .S(n305), 
        .Q(alu_i_data_B[12]) );
  OAI212 U1218 ( .A(n140), .B(n1272), .C(n657), .Q(compare_i_data_rs[13]) );
  MUX22 U1219 ( .A(compare_i_data_rt[13]), .B(i_data_immext[13]), .S(n305), 
        .Q(alu_i_data_B[13]) );
  OAI212 U1220 ( .A(n140), .B(n1273), .C(n654), .Q(compare_i_data_rs[14]) );
  MUX22 U1221 ( .A(compare_i_data_rt[14]), .B(i_data_immext[14]), .S(n305), 
        .Q(alu_i_data_B[14]) );
  OAI212 U1222 ( .A(n140), .B(n1274), .C(n651), .Q(compare_i_data_rs[15]) );
  NOR31 U1223 ( .A(n919), .B(n923), .C(n918), .Q(n1254) );
  OAI212 U1224 ( .A(i_data_immext[0]), .B(n915), .C(n1177), .Q(n923) );
  NOR31 U1225 ( .A(n912), .B(n910), .C(n911), .Q(n924) );
  OAI212 U1226 ( .A(n1261), .B(n871), .C(n1260), .Q(alu_i_con_AluCtrl[1]) );
  AOI221 U1227 ( .A(n1255), .B(n1264), .C(i_con_Ealuop[0]), .D(i_con_Ealuop[5]), .Q(n1263) );
  AOI211 U1228 ( .A(i_data_immext[2]), .B(n912), .C(n911), .Q(n921) );
  NAND22 U1229 ( .A(n909), .B(i_data_immext[1]), .Q(n911) );
  NAND22 U1230 ( .A(i_data_immext[5]), .B(n1246), .Q(n1247) );
  NAND31 U1231 ( .A(n870), .B(n909), .C(n912), .Q(n913) );
  NAND22 U1232 ( .A(n910), .B(i_data_immext[5]), .Q(n868) );
  OAI212 U1233 ( .A(n140), .B(n1285), .C(n587), .Q(compare_i_data_rs[31]) );
  NAND22 U1234 ( .A(n737), .B(n807), .Q(alu_i_data_B[31]) );
  AOI211 U1235 ( .A(n168), .B(i_data_rt[31]), .C(n735), .Q(n736) );
  OAI212 U1236 ( .A(n140), .B(n1284), .C(n590), .Q(compare_i_data_rs[30]) );
  NAND22 U1237 ( .A(n742), .B(n807), .Q(alu_i_data_B[30]) );
  OAI212 U1238 ( .A(n298), .B(n1284), .C(n741), .Q(compare_i_data_rt[30]) );
  NAND22 U1239 ( .A(n747), .B(n807), .Q(alu_i_data_B[29]) );
  AOI211 U1240 ( .A(n139), .B(i_data_rt[29]), .C(n745), .Q(n746) );
  OAI212 U1241 ( .A(n140), .B(n1283), .C(n593), .Q(compare_i_data_rs[29]) );
  NAND22 U1242 ( .A(n791), .B(n807), .Q(alu_i_data_B[20]) );
  NAND31 U1243 ( .A(n790), .B(n789), .C(n788), .Q(compare_i_data_rt[20]) );
  NAND22 U1244 ( .A(n624), .B(n623), .Q(compare_i_data_rs[20]) );
  NAND22 U1245 ( .A(n296), .B(i_data_rs[16]), .Q(n648) );
  NAND22 U1246 ( .A(n645), .B(n644), .Q(compare_i_data_rs[17]) );
  NAND22 U1247 ( .A(n638), .B(n637), .Q(compare_i_data_rs[18]) );
  NAND22 U1248 ( .A(n296), .B(i_data_rs[18]), .Q(n638) );
  OAI212 U1249 ( .A(n305), .B(n798), .C(n807), .Q(alu_i_data_B[18]) );
  NAND22 U1250 ( .A(n168), .B(i_data_rt[18]), .Q(n797) );
  NAND22 U1251 ( .A(n631), .B(n630), .Q(compare_i_data_rs[19]) );
  OAI212 U1252 ( .A(n305), .B(n935), .C(n807), .Q(alu_i_data_B[19]) );
  NAND31 U1253 ( .A(n794), .B(n793), .C(n792), .Q(compare_i_data_rt[19]) );
  OAI212 U1254 ( .A(n140), .B(n1275), .C(n617), .Q(compare_i_data_rs[21]) );
  NAND22 U1255 ( .A(n787), .B(n807), .Q(alu_i_data_B[21]) );
  OAI212 U1256 ( .A(n298), .B(n1275), .C(n786), .Q(compare_i_data_rt[21]) );
  AOI211 U1257 ( .A(n168), .B(i_data_rt[21]), .C(n785), .Q(n786) );
  OAI212 U1258 ( .A(n140), .B(n1276), .C(n614), .Q(compare_i_data_rs[22]) );
  NAND22 U1259 ( .A(n782), .B(n807), .Q(alu_i_data_B[22]) );
  NAND22 U1260 ( .A(compare_i_data_rt[22]), .B(n806), .Q(n782) );
  OAI212 U1261 ( .A(n298), .B(n1276), .C(n781), .Q(compare_i_data_rt[22]) );
  AOI211 U1262 ( .A(n168), .B(i_data_rt[22]), .C(n780), .Q(n781) );
  OAI212 U1263 ( .A(n140), .B(n1277), .C(n611), .Q(compare_i_data_rs[23]) );
  AOI211 U1264 ( .A(n720), .B(i_data_rs[23]), .C(n610), .Q(n611) );
  NAND22 U1265 ( .A(n777), .B(n807), .Q(alu_i_data_B[23]) );
  NAND22 U1266 ( .A(compare_i_data_rt[23]), .B(n806), .Q(n777) );
  OAI212 U1267 ( .A(n298), .B(n1277), .C(n776), .Q(compare_i_data_rt[23]) );
  OAI212 U1268 ( .A(n140), .B(n1278), .C(n608), .Q(compare_i_data_rs[24]) );
  NAND22 U1269 ( .A(n772), .B(n807), .Q(alu_i_data_B[24]) );
  OAI212 U1270 ( .A(n298), .B(n1278), .C(n771), .Q(compare_i_data_rt[24]) );
  AOI211 U1271 ( .A(n168), .B(i_data_rt[24]), .C(n770), .Q(n771) );
  OAI212 U1272 ( .A(n140), .B(n1279), .C(n605), .Q(compare_i_data_rs[25]) );
  NAND22 U1273 ( .A(n767), .B(n807), .Q(alu_i_data_B[25]) );
  OAI212 U1274 ( .A(n298), .B(n1279), .C(n766), .Q(compare_i_data_rt[25]) );
  OAI212 U1275 ( .A(n140), .B(n1280), .C(n602), .Q(compare_i_data_rs[26]) );
  NAND22 U1276 ( .A(n762), .B(n807), .Q(alu_i_data_B[26]) );
  OAI212 U1277 ( .A(n298), .B(n1280), .C(n761), .Q(compare_i_data_rt[26]) );
  AOI211 U1278 ( .A(n168), .B(i_data_rt[26]), .C(n760), .Q(n761) );
  OAI212 U1279 ( .A(n140), .B(n1281), .C(n599), .Q(compare_i_data_rs[27]) );
  NAND22 U1280 ( .A(n757), .B(n807), .Q(alu_i_data_B[27]) );
  NAND22 U1281 ( .A(compare_i_data_rt[27]), .B(n806), .Q(n757) );
  OAI212 U1282 ( .A(n298), .B(n1281), .C(n756), .Q(compare_i_data_rt[27]) );
  OAI212 U1283 ( .A(n140), .B(n1282), .C(n596), .Q(compare_i_data_rs[28]) );
  NOR21 U1284 ( .A(i_con_Efamux[1]), .B(n581), .Q(n582) );
  NAND22 U1285 ( .A(n752), .B(n807), .Q(alu_i_data_B[28]) );
  NOR21 U1286 ( .A(i_con_Efbmux[1]), .B(n729), .Q(n730) );
  NAND22 U1287 ( .A(i_con_Efbmux[0]), .B(i_con_Efbmux[2]), .Q(n726) );
  INV3 U1288 ( .A(i_con_Efbmux[1]), .Q(n728) );
  IMUX20 U1289 ( .A(n554), .B(n553), .S(n437), .Q(u_alu_N232) );
  IMUX20 U1290 ( .A(n515), .B(n514), .S(n440), .Q(n518) );
  IMUX20 U1291 ( .A(n538), .B(n537), .S(n437), .Q(u_alu_N229) );
  IMUX20 U1292 ( .A(n549), .B(n548), .S(n437), .Q(u_alu_N231) );
  IMUX20 U1293 ( .A(n490), .B(n526), .S(n440), .Q(n491) );
  MUX21 U1294 ( .A(n544), .B(n543), .S(n437), .Q(u_alu_N230) );
  MUX21 U1295 ( .A(n365), .B(n423), .S(n437), .Q(u_alu_N216) );
  MUX21 U1296 ( .A(n379), .B(n425), .S(n437), .Q(u_alu_N218) );
  IMUX20 U1297 ( .A(n467), .B(n470), .S(n440), .Q(n478) );
  MUX21 U1298 ( .A(n391), .B(n390), .S(n437), .Q(u_alu_N220) );
  MUX21 U1299 ( .A(n405), .B(n404), .S(n437), .Q(u_alu_N222) );
  MUX21 U1300 ( .A(n331), .B(n330), .S(n437), .Q(u_alu_N209) );
  MUX21 U1301 ( .A(n372), .B(n424), .S(n437), .Q(u_alu_N217) );
  MUX21 U1302 ( .A(n398), .B(n397), .S(n437), .Q(u_alu_N221) );
  MUX21 U1303 ( .A(n385), .B(n384), .S(n437), .Q(u_alu_N219) );
  IMUX20 U1304 ( .A(n454), .B(n453), .S(n440), .Q(n473) );
  IMUX20 U1305 ( .A(n451), .B(n454), .S(n440), .Q(n459) );
  IMUX20 U1306 ( .A(n310), .B(n309), .S(n440), .Q(n328) );
  IMUX20 U1307 ( .A(n308), .B(n307), .S(n440), .Q(n329) );
  IMUX20 U1308 ( .A(n307), .B(n310), .S(n440), .Q(n321) );
  IMUX20 U1309 ( .A(n306), .B(n308), .S(n440), .Q(n319) );
  IMUX20 U1310 ( .A(n468), .B(n467), .S(n440), .Q(n485) );
  IMUX20 U1311 ( .A(n316), .B(n315), .S(n440), .Q(n334) );
  IMUX20 U1312 ( .A(n314), .B(n313), .S(n440), .Q(n335) );
  NOR40 U1313 ( .A(n1183), .B(n874), .C(alu_i_con_AluCtrl[3]), .D(
        alu_i_con_AluCtrl[2]), .Q(n1181) );
  MUX21 U1314 ( .A(n418), .B(n417), .S(n437), .Q(u_alu_N224) );
  IMUX20 U1315 ( .A(n313), .B(n316), .S(n440), .Q(n325) );
  IMUX20 U1316 ( .A(n312), .B(n314), .S(n440), .Q(n323) );
  IMUX20 U1317 ( .A(n412), .B(n411), .S(n440), .Q(n414) );
  NAND22 U1318 ( .A(n875), .B(n873), .Q(n1078) );
  INV3 U1319 ( .A(alu_i_con_AluCtrl[2]), .Q(n873) );
  NAND22 U1320 ( .A(alu_i_con_AluCtrl[2]), .B(n1183), .Q(n881) );
  INV3 U1321 ( .A(i_data_immext[5]), .Q(n912) );
  INV3 U1322 ( .A(i_data_immext[3]), .Q(n909) );
  INV3 U1323 ( .A(i_data_immext[2]), .Q(n910) );
  INV3 U1324 ( .A(n1264), .Q(n1261) );
  NAND22 U1325 ( .A(i_con_Efamux[2]), .B(i_con_Efamux[0]), .Q(n578) );
  INV0 U1326 ( .A(u_alu_add_x_1_n14), .Q(u_alu_add_x_1_n44) );
  NAND20 U1327 ( .A(u_alu_N227), .B(n1180), .Q(n898) );
  INV0 U1328 ( .A(u_alu_add_x_1_n36), .Q(u_alu_add_x_1_n49) );
  NAND20 U1329 ( .A(u_alu_N228), .B(n1180), .Q(n895) );
  INV0 U1330 ( .A(u_alu_add_x_1_n33), .Q(u_alu_add_x_1_n48) );
  INV0 U1331 ( .A(u_alu_add_x_1_n17), .Q(u_alu_add_x_1_n45) );
  INV0 U1332 ( .A(u_alu_add_x_1_n40), .Q(u_alu_add_x_1_n50) );
  INV0 U1333 ( .A(u_alu_add_x_1_n27), .Q(u_alu_add_x_1_n47) );
  INV0 U1334 ( .A(u_alu_add_x_1_n22), .Q(u_alu_add_x_1_n46) );
  NOR30 U1335 ( .A(alu_i_data_B[15]), .B(compare_i_data_rs[15]), .C(n1144), 
        .Q(n994) );
  OAI210 U1336 ( .A(alu_i_data_B[15]), .B(n303), .C(n576), .Q(n995) );
  AOI2110 U1337 ( .A(n577), .B(compare_i_data_rs[15]), .C(n993), .D(n141), .Q(
        n997) );
  NOR20 U1338 ( .A(compare_i_data_rs[15]), .B(n303), .Q(n993) );
  NOR30 U1339 ( .A(alu_i_data_B[14]), .B(compare_i_data_rs[14]), .C(n1144), 
        .Q(n991) );
  OAI210 U1340 ( .A(alu_i_data_B[14]), .B(n303), .C(n576), .Q(n992) );
  NOR20 U1341 ( .A(compare_i_data_rs[14]), .B(n303), .Q(n990) );
  NOR30 U1342 ( .A(alu_i_data_B[9]), .B(compare_i_data_rs[9]), .C(n1144), .Q(
        n971) );
  OAI210 U1343 ( .A(alu_i_data_B[9]), .B(n303), .C(n576), .Q(n972) );
  AOI2110 U1344 ( .A(n577), .B(compare_i_data_rs[9]), .C(n970), .D(n141), .Q(
        n975) );
  NOR20 U1345 ( .A(compare_i_data_rs[9]), .B(n303), .Q(n970) );
  NAND20 U1346 ( .A(u_alu_N235), .B(n1180), .Q(n983) );
  NOR30 U1347 ( .A(u_alu_lt_x_11_B_10_), .B(compare_i_data_rs[10]), .C(n1144), 
        .Q(n981) );
  OAI210 U1348 ( .A(u_alu_lt_x_11_B_10_), .B(n303), .C(n576), .Q(n982) );
  AOI2110 U1349 ( .A(n577), .B(compare_i_data_rs[10]), .C(n980), .D(n141), .Q(
        n985) );
  NOR20 U1350 ( .A(compare_i_data_rs[10]), .B(n303), .Q(n980) );
  AOI220 U1351 ( .A(n998), .B(u_alu_N165), .C(n141), .D(alu_i_data_B[8]), .Q(
        n879) );
  INV3 U1352 ( .A(n1078), .Q(n998) );
  OAI310 U1353 ( .A(alu_i_data_B[23]), .B(compare_i_data_rs[23]), .C(n1144), 
        .D(n1065), .Q(n1066) );
  NAND20 U1354 ( .A(n1179), .B(n1064), .Q(n1065) );
  XNR21 U1355 ( .A(n159), .B(alu_i_data_B[23]), .Q(n1064) );
  OAI310 U1356 ( .A(n148), .B(n1225), .C(n1184), .D(n1063), .Q(n1067) );
  NAND20 U1357 ( .A(n1161), .B(u_alu_lt_x_11_B_7_), .Q(n1063) );
  OAI310 U1358 ( .A(alu_i_data_B[21]), .B(compare_i_data_rs[21]), .C(n1144), 
        .D(n1045), .Q(n1046) );
  NAND20 U1359 ( .A(n1179), .B(n1044), .Q(n1045) );
  XNR21 U1360 ( .A(n1043), .B(alu_i_data_B[21]), .Q(n1044) );
  OAI310 U1361 ( .A(n127), .B(n1227), .C(n1184), .D(n1042), .Q(n1047) );
  NAND20 U1362 ( .A(n1161), .B(n294), .Q(n1042) );
  AOI2110 U1363 ( .A(n141), .B(compare_i_data_rs[25]), .C(n1098), .D(n1097), 
        .Q(n1102) );
  OAI310 U1364 ( .A(alu_i_data_B[25]), .B(compare_i_data_rs[25]), .C(n1144), 
        .D(n1096), .Q(n1097) );
  NAND20 U1365 ( .A(n1179), .B(n1095), .Q(n1096) );
  XNR21 U1366 ( .A(n166), .B(alu_i_data_B[25]), .Q(n1095) );
  OAI310 U1367 ( .A(n142), .B(n1224), .C(n1184), .D(n1094), .Q(n1098) );
  NAND20 U1368 ( .A(n1161), .B(alu_i_data_B[9]), .Q(n1094) );
  AOI2110 U1369 ( .A(n141), .B(compare_i_data_rs[27]), .C(n1126), .D(n1125), 
        .Q(n1130) );
  OAI310 U1370 ( .A(alu_i_data_B[27]), .B(compare_i_data_rs[27]), .C(n1144), 
        .D(n1124), .Q(n1125) );
  NAND20 U1371 ( .A(n1179), .B(n1123), .Q(n1124) );
  XNR21 U1372 ( .A(n1122), .B(alu_i_data_B[27]), .Q(n1123) );
  OAI310 U1373 ( .A(n128), .B(n1222), .C(n1184), .D(n1121), .Q(n1126) );
  NAND20 U1374 ( .A(n1161), .B(alu_i_data_B[11]), .Q(n1121) );
  XNR21 U1375 ( .A(compare_i_data_rs[1]), .B(compare_i_data_rt[1]), .Q(n953)
         );
  XNR21 U1376 ( .A(compare_i_data_rs[18]), .B(compare_i_data_rt[18]), .Q(n954)
         );
  XNR21 U1377 ( .A(compare_i_data_rs[20]), .B(compare_i_data_rt[20]), .Q(n956)
         );
  XNR21 U1378 ( .A(compare_i_data_rs[3]), .B(compare_i_data_rt[3]), .Q(n949)
         );
  XNR21 U1379 ( .A(compare_i_data_rs[7]), .B(compare_i_data_rt[7]), .Q(n950)
         );
  XNR21 U1380 ( .A(compare_i_data_rs[6]), .B(compare_i_data_rt[6]), .Q(n951)
         );
  XNR21 U1381 ( .A(compare_i_data_rs[4]), .B(compare_i_data_rt[4]), .Q(n952)
         );
  XNR21 U1382 ( .A(compare_i_data_rt[30]), .B(compare_i_data_rs[30]), .Q(n947)
         );
  XNR21 U1383 ( .A(compare_i_data_rs[5]), .B(compare_i_data_rt[5]), .Q(n945)
         );
  XNR21 U1384 ( .A(n1122), .B(compare_i_data_rt[27]), .Q(n1294) );
  XNR21 U1385 ( .A(n1108), .B(compare_i_data_rt[26]), .Q(n1295) );
  XNR21 U1386 ( .A(n166), .B(compare_i_data_rt[25]), .Q(n1296) );
  XNR21 U1387 ( .A(n161), .B(compare_i_data_rt[24]), .Q(n1297) );
  XNR21 U1388 ( .A(compare_i_data_rt[31]), .B(compare_i_data_rs[31]), .Q(n946)
         );
  XNR21 U1389 ( .A(n157), .B(compare_i_data_rt[28]), .Q(n941) );
  XNR21 U1390 ( .A(n159), .B(compare_i_data_rt[23]), .Q(n942) );
  XNR21 U1391 ( .A(n1043), .B(compare_i_data_rt[21]), .Q(n943) );
  XNR21 U1392 ( .A(n163), .B(compare_i_data_rt[22]), .Q(n944) );
  XNR21 U1393 ( .A(n167), .B(compare_i_data_rt[9]), .Q(n937) );
  XNR21 U1394 ( .A(n151), .B(compare_i_data_rt[8]), .Q(n938) );
  XNR21 U1395 ( .A(n936), .B(compare_i_data_rt[2]), .Q(n939) );
  XNR21 U1396 ( .A(n935), .B(compare_i_data_rs[19]), .Q(n940) );
  XNR21 U1397 ( .A(n155), .B(compare_i_data_rt[11]), .Q(n931) );
  XNR21 U1398 ( .A(n930), .B(compare_i_data_rt[12]), .Q(n932) );
  XNR21 U1399 ( .A(n152), .B(compare_i_data_rt[0]), .Q(n933) );
  XNR21 U1400 ( .A(n149), .B(compare_i_data_rt[10]), .Q(n934) );
  XNR21 U1401 ( .A(n925), .B(compare_i_data_rt[15]), .Q(n926) );
  XNR21 U1402 ( .A(n154), .B(compare_i_data_rt[13]), .Q(n927) );
  XNR21 U1403 ( .A(n138), .B(compare_i_data_rt[16]), .Q(n928) );
  XNR21 U1404 ( .A(n164), .B(compare_i_data_rt[14]), .Q(n929) );
  NAND20 U1405 ( .A(u_alu_N241), .B(n1180), .Q(n1007) );
  OAI210 U1406 ( .A(n141), .B(n1003), .C(alu_i_data_B[16]), .Q(n1004) );
  IMUX20 U1407 ( .A(n1002), .B(n1001), .S(compare_i_data_rs[16]), .Q(n1005) );
  OAI210 U1408 ( .A(n303), .B(alu_i_data_B[16]), .C(n576), .Q(n1001) );
  NOR20 U1409 ( .A(alu_i_data_B[16]), .B(n1144), .Q(n1002) );
  AOI210 U1410 ( .A(n1083), .B(compare_i_data_rs[24]), .C(n1082), .Q(n1084) );
  OAI310 U1411 ( .A(alu_i_data_B[24]), .B(compare_i_data_rs[24]), .C(n1144), 
        .D(n1081), .Q(n1082) );
  NAND20 U1412 ( .A(n1161), .B(alu_i_data_B[8]), .Q(n1081) );
  OAI210 U1413 ( .A(n303), .B(alu_i_data_B[24]), .C(n576), .Q(n1083) );
  AOI2110 U1414 ( .A(n577), .B(compare_i_data_rs[24]), .C(n1080), .D(n141), 
        .Q(n1086) );
  NOR20 U1415 ( .A(compare_i_data_rs[24]), .B(n303), .Q(n1080) );
  OAI310 U1416 ( .A(alu_i_data_B[22]), .B(compare_i_data_rs[22]), .C(n1144), 
        .D(n1055), .Q(n1056) );
  NAND20 U1417 ( .A(n1179), .B(n1054), .Q(n1055) );
  XNR21 U1418 ( .A(n163), .B(alu_i_data_B[22]), .Q(n1054) );
  OAI310 U1419 ( .A(n146), .B(n1226), .C(n1184), .D(n1053), .Q(n1057) );
  NAND20 U1420 ( .A(n1161), .B(alu_i_data_B[6]), .Q(n1053) );
  OAI310 U1421 ( .A(alu_i_data_B[28]), .B(compare_i_data_rs[28]), .C(n1144), 
        .D(n1137), .Q(n1138) );
  NAND20 U1422 ( .A(n1179), .B(n1136), .Q(n1137) );
  XNR21 U1423 ( .A(n157), .B(alu_i_data_B[28]), .Q(n1136) );
  OAI310 U1424 ( .A(n143), .B(n1221), .C(n1184), .D(n1135), .Q(n1139) );
  NAND20 U1425 ( .A(n1161), .B(alu_i_data_B[12]), .Q(n1135) );
  AOI2110 U1426 ( .A(n141), .B(compare_i_data_rs[26]), .C(n1112), .D(n1111), 
        .Q(n1116) );
  OAI310 U1427 ( .A(alu_i_data_B[26]), .B(compare_i_data_rs[26]), .C(n1144), 
        .D(n1110), .Q(n1111) );
  NAND20 U1428 ( .A(n1179), .B(n1109), .Q(n1110) );
  XNR21 U1429 ( .A(n1108), .B(alu_i_data_B[26]), .Q(n1109) );
  OAI310 U1430 ( .A(n132), .B(n1223), .C(n1184), .D(n1107), .Q(n1112) );
  NAND20 U1431 ( .A(n1161), .B(u_alu_lt_x_11_B_10_), .Q(n1107) );
  NAND20 U1432 ( .A(u_alu_N245), .B(n1180), .Q(n1035) );
  AOI2110 U1433 ( .A(n141), .B(compare_i_data_rs[20]), .C(n1033), .D(n1032), 
        .Q(n1037) );
  OAI310 U1434 ( .A(alu_i_data_B[20]), .B(compare_i_data_rs[20]), .C(n1144), 
        .D(n1031), .Q(n1032) );
  NAND20 U1435 ( .A(n1179), .B(n1030), .Q(n1031) );
  XNR21 U1436 ( .A(n165), .B(alu_i_data_B[20]), .Q(n1030) );
  OAI310 U1437 ( .A(n145), .B(n1228), .C(n1184), .D(n1029), .Q(n1033) );
  NAND20 U1438 ( .A(n1161), .B(alu_i_data_B[4]), .Q(n1029) );
  OAI2110 U1439 ( .A(n158), .B(n576), .C(n1165), .D(n1164), .Q(n1166) );
  AOI220 U1440 ( .A(n1179), .B(n1163), .C(n1178), .D(n1162), .Q(n1164) );
  NOR20 U1441 ( .A(compare_i_data_rs[31]), .B(alu_i_data_B[31]), .Q(n1162) );
  XNR21 U1442 ( .A(n158), .B(alu_i_data_B[31]), .Q(n1163) );
  AOI210 U1443 ( .A(alu_i_data_B[15]), .B(n1161), .C(n1160), .Q(n1165) );
  NOR30 U1444 ( .A(n1159), .B(n1215), .C(n1184), .Q(n1160) );
  INV3 U1445 ( .A(alu_i_con_AluCtrl[0]), .Q(n874) );
  AOI220 U1446 ( .A(n301), .B(i_data_FMmemout[8]), .C(n302), .D(
        i_data_FMalures[8]), .Q(n837) );
  AOI220 U1447 ( .A(n301), .B(i_data_FMmemout[9]), .C(n302), .D(
        i_data_FMalures[9]), .Q(n833) );
  AOI220 U1448 ( .A(n301), .B(i_data_FMmemout[10]), .C(n302), .D(
        i_data_FMalures[10]), .Q(n829) );
  AOI220 U1449 ( .A(n301), .B(i_data_FMmemout[11]), .C(n302), .D(
        i_data_FMalures[11]), .Q(n825) );
  AOI220 U1450 ( .A(n301), .B(i_data_FMmemout[12]), .C(n302), .D(
        i_data_FMalures[12]), .Q(n821) );
  AOI220 U1451 ( .A(n169), .B(i_data_FMmemout[13]), .C(n721), .D(
        i_data_FMalures[13]), .Q(n655) );
  AOI220 U1452 ( .A(n301), .B(i_data_FMmemout[13]), .C(n302), .D(
        i_data_FMalures[13]), .Q(n817) );
  AOI220 U1453 ( .A(n169), .B(i_data_FMmemout[14]), .C(n721), .D(
        i_data_FMalures[14]), .Q(n652) );
  AOI220 U1454 ( .A(n301), .B(i_data_FMmemout[14]), .C(n302), .D(
        i_data_FMalures[14]), .Q(n813) );
  AOI220 U1455 ( .A(n169), .B(i_data_FMmemout[15]), .C(n721), .D(
        i_data_FMalures[15]), .Q(n649) );
  AOI220 U1456 ( .A(n301), .B(i_data_FMmemout[15]), .C(n302), .D(
        i_data_FMalures[15]), .Q(n809) );
  INV3 U1457 ( .A(alu_i_con_AluCtrl[1]), .Q(n1183) );
  AOI220 U1458 ( .A(n301), .B(i_data_FMmemout[31]), .C(n302), .D(
        i_data_FMalures[31]), .Q(n733) );
  AOI220 U1459 ( .A(n169), .B(i_data_FMmemout[30]), .C(n721), .D(
        i_data_FMalures[30]), .Q(n588) );
  AOI220 U1460 ( .A(n301), .B(i_data_FMmemout[30]), .C(n302), .D(
        i_data_FMalures[30]), .Q(n738) );
  AOI220 U1461 ( .A(n301), .B(i_data_FMmemout[29]), .C(n302), .D(
        i_data_FMalures[29]), .Q(n743) );
  AOI220 U1462 ( .A(n169), .B(i_data_FMmemout[29]), .C(n721), .D(
        i_data_FMalures[29]), .Q(n591) );
  AOI220 U1463 ( .A(n301), .B(i_data_FMmemout[20]), .C(n863), .D(
        i_data_FWmemout[20]), .Q(n788) );
  NAND20 U1464 ( .A(n169), .B(i_data_FMmemout[20]), .Q(n619) );
  AOI220 U1465 ( .A(n721), .B(i_data_FMalures[16]), .C(n573), .D(
        i_data_FEalures[16]), .Q(n647) );
  NAND20 U1466 ( .A(n169), .B(i_data_FMmemout[17]), .Q(n640) );
  NAND20 U1467 ( .A(n169), .B(i_data_FMmemout[18]), .Q(n633) );
  NAND20 U1468 ( .A(n169), .B(i_data_FMmemout[19]), .Q(n626) );
  AOI220 U1469 ( .A(n169), .B(i_data_FMmemout[21]), .C(n721), .D(
        i_data_FMalures[21]), .Q(n615) );
  AOI220 U1470 ( .A(n301), .B(i_data_FMmemout[21]), .C(n302), .D(
        i_data_FMalures[21]), .Q(n783) );
  AOI220 U1471 ( .A(n169), .B(i_data_FMmemout[22]), .C(n721), .D(
        i_data_FMalures[22]), .Q(n612) );
  AOI220 U1472 ( .A(n301), .B(i_data_FMmemout[22]), .C(n302), .D(
        i_data_FMalures[22]), .Q(n778) );
  AOI220 U1473 ( .A(n169), .B(i_data_FMmemout[23]), .C(n721), .D(
        i_data_FMalures[23]), .Q(n609) );
  AOI220 U1474 ( .A(n301), .B(i_data_FMmemout[23]), .C(n302), .D(
        i_data_FMalures[23]), .Q(n773) );
  AOI220 U1475 ( .A(n169), .B(i_data_FMmemout[24]), .C(n721), .D(
        i_data_FMalures[24]), .Q(n606) );
  AOI220 U1476 ( .A(n301), .B(i_data_FMmemout[24]), .C(n302), .D(
        i_data_FMalures[24]), .Q(n768) );
  AOI220 U1477 ( .A(n169), .B(i_data_FMmemout[25]), .C(n721), .D(
        i_data_FMalures[25]), .Q(n603) );
  AOI220 U1478 ( .A(n301), .B(i_data_FMmemout[25]), .C(n302), .D(
        i_data_FMalures[25]), .Q(n763) );
  AOI220 U1479 ( .A(n169), .B(i_data_FMmemout[26]), .C(n721), .D(
        i_data_FMalures[26]), .Q(n600) );
  AOI220 U1480 ( .A(n301), .B(i_data_FMmemout[26]), .C(n302), .D(
        i_data_FMalures[26]), .Q(n758) );
  AOI220 U1481 ( .A(n169), .B(i_data_FMmemout[27]), .C(n721), .D(
        i_data_FMalures[27]), .Q(n597) );
  AOI220 U1482 ( .A(n301), .B(i_data_FMmemout[27]), .C(n302), .D(
        i_data_FMalures[27]), .Q(n753) );
  AOI220 U1483 ( .A(n169), .B(i_data_FMmemout[28]), .C(n721), .D(
        i_data_FMalures[28]), .Q(n594) );
  INV3 U1484 ( .A(n578), .Q(n579) );
  AOI220 U1485 ( .A(n301), .B(i_data_FMmemout[28]), .C(n302), .D(
        i_data_FMalures[28]), .Q(n748) );
  INV3 U1486 ( .A(n726), .Q(n727) );
  NAND22 U1487 ( .A(n872), .B(n873), .Q(n1184) );
  INV3 U1488 ( .A(n1184), .Q(n577) );
  OAI210 U1489 ( .A(u_alu_add_x_1_n36), .B(u_alu_add_x_1_n38), .C(
        u_alu_add_x_1_n37), .Q(u_alu_add_x_1_n35) );
  AOI220 U1490 ( .A(n302), .B(i_data_FMalures[20]), .C(n300), .D(
        i_data_FEalures[20]), .Q(n789) );
  AOI220 U1491 ( .A(n302), .B(i_data_FMalures[19]), .C(n300), .D(
        i_data_FEalures[19]), .Q(n793) );
  AOI220 U1492 ( .A(n302), .B(i_data_FMalures[6]), .C(n300), .D(
        i_data_FEalures[6]), .Q(n847) );
  AOI220 U1493 ( .A(n302), .B(i_data_FMalures[18]), .C(n300), .D(
        i_data_FEalures[18]), .Q(n796) );
  XNR21 U1494 ( .A(compare_i_data_rs[17]), .B(compare_i_data_rt[17]), .Q(n955)
         );
  NOR40 U1495 ( .A(u_alu_ashr_4_SH_3_), .B(i_data_immext[8]), .C(
        u_alu_ashr_4_SH_1_), .D(n311), .Q(n330) );
  IMUX20 U1496 ( .A(n368), .B(n371), .S(u_alu_ashr_4_SH_3_), .Q(n331) );
  IMUX20 U1497 ( .A(alu_i_data_B[17]), .B(alu_i_data_B[16]), .S(
        i_data_immext[6]), .Q(n341) );
  IMUX20 U1498 ( .A(alu_i_data_B[18]), .B(alu_i_data_B[17]), .S(
        i_data_immext[6]), .Q(n346) );
  NOR20 U1499 ( .A(i_data_immext[10]), .B(n427), .Q(u_alu_N194) );
  IMUX20 U1500 ( .A(n395), .B(n348), .S(u_alu_ashr_4_SH_3_), .Q(n350) );
  IMUX20 U1501 ( .A(n402), .B(n353), .S(u_alu_ashr_4_SH_3_), .Q(n355) );
  IMUX20 U1502 ( .A(n409), .B(n358), .S(u_alu_ashr_4_SH_3_), .Q(n360) );
  IMUX20 U1503 ( .A(n415), .B(n363), .S(u_alu_ashr_4_SH_3_), .Q(n365) );
  IMUX20 U1504 ( .A(n393), .B(n367), .S(i_data_immext[8]), .Q(n369) );
  IMUX20 U1505 ( .A(n369), .B(n368), .S(u_alu_ashr_4_SH_3_), .Q(n372) );
  NAND40 U1506 ( .A(alu_i_data_B[0]), .B(n438), .C(n439), .D(n572), .Q(n370)
         );
  IMUX20 U1507 ( .A(n400), .B(n374), .S(i_data_immext[8]), .Q(n376) );
  IMUX20 U1508 ( .A(n376), .B(n375), .S(u_alu_ashr_4_SH_3_), .Q(n379) );
  IMUX20 U1509 ( .A(n408), .B(n381), .S(i_data_immext[8]), .Q(n383) );
  IMUX20 U1510 ( .A(n383), .B(n382), .S(u_alu_ashr_4_SH_3_), .Q(n385) );
  IMUX20 U1511 ( .A(n413), .B(n387), .S(i_data_immext[8]), .Q(n389) );
  IMUX20 U1512 ( .A(n389), .B(n388), .S(u_alu_ashr_4_SH_3_), .Q(n391) );
  IMUX20 U1513 ( .A(n394), .B(n393), .S(i_data_immext[8]), .Q(n396) );
  IMUX20 U1514 ( .A(n396), .B(n395), .S(u_alu_ashr_4_SH_3_), .Q(n398) );
  IMUX20 U1515 ( .A(n401), .B(n400), .S(i_data_immext[8]), .Q(n403) );
  IMUX20 U1516 ( .A(n403), .B(n402), .S(u_alu_ashr_4_SH_3_), .Q(n405) );
  NOR20 U1517 ( .A(i_data_immext[10]), .B(n428), .Q(u_alu_N195) );
  IMUX20 U1518 ( .A(n414), .B(n413), .S(i_data_immext[8]), .Q(n416) );
  IMUX20 U1519 ( .A(n416), .B(n415), .S(u_alu_ashr_4_SH_3_), .Q(n418) );
  NOR20 U1520 ( .A(i_data_immext[10]), .B(n429), .Q(u_alu_N196) );
  NOR20 U1521 ( .A(i_data_immext[10]), .B(n430), .Q(u_alu_N197) );
  NOR20 U1522 ( .A(i_data_immext[10]), .B(n431), .Q(u_alu_N198) );
  NOR20 U1523 ( .A(i_data_immext[10]), .B(n432), .Q(u_alu_N199) );
  NOR20 U1524 ( .A(i_data_immext[10]), .B(n433), .Q(u_alu_N200) );
  IMUX20 U1525 ( .A(n442), .B(n536), .S(i_data_immext[8]), .Q(n443) );
  IMUX20 U1526 ( .A(alu_i_data_B[16]), .B(alu_i_data_B[17]), .S(
        i_data_immext[6]), .Q(n447) );
  IMUX20 U1527 ( .A(n519), .B(n487), .S(u_alu_ashr_4_SH_3_), .Q(n456) );
  IMUX20 U1528 ( .A(alu_i_data_B[17]), .B(alu_i_data_B[18]), .S(
        i_data_immext[6]), .Q(n464) );
  MUX21 U1529 ( .A(n458), .B(n457), .S(i_data_immext[8]), .Q(n534) );
  MUX21 U1530 ( .A(n472), .B(n471), .S(i_data_immext[8]), .Q(n545) );
  IMUX20 U1531 ( .A(n545), .B(n504), .S(u_alu_ashr_4_SH_3_), .Q(n475) );
  MUX21 U1532 ( .A(n477), .B(n476), .S(i_data_immext[8]), .Q(n550) );
  IMUX20 U1533 ( .A(n550), .B(n507), .S(u_alu_ashr_4_SH_3_), .Q(n480) );
  NOR20 U1534 ( .A(i_data_immext[10]), .B(n566), .Q(u_alu_N241) );
  IMUX20 U1535 ( .A(n491), .B(n540), .S(i_data_immext[8]), .Q(n494) );
  IMUX20 U1536 ( .A(n494), .B(n560), .S(u_alu_ashr_4_SH_3_), .Q(n496) );
  NOR20 U1537 ( .A(i_data_immext[10]), .B(n537), .Q(u_alu_N245) );
  IMUX20 U1538 ( .A(n518), .B(n547), .S(i_data_immext[8]), .Q(n520) );
  IMUX20 U1539 ( .A(n520), .B(n519), .S(u_alu_ashr_4_SH_3_), .Q(n522) );
  NOR20 U1540 ( .A(i_data_immext[10]), .B(n524), .Q(u_alu_N256) );
  IMUX20 U1541 ( .A(n529), .B(n552), .S(i_data_immext[8]), .Q(n531) );
  IMUX20 U1542 ( .A(n531), .B(n530), .S(u_alu_ashr_4_SH_3_), .Q(n533) );
  IMUX30 U1543 ( .A(n536), .B(n535), .C(n534), .S0(i_data_immext[8]), .S1(
        u_alu_ashr_4_SH_3_), .Q(n538) );
  IMUX20 U1544 ( .A(n540), .B(n539), .S(i_data_immext[8]), .Q(n542) );
  IMUX20 U1545 ( .A(n542), .B(n541), .S(u_alu_ashr_4_SH_3_), .Q(n544) );
  IMUX30 U1546 ( .A(n547), .B(n546), .C(n545), .S0(i_data_immext[8]), .S1(
        u_alu_ashr_4_SH_3_), .Q(n549) );
  IMUX30 U1547 ( .A(n552), .B(n551), .C(n550), .S0(i_data_immext[8]), .S1(
        u_alu_ashr_4_SH_3_), .Q(n554) );
  IMUX20 U1548 ( .A(n556), .B(n555), .S(u_alu_ashr_4_SH_3_), .Q(n558) );
  OAI212 U1549 ( .A(n298), .B(n1274), .C(n812), .Q(compare_i_data_rt[15]) );
  OAI212 U1550 ( .A(n298), .B(n1273), .C(n816), .Q(compare_i_data_rt[14]) );
  OAI212 U1551 ( .A(n298), .B(n1272), .C(n820), .Q(compare_i_data_rt[13]) );
  OAI212 U1552 ( .A(n298), .B(n1271), .C(n824), .Q(compare_i_data_rt[12]) );
  OAI212 U1553 ( .A(n158), .B(n969), .C(n968), .Q(o_con_ifbranch) );
  OAI220 U1554 ( .A(n1184), .B(n1189), .C(alu_i_data_B[8]), .D(n303), .Q(n1187) );
  NOR20 U1555 ( .A(alu_i_con_AluCtrl[0]), .B(alu_i_data_B[8]), .Q(n1189) );
  IMUX20 U1556 ( .A(n303), .B(n1184), .S(u_alu_lt_x_11_B_7_), .Q(n1193) );
  IMUX20 U1557 ( .A(n1178), .B(n1179), .S(u_alu_lt_x_11_B_7_), .Q(n1190) );
  NOR20 U1558 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[31]), .Q(n1215)
         );
  NOR20 U1559 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[28]), .Q(n1221)
         );
  NOR20 U1560 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[27]), .Q(n1222)
         );
  NOR20 U1561 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[26]), .Q(n1223)
         );
  NOR20 U1562 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[25]), .Q(n1224)
         );
  NOR20 U1563 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[23]), .Q(n1225)
         );
  NOR20 U1564 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[22]), .Q(n1226)
         );
  NOR20 U1565 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[21]), .Q(n1227)
         );
  NOR20 U1566 ( .A(alu_i_con_AluCtrl[0]), .B(compare_i_data_rs[20]), .Q(n1228)
         );
  IMUX20 U1567 ( .A(n303), .B(n1184), .S(u_alu_lt_x_11_B_1_), .Q(n1232) );
  NAND20 U1568 ( .A(alu_i_con_AluCtrl[2]), .B(n1244), .Q(n1243) );
  NOR20 U1569 ( .A(alu_i_con_AluCtrl[3]), .B(n1183), .Q(n1244) );
  IMAJ30 U1570 ( .A(compare_i_data_rs[31]), .B(u_alu_N306), .C(n1159), .Q(
        n1241) );
  NOR20 U1571 ( .A(alu_i_con_AluCtrl[1]), .B(alu_i_con_AluCtrl[2]), .Q(n1245)
         );
  NOR30 U1572 ( .A(i_con_Ealuop[2]), .B(i_con_Ealuop[3]), .C(n1267), .Q(n1258)
         );
  NOR40 U1573 ( .A(n1259), .B(n1258), .C(n1257), .D(n1256), .Q(n1260) );
  IMUX20 U1574 ( .A(i_addr_rt[0]), .B(i_data_immext[11]), .S(i_con_Eregdst), 
        .Q(n1288) );
  IMUX20 U1575 ( .A(i_addr_rt[1]), .B(i_data_immext[12]), .S(i_con_Eregdst), 
        .Q(n1289) );
  IMUX20 U1576 ( .A(i_addr_rt[2]), .B(i_data_immext[13]), .S(i_con_Eregdst), 
        .Q(n1290) );
  IMUX20 U1577 ( .A(i_addr_rt[3]), .B(i_data_immext[14]), .S(i_con_Eregdst), 
        .Q(n1291) );
  IMUX20 U1578 ( .A(i_addr_rt[4]), .B(i_data_immext[15]), .S(i_con_Eregdst), 
        .Q(n1292) );
  NOR40 U1579 ( .A(n1297), .B(n1296), .C(n1295), .D(n1294), .Q(n1298) );
endmodule


module D_register_bank ( i_clk, i_rst_n, i_addr_Rs, i_con_RegWr, i_addr_Rd, 
        i_data_Rd, o_data_Rs, o_data_Rt, i_addr_Rt_4_, i_addr_Rt_3_, 
        i_addr_Rt_2_, i_addr_Rt_1_, i_addr_Rt_0_ );
  input [4:0] i_addr_Rs;
  input [4:0] i_addr_Rd;
  input [31:0] i_data_Rd;
  output [31:0] o_data_Rs;
  output [31:0] o_data_Rt;
  input i_clk, i_rst_n, i_con_RegWr, i_addr_Rt_4_, i_addr_Rt_3_, i_addr_Rt_2_,
         i_addr_Rt_1_, i_addr_Rt_0_;
  wire   n5, n6, n9, n11, n13, n15, n16, n17, n18, n20, n21, n22, n23, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n1, n2, n3, n4, n7, n8, n10, n12, n14, n19, n24,
         n33, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n232, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592;
  wire   [1023:0] regs;

  DFEC1 regs_reg_31__30_ ( .D(i_data_Rd[30]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1022]) );
  DFEC1 regs_reg_31__29_ ( .D(i_data_Rd[29]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1021]) );
  DFEC1 regs_reg_31__28_ ( .D(i_data_Rd[28]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1020]) );
  DFEC1 regs_reg_31__27_ ( .D(i_data_Rd[27]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1019]) );
  DFEC1 regs_reg_31__26_ ( .D(i_data_Rd[26]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1018]) );
  DFEC1 regs_reg_31__25_ ( .D(i_data_Rd[25]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1017]) );
  DFEC1 regs_reg_31__24_ ( .D(i_data_Rd[24]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1016]) );
  DFEC1 regs_reg_31__23_ ( .D(i_data_Rd[23]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1015]) );
  DFEC1 regs_reg_31__22_ ( .D(i_data_Rd[22]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1014]) );
  DFEC1 regs_reg_31__21_ ( .D(i_data_Rd[21]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1013]) );
  DFEC1 regs_reg_31__20_ ( .D(i_data_Rd[20]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1012]) );
  DFEC1 regs_reg_31__19_ ( .D(i_data_Rd[19]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1011]) );
  DFEC1 regs_reg_31__18_ ( .D(i_data_Rd[18]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1010]) );
  DFEC1 regs_reg_31__17_ ( .D(i_data_Rd[17]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1009]) );
  DFEC1 regs_reg_31__16_ ( .D(i_data_Rd[16]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1008]) );
  DFEC1 regs_reg_31__15_ ( .D(i_data_Rd[15]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1007]) );
  DFEC1 regs_reg_31__14_ ( .D(i_data_Rd[14]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1006]) );
  DFEC1 regs_reg_31__13_ ( .D(i_data_Rd[13]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1005]) );
  DFEC1 regs_reg_31__12_ ( .D(i_data_Rd[12]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1004]) );
  DFEC1 regs_reg_31__11_ ( .D(i_data_Rd[11]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1003]) );
  DFEC1 regs_reg_31__10_ ( .D(i_data_Rd[10]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1002]) );
  DFEC1 regs_reg_31__9_ ( .D(i_data_Rd[9]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1001]) );
  DFEC1 regs_reg_31__8_ ( .D(i_data_Rd[8]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[1000]) );
  DFEC1 regs_reg_31__7_ ( .D(i_data_Rd[7]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[999]) );
  DFEC1 regs_reg_31__6_ ( .D(i_data_Rd[6]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[998]) );
  DFEC1 regs_reg_31__5_ ( .D(i_data_Rd[5]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[997]) );
  DFEC1 regs_reg_31__4_ ( .D(i_data_Rd[4]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[996]) );
  DFEC1 regs_reg_31__3_ ( .D(i_data_Rd[3]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[995]) );
  DFEC1 regs_reg_31__2_ ( .D(i_data_Rd[2]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[994]) );
  DFEC1 regs_reg_31__1_ ( .D(i_data_Rd[1]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[993]) );
  DFEC1 regs_reg_31__0_ ( .D(i_data_Rd[0]), .E(n31), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[992]) );
  DFEC1 regs_reg_30__31_ ( .D(i_data_Rd[31]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[991]) );
  DFEC1 regs_reg_30__30_ ( .D(i_data_Rd[30]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[990]) );
  DFEC1 regs_reg_30__29_ ( .D(i_data_Rd[29]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[989]) );
  DFEC1 regs_reg_30__28_ ( .D(i_data_Rd[28]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[988]) );
  DFEC1 regs_reg_30__27_ ( .D(i_data_Rd[27]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[987]) );
  DFEC1 regs_reg_30__26_ ( .D(i_data_Rd[26]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[986]) );
  DFEC1 regs_reg_30__25_ ( .D(i_data_Rd[25]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[985]) );
  DFEC1 regs_reg_30__24_ ( .D(i_data_Rd[24]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[984]) );
  DFEC1 regs_reg_30__23_ ( .D(i_data_Rd[23]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[983]) );
  DFEC1 regs_reg_30__22_ ( .D(i_data_Rd[22]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[982]) );
  DFEC1 regs_reg_30__21_ ( .D(i_data_Rd[21]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[981]) );
  DFEC1 regs_reg_30__20_ ( .D(i_data_Rd[20]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[980]) );
  DFEC1 regs_reg_30__19_ ( .D(i_data_Rd[19]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[979]) );
  DFEC1 regs_reg_30__18_ ( .D(i_data_Rd[18]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[978]) );
  DFEC1 regs_reg_30__17_ ( .D(i_data_Rd[17]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[977]) );
  DFEC1 regs_reg_30__16_ ( .D(i_data_Rd[16]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[976]) );
  DFEC1 regs_reg_30__15_ ( .D(i_data_Rd[15]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[975]) );
  DFEC1 regs_reg_30__14_ ( .D(i_data_Rd[14]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[974]) );
  DFEC1 regs_reg_30__13_ ( .D(i_data_Rd[13]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[973]) );
  DFEC1 regs_reg_30__12_ ( .D(i_data_Rd[12]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[972]) );
  DFEC1 regs_reg_30__11_ ( .D(i_data_Rd[11]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[971]) );
  DFEC1 regs_reg_30__10_ ( .D(i_data_Rd[10]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[970]) );
  DFEC1 regs_reg_30__9_ ( .D(i_data_Rd[9]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[969]) );
  DFEC1 regs_reg_30__8_ ( .D(i_data_Rd[8]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[968]) );
  DFEC1 regs_reg_30__7_ ( .D(i_data_Rd[7]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[967]) );
  DFEC1 regs_reg_30__6_ ( .D(i_data_Rd[6]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[966]) );
  DFEC1 regs_reg_30__5_ ( .D(i_data_Rd[5]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[965]) );
  DFEC1 regs_reg_30__4_ ( .D(i_data_Rd[4]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[964]) );
  DFEC1 regs_reg_30__3_ ( .D(i_data_Rd[3]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[963]) );
  DFEC1 regs_reg_30__2_ ( .D(i_data_Rd[2]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[962]) );
  DFEC1 regs_reg_30__1_ ( .D(i_data_Rd[1]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[961]) );
  DFEC1 regs_reg_30__0_ ( .D(i_data_Rd[0]), .E(n30), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[960]) );
  DFEC1 regs_reg_29__31_ ( .D(i_data_Rd[31]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[959]) );
  DFEC1 regs_reg_29__30_ ( .D(i_data_Rd[30]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[958]) );
  DFEC1 regs_reg_29__29_ ( .D(i_data_Rd[29]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[957]) );
  DFEC1 regs_reg_29__28_ ( .D(i_data_Rd[28]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[956]) );
  DFEC1 regs_reg_29__27_ ( .D(i_data_Rd[27]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[955]) );
  DFEC1 regs_reg_29__26_ ( .D(i_data_Rd[26]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[954]) );
  DFEC1 regs_reg_29__25_ ( .D(i_data_Rd[25]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[953]) );
  DFEC1 regs_reg_29__24_ ( .D(i_data_Rd[24]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[952]) );
  DFEC1 regs_reg_29__23_ ( .D(i_data_Rd[23]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[951]) );
  DFEC1 regs_reg_29__22_ ( .D(i_data_Rd[22]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[950]) );
  DFEC1 regs_reg_29__21_ ( .D(i_data_Rd[21]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[949]) );
  DFEC1 regs_reg_29__20_ ( .D(i_data_Rd[20]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[948]) );
  DFEC1 regs_reg_29__19_ ( .D(i_data_Rd[19]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[947]) );
  DFEC1 regs_reg_29__18_ ( .D(i_data_Rd[18]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[946]) );
  DFEC1 regs_reg_29__17_ ( .D(i_data_Rd[17]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[945]) );
  DFEC1 regs_reg_29__16_ ( .D(i_data_Rd[16]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[944]) );
  DFEC1 regs_reg_29__15_ ( .D(i_data_Rd[15]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[943]) );
  DFEC1 regs_reg_29__14_ ( .D(i_data_Rd[14]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[942]) );
  DFEC1 regs_reg_29__13_ ( .D(i_data_Rd[13]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[941]) );
  DFEC1 regs_reg_29__12_ ( .D(i_data_Rd[12]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[940]) );
  DFEC1 regs_reg_29__11_ ( .D(i_data_Rd[11]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[939]) );
  DFEC1 regs_reg_29__10_ ( .D(i_data_Rd[10]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[938]) );
  DFEC1 regs_reg_29__9_ ( .D(i_data_Rd[9]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[937]) );
  DFEC1 regs_reg_29__8_ ( .D(i_data_Rd[8]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[936]) );
  DFEC1 regs_reg_29__7_ ( .D(i_data_Rd[7]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[935]) );
  DFEC1 regs_reg_29__6_ ( .D(i_data_Rd[6]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[934]) );
  DFEC1 regs_reg_29__5_ ( .D(i_data_Rd[5]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[933]) );
  DFEC1 regs_reg_29__4_ ( .D(i_data_Rd[4]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[932]) );
  DFEC1 regs_reg_29__3_ ( .D(i_data_Rd[3]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[931]) );
  DFEC1 regs_reg_29__2_ ( .D(i_data_Rd[2]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[930]) );
  DFEC1 regs_reg_29__1_ ( .D(i_data_Rd[1]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[929]) );
  DFEC1 regs_reg_29__0_ ( .D(i_data_Rd[0]), .E(n29), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[928]) );
  DFEC1 regs_reg_28__31_ ( .D(i_data_Rd[31]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[927]) );
  DFEC1 regs_reg_28__30_ ( .D(i_data_Rd[30]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[926]) );
  DFEC1 regs_reg_28__29_ ( .D(i_data_Rd[29]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[925]) );
  DFEC1 regs_reg_28__28_ ( .D(i_data_Rd[28]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[924]) );
  DFEC1 regs_reg_28__27_ ( .D(i_data_Rd[27]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[923]) );
  DFEC1 regs_reg_28__26_ ( .D(i_data_Rd[26]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[922]) );
  DFEC1 regs_reg_28__25_ ( .D(i_data_Rd[25]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[921]) );
  DFEC1 regs_reg_28__24_ ( .D(i_data_Rd[24]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[920]) );
  DFEC1 regs_reg_28__23_ ( .D(i_data_Rd[23]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[919]) );
  DFEC1 regs_reg_28__22_ ( .D(i_data_Rd[22]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[918]) );
  DFEC1 regs_reg_28__21_ ( .D(i_data_Rd[21]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[917]) );
  DFEC1 regs_reg_28__20_ ( .D(i_data_Rd[20]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[916]) );
  DFEC1 regs_reg_28__19_ ( .D(i_data_Rd[19]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[915]) );
  DFEC1 regs_reg_28__18_ ( .D(i_data_Rd[18]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[914]) );
  DFEC1 regs_reg_28__17_ ( .D(i_data_Rd[17]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[913]) );
  DFEC1 regs_reg_28__16_ ( .D(i_data_Rd[16]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[912]) );
  DFEC1 regs_reg_28__15_ ( .D(i_data_Rd[15]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[911]) );
  DFEC1 regs_reg_28__14_ ( .D(i_data_Rd[14]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[910]) );
  DFEC1 regs_reg_28__13_ ( .D(i_data_Rd[13]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[909]) );
  DFEC1 regs_reg_28__12_ ( .D(i_data_Rd[12]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[908]) );
  DFEC1 regs_reg_28__11_ ( .D(i_data_Rd[11]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[907]) );
  DFEC1 regs_reg_28__10_ ( .D(i_data_Rd[10]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[906]) );
  DFEC1 regs_reg_28__9_ ( .D(i_data_Rd[9]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[905]) );
  DFEC1 regs_reg_28__8_ ( .D(i_data_Rd[8]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[904]) );
  DFEC1 regs_reg_28__7_ ( .D(i_data_Rd[7]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[903]) );
  DFEC1 regs_reg_28__6_ ( .D(i_data_Rd[6]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[902]) );
  DFEC1 regs_reg_28__5_ ( .D(i_data_Rd[5]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[901]) );
  DFEC1 regs_reg_28__4_ ( .D(i_data_Rd[4]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[900]) );
  DFEC1 regs_reg_28__3_ ( .D(i_data_Rd[3]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[899]) );
  DFEC1 regs_reg_28__2_ ( .D(i_data_Rd[2]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[898]) );
  DFEC1 regs_reg_28__1_ ( .D(i_data_Rd[1]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[897]) );
  DFEC1 regs_reg_28__0_ ( .D(i_data_Rd[0]), .E(n28), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[896]) );
  DFEC1 regs_reg_27__31_ ( .D(i_data_Rd[31]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[895]) );
  DFEC1 regs_reg_27__30_ ( .D(i_data_Rd[30]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[894]) );
  DFEC1 regs_reg_27__29_ ( .D(i_data_Rd[29]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[893]) );
  DFEC1 regs_reg_27__28_ ( .D(i_data_Rd[28]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[892]) );
  DFEC1 regs_reg_27__27_ ( .D(i_data_Rd[27]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[891]) );
  DFEC1 regs_reg_27__26_ ( .D(i_data_Rd[26]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[890]) );
  DFEC1 regs_reg_27__25_ ( .D(i_data_Rd[25]), .E(n27), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[889]) );
  DFEC1 regs_reg_27__24_ ( .D(i_data_Rd[24]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[888]) );
  DFEC1 regs_reg_27__23_ ( .D(i_data_Rd[23]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[887]) );
  DFEC1 regs_reg_27__22_ ( .D(i_data_Rd[22]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[886]) );
  DFEC1 regs_reg_27__21_ ( .D(i_data_Rd[21]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[885]) );
  DFEC1 regs_reg_27__20_ ( .D(i_data_Rd[20]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[884]) );
  DFEC1 regs_reg_27__19_ ( .D(i_data_Rd[19]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[883]) );
  DFEC1 regs_reg_27__18_ ( .D(i_data_Rd[18]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[882]) );
  DFEC1 regs_reg_27__17_ ( .D(i_data_Rd[17]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[881]) );
  DFEC1 regs_reg_27__16_ ( .D(i_data_Rd[16]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[880]) );
  DFEC1 regs_reg_27__15_ ( .D(i_data_Rd[15]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[879]) );
  DFEC1 regs_reg_27__14_ ( .D(i_data_Rd[14]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[878]) );
  DFEC1 regs_reg_27__13_ ( .D(i_data_Rd[13]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[877]) );
  DFEC1 regs_reg_27__12_ ( .D(i_data_Rd[12]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[876]) );
  DFEC1 regs_reg_27__11_ ( .D(i_data_Rd[11]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[875]) );
  DFEC1 regs_reg_27__10_ ( .D(i_data_Rd[10]), .E(n256), .C(i_clk), .RN(i_rst_n), .Q(regs[874]) );
  DFEC1 regs_reg_27__9_ ( .D(i_data_Rd[9]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[873]) );
  DFEC1 regs_reg_27__8_ ( .D(i_data_Rd[8]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[872]) );
  DFEC1 regs_reg_27__7_ ( .D(i_data_Rd[7]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[871]) );
  DFEC1 regs_reg_27__6_ ( .D(i_data_Rd[6]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[870]) );
  DFEC1 regs_reg_27__5_ ( .D(i_data_Rd[5]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[869]) );
  DFEC1 regs_reg_27__4_ ( .D(i_data_Rd[4]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[868]) );
  DFEC1 regs_reg_27__3_ ( .D(i_data_Rd[3]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[867]) );
  DFEC1 regs_reg_27__2_ ( .D(i_data_Rd[2]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[866]) );
  DFEC1 regs_reg_27__1_ ( .D(i_data_Rd[1]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[865]) );
  DFEC1 regs_reg_27__0_ ( .D(i_data_Rd[0]), .E(n256), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[864]) );
  DFEC1 regs_reg_26__31_ ( .D(i_data_Rd[31]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[863]) );
  DFEC1 regs_reg_26__30_ ( .D(i_data_Rd[30]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[862]) );
  DFEC1 regs_reg_26__29_ ( .D(i_data_Rd[29]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[861]) );
  DFEC1 regs_reg_26__28_ ( .D(i_data_Rd[28]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[860]) );
  DFEC1 regs_reg_26__27_ ( .D(i_data_Rd[27]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[859]) );
  DFEC1 regs_reg_26__26_ ( .D(i_data_Rd[26]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[858]) );
  DFEC1 regs_reg_26__25_ ( .D(i_data_Rd[25]), .E(n26), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[857]) );
  DFEC1 regs_reg_26__24_ ( .D(i_data_Rd[24]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[856]) );
  DFEC1 regs_reg_26__23_ ( .D(i_data_Rd[23]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[855]) );
  DFEC1 regs_reg_26__22_ ( .D(i_data_Rd[22]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[854]) );
  DFEC1 regs_reg_26__21_ ( .D(i_data_Rd[21]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[853]) );
  DFEC1 regs_reg_26__20_ ( .D(i_data_Rd[20]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[852]) );
  DFEC1 regs_reg_26__19_ ( .D(i_data_Rd[19]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[851]) );
  DFEC1 regs_reg_26__18_ ( .D(i_data_Rd[18]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[850]) );
  DFEC1 regs_reg_26__17_ ( .D(i_data_Rd[17]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[849]) );
  DFEC1 regs_reg_26__16_ ( .D(i_data_Rd[16]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[848]) );
  DFEC1 regs_reg_26__15_ ( .D(i_data_Rd[15]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[847]) );
  DFEC1 regs_reg_26__14_ ( .D(i_data_Rd[14]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[846]) );
  DFEC1 regs_reg_26__13_ ( .D(i_data_Rd[13]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[845]) );
  DFEC1 regs_reg_26__12_ ( .D(i_data_Rd[12]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[844]) );
  DFEC1 regs_reg_26__11_ ( .D(i_data_Rd[11]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[843]) );
  DFEC1 regs_reg_26__10_ ( .D(i_data_Rd[10]), .E(n257), .C(i_clk), .RN(i_rst_n), .Q(regs[842]) );
  DFEC1 regs_reg_26__9_ ( .D(i_data_Rd[9]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[841]) );
  DFEC1 regs_reg_26__8_ ( .D(i_data_Rd[8]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[840]) );
  DFEC1 regs_reg_26__7_ ( .D(i_data_Rd[7]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[839]) );
  DFEC1 regs_reg_26__6_ ( .D(i_data_Rd[6]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[838]) );
  DFEC1 regs_reg_26__5_ ( .D(i_data_Rd[5]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[837]) );
  DFEC1 regs_reg_26__4_ ( .D(i_data_Rd[4]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[836]) );
  DFEC1 regs_reg_26__3_ ( .D(i_data_Rd[3]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[835]) );
  DFEC1 regs_reg_26__2_ ( .D(i_data_Rd[2]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[834]) );
  DFEC1 regs_reg_26__1_ ( .D(i_data_Rd[1]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[833]) );
  DFEC1 regs_reg_26__0_ ( .D(i_data_Rd[0]), .E(n257), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[832]) );
  DFEC1 regs_reg_25__31_ ( .D(i_data_Rd[31]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[831]) );
  DFEC1 regs_reg_25__30_ ( .D(i_data_Rd[30]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[830]) );
  DFEC1 regs_reg_25__29_ ( .D(i_data_Rd[29]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[829]) );
  DFEC1 regs_reg_25__28_ ( .D(i_data_Rd[28]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[828]) );
  DFEC1 regs_reg_25__27_ ( .D(i_data_Rd[27]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[827]) );
  DFEC1 regs_reg_25__26_ ( .D(i_data_Rd[26]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[826]) );
  DFEC1 regs_reg_25__25_ ( .D(i_data_Rd[25]), .E(n25), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[825]) );
  DFEC1 regs_reg_25__24_ ( .D(i_data_Rd[24]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[824]) );
  DFEC1 regs_reg_25__23_ ( .D(i_data_Rd[23]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[823]) );
  DFEC1 regs_reg_25__22_ ( .D(i_data_Rd[22]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[822]) );
  DFEC1 regs_reg_25__21_ ( .D(i_data_Rd[21]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[821]) );
  DFEC1 regs_reg_25__20_ ( .D(i_data_Rd[20]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[820]) );
  DFEC1 regs_reg_25__19_ ( .D(i_data_Rd[19]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[819]) );
  DFEC1 regs_reg_25__18_ ( .D(i_data_Rd[18]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[818]) );
  DFEC1 regs_reg_25__17_ ( .D(i_data_Rd[17]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[817]) );
  DFEC1 regs_reg_25__16_ ( .D(i_data_Rd[16]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[816]) );
  DFEC1 regs_reg_25__15_ ( .D(i_data_Rd[15]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[815]) );
  DFEC1 regs_reg_25__14_ ( .D(i_data_Rd[14]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[814]) );
  DFEC1 regs_reg_25__13_ ( .D(i_data_Rd[13]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[813]) );
  DFEC1 regs_reg_25__12_ ( .D(i_data_Rd[12]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[812]) );
  DFEC1 regs_reg_25__11_ ( .D(i_data_Rd[11]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[811]) );
  DFEC1 regs_reg_25__10_ ( .D(i_data_Rd[10]), .E(n258), .C(i_clk), .RN(i_rst_n), .Q(regs[810]) );
  DFEC1 regs_reg_25__9_ ( .D(i_data_Rd[9]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[809]) );
  DFEC1 regs_reg_25__8_ ( .D(i_data_Rd[8]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[808]) );
  DFEC1 regs_reg_25__7_ ( .D(i_data_Rd[7]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[807]) );
  DFEC1 regs_reg_25__6_ ( .D(i_data_Rd[6]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[806]) );
  DFEC1 regs_reg_25__5_ ( .D(i_data_Rd[5]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[805]) );
  DFEC1 regs_reg_25__4_ ( .D(i_data_Rd[4]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[804]) );
  DFEC1 regs_reg_25__3_ ( .D(i_data_Rd[3]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[803]) );
  DFEC1 regs_reg_25__2_ ( .D(i_data_Rd[2]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[802]) );
  DFEC1 regs_reg_25__1_ ( .D(i_data_Rd[1]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[801]) );
  DFEC1 regs_reg_25__0_ ( .D(i_data_Rd[0]), .E(n258), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[800]) );
  DFEC1 regs_reg_24__31_ ( .D(i_data_Rd[31]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[799]) );
  DFEC1 regs_reg_24__30_ ( .D(i_data_Rd[30]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[798]) );
  DFEC1 regs_reg_24__29_ ( .D(i_data_Rd[29]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[797]) );
  DFEC1 regs_reg_24__28_ ( .D(i_data_Rd[28]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[796]) );
  DFEC1 regs_reg_24__27_ ( .D(i_data_Rd[27]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[795]) );
  DFEC1 regs_reg_24__26_ ( .D(i_data_Rd[26]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[794]) );
  DFEC1 regs_reg_24__25_ ( .D(i_data_Rd[25]), .E(n23), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[793]) );
  DFEC1 regs_reg_24__24_ ( .D(i_data_Rd[24]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[792]) );
  DFEC1 regs_reg_24__23_ ( .D(i_data_Rd[23]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[791]) );
  DFEC1 regs_reg_24__22_ ( .D(i_data_Rd[22]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[790]) );
  DFEC1 regs_reg_24__21_ ( .D(i_data_Rd[21]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[789]) );
  DFEC1 regs_reg_24__20_ ( .D(i_data_Rd[20]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[788]) );
  DFEC1 regs_reg_24__19_ ( .D(i_data_Rd[19]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[787]) );
  DFEC1 regs_reg_24__18_ ( .D(i_data_Rd[18]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[786]) );
  DFEC1 regs_reg_24__17_ ( .D(i_data_Rd[17]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[785]) );
  DFEC1 regs_reg_24__16_ ( .D(i_data_Rd[16]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[784]) );
  DFEC1 regs_reg_24__15_ ( .D(i_data_Rd[15]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[783]) );
  DFEC1 regs_reg_24__14_ ( .D(i_data_Rd[14]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[782]) );
  DFEC1 regs_reg_24__13_ ( .D(i_data_Rd[13]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[781]) );
  DFEC1 regs_reg_24__12_ ( .D(i_data_Rd[12]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[780]) );
  DFEC1 regs_reg_24__11_ ( .D(i_data_Rd[11]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[779]) );
  DFEC1 regs_reg_24__10_ ( .D(i_data_Rd[10]), .E(n259), .C(i_clk), .RN(i_rst_n), .Q(regs[778]) );
  DFEC1 regs_reg_24__9_ ( .D(i_data_Rd[9]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[777]) );
  DFEC1 regs_reg_24__8_ ( .D(i_data_Rd[8]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[776]) );
  DFEC1 regs_reg_24__7_ ( .D(i_data_Rd[7]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[775]) );
  DFEC1 regs_reg_24__6_ ( .D(i_data_Rd[6]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[774]) );
  DFEC1 regs_reg_24__5_ ( .D(i_data_Rd[5]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[773]) );
  DFEC1 regs_reg_24__4_ ( .D(i_data_Rd[4]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[772]) );
  DFEC1 regs_reg_24__3_ ( .D(i_data_Rd[3]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[771]) );
  DFEC1 regs_reg_24__2_ ( .D(i_data_Rd[2]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[770]) );
  DFEC1 regs_reg_24__1_ ( .D(i_data_Rd[1]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[769]) );
  DFEC1 regs_reg_24__0_ ( .D(i_data_Rd[0]), .E(n259), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[768]) );
  DFEC1 regs_reg_23__31_ ( .D(i_data_Rd[31]), .E(n22), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[767]) );
  DFEC1 regs_reg_23__30_ ( .D(i_data_Rd[30]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[766]) );
  DFEC1 regs_reg_23__29_ ( .D(i_data_Rd[29]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[765]) );
  DFEC1 regs_reg_23__28_ ( .D(i_data_Rd[28]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[764]) );
  DFEC1 regs_reg_23__27_ ( .D(i_data_Rd[27]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[763]) );
  DFEC1 regs_reg_23__26_ ( .D(i_data_Rd[26]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[762]) );
  DFEC1 regs_reg_23__25_ ( .D(i_data_Rd[25]), .E(n22), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[761]) );
  DFEC1 regs_reg_23__24_ ( .D(i_data_Rd[24]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[760]) );
  DFEC1 regs_reg_23__23_ ( .D(i_data_Rd[23]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[759]) );
  DFEC1 regs_reg_23__22_ ( .D(i_data_Rd[22]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[758]) );
  DFEC1 regs_reg_23__21_ ( .D(i_data_Rd[21]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[757]) );
  DFEC1 regs_reg_23__20_ ( .D(i_data_Rd[20]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[756]) );
  DFEC1 regs_reg_23__19_ ( .D(i_data_Rd[19]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[755]) );
  DFEC1 regs_reg_23__18_ ( .D(i_data_Rd[18]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[754]) );
  DFEC1 regs_reg_23__17_ ( .D(i_data_Rd[17]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[753]) );
  DFEC1 regs_reg_23__16_ ( .D(i_data_Rd[16]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[752]) );
  DFEC1 regs_reg_23__15_ ( .D(i_data_Rd[15]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[751]) );
  DFEC1 regs_reg_23__14_ ( .D(i_data_Rd[14]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[750]) );
  DFEC1 regs_reg_23__13_ ( .D(i_data_Rd[13]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[749]) );
  DFEC1 regs_reg_23__12_ ( .D(i_data_Rd[12]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[748]) );
  DFEC1 regs_reg_23__11_ ( .D(i_data_Rd[11]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[747]) );
  DFEC1 regs_reg_23__10_ ( .D(i_data_Rd[10]), .E(n260), .C(i_clk), .RN(i_rst_n), .Q(regs[746]) );
  DFEC1 regs_reg_23__9_ ( .D(i_data_Rd[9]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[745]) );
  DFEC1 regs_reg_23__8_ ( .D(i_data_Rd[8]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[744]) );
  DFEC1 regs_reg_23__7_ ( .D(i_data_Rd[7]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[743]) );
  DFEC1 regs_reg_23__6_ ( .D(i_data_Rd[6]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[742]) );
  DFEC1 regs_reg_23__5_ ( .D(i_data_Rd[5]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[741]) );
  DFEC1 regs_reg_23__4_ ( .D(i_data_Rd[4]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[740]) );
  DFEC1 regs_reg_23__3_ ( .D(i_data_Rd[3]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[739]) );
  DFEC1 regs_reg_23__2_ ( .D(i_data_Rd[2]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[738]) );
  DFEC1 regs_reg_23__1_ ( .D(i_data_Rd[1]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[737]) );
  DFEC1 regs_reg_23__0_ ( .D(i_data_Rd[0]), .E(n260), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[736]) );
  DFEC1 regs_reg_22__31_ ( .D(i_data_Rd[31]), .E(n21), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[735]) );
  DFEC1 regs_reg_22__30_ ( .D(i_data_Rd[30]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[734]) );
  DFEC1 regs_reg_22__29_ ( .D(i_data_Rd[29]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[733]) );
  DFEC1 regs_reg_22__28_ ( .D(i_data_Rd[28]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[732]) );
  DFEC1 regs_reg_22__27_ ( .D(i_data_Rd[27]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[731]) );
  DFEC1 regs_reg_22__26_ ( .D(i_data_Rd[26]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[730]) );
  DFEC1 regs_reg_22__25_ ( .D(i_data_Rd[25]), .E(n21), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[729]) );
  DFEC1 regs_reg_22__24_ ( .D(i_data_Rd[24]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[728]) );
  DFEC1 regs_reg_22__23_ ( .D(i_data_Rd[23]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[727]) );
  DFEC1 regs_reg_22__22_ ( .D(i_data_Rd[22]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[726]) );
  DFEC1 regs_reg_22__21_ ( .D(i_data_Rd[21]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[725]) );
  DFEC1 regs_reg_22__20_ ( .D(i_data_Rd[20]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[724]) );
  DFEC1 regs_reg_22__19_ ( .D(i_data_Rd[19]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[723]) );
  DFEC1 regs_reg_22__18_ ( .D(i_data_Rd[18]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[722]) );
  DFEC1 regs_reg_22__17_ ( .D(i_data_Rd[17]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[721]) );
  DFEC1 regs_reg_22__16_ ( .D(i_data_Rd[16]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[720]) );
  DFEC1 regs_reg_22__15_ ( .D(i_data_Rd[15]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[719]) );
  DFEC1 regs_reg_22__14_ ( .D(i_data_Rd[14]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[718]) );
  DFEC1 regs_reg_22__13_ ( .D(i_data_Rd[13]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[717]) );
  DFEC1 regs_reg_22__12_ ( .D(i_data_Rd[12]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[716]) );
  DFEC1 regs_reg_22__11_ ( .D(i_data_Rd[11]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[715]) );
  DFEC1 regs_reg_22__10_ ( .D(i_data_Rd[10]), .E(n261), .C(i_clk), .RN(i_rst_n), .Q(regs[714]) );
  DFEC1 regs_reg_22__9_ ( .D(i_data_Rd[9]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[713]) );
  DFEC1 regs_reg_22__8_ ( .D(i_data_Rd[8]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[712]) );
  DFEC1 regs_reg_22__7_ ( .D(i_data_Rd[7]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[711]) );
  DFEC1 regs_reg_22__6_ ( .D(i_data_Rd[6]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[710]) );
  DFEC1 regs_reg_22__5_ ( .D(i_data_Rd[5]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[709]) );
  DFEC1 regs_reg_22__4_ ( .D(i_data_Rd[4]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[708]) );
  DFEC1 regs_reg_22__3_ ( .D(i_data_Rd[3]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[707]) );
  DFEC1 regs_reg_22__2_ ( .D(i_data_Rd[2]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[706]) );
  DFEC1 regs_reg_22__1_ ( .D(i_data_Rd[1]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[705]) );
  DFEC1 regs_reg_22__0_ ( .D(i_data_Rd[0]), .E(n261), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[704]) );
  DFEC1 regs_reg_21__31_ ( .D(i_data_Rd[31]), .E(n20), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[703]) );
  DFEC1 regs_reg_21__30_ ( .D(i_data_Rd[30]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[702]) );
  DFEC1 regs_reg_21__29_ ( .D(i_data_Rd[29]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[701]) );
  DFEC1 regs_reg_21__28_ ( .D(i_data_Rd[28]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[700]) );
  DFEC1 regs_reg_21__27_ ( .D(i_data_Rd[27]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[699]) );
  DFEC1 regs_reg_21__26_ ( .D(i_data_Rd[26]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[698]) );
  DFEC1 regs_reg_21__25_ ( .D(i_data_Rd[25]), .E(n20), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[697]) );
  DFEC1 regs_reg_21__24_ ( .D(i_data_Rd[24]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[696]) );
  DFEC1 regs_reg_21__23_ ( .D(i_data_Rd[23]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[695]) );
  DFEC1 regs_reg_21__22_ ( .D(i_data_Rd[22]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[694]) );
  DFEC1 regs_reg_21__21_ ( .D(i_data_Rd[21]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[693]) );
  DFEC1 regs_reg_21__20_ ( .D(i_data_Rd[20]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[692]) );
  DFEC1 regs_reg_21__19_ ( .D(i_data_Rd[19]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[691]) );
  DFEC1 regs_reg_21__18_ ( .D(i_data_Rd[18]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[690]) );
  DFEC1 regs_reg_21__17_ ( .D(i_data_Rd[17]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[689]) );
  DFEC1 regs_reg_21__16_ ( .D(i_data_Rd[16]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[688]) );
  DFEC1 regs_reg_21__15_ ( .D(i_data_Rd[15]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[687]) );
  DFEC1 regs_reg_21__14_ ( .D(i_data_Rd[14]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[686]) );
  DFEC1 regs_reg_21__13_ ( .D(i_data_Rd[13]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[685]) );
  DFEC1 regs_reg_21__12_ ( .D(i_data_Rd[12]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[684]) );
  DFEC1 regs_reg_21__11_ ( .D(i_data_Rd[11]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[683]) );
  DFEC1 regs_reg_21__10_ ( .D(i_data_Rd[10]), .E(n262), .C(i_clk), .RN(i_rst_n), .Q(regs[682]) );
  DFEC1 regs_reg_21__9_ ( .D(i_data_Rd[9]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[681]) );
  DFEC1 regs_reg_21__8_ ( .D(i_data_Rd[8]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[680]) );
  DFEC1 regs_reg_21__7_ ( .D(i_data_Rd[7]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[679]) );
  DFEC1 regs_reg_21__6_ ( .D(i_data_Rd[6]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[678]) );
  DFEC1 regs_reg_21__5_ ( .D(i_data_Rd[5]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[677]) );
  DFEC1 regs_reg_21__4_ ( .D(i_data_Rd[4]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[676]) );
  DFEC1 regs_reg_21__3_ ( .D(i_data_Rd[3]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[675]) );
  DFEC1 regs_reg_21__2_ ( .D(i_data_Rd[2]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[674]) );
  DFEC1 regs_reg_21__1_ ( .D(i_data_Rd[1]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[673]) );
  DFEC1 regs_reg_21__0_ ( .D(i_data_Rd[0]), .E(n262), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[672]) );
  DFEC1 regs_reg_20__31_ ( .D(i_data_Rd[31]), .E(n18), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[671]) );
  DFEC1 regs_reg_20__30_ ( .D(i_data_Rd[30]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[670]) );
  DFEC1 regs_reg_20__29_ ( .D(i_data_Rd[29]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[669]) );
  DFEC1 regs_reg_20__28_ ( .D(i_data_Rd[28]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[668]) );
  DFEC1 regs_reg_20__27_ ( .D(i_data_Rd[27]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[667]) );
  DFEC1 regs_reg_20__26_ ( .D(i_data_Rd[26]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[666]) );
  DFEC1 regs_reg_20__25_ ( .D(i_data_Rd[25]), .E(n18), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[665]) );
  DFEC1 regs_reg_20__24_ ( .D(i_data_Rd[24]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[664]) );
  DFEC1 regs_reg_20__23_ ( .D(i_data_Rd[23]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[663]) );
  DFEC1 regs_reg_20__22_ ( .D(i_data_Rd[22]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[662]) );
  DFEC1 regs_reg_20__21_ ( .D(i_data_Rd[21]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[661]) );
  DFEC1 regs_reg_20__20_ ( .D(i_data_Rd[20]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[660]) );
  DFEC1 regs_reg_20__19_ ( .D(i_data_Rd[19]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[659]) );
  DFEC1 regs_reg_20__18_ ( .D(i_data_Rd[18]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[658]) );
  DFEC1 regs_reg_20__17_ ( .D(i_data_Rd[17]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[657]) );
  DFEC1 regs_reg_20__16_ ( .D(i_data_Rd[16]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[656]) );
  DFEC1 regs_reg_20__15_ ( .D(i_data_Rd[15]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[655]) );
  DFEC1 regs_reg_20__14_ ( .D(i_data_Rd[14]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[654]) );
  DFEC1 regs_reg_20__13_ ( .D(i_data_Rd[13]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[653]) );
  DFEC1 regs_reg_20__12_ ( .D(i_data_Rd[12]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[652]) );
  DFEC1 regs_reg_20__11_ ( .D(i_data_Rd[11]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[651]) );
  DFEC1 regs_reg_20__10_ ( .D(i_data_Rd[10]), .E(n263), .C(i_clk), .RN(i_rst_n), .Q(regs[650]) );
  DFEC1 regs_reg_20__9_ ( .D(i_data_Rd[9]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[649]) );
  DFEC1 regs_reg_20__8_ ( .D(i_data_Rd[8]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[648]) );
  DFEC1 regs_reg_20__7_ ( .D(i_data_Rd[7]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[647]) );
  DFEC1 regs_reg_20__6_ ( .D(i_data_Rd[6]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[646]) );
  DFEC1 regs_reg_20__5_ ( .D(i_data_Rd[5]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[645]) );
  DFEC1 regs_reg_20__4_ ( .D(i_data_Rd[4]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[644]) );
  DFEC1 regs_reg_20__3_ ( .D(i_data_Rd[3]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[643]) );
  DFEC1 regs_reg_20__2_ ( .D(i_data_Rd[2]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[642]) );
  DFEC1 regs_reg_20__1_ ( .D(i_data_Rd[1]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[641]) );
  DFEC1 regs_reg_20__0_ ( .D(i_data_Rd[0]), .E(n263), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[640]) );
  DFEC1 regs_reg_19__31_ ( .D(i_data_Rd[31]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[639]) );
  DFEC1 regs_reg_19__30_ ( .D(i_data_Rd[30]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[638]) );
  DFEC1 regs_reg_19__29_ ( .D(i_data_Rd[29]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[637]) );
  DFEC1 regs_reg_19__28_ ( .D(i_data_Rd[28]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[636]) );
  DFEC1 regs_reg_19__27_ ( .D(i_data_Rd[27]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[635]) );
  DFEC1 regs_reg_19__26_ ( .D(i_data_Rd[26]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[634]) );
  DFEC1 regs_reg_19__25_ ( .D(i_data_Rd[25]), .E(n17), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[633]) );
  DFEC1 regs_reg_19__24_ ( .D(i_data_Rd[24]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[632]) );
  DFEC1 regs_reg_19__23_ ( .D(i_data_Rd[23]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[631]) );
  DFEC1 regs_reg_19__22_ ( .D(i_data_Rd[22]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[630]) );
  DFEC1 regs_reg_19__21_ ( .D(i_data_Rd[21]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[629]) );
  DFEC1 regs_reg_19__20_ ( .D(i_data_Rd[20]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[628]) );
  DFEC1 regs_reg_19__19_ ( .D(i_data_Rd[19]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[627]) );
  DFEC1 regs_reg_19__18_ ( .D(i_data_Rd[18]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[626]) );
  DFEC1 regs_reg_19__17_ ( .D(i_data_Rd[17]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[625]) );
  DFEC1 regs_reg_19__16_ ( .D(i_data_Rd[16]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[624]) );
  DFEC1 regs_reg_19__15_ ( .D(i_data_Rd[15]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[623]) );
  DFEC1 regs_reg_19__14_ ( .D(i_data_Rd[14]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[622]) );
  DFEC1 regs_reg_19__13_ ( .D(i_data_Rd[13]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[621]) );
  DFEC1 regs_reg_19__12_ ( .D(i_data_Rd[12]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[620]) );
  DFEC1 regs_reg_19__11_ ( .D(i_data_Rd[11]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[619]) );
  DFEC1 regs_reg_19__10_ ( .D(i_data_Rd[10]), .E(n264), .C(i_clk), .RN(i_rst_n), .Q(regs[618]) );
  DFEC1 regs_reg_19__9_ ( .D(i_data_Rd[9]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[617]) );
  DFEC1 regs_reg_19__8_ ( .D(i_data_Rd[8]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[616]) );
  DFEC1 regs_reg_19__7_ ( .D(i_data_Rd[7]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[615]) );
  DFEC1 regs_reg_19__6_ ( .D(i_data_Rd[6]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[614]) );
  DFEC1 regs_reg_19__5_ ( .D(i_data_Rd[5]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[613]) );
  DFEC1 regs_reg_19__4_ ( .D(i_data_Rd[4]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[612]) );
  DFEC1 regs_reg_19__3_ ( .D(i_data_Rd[3]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[611]) );
  DFEC1 regs_reg_19__2_ ( .D(i_data_Rd[2]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[610]) );
  DFEC1 regs_reg_19__1_ ( .D(i_data_Rd[1]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[609]) );
  DFEC1 regs_reg_19__0_ ( .D(i_data_Rd[0]), .E(n264), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[608]) );
  DFEC1 regs_reg_18__31_ ( .D(i_data_Rd[31]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[607]) );
  DFEC1 regs_reg_18__30_ ( .D(i_data_Rd[30]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[606]) );
  DFEC1 regs_reg_18__29_ ( .D(i_data_Rd[29]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[605]) );
  DFEC1 regs_reg_18__28_ ( .D(i_data_Rd[28]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[604]) );
  DFEC1 regs_reg_18__27_ ( .D(i_data_Rd[27]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[603]) );
  DFEC1 regs_reg_18__26_ ( .D(i_data_Rd[26]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[602]) );
  DFEC1 regs_reg_18__25_ ( .D(i_data_Rd[25]), .E(n16), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[601]) );
  DFEC1 regs_reg_18__24_ ( .D(i_data_Rd[24]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[600]) );
  DFEC1 regs_reg_18__23_ ( .D(i_data_Rd[23]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[599]) );
  DFEC1 regs_reg_18__22_ ( .D(i_data_Rd[22]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[598]) );
  DFEC1 regs_reg_18__21_ ( .D(i_data_Rd[21]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[597]) );
  DFEC1 regs_reg_18__20_ ( .D(i_data_Rd[20]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[596]) );
  DFEC1 regs_reg_18__19_ ( .D(i_data_Rd[19]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[595]) );
  DFEC1 regs_reg_18__18_ ( .D(i_data_Rd[18]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[594]) );
  DFEC1 regs_reg_18__17_ ( .D(i_data_Rd[17]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[593]) );
  DFEC1 regs_reg_18__16_ ( .D(i_data_Rd[16]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[592]) );
  DFEC1 regs_reg_18__15_ ( .D(i_data_Rd[15]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[591]) );
  DFEC1 regs_reg_18__14_ ( .D(i_data_Rd[14]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[590]) );
  DFEC1 regs_reg_18__13_ ( .D(i_data_Rd[13]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[589]) );
  DFEC1 regs_reg_18__12_ ( .D(i_data_Rd[12]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[588]) );
  DFEC1 regs_reg_18__11_ ( .D(i_data_Rd[11]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[587]) );
  DFEC1 regs_reg_18__10_ ( .D(i_data_Rd[10]), .E(n265), .C(i_clk), .RN(i_rst_n), .Q(regs[586]) );
  DFEC1 regs_reg_18__9_ ( .D(i_data_Rd[9]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[585]) );
  DFEC1 regs_reg_18__8_ ( .D(i_data_Rd[8]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[584]) );
  DFEC1 regs_reg_18__7_ ( .D(i_data_Rd[7]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[583]) );
  DFEC1 regs_reg_18__6_ ( .D(i_data_Rd[6]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[582]) );
  DFEC1 regs_reg_18__5_ ( .D(i_data_Rd[5]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[581]) );
  DFEC1 regs_reg_18__4_ ( .D(i_data_Rd[4]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[580]) );
  DFEC1 regs_reg_18__3_ ( .D(i_data_Rd[3]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[579]) );
  DFEC1 regs_reg_18__2_ ( .D(i_data_Rd[2]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[578]) );
  DFEC1 regs_reg_18__1_ ( .D(i_data_Rd[1]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[577]) );
  DFEC1 regs_reg_18__0_ ( .D(i_data_Rd[0]), .E(n265), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[576]) );
  DFEC1 regs_reg_17__31_ ( .D(i_data_Rd[31]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[575]) );
  DFEC1 regs_reg_17__30_ ( .D(i_data_Rd[30]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[574]) );
  DFEC1 regs_reg_17__29_ ( .D(i_data_Rd[29]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[573]) );
  DFEC1 regs_reg_17__28_ ( .D(i_data_Rd[28]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[572]) );
  DFEC1 regs_reg_17__27_ ( .D(i_data_Rd[27]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[571]) );
  DFEC1 regs_reg_17__26_ ( .D(i_data_Rd[26]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[570]) );
  DFEC1 regs_reg_17__25_ ( .D(i_data_Rd[25]), .E(n15), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[569]) );
  DFEC1 regs_reg_17__24_ ( .D(i_data_Rd[24]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[568]) );
  DFEC1 regs_reg_17__23_ ( .D(i_data_Rd[23]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[567]) );
  DFEC1 regs_reg_17__22_ ( .D(i_data_Rd[22]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[566]) );
  DFEC1 regs_reg_17__21_ ( .D(i_data_Rd[21]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[565]) );
  DFEC1 regs_reg_17__20_ ( .D(i_data_Rd[20]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[564]) );
  DFEC1 regs_reg_17__19_ ( .D(i_data_Rd[19]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[563]) );
  DFEC1 regs_reg_17__18_ ( .D(i_data_Rd[18]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[562]) );
  DFEC1 regs_reg_17__17_ ( .D(i_data_Rd[17]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[561]) );
  DFEC1 regs_reg_17__16_ ( .D(i_data_Rd[16]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[560]) );
  DFEC1 regs_reg_17__15_ ( .D(i_data_Rd[15]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[559]) );
  DFEC1 regs_reg_17__14_ ( .D(i_data_Rd[14]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[558]) );
  DFEC1 regs_reg_17__13_ ( .D(i_data_Rd[13]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[557]) );
  DFEC1 regs_reg_17__12_ ( .D(i_data_Rd[12]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[556]) );
  DFEC1 regs_reg_17__11_ ( .D(i_data_Rd[11]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[555]) );
  DFEC1 regs_reg_17__10_ ( .D(i_data_Rd[10]), .E(n266), .C(i_clk), .RN(i_rst_n), .Q(regs[554]) );
  DFEC1 regs_reg_17__9_ ( .D(i_data_Rd[9]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[553]) );
  DFEC1 regs_reg_17__8_ ( .D(i_data_Rd[8]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[552]) );
  DFEC1 regs_reg_17__7_ ( .D(i_data_Rd[7]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[551]) );
  DFEC1 regs_reg_17__6_ ( .D(i_data_Rd[6]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[550]) );
  DFEC1 regs_reg_17__5_ ( .D(i_data_Rd[5]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[549]) );
  DFEC1 regs_reg_17__4_ ( .D(i_data_Rd[4]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[548]) );
  DFEC1 regs_reg_17__3_ ( .D(i_data_Rd[3]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[547]) );
  DFEC1 regs_reg_17__2_ ( .D(i_data_Rd[2]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[546]) );
  DFEC1 regs_reg_17__1_ ( .D(i_data_Rd[1]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[545]) );
  DFEC1 regs_reg_17__0_ ( .D(i_data_Rd[0]), .E(n266), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[544]) );
  DFEC1 regs_reg_16__31_ ( .D(i_data_Rd[31]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[543]) );
  DFEC1 regs_reg_16__30_ ( .D(i_data_Rd[30]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[542]) );
  DFEC1 regs_reg_16__29_ ( .D(i_data_Rd[29]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[541]) );
  DFEC1 regs_reg_16__28_ ( .D(i_data_Rd[28]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[540]) );
  DFEC1 regs_reg_16__27_ ( .D(i_data_Rd[27]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[539]) );
  DFEC1 regs_reg_16__26_ ( .D(i_data_Rd[26]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[538]) );
  DFEC1 regs_reg_16__25_ ( .D(i_data_Rd[25]), .E(n13), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[537]) );
  DFEC1 regs_reg_16__24_ ( .D(i_data_Rd[24]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[536]) );
  DFEC1 regs_reg_16__23_ ( .D(i_data_Rd[23]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[535]) );
  DFEC1 regs_reg_16__22_ ( .D(i_data_Rd[22]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[534]) );
  DFEC1 regs_reg_16__21_ ( .D(i_data_Rd[21]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[533]) );
  DFEC1 regs_reg_16__20_ ( .D(i_data_Rd[20]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[532]) );
  DFEC1 regs_reg_16__19_ ( .D(i_data_Rd[19]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[531]) );
  DFEC1 regs_reg_16__18_ ( .D(i_data_Rd[18]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[530]) );
  DFEC1 regs_reg_16__17_ ( .D(i_data_Rd[17]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[529]) );
  DFEC1 regs_reg_16__16_ ( .D(i_data_Rd[16]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[528]) );
  DFEC1 regs_reg_16__15_ ( .D(i_data_Rd[15]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[527]) );
  DFEC1 regs_reg_16__14_ ( .D(i_data_Rd[14]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[526]) );
  DFEC1 regs_reg_16__13_ ( .D(i_data_Rd[13]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[525]) );
  DFEC1 regs_reg_16__12_ ( .D(i_data_Rd[12]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[524]) );
  DFEC1 regs_reg_16__11_ ( .D(i_data_Rd[11]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[523]) );
  DFEC1 regs_reg_16__10_ ( .D(i_data_Rd[10]), .E(n267), .C(i_clk), .RN(i_rst_n), .Q(regs[522]) );
  DFEC1 regs_reg_16__9_ ( .D(i_data_Rd[9]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[521]) );
  DFEC1 regs_reg_16__8_ ( .D(i_data_Rd[8]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[520]) );
  DFEC1 regs_reg_16__7_ ( .D(i_data_Rd[7]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[519]) );
  DFEC1 regs_reg_16__6_ ( .D(i_data_Rd[6]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[518]) );
  DFEC1 regs_reg_16__5_ ( .D(i_data_Rd[5]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[517]) );
  DFEC1 regs_reg_16__4_ ( .D(i_data_Rd[4]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[516]) );
  DFEC1 regs_reg_16__3_ ( .D(i_data_Rd[3]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[515]) );
  DFEC1 regs_reg_16__2_ ( .D(i_data_Rd[2]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[514]) );
  DFEC1 regs_reg_16__1_ ( .D(i_data_Rd[1]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[513]) );
  DFEC1 regs_reg_16__0_ ( .D(i_data_Rd[0]), .E(n267), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[512]) );
  DFEC1 regs_reg_15__31_ ( .D(i_data_Rd[31]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[511]) );
  DFEC1 regs_reg_15__30_ ( .D(i_data_Rd[30]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[510]) );
  DFEC1 regs_reg_15__29_ ( .D(i_data_Rd[29]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[509]) );
  DFEC1 regs_reg_15__28_ ( .D(i_data_Rd[28]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[508]) );
  DFEC1 regs_reg_15__27_ ( .D(i_data_Rd[27]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[507]) );
  DFEC1 regs_reg_15__26_ ( .D(i_data_Rd[26]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[506]) );
  DFEC1 regs_reg_15__25_ ( .D(i_data_Rd[25]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[505]) );
  DFEC1 regs_reg_15__24_ ( .D(i_data_Rd[24]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[504]) );
  DFEC1 regs_reg_15__23_ ( .D(i_data_Rd[23]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[503]) );
  DFEC1 regs_reg_15__22_ ( .D(i_data_Rd[22]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[502]) );
  DFEC1 regs_reg_15__21_ ( .D(i_data_Rd[21]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[501]) );
  DFEC1 regs_reg_15__20_ ( .D(i_data_Rd[20]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[500]) );
  DFEC1 regs_reg_15__19_ ( .D(i_data_Rd[19]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[499]) );
  DFEC1 regs_reg_15__18_ ( .D(i_data_Rd[18]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[498]) );
  DFEC1 regs_reg_15__17_ ( .D(i_data_Rd[17]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[497]) );
  DFEC1 regs_reg_15__16_ ( .D(i_data_Rd[16]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[496]) );
  DFEC1 regs_reg_15__15_ ( .D(i_data_Rd[15]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[495]) );
  DFEC1 regs_reg_15__14_ ( .D(i_data_Rd[14]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[494]) );
  DFEC1 regs_reg_15__13_ ( .D(i_data_Rd[13]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[493]) );
  DFEC1 regs_reg_15__12_ ( .D(i_data_Rd[12]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[492]) );
  DFEC1 regs_reg_15__11_ ( .D(i_data_Rd[11]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[491]) );
  DFEC1 regs_reg_15__10_ ( .D(i_data_Rd[10]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[490]) );
  DFEC1 regs_reg_15__9_ ( .D(i_data_Rd[9]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[489]) );
  DFEC1 regs_reg_15__8_ ( .D(i_data_Rd[8]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[488]) );
  DFEC1 regs_reg_15__7_ ( .D(i_data_Rd[7]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[487]) );
  DFEC1 regs_reg_15__6_ ( .D(i_data_Rd[6]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[486]) );
  DFEC1 regs_reg_15__5_ ( .D(i_data_Rd[5]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[485]) );
  DFEC1 regs_reg_15__4_ ( .D(i_data_Rd[4]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[484]) );
  DFEC1 regs_reg_15__3_ ( .D(i_data_Rd[3]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[483]) );
  DFEC1 regs_reg_15__2_ ( .D(i_data_Rd[2]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[482]) );
  DFEC1 regs_reg_15__1_ ( .D(i_data_Rd[1]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[481]) );
  DFEC1 regs_reg_15__0_ ( .D(i_data_Rd[0]), .E(n11), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[480]) );
  DFEC1 regs_reg_14__31_ ( .D(i_data_Rd[31]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[479]) );
  DFEC1 regs_reg_14__30_ ( .D(i_data_Rd[30]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[478]) );
  DFEC1 regs_reg_14__29_ ( .D(i_data_Rd[29]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[477]) );
  DFEC1 regs_reg_14__28_ ( .D(i_data_Rd[28]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[476]) );
  DFEC1 regs_reg_14__27_ ( .D(i_data_Rd[27]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[475]) );
  DFEC1 regs_reg_14__26_ ( .D(i_data_Rd[26]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[474]) );
  DFEC1 regs_reg_14__25_ ( .D(i_data_Rd[25]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[473]) );
  DFEC1 regs_reg_14__24_ ( .D(i_data_Rd[24]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[472]) );
  DFEC1 regs_reg_14__23_ ( .D(i_data_Rd[23]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[471]) );
  DFEC1 regs_reg_14__22_ ( .D(i_data_Rd[22]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[470]) );
  DFEC1 regs_reg_14__21_ ( .D(i_data_Rd[21]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[469]) );
  DFEC1 regs_reg_14__20_ ( .D(i_data_Rd[20]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[468]) );
  DFEC1 regs_reg_14__19_ ( .D(i_data_Rd[19]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[467]) );
  DFEC1 regs_reg_14__18_ ( .D(i_data_Rd[18]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[466]) );
  DFEC1 regs_reg_14__17_ ( .D(i_data_Rd[17]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[465]) );
  DFEC1 regs_reg_14__16_ ( .D(i_data_Rd[16]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[464]) );
  DFEC1 regs_reg_14__15_ ( .D(i_data_Rd[15]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[463]) );
  DFEC1 regs_reg_14__14_ ( .D(i_data_Rd[14]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[462]) );
  DFEC1 regs_reg_14__13_ ( .D(i_data_Rd[13]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[461]) );
  DFEC1 regs_reg_14__12_ ( .D(i_data_Rd[12]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[460]) );
  DFEC1 regs_reg_14__11_ ( .D(i_data_Rd[11]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[459]) );
  DFEC1 regs_reg_14__10_ ( .D(i_data_Rd[10]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[458]) );
  DFEC1 regs_reg_14__9_ ( .D(i_data_Rd[9]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[457]) );
  DFEC1 regs_reg_14__8_ ( .D(i_data_Rd[8]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[456]) );
  DFEC1 regs_reg_14__7_ ( .D(i_data_Rd[7]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[455]) );
  DFEC1 regs_reg_14__6_ ( .D(i_data_Rd[6]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[454]) );
  DFEC1 regs_reg_14__5_ ( .D(i_data_Rd[5]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[453]) );
  DFEC1 regs_reg_14__4_ ( .D(i_data_Rd[4]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[452]) );
  DFEC1 regs_reg_14__3_ ( .D(i_data_Rd[3]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[451]) );
  DFEC1 regs_reg_14__2_ ( .D(i_data_Rd[2]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[450]) );
  DFEC1 regs_reg_14__1_ ( .D(i_data_Rd[1]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[449]) );
  DFEC1 regs_reg_14__0_ ( .D(i_data_Rd[0]), .E(n9), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[448]) );
  DFEC1 regs_reg_13__31_ ( .D(i_data_Rd[31]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[447]) );
  DFEC1 regs_reg_13__30_ ( .D(i_data_Rd[30]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[446]) );
  DFEC1 regs_reg_13__29_ ( .D(i_data_Rd[29]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[445]) );
  DFEC1 regs_reg_13__28_ ( .D(i_data_Rd[28]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[444]) );
  DFEC1 regs_reg_13__27_ ( .D(i_data_Rd[27]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[443]) );
  DFEC1 regs_reg_13__26_ ( .D(i_data_Rd[26]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[442]) );
  DFEC1 regs_reg_13__25_ ( .D(i_data_Rd[25]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[441]) );
  DFEC1 regs_reg_13__24_ ( .D(i_data_Rd[24]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[440]) );
  DFEC1 regs_reg_13__23_ ( .D(i_data_Rd[23]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[439]) );
  DFEC1 regs_reg_13__22_ ( .D(i_data_Rd[22]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[438]) );
  DFEC1 regs_reg_13__21_ ( .D(i_data_Rd[21]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[437]) );
  DFEC1 regs_reg_13__20_ ( .D(i_data_Rd[20]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[436]) );
  DFEC1 regs_reg_13__19_ ( .D(i_data_Rd[19]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[435]) );
  DFEC1 regs_reg_13__18_ ( .D(i_data_Rd[18]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[434]) );
  DFEC1 regs_reg_13__17_ ( .D(i_data_Rd[17]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[433]) );
  DFEC1 regs_reg_13__16_ ( .D(i_data_Rd[16]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[432]) );
  DFEC1 regs_reg_13__15_ ( .D(i_data_Rd[15]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[431]) );
  DFEC1 regs_reg_13__14_ ( .D(i_data_Rd[14]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[430]) );
  DFEC1 regs_reg_13__13_ ( .D(i_data_Rd[13]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[429]) );
  DFEC1 regs_reg_13__12_ ( .D(i_data_Rd[12]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[428]) );
  DFEC1 regs_reg_13__11_ ( .D(i_data_Rd[11]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[427]) );
  DFEC1 regs_reg_13__10_ ( .D(i_data_Rd[10]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[426]) );
  DFEC1 regs_reg_13__9_ ( .D(i_data_Rd[9]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[425]) );
  DFEC1 regs_reg_13__8_ ( .D(i_data_Rd[8]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[424]) );
  DFEC1 regs_reg_13__7_ ( .D(i_data_Rd[7]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[423]) );
  DFEC1 regs_reg_13__6_ ( .D(i_data_Rd[6]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[422]) );
  DFEC1 regs_reg_13__5_ ( .D(i_data_Rd[5]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[421]) );
  DFEC1 regs_reg_13__4_ ( .D(i_data_Rd[4]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[420]) );
  DFEC1 regs_reg_13__3_ ( .D(i_data_Rd[3]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[419]) );
  DFEC1 regs_reg_13__2_ ( .D(i_data_Rd[2]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[418]) );
  DFEC1 regs_reg_13__1_ ( .D(i_data_Rd[1]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[417]) );
  DFEC1 regs_reg_13__0_ ( .D(i_data_Rd[0]), .E(n6), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[416]) );
  DFEC1 regs_reg_12__31_ ( .D(i_data_Rd[31]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[415]) );
  DFEC1 regs_reg_12__30_ ( .D(i_data_Rd[30]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[414]) );
  DFEC1 regs_reg_12__29_ ( .D(i_data_Rd[29]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[413]) );
  DFEC1 regs_reg_12__28_ ( .D(i_data_Rd[28]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[412]) );
  DFEC1 regs_reg_12__27_ ( .D(i_data_Rd[27]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[411]) );
  DFEC1 regs_reg_12__26_ ( .D(i_data_Rd[26]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[410]) );
  DFEC1 regs_reg_12__25_ ( .D(i_data_Rd[25]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[409]) );
  DFEC1 regs_reg_12__24_ ( .D(i_data_Rd[24]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[408]) );
  DFEC1 regs_reg_12__23_ ( .D(i_data_Rd[23]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[407]) );
  DFEC1 regs_reg_12__22_ ( .D(i_data_Rd[22]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[406]) );
  DFEC1 regs_reg_12__21_ ( .D(i_data_Rd[21]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[405]) );
  DFEC1 regs_reg_12__20_ ( .D(i_data_Rd[20]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[404]) );
  DFEC1 regs_reg_12__19_ ( .D(i_data_Rd[19]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[403]) );
  DFEC1 regs_reg_12__18_ ( .D(i_data_Rd[18]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[402]) );
  DFEC1 regs_reg_12__17_ ( .D(i_data_Rd[17]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[401]) );
  DFEC1 regs_reg_12__16_ ( .D(i_data_Rd[16]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[400]) );
  DFEC1 regs_reg_12__15_ ( .D(i_data_Rd[15]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[399]) );
  DFEC1 regs_reg_12__14_ ( .D(i_data_Rd[14]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[398]) );
  DFEC1 regs_reg_12__13_ ( .D(i_data_Rd[13]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[397]) );
  DFEC1 regs_reg_12__12_ ( .D(i_data_Rd[12]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[396]) );
  DFEC1 regs_reg_12__11_ ( .D(i_data_Rd[11]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[395]) );
  DFEC1 regs_reg_12__10_ ( .D(i_data_Rd[10]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[394]) );
  DFEC1 regs_reg_12__9_ ( .D(i_data_Rd[9]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[393]) );
  DFEC1 regs_reg_12__8_ ( .D(i_data_Rd[8]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[392]) );
  DFEC1 regs_reg_12__7_ ( .D(i_data_Rd[7]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[391]) );
  DFEC1 regs_reg_12__6_ ( .D(i_data_Rd[6]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[390]) );
  DFEC1 regs_reg_12__5_ ( .D(i_data_Rd[5]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[389]) );
  DFEC1 regs_reg_12__4_ ( .D(i_data_Rd[4]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[388]) );
  DFEC1 regs_reg_12__3_ ( .D(i_data_Rd[3]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[387]) );
  DFEC1 regs_reg_12__2_ ( .D(i_data_Rd[2]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[386]) );
  DFEC1 regs_reg_12__1_ ( .D(i_data_Rd[1]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[385]) );
  DFEC1 regs_reg_12__0_ ( .D(i_data_Rd[0]), .E(n5), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[384]) );
  DFEC1 regs_reg_11__31_ ( .D(i_data_Rd[31]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[383]) );
  DFEC1 regs_reg_11__30_ ( .D(i_data_Rd[30]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[382]) );
  DFEC1 regs_reg_11__29_ ( .D(i_data_Rd[29]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[381]) );
  DFEC1 regs_reg_11__28_ ( .D(i_data_Rd[28]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[380]) );
  DFEC1 regs_reg_11__27_ ( .D(i_data_Rd[27]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[379]) );
  DFEC1 regs_reg_11__26_ ( .D(i_data_Rd[26]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[378]) );
  DFEC1 regs_reg_11__25_ ( .D(i_data_Rd[25]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[377]) );
  DFEC1 regs_reg_11__24_ ( .D(i_data_Rd[24]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[376]) );
  DFEC1 regs_reg_11__23_ ( .D(i_data_Rd[23]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[375]) );
  DFEC1 regs_reg_11__22_ ( .D(i_data_Rd[22]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[374]) );
  DFEC1 regs_reg_11__21_ ( .D(i_data_Rd[21]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[373]) );
  DFEC1 regs_reg_11__20_ ( .D(i_data_Rd[20]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[372]) );
  DFEC1 regs_reg_11__19_ ( .D(i_data_Rd[19]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[371]) );
  DFEC1 regs_reg_11__18_ ( .D(i_data_Rd[18]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[370]) );
  DFEC1 regs_reg_11__17_ ( .D(i_data_Rd[17]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[369]) );
  DFEC1 regs_reg_11__16_ ( .D(i_data_Rd[16]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[368]) );
  DFEC1 regs_reg_11__15_ ( .D(i_data_Rd[15]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[367]) );
  DFEC1 regs_reg_11__14_ ( .D(i_data_Rd[14]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[366]) );
  DFEC1 regs_reg_11__13_ ( .D(i_data_Rd[13]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[365]) );
  DFEC1 regs_reg_11__12_ ( .D(i_data_Rd[12]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[364]) );
  DFEC1 regs_reg_11__11_ ( .D(i_data_Rd[11]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[363]) );
  DFEC1 regs_reg_11__10_ ( .D(i_data_Rd[10]), .E(n248), .C(i_clk), .RN(i_rst_n), .Q(regs[362]) );
  DFEC1 regs_reg_11__9_ ( .D(i_data_Rd[9]), .E(n248), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[361]) );
  DFEC1 regs_reg_11__8_ ( .D(i_data_Rd[8]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[360]) );
  DFEC1 regs_reg_11__7_ ( .D(i_data_Rd[7]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[359]) );
  DFEC1 regs_reg_11__6_ ( .D(i_data_Rd[6]), .E(n248), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[358]) );
  DFEC1 regs_reg_11__5_ ( .D(i_data_Rd[5]), .E(n248), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[357]) );
  DFEC1 regs_reg_11__4_ ( .D(i_data_Rd[4]), .E(n248), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[356]) );
  DFEC1 regs_reg_11__3_ ( .D(i_data_Rd[3]), .E(n248), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[355]) );
  DFEC1 regs_reg_11__2_ ( .D(i_data_Rd[2]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[354]) );
  DFEC1 regs_reg_11__1_ ( .D(i_data_Rd[1]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[353]) );
  DFEC1 regs_reg_11__0_ ( .D(i_data_Rd[0]), .E(n44), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[352]) );
  DFEC1 regs_reg_10__31_ ( .D(i_data_Rd[31]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[351]) );
  DFEC1 regs_reg_10__30_ ( .D(i_data_Rd[30]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[350]) );
  DFEC1 regs_reg_10__29_ ( .D(i_data_Rd[29]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[349]) );
  DFEC1 regs_reg_10__28_ ( .D(i_data_Rd[28]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[348]) );
  DFEC1 regs_reg_10__27_ ( .D(i_data_Rd[27]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[347]) );
  DFEC1 regs_reg_10__26_ ( .D(i_data_Rd[26]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[346]) );
  DFEC1 regs_reg_10__25_ ( .D(i_data_Rd[25]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[345]) );
  DFEC1 regs_reg_10__24_ ( .D(i_data_Rd[24]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[344]) );
  DFEC1 regs_reg_10__23_ ( .D(i_data_Rd[23]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[343]) );
  DFEC1 regs_reg_10__22_ ( .D(i_data_Rd[22]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[342]) );
  DFEC1 regs_reg_10__21_ ( .D(i_data_Rd[21]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[341]) );
  DFEC1 regs_reg_10__20_ ( .D(i_data_Rd[20]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[340]) );
  DFEC1 regs_reg_10__19_ ( .D(i_data_Rd[19]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[339]) );
  DFEC1 regs_reg_10__18_ ( .D(i_data_Rd[18]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[338]) );
  DFEC1 regs_reg_10__17_ ( .D(i_data_Rd[17]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[337]) );
  DFEC1 regs_reg_10__16_ ( .D(i_data_Rd[16]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[336]) );
  DFEC1 regs_reg_10__15_ ( .D(i_data_Rd[15]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[335]) );
  DFEC1 regs_reg_10__14_ ( .D(i_data_Rd[14]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[334]) );
  DFEC1 regs_reg_10__13_ ( .D(i_data_Rd[13]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[333]) );
  DFEC1 regs_reg_10__12_ ( .D(i_data_Rd[12]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[332]) );
  DFEC1 regs_reg_10__11_ ( .D(i_data_Rd[11]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[331]) );
  DFEC1 regs_reg_10__10_ ( .D(i_data_Rd[10]), .E(n249), .C(i_clk), .RN(i_rst_n), .Q(regs[330]) );
  DFEC1 regs_reg_10__9_ ( .D(i_data_Rd[9]), .E(n249), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[329]) );
  DFEC1 regs_reg_10__8_ ( .D(i_data_Rd[8]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[328]) );
  DFEC1 regs_reg_10__7_ ( .D(i_data_Rd[7]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[327]) );
  DFEC1 regs_reg_10__6_ ( .D(i_data_Rd[6]), .E(n249), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[326]) );
  DFEC1 regs_reg_10__5_ ( .D(i_data_Rd[5]), .E(n249), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[325]) );
  DFEC1 regs_reg_10__4_ ( .D(i_data_Rd[4]), .E(n249), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[324]) );
  DFEC1 regs_reg_10__3_ ( .D(i_data_Rd[3]), .E(n249), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[323]) );
  DFEC1 regs_reg_10__2_ ( .D(i_data_Rd[2]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[322]) );
  DFEC1 regs_reg_10__1_ ( .D(i_data_Rd[1]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[321]) );
  DFEC1 regs_reg_10__0_ ( .D(i_data_Rd[0]), .E(n43), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[320]) );
  DFEC1 regs_reg_9__31_ ( .D(i_data_Rd[31]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[319]) );
  DFEC1 regs_reg_9__30_ ( .D(i_data_Rd[30]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[318]) );
  DFEC1 regs_reg_9__29_ ( .D(i_data_Rd[29]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[317]) );
  DFEC1 regs_reg_9__28_ ( .D(i_data_Rd[28]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[316]) );
  DFEC1 regs_reg_9__27_ ( .D(i_data_Rd[27]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[315]) );
  DFEC1 regs_reg_9__26_ ( .D(i_data_Rd[26]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[314]) );
  DFEC1 regs_reg_9__25_ ( .D(i_data_Rd[25]), .E(n42), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[313]) );
  DFEC1 regs_reg_9__24_ ( .D(i_data_Rd[24]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[312]) );
  DFEC1 regs_reg_9__23_ ( .D(i_data_Rd[23]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[311]) );
  DFEC1 regs_reg_9__22_ ( .D(i_data_Rd[22]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[310]) );
  DFEC1 regs_reg_9__21_ ( .D(i_data_Rd[21]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[309]) );
  DFEC1 regs_reg_9__20_ ( .D(i_data_Rd[20]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[308]) );
  DFEC1 regs_reg_9__19_ ( .D(i_data_Rd[19]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[307]) );
  DFEC1 regs_reg_9__18_ ( .D(i_data_Rd[18]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[306]) );
  DFEC1 regs_reg_9__17_ ( .D(i_data_Rd[17]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[305]) );
  DFEC1 regs_reg_9__16_ ( .D(i_data_Rd[16]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[304]) );
  DFEC1 regs_reg_9__15_ ( .D(i_data_Rd[15]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[303]) );
  DFEC1 regs_reg_9__14_ ( .D(i_data_Rd[14]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[302]) );
  DFEC1 regs_reg_9__13_ ( .D(i_data_Rd[13]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[301]) );
  DFEC1 regs_reg_9__12_ ( .D(i_data_Rd[12]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[300]) );
  DFEC1 regs_reg_9__11_ ( .D(i_data_Rd[11]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[299]) );
  DFEC1 regs_reg_9__10_ ( .D(i_data_Rd[10]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[298]) );
  DFEC1 regs_reg_9__9_ ( .D(i_data_Rd[9]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[297]) );
  DFEC1 regs_reg_9__8_ ( .D(i_data_Rd[8]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[296]) );
  DFEC1 regs_reg_9__7_ ( .D(i_data_Rd[7]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[295]) );
  DFEC1 regs_reg_9__6_ ( .D(i_data_Rd[6]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[294]) );
  DFEC1 regs_reg_9__5_ ( .D(i_data_Rd[5]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[293]) );
  DFEC1 regs_reg_9__4_ ( .D(i_data_Rd[4]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[292]) );
  DFEC1 regs_reg_9__3_ ( .D(i_data_Rd[3]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[291]) );
  DFEC1 regs_reg_9__2_ ( .D(i_data_Rd[2]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[290]) );
  DFEC1 regs_reg_9__1_ ( .D(i_data_Rd[1]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[289]) );
  DFEC1 regs_reg_9__0_ ( .D(i_data_Rd[0]), .E(n250), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[288]) );
  DFEC1 regs_reg_8__31_ ( .D(i_data_Rd[31]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[287]) );
  DFEC1 regs_reg_8__30_ ( .D(i_data_Rd[30]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[286]) );
  DFEC1 regs_reg_8__29_ ( .D(i_data_Rd[29]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[285]) );
  DFEC1 regs_reg_8__28_ ( .D(i_data_Rd[28]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[284]) );
  DFEC1 regs_reg_8__27_ ( .D(i_data_Rd[27]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[283]) );
  DFEC1 regs_reg_8__26_ ( .D(i_data_Rd[26]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[282]) );
  DFEC1 regs_reg_8__25_ ( .D(i_data_Rd[25]), .E(n41), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[281]) );
  DFEC1 regs_reg_8__24_ ( .D(i_data_Rd[24]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[280]) );
  DFEC1 regs_reg_8__23_ ( .D(i_data_Rd[23]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[279]) );
  DFEC1 regs_reg_8__22_ ( .D(i_data_Rd[22]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[278]) );
  DFEC1 regs_reg_8__21_ ( .D(i_data_Rd[21]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[277]) );
  DFEC1 regs_reg_8__20_ ( .D(i_data_Rd[20]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[276]) );
  DFEC1 regs_reg_8__19_ ( .D(i_data_Rd[19]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[275]) );
  DFEC1 regs_reg_8__18_ ( .D(i_data_Rd[18]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[274]) );
  DFEC1 regs_reg_8__17_ ( .D(i_data_Rd[17]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[273]) );
  DFEC1 regs_reg_8__16_ ( .D(i_data_Rd[16]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[272]) );
  DFEC1 regs_reg_8__15_ ( .D(i_data_Rd[15]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[271]) );
  DFEC1 regs_reg_8__14_ ( .D(i_data_Rd[14]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[270]) );
  DFEC1 regs_reg_8__13_ ( .D(i_data_Rd[13]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[269]) );
  DFEC1 regs_reg_8__12_ ( .D(i_data_Rd[12]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[268]) );
  DFEC1 regs_reg_8__11_ ( .D(i_data_Rd[11]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[267]) );
  DFEC1 regs_reg_8__10_ ( .D(i_data_Rd[10]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[266]) );
  DFEC1 regs_reg_8__9_ ( .D(i_data_Rd[9]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[265]) );
  DFEC1 regs_reg_8__8_ ( .D(i_data_Rd[8]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[264]) );
  DFEC1 regs_reg_8__7_ ( .D(i_data_Rd[7]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[263]) );
  DFEC1 regs_reg_8__6_ ( .D(i_data_Rd[6]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[262]) );
  DFEC1 regs_reg_8__5_ ( .D(i_data_Rd[5]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[261]) );
  DFEC1 regs_reg_8__4_ ( .D(i_data_Rd[4]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[260]) );
  DFEC1 regs_reg_8__3_ ( .D(i_data_Rd[3]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[259]) );
  DFEC1 regs_reg_8__2_ ( .D(i_data_Rd[2]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[258]) );
  DFEC1 regs_reg_8__1_ ( .D(i_data_Rd[1]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[257]) );
  DFEC1 regs_reg_8__0_ ( .D(i_data_Rd[0]), .E(n251), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[256]) );
  DFEC1 regs_reg_7__31_ ( .D(i_data_Rd[31]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[255]) );
  DFEC1 regs_reg_7__30_ ( .D(i_data_Rd[30]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[254]) );
  DFEC1 regs_reg_7__29_ ( .D(i_data_Rd[29]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[253]) );
  DFEC1 regs_reg_7__28_ ( .D(i_data_Rd[28]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[252]) );
  DFEC1 regs_reg_7__27_ ( .D(i_data_Rd[27]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[251]) );
  DFEC1 regs_reg_7__26_ ( .D(i_data_Rd[26]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[250]) );
  DFEC1 regs_reg_7__25_ ( .D(i_data_Rd[25]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[249]) );
  DFEC1 regs_reg_7__24_ ( .D(i_data_Rd[24]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[248]) );
  DFEC1 regs_reg_7__23_ ( .D(i_data_Rd[23]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[247]) );
  DFEC1 regs_reg_7__22_ ( .D(i_data_Rd[22]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[246]) );
  DFEC1 regs_reg_7__21_ ( .D(i_data_Rd[21]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[245]) );
  DFEC1 regs_reg_7__20_ ( .D(i_data_Rd[20]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[244]) );
  DFEC1 regs_reg_7__19_ ( .D(i_data_Rd[19]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[243]) );
  DFEC1 regs_reg_7__18_ ( .D(i_data_Rd[18]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[242]) );
  DFEC1 regs_reg_7__17_ ( .D(i_data_Rd[17]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[241]) );
  DFEC1 regs_reg_7__16_ ( .D(i_data_Rd[16]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[240]) );
  DFEC1 regs_reg_7__15_ ( .D(i_data_Rd[15]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[239]) );
  DFEC1 regs_reg_7__14_ ( .D(i_data_Rd[14]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[238]) );
  DFEC1 regs_reg_7__13_ ( .D(i_data_Rd[13]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[237]) );
  DFEC1 regs_reg_7__12_ ( .D(i_data_Rd[12]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[236]) );
  DFEC1 regs_reg_7__11_ ( .D(i_data_Rd[11]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[235]) );
  DFEC1 regs_reg_7__10_ ( .D(i_data_Rd[10]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[234]) );
  DFEC1 regs_reg_7__9_ ( .D(i_data_Rd[9]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[233]) );
  DFEC1 regs_reg_7__8_ ( .D(i_data_Rd[8]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[232]) );
  DFEC1 regs_reg_7__7_ ( .D(i_data_Rd[7]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[231]) );
  DFEC1 regs_reg_7__6_ ( .D(i_data_Rd[6]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[230]) );
  DFEC1 regs_reg_7__5_ ( .D(i_data_Rd[5]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[229]) );
  DFEC1 regs_reg_7__4_ ( .D(i_data_Rd[4]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[228]) );
  DFEC1 regs_reg_7__3_ ( .D(i_data_Rd[3]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[227]) );
  DFEC1 regs_reg_7__2_ ( .D(i_data_Rd[2]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[226]) );
  DFEC1 regs_reg_7__1_ ( .D(i_data_Rd[1]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[225]) );
  DFEC1 regs_reg_7__0_ ( .D(i_data_Rd[0]), .E(n40), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[224]) );
  DFEC1 regs_reg_6__31_ ( .D(i_data_Rd[31]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[223]) );
  DFEC1 regs_reg_6__30_ ( .D(i_data_Rd[30]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[222]) );
  DFEC1 regs_reg_6__29_ ( .D(i_data_Rd[29]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[221]) );
  DFEC1 regs_reg_6__28_ ( .D(i_data_Rd[28]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[220]) );
  DFEC1 regs_reg_6__27_ ( .D(i_data_Rd[27]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[219]) );
  DFEC1 regs_reg_6__26_ ( .D(i_data_Rd[26]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[218]) );
  DFEC1 regs_reg_6__25_ ( .D(i_data_Rd[25]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[217]) );
  DFEC1 regs_reg_6__24_ ( .D(i_data_Rd[24]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[216]) );
  DFEC1 regs_reg_6__23_ ( .D(i_data_Rd[23]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[215]) );
  DFEC1 regs_reg_6__22_ ( .D(i_data_Rd[22]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[214]) );
  DFEC1 regs_reg_6__21_ ( .D(i_data_Rd[21]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[213]) );
  DFEC1 regs_reg_6__20_ ( .D(i_data_Rd[20]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[212]) );
  DFEC1 regs_reg_6__19_ ( .D(i_data_Rd[19]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[211]) );
  DFEC1 regs_reg_6__18_ ( .D(i_data_Rd[18]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[210]) );
  DFEC1 regs_reg_6__17_ ( .D(i_data_Rd[17]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[209]) );
  DFEC1 regs_reg_6__16_ ( .D(i_data_Rd[16]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[208]) );
  DFEC1 regs_reg_6__15_ ( .D(i_data_Rd[15]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[207]) );
  DFEC1 regs_reg_6__14_ ( .D(i_data_Rd[14]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[206]) );
  DFEC1 regs_reg_6__13_ ( .D(i_data_Rd[13]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[205]) );
  DFEC1 regs_reg_6__12_ ( .D(i_data_Rd[12]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[204]) );
  DFEC1 regs_reg_6__11_ ( .D(i_data_Rd[11]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[203]) );
  DFEC1 regs_reg_6__10_ ( .D(i_data_Rd[10]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[202]) );
  DFEC1 regs_reg_6__9_ ( .D(i_data_Rd[9]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[201]) );
  DFEC1 regs_reg_6__8_ ( .D(i_data_Rd[8]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[200]) );
  DFEC1 regs_reg_6__7_ ( .D(i_data_Rd[7]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[199]) );
  DFEC1 regs_reg_6__6_ ( .D(i_data_Rd[6]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[198]) );
  DFEC1 regs_reg_6__5_ ( .D(i_data_Rd[5]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[197]) );
  DFEC1 regs_reg_6__4_ ( .D(i_data_Rd[4]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[196]) );
  DFEC1 regs_reg_6__3_ ( .D(i_data_Rd[3]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[195]) );
  DFEC1 regs_reg_6__2_ ( .D(i_data_Rd[2]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[194]) );
  DFEC1 regs_reg_6__1_ ( .D(i_data_Rd[1]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[193]) );
  DFEC1 regs_reg_6__0_ ( .D(i_data_Rd[0]), .E(n39), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[192]) );
  DFEC1 regs_reg_5__31_ ( .D(i_data_Rd[31]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[191]) );
  DFEC1 regs_reg_5__30_ ( .D(i_data_Rd[30]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[190]) );
  DFEC1 regs_reg_5__29_ ( .D(i_data_Rd[29]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[189]) );
  DFEC1 regs_reg_5__28_ ( .D(i_data_Rd[28]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[188]) );
  DFEC1 regs_reg_5__27_ ( .D(i_data_Rd[27]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[187]) );
  DFEC1 regs_reg_5__26_ ( .D(i_data_Rd[26]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[186]) );
  DFEC1 regs_reg_5__25_ ( .D(i_data_Rd[25]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[185]) );
  DFEC1 regs_reg_5__24_ ( .D(i_data_Rd[24]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[184]) );
  DFEC1 regs_reg_5__23_ ( .D(i_data_Rd[23]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[183]) );
  DFEC1 regs_reg_5__22_ ( .D(i_data_Rd[22]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[182]) );
  DFEC1 regs_reg_5__21_ ( .D(i_data_Rd[21]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[181]) );
  DFEC1 regs_reg_5__20_ ( .D(i_data_Rd[20]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[180]) );
  DFEC1 regs_reg_5__19_ ( .D(i_data_Rd[19]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[179]) );
  DFEC1 regs_reg_5__18_ ( .D(i_data_Rd[18]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[178]) );
  DFEC1 regs_reg_5__17_ ( .D(i_data_Rd[17]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[177]) );
  DFEC1 regs_reg_5__16_ ( .D(i_data_Rd[16]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[176]) );
  DFEC1 regs_reg_5__15_ ( .D(i_data_Rd[15]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[175]) );
  DFEC1 regs_reg_5__14_ ( .D(i_data_Rd[14]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[174]) );
  DFEC1 regs_reg_5__13_ ( .D(i_data_Rd[13]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[173]) );
  DFEC1 regs_reg_5__12_ ( .D(i_data_Rd[12]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[172]) );
  DFEC1 regs_reg_5__11_ ( .D(i_data_Rd[11]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[171]) );
  DFEC1 regs_reg_5__10_ ( .D(i_data_Rd[10]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[170]) );
  DFEC1 regs_reg_5__9_ ( .D(i_data_Rd[9]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[169]) );
  DFEC1 regs_reg_5__8_ ( .D(i_data_Rd[8]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[168]) );
  DFEC1 regs_reg_5__7_ ( .D(i_data_Rd[7]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[167]) );
  DFEC1 regs_reg_5__6_ ( .D(i_data_Rd[6]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[166]) );
  DFEC1 regs_reg_5__5_ ( .D(i_data_Rd[5]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[165]) );
  DFEC1 regs_reg_5__4_ ( .D(i_data_Rd[4]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[164]) );
  DFEC1 regs_reg_5__3_ ( .D(i_data_Rd[3]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[163]) );
  DFEC1 regs_reg_5__2_ ( .D(i_data_Rd[2]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[162]) );
  DFEC1 regs_reg_5__1_ ( .D(i_data_Rd[1]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[161]) );
  DFEC1 regs_reg_5__0_ ( .D(i_data_Rd[0]), .E(n38), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[160]) );
  DFEC1 regs_reg_4__31_ ( .D(i_data_Rd[31]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[159]) );
  DFEC1 regs_reg_4__30_ ( .D(i_data_Rd[30]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[158]) );
  DFEC1 regs_reg_4__29_ ( .D(i_data_Rd[29]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[157]) );
  DFEC1 regs_reg_4__28_ ( .D(i_data_Rd[28]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[156]) );
  DFEC1 regs_reg_4__27_ ( .D(i_data_Rd[27]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[155]) );
  DFEC1 regs_reg_4__26_ ( .D(i_data_Rd[26]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[154]) );
  DFEC1 regs_reg_4__25_ ( .D(i_data_Rd[25]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[153]) );
  DFEC1 regs_reg_4__24_ ( .D(i_data_Rd[24]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[152]) );
  DFEC1 regs_reg_4__23_ ( .D(i_data_Rd[23]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[151]) );
  DFEC1 regs_reg_4__22_ ( .D(i_data_Rd[22]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[150]) );
  DFEC1 regs_reg_4__21_ ( .D(i_data_Rd[21]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[149]) );
  DFEC1 regs_reg_4__20_ ( .D(i_data_Rd[20]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[148]) );
  DFEC1 regs_reg_4__19_ ( .D(i_data_Rd[19]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[147]) );
  DFEC1 regs_reg_4__18_ ( .D(i_data_Rd[18]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[146]) );
  DFEC1 regs_reg_4__17_ ( .D(i_data_Rd[17]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[145]) );
  DFEC1 regs_reg_4__16_ ( .D(i_data_Rd[16]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[144]) );
  DFEC1 regs_reg_4__15_ ( .D(i_data_Rd[15]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[143]) );
  DFEC1 regs_reg_4__14_ ( .D(i_data_Rd[14]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[142]) );
  DFEC1 regs_reg_4__13_ ( .D(i_data_Rd[13]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[141]) );
  DFEC1 regs_reg_4__12_ ( .D(i_data_Rd[12]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[140]) );
  DFEC1 regs_reg_4__11_ ( .D(i_data_Rd[11]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[139]) );
  DFEC1 regs_reg_4__10_ ( .D(i_data_Rd[10]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[138]) );
  DFEC1 regs_reg_4__9_ ( .D(i_data_Rd[9]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[137]) );
  DFEC1 regs_reg_4__8_ ( .D(i_data_Rd[8]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[136]) );
  DFEC1 regs_reg_4__7_ ( .D(i_data_Rd[7]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[135]) );
  DFEC1 regs_reg_4__6_ ( .D(i_data_Rd[6]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[134]) );
  DFEC1 regs_reg_4__5_ ( .D(i_data_Rd[5]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[133]) );
  DFEC1 regs_reg_4__4_ ( .D(i_data_Rd[4]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[132]) );
  DFEC1 regs_reg_4__3_ ( .D(i_data_Rd[3]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[131]) );
  DFEC1 regs_reg_4__2_ ( .D(i_data_Rd[2]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[130]) );
  DFEC1 regs_reg_4__1_ ( .D(i_data_Rd[1]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[129]) );
  DFEC1 regs_reg_4__0_ ( .D(i_data_Rd[0]), .E(n37), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[128]) );
  DFEC1 regs_reg_3__31_ ( .D(i_data_Rd[31]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[127]) );
  DFEC1 regs_reg_3__30_ ( .D(i_data_Rd[30]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[126]) );
  DFEC1 regs_reg_3__29_ ( .D(i_data_Rd[29]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[125]) );
  DFEC1 regs_reg_3__28_ ( .D(i_data_Rd[28]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[124]) );
  DFEC1 regs_reg_3__27_ ( .D(i_data_Rd[27]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[123]) );
  DFEC1 regs_reg_3__26_ ( .D(i_data_Rd[26]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[122]) );
  DFEC1 regs_reg_3__25_ ( .D(i_data_Rd[25]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[121]) );
  DFEC1 regs_reg_3__24_ ( .D(i_data_Rd[24]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[120]) );
  DFEC1 regs_reg_3__23_ ( .D(i_data_Rd[23]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[119]) );
  DFEC1 regs_reg_3__22_ ( .D(i_data_Rd[22]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[118]) );
  DFEC1 regs_reg_3__21_ ( .D(i_data_Rd[21]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[117]) );
  DFEC1 regs_reg_3__20_ ( .D(i_data_Rd[20]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[116]) );
  DFEC1 regs_reg_3__19_ ( .D(i_data_Rd[19]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[115]) );
  DFEC1 regs_reg_3__18_ ( .D(i_data_Rd[18]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[114]) );
  DFEC1 regs_reg_3__17_ ( .D(i_data_Rd[17]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[113]) );
  DFEC1 regs_reg_3__16_ ( .D(i_data_Rd[16]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[112]) );
  DFEC1 regs_reg_3__15_ ( .D(i_data_Rd[15]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[111]) );
  DFEC1 regs_reg_3__14_ ( .D(i_data_Rd[14]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[110]) );
  DFEC1 regs_reg_3__13_ ( .D(i_data_Rd[13]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[109]) );
  DFEC1 regs_reg_3__12_ ( .D(i_data_Rd[12]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[108]) );
  DFEC1 regs_reg_3__11_ ( .D(i_data_Rd[11]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[107]) );
  DFEC1 regs_reg_3__10_ ( .D(i_data_Rd[10]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[106]) );
  DFEC1 regs_reg_3__9_ ( .D(i_data_Rd[9]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[105]) );
  DFEC1 regs_reg_3__8_ ( .D(i_data_Rd[8]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[104]) );
  DFEC1 regs_reg_3__7_ ( .D(i_data_Rd[7]), .E(n36), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[103]) );
  DFEC1 regs_reg_3__6_ ( .D(i_data_Rd[6]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[102]) );
  DFEC1 regs_reg_3__5_ ( .D(i_data_Rd[5]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[101]) );
  DFEC1 regs_reg_3__4_ ( .D(i_data_Rd[4]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[100]) );
  DFEC1 regs_reg_3__3_ ( .D(i_data_Rd[3]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[99]) );
  DFEC1 regs_reg_3__2_ ( .D(i_data_Rd[2]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[98]) );
  DFEC1 regs_reg_3__1_ ( .D(i_data_Rd[1]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[97]) );
  DFEC1 regs_reg_3__0_ ( .D(i_data_Rd[0]), .E(n252), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[96]) );
  DFEC1 regs_reg_2__31_ ( .D(i_data_Rd[31]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[95]) );
  DFEC1 regs_reg_2__30_ ( .D(i_data_Rd[30]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[94]) );
  DFEC1 regs_reg_2__29_ ( .D(i_data_Rd[29]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[93]) );
  DFEC1 regs_reg_2__28_ ( .D(i_data_Rd[28]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[92]) );
  DFEC1 regs_reg_2__27_ ( .D(i_data_Rd[27]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[91]) );
  DFEC1 regs_reg_2__26_ ( .D(i_data_Rd[26]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[90]) );
  DFEC1 regs_reg_2__25_ ( .D(i_data_Rd[25]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[89]) );
  DFEC1 regs_reg_2__24_ ( .D(i_data_Rd[24]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[88]) );
  DFEC1 regs_reg_2__23_ ( .D(i_data_Rd[23]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[87]) );
  DFEC1 regs_reg_2__22_ ( .D(i_data_Rd[22]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[86]) );
  DFEC1 regs_reg_2__21_ ( .D(i_data_Rd[21]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[85]) );
  DFEC1 regs_reg_2__20_ ( .D(i_data_Rd[20]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[84]) );
  DFEC1 regs_reg_2__19_ ( .D(i_data_Rd[19]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[83]) );
  DFEC1 regs_reg_2__18_ ( .D(i_data_Rd[18]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[82]) );
  DFEC1 regs_reg_2__17_ ( .D(i_data_Rd[17]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[81]) );
  DFEC1 regs_reg_2__16_ ( .D(i_data_Rd[16]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[80]) );
  DFEC1 regs_reg_2__15_ ( .D(i_data_Rd[15]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[79]) );
  DFEC1 regs_reg_2__14_ ( .D(i_data_Rd[14]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[78]) );
  DFEC1 regs_reg_2__13_ ( .D(i_data_Rd[13]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[77]) );
  DFEC1 regs_reg_2__12_ ( .D(i_data_Rd[12]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[76]) );
  DFEC1 regs_reg_2__11_ ( .D(i_data_Rd[11]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[75]) );
  DFEC1 regs_reg_2__10_ ( .D(i_data_Rd[10]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[74]) );
  DFEC1 regs_reg_2__9_ ( .D(i_data_Rd[9]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[73]) );
  DFEC1 regs_reg_2__8_ ( .D(i_data_Rd[8]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[72]) );
  DFEC1 regs_reg_2__7_ ( .D(i_data_Rd[7]), .E(n35), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[71]) );
  DFEC1 regs_reg_2__6_ ( .D(i_data_Rd[6]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[70]) );
  DFEC1 regs_reg_2__5_ ( .D(i_data_Rd[5]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[69]) );
  DFEC1 regs_reg_2__4_ ( .D(i_data_Rd[4]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[68]) );
  DFEC1 regs_reg_2__3_ ( .D(i_data_Rd[3]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[67]) );
  DFEC1 regs_reg_2__2_ ( .D(i_data_Rd[2]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[66]) );
  DFEC1 regs_reg_2__1_ ( .D(i_data_Rd[1]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[65]) );
  DFEC1 regs_reg_2__0_ ( .D(i_data_Rd[0]), .E(n253), .C(i_clk), .RN(i_rst_n), 
        .Q(regs[64]) );
  DFEC1 regs_reg_1__31_ ( .D(n165), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[63]) );
  DFEC1 regs_reg_1__30_ ( .D(n196), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[62]) );
  DFEC1 regs_reg_1__29_ ( .D(n195), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[61]) );
  DFEC1 regs_reg_1__28_ ( .D(n194), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[60]) );
  DFEC1 regs_reg_1__27_ ( .D(n193), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[59]) );
  DFEC1 regs_reg_1__26_ ( .D(n192), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[58]) );
  DFEC1 regs_reg_1__25_ ( .D(n191), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[57]) );
  DFEC1 regs_reg_1__24_ ( .D(n190), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[56]) );
  DFEC1 regs_reg_1__23_ ( .D(n189), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[55]) );
  DFEC1 regs_reg_1__22_ ( .D(n188), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[54]) );
  DFEC1 regs_reg_1__21_ ( .D(n187), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[53]) );
  DFEC1 regs_reg_1__20_ ( .D(n186), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[52]) );
  DFEC1 regs_reg_1__19_ ( .D(n185), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[51]) );
  DFEC1 regs_reg_1__18_ ( .D(n184), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[50]) );
  DFEC1 regs_reg_1__17_ ( .D(n183), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[49]) );
  DFEC1 regs_reg_1__16_ ( .D(n182), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[48]) );
  DFEC1 regs_reg_1__15_ ( .D(n181), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[47]) );
  DFEC1 regs_reg_1__14_ ( .D(n180), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[46]) );
  DFEC1 regs_reg_1__13_ ( .D(n179), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[45]) );
  DFEC1 regs_reg_1__12_ ( .D(n178), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[44]) );
  DFEC1 regs_reg_1__11_ ( .D(n177), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[43]) );
  DFEC1 regs_reg_1__10_ ( .D(n176), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[42]) );
  DFEC1 regs_reg_1__9_ ( .D(n175), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[41]) );
  DFEC1 regs_reg_1__8_ ( .D(n174), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[40]) );
  DFEC1 regs_reg_1__7_ ( .D(n173), .E(n34), .C(i_clk), .RN(i_rst_n), .Q(
        regs[39]) );
  DFEC1 regs_reg_1__6_ ( .D(n172), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[38]) );
  DFEC1 regs_reg_1__5_ ( .D(n171), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[37]) );
  DFEC1 regs_reg_1__4_ ( .D(n170), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[36]) );
  DFEC1 regs_reg_1__3_ ( .D(n169), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[35]) );
  DFEC1 regs_reg_1__2_ ( .D(n168), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[34]) );
  DFEC1 regs_reg_1__1_ ( .D(n167), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[33]) );
  DFEC1 regs_reg_1__0_ ( .D(n166), .E(n254), .C(i_clk), .RN(i_rst_n), .Q(
        regs[32]) );
  DFEC1 regs_reg_0__31_ ( .D(n165), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[31]) );
  DFEC1 regs_reg_0__30_ ( .D(n196), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[30]) );
  DFEC1 regs_reg_0__29_ ( .D(n195), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[29]) );
  DFEC1 regs_reg_0__28_ ( .D(n194), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[28]) );
  DFEC1 regs_reg_0__27_ ( .D(n193), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[27]) );
  DFEC1 regs_reg_0__26_ ( .D(n192), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[26]) );
  DFEC1 regs_reg_0__25_ ( .D(n191), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[25]) );
  DFEC1 regs_reg_0__24_ ( .D(n190), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[24]) );
  DFEC1 regs_reg_0__23_ ( .D(n189), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[23]) );
  DFEC1 regs_reg_0__22_ ( .D(n188), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[22]) );
  DFEC1 regs_reg_0__21_ ( .D(n187), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[21]) );
  DFEC1 regs_reg_0__20_ ( .D(n186), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[20]) );
  DFEC1 regs_reg_0__19_ ( .D(n185), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[19]) );
  DFEC1 regs_reg_0__18_ ( .D(n184), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[18]) );
  DFEC1 regs_reg_0__17_ ( .D(n183), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[17]) );
  DFEC1 regs_reg_0__16_ ( .D(n182), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[16]) );
  DFEC1 regs_reg_0__15_ ( .D(n181), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[15]) );
  DFEC1 regs_reg_0__14_ ( .D(n180), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[14]) );
  DFEC1 regs_reg_0__13_ ( .D(n179), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[13]) );
  DFEC1 regs_reg_0__12_ ( .D(n178), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[12]) );
  DFEC1 regs_reg_0__11_ ( .D(n177), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[11]) );
  DFEC1 regs_reg_0__10_ ( .D(n176), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[10]) );
  DFEC1 regs_reg_0__9_ ( .D(n175), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[9]) );
  DFEC1 regs_reg_0__8_ ( .D(n174), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[8]) );
  DFEC1 regs_reg_0__7_ ( .D(n173), .E(n32), .C(i_clk), .RN(i_rst_n), .Q(
        regs[7]) );
  DFEC1 regs_reg_0__6_ ( .D(n172), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[6]) );
  DFEC1 regs_reg_0__5_ ( .D(n171), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[5]) );
  DFEC1 regs_reg_0__4_ ( .D(n170), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[4]) );
  DFEC1 regs_reg_0__3_ ( .D(n169), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[3]) );
  DFEC1 regs_reg_0__2_ ( .D(n168), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[2]) );
  DFEC1 regs_reg_0__1_ ( .D(n167), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[1]) );
  DFEC1 regs_reg_0__0_ ( .D(n166), .E(n255), .C(i_clk), .RN(i_rst_n), .Q(
        regs[0]) );
  MUX21 regs_reg_31__31__U4 ( .A(regs[1023]), .B(i_data_Rd[31]), .S(n31), .Q(
        n197) );
  DFC1 regs_reg_31__31_ ( .D(n197), .C(i_clk), .RN(i_rst_n), .Q(regs[1023]) );
  BUF6 U2 ( .A(n1565), .Q(n246) );
  BUF6 U3 ( .A(n1563), .Q(n245) );
  BUF6 U4 ( .A(n973), .Q(n201) );
  BUF6 U5 ( .A(n976), .Q(n206) );
  BUF8 U6 ( .A(n979), .Q(n244) );
  BUF8 U7 ( .A(n978), .Q(n232) );
  AOI220 U8 ( .A(n1562), .B(regs[673]), .C(n245), .D(regs[737]), .Q(n1) );
  AOI220 U9 ( .A(n1565), .B(regs[705]), .C(n200), .D(regs[641]), .Q(n2) );
  AOI220 U10 ( .A(n1566), .B(regs[545]), .C(n247), .D(regs[609]), .Q(n3) );
  AOI220 U11 ( .A(n203), .B(regs[577]), .C(n204), .D(regs[513]), .Q(n4) );
  NAND40 U12 ( .A(n1), .B(n2), .C(n3), .D(n4), .Q(n7) );
  AOI220 U13 ( .A(n199), .B(regs[161]), .C(n245), .D(regs[225]), .Q(n8) );
  AOI220 U14 ( .A(n200), .B(regs[129]), .C(n246), .D(regs[193]), .Q(n10) );
  AOI220 U15 ( .A(n205), .B(regs[33]), .C(n247), .D(regs[97]), .Q(n12) );
  AOI220 U16 ( .A(n203), .B(regs[65]), .C(n204), .D(regs[1]), .Q(n14) );
  NAND40 U17 ( .A(n8), .B(n10), .C(n12), .D(n14), .Q(n19) );
  AOI220 U18 ( .A(n1577), .B(n7), .C(n1575), .D(n19), .Q(n24) );
  AOI220 U19 ( .A(n199), .B(regs[929]), .C(n245), .D(regs[993]), .Q(n33) );
  AOI220 U20 ( .A(n200), .B(regs[897]), .C(n246), .D(regs[961]), .Q(n45) );
  AOI220 U21 ( .A(n205), .B(regs[801]), .C(n247), .D(regs[865]), .Q(n46) );
  AOI220 U22 ( .A(n1569), .B(regs[833]), .C(n204), .D(regs[769]), .Q(n47) );
  NAND40 U23 ( .A(n33), .B(n45), .C(n46), .D(n47), .Q(n48) );
  AOI220 U24 ( .A(n199), .B(regs[417]), .C(n245), .D(regs[481]), .Q(n49) );
  AOI220 U25 ( .A(n200), .B(regs[385]), .C(n246), .D(regs[449]), .Q(n50) );
  AOI220 U26 ( .A(n205), .B(regs[289]), .C(n247), .D(regs[353]), .Q(n51) );
  AOI220 U27 ( .A(n203), .B(regs[321]), .C(n204), .D(regs[257]), .Q(n52) );
  NAND40 U28 ( .A(n49), .B(n50), .C(n51), .D(n52), .Q(n53) );
  AOI220 U29 ( .A(n1557), .B(n48), .C(n1555), .D(n53), .Q(n54) );
  NAND20 U30 ( .A(n24), .B(n54), .Q(o_data_Rs[1]) );
  AOI220 U31 ( .A(n199), .B(regs[693]), .C(n245), .D(regs[757]), .Q(n55) );
  AOI220 U32 ( .A(n200), .B(regs[661]), .C(n246), .D(regs[725]), .Q(n56) );
  AOI220 U33 ( .A(n205), .B(regs[565]), .C(n247), .D(regs[629]), .Q(n57) );
  AOI220 U34 ( .A(n203), .B(regs[597]), .C(n1568), .D(regs[533]), .Q(n58) );
  NAND40 U35 ( .A(n55), .B(n56), .C(n57), .D(n58), .Q(n59) );
  AOI220 U36 ( .A(n199), .B(regs[181]), .C(n245), .D(regs[245]), .Q(n60) );
  AOI220 U37 ( .A(n200), .B(regs[149]), .C(n246), .D(regs[213]), .Q(n61) );
  AOI220 U38 ( .A(n205), .B(regs[53]), .C(n247), .D(regs[117]), .Q(n62) );
  AOI220 U39 ( .A(n203), .B(regs[85]), .C(n1568), .D(regs[21]), .Q(n63) );
  NAND40 U40 ( .A(n60), .B(n61), .C(n62), .D(n63), .Q(n64) );
  AOI220 U41 ( .A(n1577), .B(n59), .C(n1575), .D(n64), .Q(n65) );
  AOI220 U42 ( .A(n199), .B(regs[949]), .C(n245), .D(regs[1013]), .Q(n66) );
  AOI220 U43 ( .A(n200), .B(regs[917]), .C(n246), .D(regs[981]), .Q(n67) );
  AOI220 U44 ( .A(n205), .B(regs[821]), .C(n247), .D(regs[885]), .Q(n68) );
  AOI220 U45 ( .A(n203), .B(regs[853]), .C(n1568), .D(regs[789]), .Q(n69) );
  NAND40 U46 ( .A(n66), .B(n67), .C(n68), .D(n69), .Q(n70) );
  AOI220 U47 ( .A(n199), .B(regs[437]), .C(n245), .D(regs[501]), .Q(n71) );
  AOI220 U48 ( .A(n200), .B(regs[405]), .C(n246), .D(regs[469]), .Q(n72) );
  AOI220 U49 ( .A(n205), .B(regs[309]), .C(n247), .D(regs[373]), .Q(n73) );
  AOI220 U50 ( .A(n203), .B(regs[341]), .C(n1568), .D(regs[277]), .Q(n74) );
  NAND40 U51 ( .A(n71), .B(n72), .C(n73), .D(n74), .Q(n75) );
  AOI220 U52 ( .A(n1557), .B(n70), .C(n1555), .D(n75), .Q(n76) );
  NAND20 U53 ( .A(n65), .B(n76), .Q(o_data_Rs[21]) );
  AOI220 U54 ( .A(n199), .B(regs[686]), .C(n245), .D(regs[750]), .Q(n77) );
  AOI220 U55 ( .A(n200), .B(regs[654]), .C(n246), .D(regs[718]), .Q(n78) );
  AOI220 U56 ( .A(n205), .B(regs[558]), .C(n247), .D(regs[622]), .Q(n79) );
  AOI220 U57 ( .A(n203), .B(regs[590]), .C(n204), .D(regs[526]), .Q(n80) );
  NAND40 U58 ( .A(n77), .B(n78), .C(n79), .D(n80), .Q(n81) );
  AOI220 U59 ( .A(n199), .B(regs[174]), .C(n245), .D(regs[238]), .Q(n82) );
  AOI220 U60 ( .A(n200), .B(regs[142]), .C(n246), .D(regs[206]), .Q(n83) );
  AOI220 U61 ( .A(n205), .B(regs[46]), .C(n247), .D(regs[110]), .Q(n84) );
  AOI220 U62 ( .A(n1568), .B(regs[14]), .C(n203), .D(regs[78]), .Q(n85) );
  NAND40 U63 ( .A(n82), .B(n83), .C(n84), .D(n85), .Q(n86) );
  AOI220 U64 ( .A(n1577), .B(n81), .C(n1575), .D(n86), .Q(n87) );
  AOI220 U65 ( .A(n199), .B(regs[942]), .C(n245), .D(regs[1006]), .Q(n88) );
  AOI220 U66 ( .A(n200), .B(regs[910]), .C(n246), .D(regs[974]), .Q(n89) );
  AOI220 U67 ( .A(n205), .B(regs[814]), .C(n247), .D(regs[878]), .Q(n90) );
  AOI220 U68 ( .A(n1568), .B(regs[782]), .C(n203), .D(regs[846]), .Q(n91) );
  NAND40 U69 ( .A(n88), .B(n89), .C(n90), .D(n91), .Q(n92) );
  AOI220 U70 ( .A(n199), .B(regs[430]), .C(n245), .D(regs[494]), .Q(n93) );
  AOI220 U71 ( .A(n200), .B(regs[398]), .C(n246), .D(regs[462]), .Q(n94) );
  AOI220 U72 ( .A(n205), .B(regs[302]), .C(n247), .D(regs[366]), .Q(n95) );
  AOI220 U73 ( .A(n1568), .B(regs[270]), .C(n203), .D(regs[334]), .Q(n96) );
  NAND40 U74 ( .A(n93), .B(n94), .C(n95), .D(n96), .Q(n97) );
  AOI220 U75 ( .A(n1557), .B(n92), .C(n1555), .D(n97), .Q(n98) );
  NAND20 U76 ( .A(n87), .B(n98), .Q(o_data_Rs[14]) );
  AOI220 U77 ( .A(n199), .B(regs[682]), .C(n245), .D(regs[746]), .Q(n99) );
  AOI220 U78 ( .A(n200), .B(regs[650]), .C(n246), .D(regs[714]), .Q(n100) );
  AOI220 U79 ( .A(n205), .B(regs[554]), .C(n247), .D(regs[618]), .Q(n101) );
  AOI220 U80 ( .A(n203), .B(regs[586]), .C(n204), .D(regs[522]), .Q(n102) );
  NAND40 U81 ( .A(n99), .B(n100), .C(n101), .D(n102), .Q(n103) );
  AOI220 U82 ( .A(n199), .B(regs[170]), .C(n245), .D(regs[234]), .Q(n104) );
  AOI220 U83 ( .A(n200), .B(regs[138]), .C(n246), .D(regs[202]), .Q(n105) );
  AOI220 U84 ( .A(n205), .B(regs[42]), .C(n247), .D(regs[106]), .Q(n106) );
  AOI220 U85 ( .A(n1568), .B(regs[10]), .C(n203), .D(regs[74]), .Q(n107) );
  NAND40 U86 ( .A(n104), .B(n105), .C(n106), .D(n107), .Q(n108) );
  AOI220 U87 ( .A(n1577), .B(n103), .C(n1575), .D(n108), .Q(n109) );
  AOI220 U88 ( .A(n199), .B(regs[938]), .C(n245), .D(regs[1002]), .Q(n110) );
  AOI220 U89 ( .A(n200), .B(regs[906]), .C(n246), .D(regs[970]), .Q(n111) );
  AOI220 U90 ( .A(n205), .B(regs[810]), .C(n247), .D(regs[874]), .Q(n112) );
  AOI220 U91 ( .A(n203), .B(regs[842]), .C(n204), .D(regs[778]), .Q(n113) );
  NAND40 U92 ( .A(n110), .B(n111), .C(n112), .D(n113), .Q(n114) );
  AOI220 U93 ( .A(n199), .B(regs[426]), .C(n245), .D(regs[490]), .Q(n115) );
  AOI220 U94 ( .A(n200), .B(regs[394]), .C(n246), .D(regs[458]), .Q(n116) );
  AOI220 U95 ( .A(n205), .B(regs[298]), .C(n247), .D(regs[362]), .Q(n117) );
  AOI220 U96 ( .A(n203), .B(regs[330]), .C(n204), .D(regs[266]), .Q(n118) );
  NAND40 U97 ( .A(n115), .B(n116), .C(n117), .D(n118), .Q(n119) );
  AOI220 U98 ( .A(n1557), .B(n114), .C(n1555), .D(n119), .Q(n120) );
  NAND20 U99 ( .A(n109), .B(n120), .Q(o_data_Rs[10]) );
  AOI220 U100 ( .A(n199), .B(regs[675]), .C(n245), .D(regs[739]), .Q(n121) );
  AOI220 U101 ( .A(n200), .B(regs[643]), .C(n246), .D(regs[707]), .Q(n122) );
  AOI220 U102 ( .A(n205), .B(regs[547]), .C(n247), .D(regs[611]), .Q(n123) );
  AOI220 U103 ( .A(n203), .B(regs[579]), .C(n204), .D(regs[515]), .Q(n124) );
  NAND40 U104 ( .A(n121), .B(n122), .C(n123), .D(n124), .Q(n125) );
  AOI220 U105 ( .A(n199), .B(regs[163]), .C(n245), .D(regs[227]), .Q(n126) );
  AOI220 U106 ( .A(n200), .B(regs[131]), .C(n246), .D(regs[195]), .Q(n127) );
  AOI220 U107 ( .A(n205), .B(regs[35]), .C(n247), .D(regs[99]), .Q(n128) );
  AOI220 U108 ( .A(n203), .B(regs[67]), .C(n204), .D(regs[3]), .Q(n129) );
  NAND40 U109 ( .A(n126), .B(n127), .C(n128), .D(n129), .Q(n130) );
  AOI220 U110 ( .A(n1577), .B(n125), .C(n1575), .D(n130), .Q(n131) );
  AOI220 U111 ( .A(n199), .B(regs[931]), .C(n245), .D(regs[995]), .Q(n132) );
  AOI220 U112 ( .A(n200), .B(regs[899]), .C(n246), .D(regs[963]), .Q(n133) );
  AOI220 U113 ( .A(n205), .B(regs[803]), .C(n247), .D(regs[867]), .Q(n134) );
  AOI220 U114 ( .A(n203), .B(regs[835]), .C(n204), .D(regs[771]), .Q(n135) );
  NAND40 U115 ( .A(n132), .B(n133), .C(n134), .D(n135), .Q(n136) );
  AOI220 U116 ( .A(n199), .B(regs[419]), .C(n245), .D(regs[483]), .Q(n137) );
  AOI220 U117 ( .A(n200), .B(regs[387]), .C(n246), .D(regs[451]), .Q(n138) );
  AOI220 U118 ( .A(n205), .B(regs[291]), .C(n247), .D(regs[355]), .Q(n139) );
  AOI220 U119 ( .A(n203), .B(regs[323]), .C(n204), .D(regs[259]), .Q(n140) );
  NAND40 U120 ( .A(n137), .B(n138), .C(n139), .D(n140), .Q(n141) );
  AOI220 U121 ( .A(n1557), .B(n136), .C(n1555), .D(n141), .Q(n142) );
  NAND20 U122 ( .A(n131), .B(n142), .Q(o_data_Rs[3]) );
  AOI220 U123 ( .A(n199), .B(regs[672]), .C(n245), .D(regs[736]), .Q(n143) );
  AOI220 U124 ( .A(n1564), .B(regs[640]), .C(n246), .D(regs[704]), .Q(n144) );
  AOI220 U125 ( .A(n1566), .B(regs[544]), .C(n247), .D(regs[608]), .Q(n145) );
  AOI220 U126 ( .A(n1568), .B(regs[512]), .C(n1569), .D(regs[576]), .Q(n146)
         );
  NAND40 U127 ( .A(n143), .B(n144), .C(n145), .D(n146), .Q(n147) );
  AOI220 U128 ( .A(n199), .B(regs[160]), .C(n245), .D(regs[224]), .Q(n148) );
  AOI220 U129 ( .A(n200), .B(regs[128]), .C(n246), .D(regs[192]), .Q(n149) );
  AOI220 U130 ( .A(n205), .B(regs[32]), .C(n247), .D(regs[96]), .Q(n150) );
  AOI220 U131 ( .A(n203), .B(regs[64]), .C(n204), .D(regs[0]), .Q(n151) );
  NAND40 U132 ( .A(n148), .B(n149), .C(n150), .D(n151), .Q(n152) );
  AOI220 U133 ( .A(n1577), .B(n147), .C(n1575), .D(n152), .Q(n153) );
  AOI220 U134 ( .A(n199), .B(regs[928]), .C(n245), .D(regs[992]), .Q(n154) );
  AOI220 U135 ( .A(n200), .B(regs[896]), .C(n246), .D(regs[960]), .Q(n155) );
  AOI220 U136 ( .A(n205), .B(regs[800]), .C(n247), .D(regs[864]), .Q(n156) );
  AOI220 U137 ( .A(n203), .B(regs[832]), .C(n204), .D(regs[768]), .Q(n157) );
  NAND40 U138 ( .A(n154), .B(n155), .C(n156), .D(n157), .Q(n158) );
  AOI220 U139 ( .A(n199), .B(regs[416]), .C(n245), .D(regs[480]), .Q(n159) );
  AOI220 U140 ( .A(n200), .B(regs[384]), .C(n246), .D(regs[448]), .Q(n160) );
  AOI220 U141 ( .A(n205), .B(regs[288]), .C(n247), .D(regs[352]), .Q(n161) );
  AOI220 U142 ( .A(n203), .B(regs[320]), .C(n204), .D(regs[256]), .Q(n162) );
  NAND40 U143 ( .A(n159), .B(n160), .C(n161), .D(n162), .Q(n163) );
  AOI220 U144 ( .A(n1557), .B(n158), .C(n1555), .D(n163), .Q(n164) );
  NAND20 U145 ( .A(n153), .B(n164), .Q(o_data_Rs[0]) );
  BUF6 U146 ( .A(n1566), .Q(n205) );
  BUF6 U147 ( .A(n977), .Q(n243) );
  BUF6 U148 ( .A(n972), .Q(n198) );
  BUF2 U149 ( .A(i_data_Rd[31]), .Q(n165) );
  BUF2 U150 ( .A(i_data_Rd[0]), .Q(n166) );
  BUF2 U151 ( .A(i_data_Rd[1]), .Q(n167) );
  BUF2 U152 ( .A(i_data_Rd[2]), .Q(n168) );
  BUF2 U153 ( .A(i_data_Rd[3]), .Q(n169) );
  BUF2 U154 ( .A(i_data_Rd[4]), .Q(n170) );
  BUF2 U155 ( .A(i_data_Rd[5]), .Q(n171) );
  BUF2 U156 ( .A(i_data_Rd[6]), .Q(n172) );
  BUF2 U157 ( .A(i_data_Rd[7]), .Q(n173) );
  BUF2 U158 ( .A(i_data_Rd[8]), .Q(n174) );
  BUF2 U159 ( .A(i_data_Rd[9]), .Q(n175) );
  BUF2 U160 ( .A(i_data_Rd[10]), .Q(n176) );
  BUF2 U161 ( .A(i_data_Rd[11]), .Q(n177) );
  BUF2 U162 ( .A(i_data_Rd[12]), .Q(n178) );
  BUF2 U163 ( .A(i_data_Rd[13]), .Q(n179) );
  BUF2 U164 ( .A(i_data_Rd[14]), .Q(n180) );
  BUF2 U165 ( .A(i_data_Rd[15]), .Q(n181) );
  BUF2 U166 ( .A(i_data_Rd[16]), .Q(n182) );
  BUF2 U167 ( .A(i_data_Rd[17]), .Q(n183) );
  BUF2 U168 ( .A(i_data_Rd[18]), .Q(n184) );
  BUF2 U169 ( .A(i_data_Rd[19]), .Q(n185) );
  BUF2 U170 ( .A(i_data_Rd[20]), .Q(n186) );
  BUF2 U171 ( .A(i_data_Rd[21]), .Q(n187) );
  BUF2 U172 ( .A(i_data_Rd[22]), .Q(n188) );
  BUF2 U173 ( .A(i_data_Rd[23]), .Q(n189) );
  BUF2 U174 ( .A(i_data_Rd[24]), .Q(n190) );
  BUF2 U175 ( .A(i_data_Rd[25]), .Q(n191) );
  BUF2 U176 ( .A(i_data_Rd[26]), .Q(n192) );
  BUF2 U177 ( .A(i_data_Rd[27]), .Q(n193) );
  BUF2 U178 ( .A(i_data_Rd[28]), .Q(n194) );
  BUF2 U179 ( .A(i_data_Rd[29]), .Q(n195) );
  BUF2 U180 ( .A(i_data_Rd[30]), .Q(n196) );
  AOI220 U181 ( .A(n967), .B(n679), .C(n965), .D(n678), .Q(n691) );
  AOI221 U182 ( .A(n967), .B(n767), .C(n965), .D(n766), .Q(n779) );
  NAND21 U183 ( .A(n989), .B(n988), .Q(o_data_Rt[31]) );
  AOI221 U184 ( .A(n967), .B(n921), .C(n965), .D(n920), .Q(n933) );
  AOI220 U185 ( .A(n967), .B(n327), .C(n965), .D(n326), .Q(n339) );
  AOI220 U186 ( .A(n967), .B(n371), .C(n965), .D(n370), .Q(n383) );
  AOI220 U187 ( .A(n967), .B(n415), .C(n965), .D(n414), .Q(n427) );
  AOI221 U188 ( .A(n1557), .B(n1203), .C(n1555), .D(n1202), .Q(n1215) );
  AOI220 U189 ( .A(n987), .B(n469), .C(n985), .D(n468), .Q(n470) );
  AOI220 U190 ( .A(n987), .B(n909), .C(n985), .D(n908), .Q(n910) );
  AOI220 U191 ( .A(n967), .B(n525), .C(n965), .D(n524), .Q(n537) );
  AOI220 U192 ( .A(n967), .B(n943), .C(n965), .D(n942), .Q(n955) );
  AOI220 U193 ( .A(n967), .B(n393), .C(n965), .D(n392), .Q(n405) );
  AOI220 U194 ( .A(n967), .B(n899), .C(n965), .D(n898), .Q(n911) );
  AOI220 U195 ( .A(n967), .B(n745), .C(n965), .D(n744), .Q(n757) );
  AOI220 U196 ( .A(n967), .B(n547), .C(n965), .D(n546), .Q(n559) );
  AOI220 U197 ( .A(n987), .B(n986), .C(n985), .D(n984), .Q(n988) );
  AOI220 U198 ( .A(n243), .B(regs[627]), .C(n206), .D(regs[563]), .Q(n703) );
  AOI221 U199 ( .A(n243), .B(regs[891]), .C(n206), .D(regs[827]), .Q(n869) );
  AOI221 U200 ( .A(n243), .B(regs[622]), .C(n206), .D(regs[558]), .Q(n593) );
  AOI220 U201 ( .A(n243), .B(regs[369]), .C(n206), .D(regs[305]), .Q(n653) );
  AOI221 U202 ( .A(n243), .B(regs[374]), .C(n206), .D(regs[310]), .Q(n763) );
  AOI220 U203 ( .A(n243), .B(regs[371]), .C(n206), .D(regs[307]), .Q(n697) );
  AOI221 U204 ( .A(n977), .B(regs[120]), .C(n206), .D(regs[56]), .Q(n817) );
  AOI221 U205 ( .A(n243), .B(regs[381]), .C(n206), .D(regs[317]), .Q(n917) );
  AOI221 U206 ( .A(n977), .B(regs[365]), .C(n206), .D(regs[301]), .Q(n565) );
  AOI220 U207 ( .A(n243), .B(regs[370]), .C(n206), .D(regs[306]), .Q(n675) );
  AOI220 U208 ( .A(n243), .B(regs[626]), .C(n206), .D(regs[562]), .Q(n681) );
  AOI220 U209 ( .A(n243), .B(regs[884]), .C(n206), .D(regs[820]), .Q(n715) );
  AOI220 U210 ( .A(n243), .B(regs[114]), .C(n206), .D(regs[50]), .Q(n685) );
  AOI221 U211 ( .A(n243), .B(regs[614]), .C(n206), .D(regs[550]), .Q(n417) );
  AOI220 U212 ( .A(n243), .B(regs[115]), .C(n206), .D(regs[51]), .Q(n707) );
  AOI221 U213 ( .A(n243), .B(regs[632]), .C(n206), .D(regs[568]), .Q(n813) );
  AOI221 U214 ( .A(n977), .B(regs[880]), .C(n206), .D(regs[816]), .Q(n627) );
  AOI221 U215 ( .A(n243), .B(regs[889]), .C(n206), .D(regs[825]), .Q(n825) );
  AOI221 U216 ( .A(n977), .B(regs[623]), .C(n206), .D(regs[559]), .Q(n615) );
  AOI221 U217 ( .A(n243), .B(regs[864]), .C(n206), .D(regs[800]), .Q(n273) );
  AOI220 U218 ( .A(n201), .B(regs[253]), .C(n198), .D(regs[189]), .Q(n929) );
  AOI220 U219 ( .A(regs[987]), .B(n246), .C(regs[923]), .D(n200), .Q(n1460) );
  AOI220 U220 ( .A(n201), .B(regs[756]), .C(n198), .D(regs[692]), .Q(n727) );
  AOI220 U221 ( .A(n201), .B(regs[233]), .C(n198), .D(regs[169]), .Q(n489) );
  AOI220 U222 ( .A(regs[1020]), .B(n245), .C(regs[956]), .D(n199), .Q(n1483)
         );
  AOI220 U223 ( .A(n201), .B(regs[765]), .C(n198), .D(regs[701]), .Q(n925) );
  AOI221 U224 ( .A(n244), .B(regs[80]), .C(n232), .D(regs[16]), .Q(n640) );
  AOI220 U225 ( .A(n201), .B(regs[754]), .C(n198), .D(regs[690]), .Q(n683) );
  AOI221 U226 ( .A(n975), .B(regs[477]), .C(n202), .D(regs[413]), .Q(n918) );
  AOI220 U227 ( .A(n241), .B(regs[711]), .C(n202), .D(regs[647]), .Q(n440) );
  AOI220 U228 ( .A(n201), .B(regs[1012]), .C(n198), .D(regs[948]), .Q(n717) );
  AOI220 U229 ( .A(regs[764]), .B(n245), .C(regs[700]), .D(n199), .Q(n1493) );
  AOI220 U230 ( .A(n241), .B(regs[199]), .C(n202), .D(regs[135]), .Q(n444) );
  AOI220 U231 ( .A(regs[732]), .B(n246), .C(regs[668]), .D(n200), .Q(n1492) );
  AOI220 U232 ( .A(n201), .B(regs[745]), .C(n198), .D(regs[681]), .Q(n485) );
  AOI220 U233 ( .A(n201), .B(regs[498]), .C(n198), .D(regs[434]), .Q(n677) );
  AOI220 U234 ( .A(n243), .B(regs[617]), .C(n206), .D(regs[553]), .Q(n483) );
  AOI220 U235 ( .A(regs[220]), .B(n246), .C(regs[156]), .D(n200), .Q(n1496) );
  AOI220 U236 ( .A(n201), .B(regs[1016]), .C(n198), .D(regs[952]), .Q(n805) );
  AOI220 U237 ( .A(n201), .B(regs[1011]), .C(n198), .D(regs[947]), .Q(n695) );
  AOI221 U238 ( .A(n244), .B(regs[323]), .C(n232), .D(regs[259]), .Q(n344) );
  AOI220 U239 ( .A(n243), .B(regs[881]), .C(n206), .D(regs[817]), .Q(n649) );
  AOI220 U240 ( .A(n201), .B(regs[243]), .C(n972), .D(regs[179]), .Q(n709) );
  AOI221 U241 ( .A(n244), .B(regs[835]), .C(n232), .D(regs[771]), .Q(n340) );
  AOI220 U242 ( .A(regs[477]), .B(n246), .C(regs[413]), .D(n200), .Q(n1508) );
  AOI220 U243 ( .A(n201), .B(regs[232]), .C(n198), .D(regs[168]), .Q(n467) );
  AOI220 U244 ( .A(regs[733]), .B(n246), .C(regs[669]), .D(n200), .Q(n1514) );
  AOI220 U245 ( .A(n243), .B(regs[100]), .C(n206), .D(regs[36]), .Q(n377) );
  AOI220 U246 ( .A(n201), .B(regs[499]), .C(n198), .D(regs[435]), .Q(n699) );
  AOI221 U247 ( .A(n201), .B(regs[753]), .C(n198), .D(regs[689]), .Q(n661) );
  AOI220 U248 ( .A(n243), .B(regs[356]), .C(n206), .D(regs[292]), .Q(n367) );
  AOI220 U249 ( .A(n201), .B(regs[755]), .C(n198), .D(regs[691]), .Q(n705) );
  AOI220 U250 ( .A(n201), .B(regs[508]), .C(n198), .D(regs[444]), .Q(n897) );
  AOI220 U251 ( .A(regs[765]), .B(n245), .C(regs[701]), .D(n199), .Q(n1515) );
  AOI220 U252 ( .A(n243), .B(regs[105]), .C(n206), .D(regs[41]), .Q(n487) );
  AOI221 U253 ( .A(n201), .B(regs[742]), .C(n198), .D(regs[678]), .Q(n419) );
  AOI220 U254 ( .A(regs[763]), .B(n245), .C(regs[699]), .D(n199), .Q(n1471) );
  AOI221 U255 ( .A(n244), .B(regs[578]), .C(n232), .D(regs[514]), .Q(n328) );
  AOI220 U256 ( .A(regs[731]), .B(n246), .C(regs[667]), .D(n200), .Q(n1470) );
  AOI220 U257 ( .A(regs[989]), .B(n246), .C(regs[925]), .D(n200), .Q(n1504) );
  AOI220 U258 ( .A(n201), .B(regs[1022]), .C(n198), .D(regs[958]), .Q(n937) );
  AOI220 U259 ( .A(n243), .B(regs[104]), .C(n206), .D(regs[40]), .Q(n465) );
  AOI220 U260 ( .A(n201), .B(regs[1000]), .C(n198), .D(regs[936]), .Q(n453) );
  AOI220 U261 ( .A(n241), .B(regs[968]), .C(n202), .D(regs[904]), .Q(n452) );
  AOI220 U262 ( .A(regs[982]), .B(n246), .C(regs[918]), .D(n200), .Q(n1350) );
  AOI220 U263 ( .A(n243), .B(regs[872]), .C(n206), .D(regs[808]), .Q(n451) );
  AOI221 U264 ( .A(n244), .B(regs[857]), .C(n232), .D(regs[793]), .Q(n824) );
  AOI220 U265 ( .A(regs[712]), .B(n246), .C(regs[648]), .D(n200), .Q(n1118) );
  AOI220 U266 ( .A(regs[744]), .B(n245), .C(regs[680]), .D(n199), .Q(n1119) );
  AOI221 U267 ( .A(n244), .B(regs[855]), .C(n232), .D(regs[791]), .Q(n780) );
  AOI220 U268 ( .A(regs[488]), .B(n245), .C(regs[424]), .D(n199), .Q(n1113) );
  AOI220 U269 ( .A(n201), .B(regs[503]), .C(n198), .D(regs[439]), .Q(n787) );
  AOI220 U270 ( .A(regs[968]), .B(n246), .C(regs[904]), .D(n200), .Q(n1108) );
  AOI220 U271 ( .A(n201), .B(regs[1017]), .C(n198), .D(regs[953]), .Q(n827) );
  AOI221 U272 ( .A(n244), .B(regs[343]), .C(n232), .D(regs[279]), .Q(n784) );
  AOI220 U273 ( .A(n201), .B(regs[759]), .C(n198), .D(regs[695]), .Q(n793) );
  AOI220 U274 ( .A(n243), .B(regs[107]), .C(n206), .D(regs[43]), .Q(n531) );
  AOI221 U275 ( .A(n244), .B(regs[333]), .C(n232), .D(regs[269]), .Q(n564) );
  AOI220 U276 ( .A(regs[223]), .B(n246), .C(regs[159]), .D(n200), .Q(n1572) );
  AOI221 U277 ( .A(n244), .B(regs[599]), .C(n232), .D(regs[535]), .Q(n790) );
  AOI220 U278 ( .A(n201), .B(regs[247]), .C(n972), .D(regs[183]), .Q(n797) );
  AOI220 U279 ( .A(n201), .B(regs[250]), .C(n198), .D(regs[186]), .Q(n863) );
  AOI220 U280 ( .A(n201), .B(regs[1014]), .C(n198), .D(regs[950]), .Q(n761) );
  AOI220 U281 ( .A(n201), .B(regs[504]), .C(n198), .D(regs[440]), .Q(n809) );
  AOI220 U282 ( .A(n201), .B(regs[249]), .C(n198), .D(regs[185]), .Q(n841) );
  AOI221 U283 ( .A(n244), .B(regs[601]), .C(n232), .D(regs[537]), .Q(n834) );
  AOI220 U284 ( .A(regs[741]), .B(n245), .C(regs[677]), .D(n199), .Q(n1053) );
  AOI220 U285 ( .A(n201), .B(regs[760]), .C(n198), .D(regs[696]), .Q(n815) );
  AOI220 U286 ( .A(n201), .B(regs[761]), .C(n972), .D(regs[697]), .Q(n837) );
  AOI221 U287 ( .A(n244), .B(regs[345]), .C(n232), .D(regs[281]), .Q(n828) );
  AOI221 U288 ( .A(n244), .B(regs[600]), .C(n232), .D(regs[536]), .Q(n812) );
  AOI220 U289 ( .A(n201), .B(regs[248]), .C(n198), .D(regs[184]), .Q(n819) );
  AOI220 U290 ( .A(regs[998]), .B(n245), .C(regs[934]), .D(n199), .Q(n1065) );
  AOI220 U291 ( .A(regs[199]), .B(n246), .C(regs[135]), .D(n200), .Q(n1100) );
  AOI220 U292 ( .A(n201), .B(regs[505]), .C(n198), .D(regs[441]), .Q(n831) );
  AOI220 U293 ( .A(n201), .B(regs[1015]), .C(n972), .D(regs[951]), .Q(n783) );
  AOI220 U294 ( .A(n201), .B(regs[246]), .C(n198), .D(regs[182]), .Q(n775) );
  AOI220 U295 ( .A(n201), .B(regs[1018]), .C(n198), .D(regs[954]), .Q(n849) );
  AOI220 U296 ( .A(regs[766]), .B(n245), .C(regs[702]), .D(n199), .Q(n1537) );
  AOI220 U297 ( .A(regs[751]), .B(n245), .C(regs[687]), .D(n199), .Q(n1229) );
  AOI220 U298 ( .A(n201), .B(regs[1013]), .C(n972), .D(regs[949]), .Q(n739) );
  AOI220 U299 ( .A(n241), .B(regs[202]), .C(n202), .D(regs[138]), .Q(n510) );
  AOI220 U300 ( .A(n243), .B(regs[106]), .C(n206), .D(regs[42]), .Q(n509) );
  AOI221 U301 ( .A(n244), .B(regs[591]), .C(n232), .D(regs[527]), .Q(n614) );
  AOI220 U302 ( .A(regs[208]), .B(n246), .C(regs[144]), .D(n200), .Q(n1254) );
  AOI220 U303 ( .A(regs[752]), .B(n245), .C(regs[688]), .D(n199), .Q(n1251) );
  AOI220 U304 ( .A(regs[496]), .B(n245), .C(regs[432]), .D(n199), .Q(n1245) );
  AOI220 U305 ( .A(regs[976]), .B(n246), .C(regs[912]), .D(n200), .Q(n1240) );
  AOI221 U306 ( .A(n244), .B(regs[335]), .C(n232), .D(regs[271]), .Q(n608) );
  AOI220 U307 ( .A(regs[1008]), .B(n245), .C(regs[944]), .D(n199), .Q(n1241)
         );
  AOI220 U308 ( .A(regs[209]), .B(n246), .C(regs[145]), .D(n200), .Q(n1276) );
  AOI220 U309 ( .A(regs[254]), .B(n245), .C(regs[190]), .D(n199), .Q(n1541) );
  AOI220 U310 ( .A(regs[241]), .B(n245), .C(regs[177]), .D(n199), .Q(n1277) );
  AOI220 U311 ( .A(n201), .B(regs[757]), .C(n972), .D(regs[693]), .Q(n749) );
  AOI220 U312 ( .A(regs[497]), .B(n245), .C(regs[433]), .D(n199), .Q(n1267) );
  NOR22 U313 ( .A(n1585), .B(n1582), .Q(n37) );
  AOI220 U314 ( .A(regs[210]), .B(n246), .C(regs[146]), .D(n200), .Q(n1298) );
  AOI220 U315 ( .A(regs[749]), .B(n245), .C(regs[685]), .D(n199), .Q(n1207) );
  AOI220 U316 ( .A(n201), .B(regs[758]), .C(n972), .D(regs[694]), .Q(n771) );
  AOI220 U317 ( .A(n975), .B(regs[474]), .C(n202), .D(regs[410]), .Q(n852) );
  AOI220 U318 ( .A(regs[237]), .B(n245), .C(regs[173]), .D(n199), .Q(n1211) );
  AOI220 U319 ( .A(n201), .B(regs[506]), .C(n198), .D(regs[442]), .Q(n853) );
  AOI221 U320 ( .A(n244), .B(regs[342]), .C(n232), .D(regs[278]), .Q(n762) );
  AOI220 U321 ( .A(n243), .B(regs[366]), .C(n206), .D(regs[302]), .Q(n587) );
  AOI221 U322 ( .A(n201), .B(regs[750]), .C(n198), .D(regs[686]), .Q(n595) );
  AOI220 U323 ( .A(regs[1005]), .B(n245), .C(regs[941]), .D(n199), .Q(n1197)
         );
  AOI221 U324 ( .A(n244), .B(regs[858]), .C(n232), .D(regs[794]), .Q(n846) );
  NOR22 U325 ( .A(n1589), .B(n1582), .Q(n40) );
  AOI221 U326 ( .A(n244), .B(regs[598]), .C(n232), .D(regs[534]), .Q(n768) );
  AOI220 U327 ( .A(regs[990]), .B(n246), .C(regs[926]), .D(n200), .Q(n1526) );
  AOI221 U328 ( .A(n244), .B(regs[346]), .C(n232), .D(regs[282]), .Q(n850) );
  NOR22 U329 ( .A(n1591), .B(n1583), .Q(n29) );
  NOR22 U330 ( .A(n1590), .B(n1583), .Q(n30) );
  BUF6 U331 ( .A(n1569), .Q(n203) );
  BUF6 U332 ( .A(n1567), .Q(n247) );
  BUF8 U333 ( .A(n1564), .Q(n200) );
  BUF12 U334 ( .A(n1562), .Q(n199) );
  NOR22 U335 ( .A(n1589), .B(n1583), .Q(n31) );
  BUF6 U336 ( .A(n974), .Q(n202) );
  NOR22 U337 ( .A(n1585), .B(n1583), .Q(n28) );
  NOR31 U338 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[1]), .C(n990), .Q(n1564) );
  AOI220 U339 ( .A(n967), .B(n459), .C(n965), .D(n458), .Q(n471) );
  AOI220 U340 ( .A(n967), .B(n789), .C(n965), .D(n788), .Q(n801) );
  AOI220 U341 ( .A(n967), .B(n811), .C(n965), .D(n810), .Q(n823) );
  AOI220 U342 ( .A(n967), .B(n966), .C(n965), .D(n964), .Q(n989) );
  AOI220 U343 ( .A(n967), .B(n569), .C(n965), .D(n568), .Q(n581) );
  AOI221 U344 ( .A(n244), .B(regs[337]), .C(n232), .D(regs[273]), .Q(n652) );
  AOI221 U345 ( .A(n244), .B(regs[594]), .C(n232), .D(regs[530]), .Q(n680) );
  AOI221 U346 ( .A(n244), .B(regs[75]), .C(n232), .D(regs[11]), .Q(n530) );
  AOI220 U347 ( .A(n967), .B(n503), .C(n965), .D(n502), .Q(n515) );
  AOI221 U348 ( .A(n244), .B(regs[68]), .C(n232), .D(regs[4]), .Q(n376) );
  AOI220 U349 ( .A(n967), .B(n437), .C(n965), .D(n436), .Q(n449) );
  AOI220 U350 ( .A(n967), .B(n481), .C(n965), .D(n480), .Q(n493) );
  AOI221 U351 ( .A(n244), .B(regs[339]), .C(n232), .D(regs[275]), .Q(n696) );
  AOI221 U352 ( .A(n244), .B(regs[83]), .C(n232), .D(regs[19]), .Q(n706) );
  AOI221 U353 ( .A(n244), .B(regs[86]), .C(n232), .D(regs[22]), .Q(n772) );
  AOI221 U354 ( .A(n244), .B(regs[586]), .C(n232), .D(regs[522]), .Q(n504) );
  AOI221 U355 ( .A(n977), .B(regs[618]), .C(n206), .D(regs[554]), .Q(n505) );
  AOI221 U356 ( .A(n243), .B(regs[633]), .C(n206), .D(regs[569]), .Q(n835) );
  AOI221 U357 ( .A(n244), .B(regs[74]), .C(n232), .D(regs[10]), .Q(n508) );
  AOI221 U358 ( .A(n244), .B(regs[847]), .C(n232), .D(regs[783]), .Q(n604) );
  AOI221 U359 ( .A(n244), .B(regs[592]), .C(n232), .D(regs[528]), .Q(n636) );
  AOI221 U360 ( .A(n244), .B(regs[79]), .C(n232), .D(regs[15]), .Q(n618) );
  AOI221 U361 ( .A(n244), .B(regs[590]), .C(n232), .D(regs[526]), .Q(n592) );
  AOI221 U362 ( .A(n244), .B(regs[848]), .C(n232), .D(regs[784]), .Q(n626) );
  AOI221 U363 ( .A(n244), .B(regs[78]), .C(n232), .D(regs[14]), .Q(n596) );
  AOI221 U364 ( .A(n244), .B(regs[81]), .C(n232), .D(regs[17]), .Q(n662) );
  AOI221 U365 ( .A(n243), .B(regs[621]), .C(n206), .D(regs[557]), .Q(n571) );
  AOI221 U366 ( .A(n244), .B(regs[593]), .C(n232), .D(regs[529]), .Q(n658) );
  AOI221 U367 ( .A(n244), .B(regs[849]), .C(n232), .D(regs[785]), .Q(n648) );
  AOI221 U368 ( .A(n244), .B(regs[844]), .C(n232), .D(regs[780]), .Q(n538) );
  AOI221 U369 ( .A(n244), .B(regs[332]), .C(n232), .D(regs[268]), .Q(n542) );
  AOI221 U370 ( .A(n244), .B(regs[850]), .C(n232), .D(regs[786]), .Q(n670) );
  AOI221 U371 ( .A(n244), .B(regs[843]), .C(n232), .D(regs[779]), .Q(n516) );
  AOI220 U372 ( .A(n243), .B(regs[883]), .C(n206), .D(regs[819]), .Q(n693) );
  AOI221 U373 ( .A(n244), .B(regs[331]), .C(n232), .D(regs[267]), .Q(n520) );
  AOI221 U374 ( .A(n244), .B(regs[596]), .C(n232), .D(regs[532]), .Q(n724) );
  AOI221 U375 ( .A(n244), .B(regs[587]), .C(n232), .D(regs[523]), .Q(n526) );
  AOI221 U376 ( .A(n244), .B(regs[597]), .C(n232), .D(regs[533]), .Q(n746) );
  AOI221 U377 ( .A(n244), .B(regs[325]), .C(n232), .D(regs[261]), .Q(n388) );
  AOI221 U378 ( .A(n244), .B(regs[859]), .C(n232), .D(regs[795]), .Q(n868) );
  AOI221 U379 ( .A(n244), .B(regs[92]), .C(n232), .D(regs[28]), .Q(n904) );
  AOI221 U380 ( .A(n244), .B(regs[604]), .C(n232), .D(regs[540]), .Q(n900) );
  AOI221 U381 ( .A(n244), .B(regs[836]), .C(n232), .D(regs[772]), .Q(n362) );
  AOI221 U382 ( .A(n244), .B(regs[348]), .C(n232), .D(regs[284]), .Q(n894) );
  AOI220 U383 ( .A(n243), .B(regs[637]), .C(n206), .D(regs[573]), .Q(n923) );
  AOI221 U384 ( .A(n244), .B(regs[862]), .C(n232), .D(regs[798]), .Q(n934) );
  AOI221 U385 ( .A(n243), .B(regs[866]), .C(n206), .D(regs[802]), .Q(n319) );
  AOI221 U386 ( .A(n244), .B(regs[834]), .C(n232), .D(regs[770]), .Q(n318) );
  AOI221 U387 ( .A(n243), .B(regs[354]), .C(n206), .D(regs[290]), .Q(n323) );
  AOI221 U388 ( .A(n244), .B(regs[64]), .C(n232), .D(regs[0]), .Q(n288) );
  AOI221 U389 ( .A(n244), .B(regs[322]), .C(n232), .D(regs[258]), .Q(n322) );
  AOI221 U390 ( .A(n243), .B(regs[96]), .C(n206), .D(regs[32]), .Q(n289) );
  AOI221 U391 ( .A(n244), .B(regs[320]), .C(n232), .D(regs[256]), .Q(n277) );
  AOI221 U392 ( .A(n243), .B(regs[352]), .C(n206), .D(regs[288]), .Q(n278) );
  AOI221 U393 ( .A(n244), .B(regs[65]), .C(n232), .D(regs[1]), .Q(n310) );
  AOI221 U394 ( .A(n243), .B(regs[97]), .C(n206), .D(regs[33]), .Q(n311) );
  AOI221 U395 ( .A(n244), .B(regs[577]), .C(n232), .D(regs[513]), .Q(n306) );
  AOI221 U396 ( .A(n243), .B(regs[609]), .C(n206), .D(regs[545]), .Q(n307) );
  AOI221 U397 ( .A(n243), .B(regs[865]), .C(n206), .D(regs[801]), .Q(n297) );
  AOI221 U398 ( .A(n244), .B(regs[321]), .C(n232), .D(regs[257]), .Q(n300) );
  AOI221 U399 ( .A(n243), .B(regs[353]), .C(n206), .D(regs[289]), .Q(n301) );
  AOI221 U400 ( .A(n244), .B(regs[833]), .C(n232), .D(regs[769]), .Q(n296) );
  AOI221 U401 ( .A(n244), .B(regs[90]), .C(n232), .D(regs[26]), .Q(n860) );
  AOI221 U402 ( .A(n243), .B(regs[615]), .C(n206), .D(regs[551]), .Q(n439) );
  AOI220 U403 ( .A(n243), .B(regs[874]), .C(n206), .D(regs[810]), .Q(n495) );
  AOI220 U404 ( .A(n244), .B(regs[842]), .C(n232), .D(regs[778]), .Q(n494) );
  AOI220 U405 ( .A(n244), .B(regs[330]), .C(n232), .D(regs[266]), .Q(n498) );
  AOI221 U406 ( .A(n244), .B(regs[347]), .C(n232), .D(regs[283]), .Q(n872) );
  NOR22 U407 ( .A(n1592), .B(n1591), .Q(n6) );
  AOI220 U408 ( .A(n244), .B(regs[76]), .C(n232), .D(regs[12]), .Q(n552) );
  AOI221 U409 ( .A(n244), .B(regs[344]), .C(n232), .D(regs[280]), .Q(n806) );
  AOI220 U410 ( .A(n244), .B(regs[66]), .C(n232), .D(regs[2]), .Q(n332) );
  AOI220 U411 ( .A(n244), .B(regs[73]), .C(n232), .D(regs[9]), .Q(n486) );
  AOI221 U412 ( .A(n244), .B(regs[832]), .C(n232), .D(regs[768]), .Q(n272) );
  AOI221 U413 ( .A(n244), .B(regs[350]), .C(n232), .D(regs[286]), .Q(n938) );
  AOI221 U414 ( .A(n244), .B(regs[606]), .C(n232), .D(regs[542]), .Q(n944) );
  AOI221 U415 ( .A(n244), .B(regs[94]), .C(n232), .D(regs[30]), .Q(n948) );
  AOI221 U416 ( .A(n244), .B(regs[93]), .C(n232), .D(regs[29]), .Q(n926) );
  AOI220 U417 ( .A(n243), .B(regs[125]), .C(n206), .D(regs[61]), .Q(n927) );
  AOI221 U418 ( .A(n244), .B(regs[861]), .C(n232), .D(regs[797]), .Q(n912) );
  AOI220 U419 ( .A(n244), .B(regs[584]), .C(n232), .D(regs[520]), .Q(n460) );
  AOI221 U420 ( .A(n244), .B(regs[349]), .C(n232), .D(regs[285]), .Q(n916) );
  AOI220 U421 ( .A(n244), .B(regs[72]), .C(n232), .D(regs[8]), .Q(n464) );
  AOI221 U422 ( .A(n244), .B(regs[863]), .C(n232), .D(regs[799]), .Q(n956) );
  AOI221 U423 ( .A(n244), .B(regs[351]), .C(n232), .D(regs[287]), .Q(n960) );
  NOR22 U424 ( .A(n1592), .B(n1585), .Q(n5) );
  AOI220 U425 ( .A(n244), .B(regs[841]), .C(n232), .D(regs[777]), .Q(n472) );
  AOI221 U426 ( .A(n244), .B(regs[607]), .C(n232), .D(regs[543]), .Q(n968) );
  NOR22 U427 ( .A(n1582), .B(n1591), .Q(n38) );
  AOI220 U428 ( .A(n244), .B(regs[329]), .C(n232), .D(regs[265]), .Q(n476) );
  AOI220 U429 ( .A(n243), .B(regs[894]), .C(n206), .D(regs[830]), .Q(n935) );
  AOI220 U430 ( .A(n244), .B(regs[585]), .C(n232), .D(regs[521]), .Q(n482) );
  AOI221 U431 ( .A(n244), .B(regs[88]), .C(n232), .D(regs[24]), .Q(n816) );
  AOI220 U432 ( .A(n243), .B(regs[882]), .C(n206), .D(regs[818]), .Q(n671) );
  AOI220 U433 ( .A(n243), .B(regs[624]), .C(n206), .D(regs[560]), .Q(n637) );
  AOI220 U434 ( .A(n244), .B(regs[324]), .C(n232), .D(regs[260]), .Q(n366) );
  NOR22 U435 ( .A(n1582), .B(n1590), .Q(n39) );
  NOR22 U436 ( .A(n1592), .B(n1589), .Q(n11) );
  AOI220 U437 ( .A(n243), .B(regs[368]), .C(n206), .D(regs[304]), .Q(n631) );
  AOI221 U438 ( .A(n244), .B(regs[91]), .C(n232), .D(regs[27]), .Q(n882) );
  AOI220 U439 ( .A(n244), .B(regs[579]), .C(n232), .D(regs[515]), .Q(n350) );
  AOI221 U440 ( .A(n244), .B(regs[326]), .C(n232), .D(regs[262]), .Q(n410) );
  AOI220 U441 ( .A(n244), .B(regs[67]), .C(n232), .D(regs[3]), .Q(n354) );
  NOR22 U442 ( .A(n1592), .B(n1590), .Q(n9) );
  AOI221 U443 ( .A(n244), .B(regs[89]), .C(n232), .D(regs[25]), .Q(n838) );
  NOR22 U444 ( .A(i_addr_Rt_4_), .B(n276), .Q(n965) );
  NOR22 U445 ( .A(n994), .B(n995), .Q(n1557) );
  NOR22 U446 ( .A(n276), .B(n283), .Q(n967) );
  NOR31 U447 ( .A(i_addr_Rs[1]), .B(i_addr_Rs[2]), .C(n992), .Q(n1566) );
  BUF6 U448 ( .A(n1568), .Q(n204) );
  NOR22 U449 ( .A(i_addr_Rs[3]), .B(i_addr_Rs[4]), .Q(n1575) );
  NOR22 U450 ( .A(i_addr_Rt_3_), .B(i_addr_Rt_4_), .Q(n985) );
  AOI220 U451 ( .A(n241), .B(regs[991]), .C(n974), .D(regs[927]), .Q(n958) );
  AOI220 U452 ( .A(n242), .B(regs[990]), .C(n202), .D(regs[926]), .Q(n936) );
  AOI220 U453 ( .A(n241), .B(regs[479]), .C(n202), .D(regs[415]), .Q(n962) );
  AOI220 U454 ( .A(n975), .B(regs[735]), .C(n974), .D(regs[671]), .Q(n970) );
  AOI220 U455 ( .A(n242), .B(regs[709]), .C(n202), .D(regs[645]), .Q(n396) );
  AOI220 U456 ( .A(regs[873]), .B(n247), .C(regs[809]), .D(n205), .Q(n1129) );
  AOI220 U457 ( .A(n242), .B(regs[965]), .C(n202), .D(regs[901]), .Q(n386) );
  AOI220 U458 ( .A(regs[361]), .B(n247), .C(regs[297]), .D(n205), .Q(n1133) );
  AOI220 U459 ( .A(n241), .B(regs[198]), .C(n202), .D(regs[134]), .Q(n422) );
  AOI220 U460 ( .A(n241), .B(regs[710]), .C(n202), .D(regs[646]), .Q(n418) );
  AOI220 U461 ( .A(regs[617]), .B(n247), .C(regs[553]), .D(n205), .Q(n1139) );
  AOI220 U462 ( .A(n242), .B(regs[454]), .C(n202), .D(regs[390]), .Q(n412) );
  AOI220 U463 ( .A(regs[105]), .B(n247), .C(regs[41]), .D(n205), .Q(n1143) );
  AOI220 U464 ( .A(n242), .B(regs[966]), .C(n202), .D(regs[902]), .Q(n408) );
  AOI220 U465 ( .A(regs[1000]), .B(n245), .C(regs[936]), .D(n199), .Q(n1109)
         );
  AOI220 U466 ( .A(regs[872]), .B(n247), .C(regs[808]), .D(n205), .Q(n1107) );
  AOI220 U467 ( .A(n241), .B(regs[455]), .C(n202), .D(regs[391]), .Q(n434) );
  AOI220 U468 ( .A(regs[456]), .B(n246), .C(regs[392]), .D(n200), .Q(n1112) );
  AOI220 U469 ( .A(regs[360]), .B(n247), .C(regs[296]), .D(n205), .Q(n1111) );
  AOI220 U470 ( .A(n241), .B(regs[967]), .C(n202), .D(regs[903]), .Q(n430) );
  AOI220 U471 ( .A(regs[616]), .B(n247), .C(regs[552]), .D(n205), .Q(n1117) );
  AOI220 U472 ( .A(n242), .B(regs[200]), .C(n202), .D(regs[136]), .Q(n466) );
  AOI220 U473 ( .A(n975), .B(regs[712]), .C(n974), .D(regs[648]), .Q(n462) );
  AOI220 U474 ( .A(regs[104]), .B(n247), .C(regs[40]), .D(n205), .Q(n1121) );
  AOI220 U475 ( .A(n241), .B(regs[456]), .C(n202), .D(regs[392]), .Q(n456) );
  AOI220 U476 ( .A(regs[999]), .B(n245), .C(regs[935]), .D(n199), .Q(n1087) );
  AOI220 U477 ( .A(regs[967]), .B(n246), .C(regs[903]), .D(n200), .Q(n1086) );
  AOI220 U478 ( .A(regs[871]), .B(n247), .C(regs[807]), .D(n205), .Q(n1085) );
  AOI220 U479 ( .A(regs[487]), .B(n245), .C(regs[423]), .D(n199), .Q(n1091) );
  AOI220 U480 ( .A(regs[455]), .B(n246), .C(regs[391]), .D(n200), .Q(n1090) );
  AOI220 U481 ( .A(regs[743]), .B(n245), .C(regs[679]), .D(n199), .Q(n1097) );
  AOI220 U482 ( .A(regs[711]), .B(n246), .C(regs[647]), .D(n200), .Q(n1096) );
  AOI220 U483 ( .A(n241), .B(regs[457]), .C(n202), .D(regs[393]), .Q(n478) );
  AOI220 U484 ( .A(regs[615]), .B(n247), .C(regs[551]), .D(n205), .Q(n1095) );
  AOI220 U485 ( .A(n241), .B(regs[969]), .C(n202), .D(regs[905]), .Q(n474) );
  AOI220 U486 ( .A(regs[231]), .B(n245), .C(regs[167]), .D(n199), .Q(n1101) );
  AOI220 U487 ( .A(regs[103]), .B(n247), .C(regs[39]), .D(n205), .Q(n1099) );
  AOI220 U488 ( .A(n241), .B(regs[714]), .C(n202), .D(regs[650]), .Q(n506) );
  AOI220 U489 ( .A(n241), .B(regs[970]), .C(n202), .D(regs[906]), .Q(n496) );
  AOI220 U490 ( .A(regs[742]), .B(n245), .C(regs[678]), .D(n199), .Q(n1075) );
  AOI220 U491 ( .A(regs[710]), .B(n246), .C(regs[646]), .D(n200), .Q(n1074) );
  AOI220 U492 ( .A(n242), .B(regs[203]), .C(n202), .D(regs[139]), .Q(n532) );
  AOI220 U493 ( .A(n241), .B(regs[715]), .C(n974), .D(regs[651]), .Q(n528) );
  AOI220 U494 ( .A(n242), .B(regs[197]), .C(n202), .D(regs[133]), .Q(n400) );
  AOI220 U495 ( .A(n975), .B(regs[459]), .C(n202), .D(regs[395]), .Q(n522) );
  AOI220 U496 ( .A(regs[997]), .B(n245), .C(regs[933]), .D(n199), .Q(n1043) );
  AOI220 U497 ( .A(regs[965]), .B(n246), .C(regs[901]), .D(n200), .Q(n1042) );
  AOI220 U498 ( .A(n241), .B(regs[971]), .C(n202), .D(regs[907]), .Q(n518) );
  AOI220 U499 ( .A(n242), .B(regs[204]), .C(n974), .D(regs[140]), .Q(n554) );
  AOI220 U500 ( .A(n241), .B(regs[716]), .C(n202), .D(regs[652]), .Q(n550) );
  AOI220 U501 ( .A(n201), .B(regs[748]), .C(n198), .D(regs[684]), .Q(n551) );
  AOI220 U502 ( .A(n243), .B(regs[364]), .C(n206), .D(regs[300]), .Q(n543) );
  AOI220 U503 ( .A(n242), .B(regs[460]), .C(n202), .D(regs[396]), .Q(n544) );
  AOI220 U504 ( .A(n242), .B(regs[972]), .C(n202), .D(regs[908]), .Q(n540) );
  AOI220 U505 ( .A(regs[996]), .B(n245), .C(regs[932]), .D(n199), .Q(n1021) );
  AOI220 U506 ( .A(regs[964]), .B(n246), .C(regs[900]), .D(n200), .Q(n1020) );
  AOI220 U507 ( .A(n242), .B(regs[205]), .C(n202), .D(regs[141]), .Q(n576) );
  AOI220 U508 ( .A(n201), .B(regs[237]), .C(n198), .D(regs[173]), .Q(n577) );
  AOI220 U509 ( .A(regs[484]), .B(n245), .C(regs[420]), .D(n199), .Q(n1025) );
  AOI220 U510 ( .A(n242), .B(regs[717]), .C(n202), .D(regs[653]), .Q(n572) );
  AOI220 U511 ( .A(regs[452]), .B(n246), .C(regs[388]), .D(n200), .Q(n1024) );
  AOI220 U512 ( .A(n241), .B(regs[461]), .C(n202), .D(regs[397]), .Q(n566) );
  AOI220 U513 ( .A(n201), .B(regs[493]), .C(n198), .D(regs[429]), .Q(n567) );
  AOI220 U514 ( .A(regs[740]), .B(n245), .C(regs[676]), .D(n199), .Q(n1031) );
  AOI220 U515 ( .A(regs[708]), .B(n246), .C(regs[644]), .D(n200), .Q(n1030) );
  AOI220 U516 ( .A(n241), .B(regs[973]), .C(n974), .D(regs[909]), .Q(n562) );
  AOI220 U517 ( .A(regs[612]), .B(n247), .C(regs[548]), .D(n1566), .Q(n1029)
         );
  AOI220 U518 ( .A(regs[228]), .B(n245), .C(regs[164]), .D(n199), .Q(n1035) );
  AOI220 U519 ( .A(regs[196]), .B(n246), .C(regs[132]), .D(n200), .Q(n1034) );
  AOI220 U520 ( .A(n242), .B(regs[462]), .C(n974), .D(regs[398]), .Q(n588) );
  AOI220 U521 ( .A(n242), .B(regs[974]), .C(n202), .D(regs[910]), .Q(n584) );
  AOI220 U522 ( .A(n242), .B(regs[207]), .C(n974), .D(regs[143]), .Q(n620) );
  AOI220 U523 ( .A(n201), .B(regs[239]), .C(n198), .D(regs[175]), .Q(n621) );
  AOI220 U524 ( .A(n201), .B(regs[751]), .C(n972), .D(regs[687]), .Q(n617) );
  AOI220 U525 ( .A(n975), .B(regs[975]), .C(n202), .D(regs[911]), .Q(n606) );
  AOI220 U526 ( .A(n201), .B(regs[240]), .C(n198), .D(regs[176]), .Q(n643) );
  AOI220 U527 ( .A(n201), .B(regs[752]), .C(n198), .D(regs[688]), .Q(n639) );
  AOI220 U528 ( .A(n975), .B(regs[464]), .C(n202), .D(regs[400]), .Q(n632) );
  AOI220 U529 ( .A(regs[375]), .B(n247), .C(regs[311]), .D(n1566), .Q(n1375)
         );
  AOI220 U530 ( .A(regs[887]), .B(n247), .C(regs[823]), .D(n205), .Q(n1371) );
  AOI220 U531 ( .A(regs[119]), .B(n247), .C(regs[55]), .D(n205), .Q(n1385) );
  AOI220 U532 ( .A(regs[120]), .B(n247), .C(regs[56]), .D(n205), .Q(n1407) );
  AOI220 U533 ( .A(regs[632]), .B(n247), .C(regs[568]), .D(n205), .Q(n1403) );
  AOI220 U534 ( .A(regs[728]), .B(n246), .C(regs[664]), .D(n200), .Q(n1404) );
  AOI220 U535 ( .A(regs[760]), .B(n245), .C(regs[696]), .D(n199), .Q(n1405) );
  AOI220 U536 ( .A(regs[376]), .B(n247), .C(regs[312]), .D(n1566), .Q(n1397)
         );
  AOI220 U537 ( .A(regs[888]), .B(n247), .C(regs[824]), .D(n205), .Q(n1393) );
  AOI220 U538 ( .A(regs[118]), .B(n247), .C(regs[54]), .D(n205), .Q(n1363) );
  AOI220 U539 ( .A(regs[121]), .B(n247), .C(regs[57]), .D(n205), .Q(n1429) );
  AOI220 U540 ( .A(regs[633]), .B(n247), .C(regs[569]), .D(n205), .Q(n1425) );
  AOI220 U541 ( .A(regs[377]), .B(n247), .C(regs[313]), .D(n1566), .Q(n1419)
         );
  AOI220 U542 ( .A(regs[889]), .B(n247), .C(regs[825]), .D(n1566), .Q(n1415)
         );
  AOI220 U543 ( .A(regs[730]), .B(n246), .C(regs[666]), .D(n200), .Q(n1448) );
  AOI220 U544 ( .A(regs[762]), .B(n245), .C(regs[698]), .D(n199), .Q(n1449) );
  AOI220 U545 ( .A(regs[890]), .B(n247), .C(regs[826]), .D(n1566), .Q(n1437)
         );
  AOI220 U546 ( .A(regs[475]), .B(n246), .C(regs[411]), .D(n200), .Q(n1464) );
  AOI220 U547 ( .A(regs[507]), .B(n245), .C(regs[443]), .D(n199), .Q(n1465) );
  AOI220 U548 ( .A(regs[252]), .B(n245), .C(regs[188]), .D(n199), .Q(n1497) );
  AOI220 U549 ( .A(regs[627]), .B(n247), .C(regs[563]), .D(n205), .Q(n1315) );
  AOI220 U550 ( .A(regs[242]), .B(n245), .C(regs[178]), .D(n199), .Q(n1299) );
  AOI220 U551 ( .A(regs[1022]), .B(n245), .C(regs[958]), .D(n199), .Q(n1527)
         );
  AOI220 U552 ( .A(regs[383]), .B(n247), .C(regs[319]), .D(n205), .Q(n1551) );
  AOI220 U553 ( .A(regs[240]), .B(n245), .C(regs[176]), .D(n199), .Q(n1255) );
  AOI220 U554 ( .A(regs[631]), .B(n247), .C(regs[567]), .D(n205), .Q(n1381) );
  AOI220 U555 ( .A(regs[610]), .B(n247), .C(regs[546]), .D(n205), .Q(n1007) );
  AOI220 U556 ( .A(regs[704]), .B(n242), .C(regs[640]), .D(n202), .Q(n286) );
  AOI220 U557 ( .A(n242), .B(regs[960]), .C(n202), .D(regs[896]), .Q(n274) );
  AOI220 U558 ( .A(n241), .B(regs[194]), .C(n202), .D(regs[130]), .Q(n334) );
  AOI220 U559 ( .A(n242), .B(regs[706]), .C(n202), .D(regs[642]), .Q(n330) );
  AOI220 U560 ( .A(n201), .B(regs[738]), .C(n972), .D(regs[674]), .Q(n331) );
  AOI220 U561 ( .A(regs[1003]), .B(n245), .C(regs[939]), .D(n199), .Q(n1153)
         );
  AOI220 U562 ( .A(regs[971]), .B(n246), .C(regs[907]), .D(n200), .Q(n1152) );
  AOI220 U563 ( .A(n242), .B(regs[195]), .C(n202), .D(regs[131]), .Q(n356) );
  AOI220 U564 ( .A(n201), .B(regs[227]), .C(n198), .D(regs[163]), .Q(n357) );
  AOI220 U565 ( .A(n241), .B(regs[451]), .C(n974), .D(regs[387]), .Q(n346) );
  AOI220 U566 ( .A(n241), .B(regs[963]), .C(n202), .D(regs[899]), .Q(n342) );
  AOI220 U567 ( .A(n242), .B(regs[708]), .C(n974), .D(regs[644]), .Q(n374) );
  AOI220 U568 ( .A(n242), .B(regs[964]), .C(n202), .D(regs[900]), .Q(n364) );
  AOI220 U569 ( .A(n241), .B(regs[221]), .C(n202), .D(regs[157]), .Q(n928) );
  AOI220 U570 ( .A(n241), .B(regs[980]), .C(n202), .D(regs[916]), .Q(n716) );
  AOI220 U571 ( .A(n243), .B(regs[892]), .C(n206), .D(regs[828]), .Q(n891) );
  AOI220 U572 ( .A(n242), .B(regs[725]), .C(n202), .D(regs[661]), .Q(n748) );
  AOI220 U573 ( .A(n241), .B(regs[476]), .C(n974), .D(regs[412]), .Q(n896) );
  AOI220 U574 ( .A(n242), .B(regs[981]), .C(n202), .D(regs[917]), .Q(n738) );
  AOI220 U575 ( .A(n242), .B(regs[214]), .C(n202), .D(regs[150]), .Q(n774) );
  AOI220 U576 ( .A(n241), .B(regs[726]), .C(n202), .D(regs[662]), .Q(n770) );
  AOI220 U577 ( .A(n241), .B(regs[470]), .C(n202), .D(regs[406]), .Q(n764) );
  AOI220 U578 ( .A(n975), .B(regs[220]), .C(n202), .D(regs[156]), .Q(n906) );
  AOI220 U579 ( .A(n241), .B(regs[982]), .C(n202), .D(regs[918]), .Q(n760) );
  AOI220 U580 ( .A(n242), .B(regs[215]), .C(n202), .D(regs[151]), .Q(n796) );
  AOI220 U581 ( .A(n242), .B(regs[727]), .C(n202), .D(regs[663]), .Q(n792) );
  AOI220 U582 ( .A(n241), .B(regs[471]), .C(n202), .D(regs[407]), .Q(n786) );
  AOI220 U583 ( .A(n242), .B(regs[983]), .C(n202), .D(regs[919]), .Q(n782) );
  AOI220 U584 ( .A(n243), .B(regs[635]), .C(n206), .D(regs[571]), .Q(n879) );
  AOI220 U585 ( .A(n242), .B(regs[216]), .C(n202), .D(regs[152]), .Q(n818) );
  AOI220 U586 ( .A(n241), .B(regs[728]), .C(n202), .D(regs[664]), .Q(n814) );
  AOI220 U587 ( .A(n242), .B(regs[472]), .C(n202), .D(regs[408]), .Q(n808) );
  AOI220 U588 ( .A(n241), .B(regs[986]), .C(n202), .D(regs[922]), .Q(n848) );
  AOI220 U589 ( .A(n241), .B(regs[984]), .C(n202), .D(regs[920]), .Q(n804) );
  AOI220 U590 ( .A(n241), .B(regs[217]), .C(n202), .D(regs[153]), .Q(n840) );
  AOI220 U591 ( .A(n243), .B(regs[378]), .C(n206), .D(regs[314]), .Q(n851) );
  AOI220 U592 ( .A(n241), .B(regs[473]), .C(n202), .D(regs[409]), .Q(n830) );
  AOI220 U593 ( .A(n242), .B(regs[730]), .C(n974), .D(regs[666]), .Q(n858) );
  AOI220 U594 ( .A(n243), .B(regs[634]), .C(n206), .D(regs[570]), .Q(n857) );
  AOI220 U595 ( .A(n242), .B(regs[985]), .C(n202), .D(regs[921]), .Q(n826) );
  AOI220 U596 ( .A(n241), .B(regs[979]), .C(n974), .D(regs[915]), .Q(n694) );
  AOI220 U597 ( .A(n242), .B(regs[466]), .C(n202), .D(regs[402]), .Q(n676) );
  AOI220 U598 ( .A(n241), .B(regs[222]), .C(n974), .D(regs[158]), .Q(n950) );
  AOI220 U599 ( .A(n242), .B(regs[722]), .C(n202), .D(regs[658]), .Q(n682) );
  AOI220 U600 ( .A(n975), .B(regs[734]), .C(n202), .D(regs[670]), .Q(n946) );
  AOI220 U601 ( .A(n241), .B(regs[211]), .C(n974), .D(regs[147]), .Q(n708) );
  AOI220 U602 ( .A(n975), .B(regs[989]), .C(n974), .D(regs[925]), .Q(n914) );
  AOI220 U603 ( .A(n242), .B(regs[210]), .C(n974), .D(regs[146]), .Q(n686) );
  AOI220 U604 ( .A(n975), .B(regs[723]), .C(n202), .D(regs[659]), .Q(n704) );
  AOI220 U605 ( .A(n242), .B(regs[467]), .C(n974), .D(regs[403]), .Q(n698) );
  AOI220 U606 ( .A(n242), .B(regs[478]), .C(n974), .D(regs[414]), .Q(n940) );
  AOI220 U607 ( .A(n975), .B(regs[724]), .C(n202), .D(regs[660]), .Q(n726) );
  AOI220 U608 ( .A(n242), .B(regs[733]), .C(n202), .D(regs[669]), .Q(n924) );
  AOI220 U609 ( .A(n241), .B(regs[458]), .C(n202), .D(regs[394]), .Q(n500) );
  AOI220 U610 ( .A(n975), .B(regs[465]), .C(n202), .D(regs[401]), .Q(n654) );
  AOI220 U611 ( .A(n241), .B(regs[212]), .C(n202), .D(regs[148]), .Q(n730) );
  AOI220 U612 ( .A(regs[1021]), .B(n245), .C(regs[957]), .D(n199), .Q(n1505)
         );
  AOI220 U613 ( .A(regs[509]), .B(n245), .C(regs[445]), .D(n199), .Q(n1509) );
  AOI220 U614 ( .A(regs[510]), .B(n245), .C(regs[446]), .D(n199), .Q(n1531) );
  AOI220 U615 ( .A(regs[255]), .B(n245), .C(regs[191]), .D(n199), .Q(n1573) );
  AOI220 U616 ( .A(regs[495]), .B(n245), .C(regs[431]), .D(n199), .Q(n1223) );
  AOI220 U617 ( .A(regs[1016]), .B(n245), .C(regs[952]), .D(n199), .Q(n1395)
         );
  AOI220 U618 ( .A(regs[489]), .B(n245), .C(regs[425]), .D(n199), .Q(n1135) );
  AOI220 U619 ( .A(regs[251]), .B(n245), .C(regs[187]), .D(n199), .Q(n1475) );
  AOI220 U620 ( .A(regs[508]), .B(n245), .C(regs[444]), .D(n199), .Q(n1487) );
  AOI220 U621 ( .A(n201), .B(regs[226]), .C(n198), .D(regs[162]), .Q(n335) );
  AOI220 U622 ( .A(n201), .B(regs[739]), .C(n198), .D(regs[675]), .Q(n353) );
  AOI220 U623 ( .A(n201), .B(regs[483]), .C(n198), .D(regs[419]), .Q(n347) );
  AOI220 U624 ( .A(n201), .B(regs[995]), .C(n198), .D(regs[931]), .Q(n343) );
  AOI220 U625 ( .A(n201), .B(regs[497]), .C(n198), .D(regs[433]), .Q(n655) );
  AOI220 U626 ( .A(n201), .B(regs[484]), .C(n198), .D(regs[420]), .Q(n369) );
  AOI220 U627 ( .A(n201), .B(regs[996]), .C(n198), .D(regs[932]), .Q(n365) );
  AOI220 U628 ( .A(n201), .B(regs[487]), .C(n198), .D(regs[423]), .Q(n435) );
  AOI220 U629 ( .A(n201), .B(regs[744]), .C(n198), .D(regs[680]), .Q(n463) );
  AOI220 U630 ( .A(n201), .B(regs[488]), .C(n198), .D(regs[424]), .Q(n457) );
  AOI220 U631 ( .A(n201), .B(regs[495]), .C(n198), .D(regs[431]), .Q(n611) );
  AOI220 U632 ( .A(n201), .B(regs[489]), .C(n198), .D(regs[425]), .Q(n479) );
  AOI220 U633 ( .A(n201), .B(regs[1001]), .C(n198), .D(regs[937]), .Q(n475) );
  AOI220 U634 ( .A(n201), .B(regs[234]), .C(n198), .D(regs[170]), .Q(n511) );
  AOI220 U635 ( .A(n201), .B(regs[746]), .C(n198), .D(regs[682]), .Q(n507) );
  AOI220 U636 ( .A(n201), .B(regs[490]), .C(n198), .D(regs[426]), .Q(n501) );
  AOI220 U637 ( .A(n201), .B(regs[1002]), .C(n198), .D(regs[938]), .Q(n497) );
  AOI220 U638 ( .A(n201), .B(regs[235]), .C(n198), .D(regs[171]), .Q(n533) );
  AOI220 U639 ( .A(n201), .B(regs[747]), .C(n198), .D(regs[683]), .Q(n529) );
  AOI220 U640 ( .A(n201), .B(regs[491]), .C(n198), .D(regs[427]), .Q(n523) );
  AOI220 U641 ( .A(n201), .B(regs[1003]), .C(n198), .D(regs[939]), .Q(n519) );
  AOI220 U642 ( .A(n201), .B(regs[494]), .C(n198), .D(regs[430]), .Q(n589) );
  AOI220 U643 ( .A(regs[748]), .B(n245), .C(regs[684]), .D(n199), .Q(n1185) );
  AOI220 U644 ( .A(n201), .B(regs[1004]), .C(n198), .D(regs[940]), .Q(n541) );
  AOI220 U645 ( .A(n201), .B(regs[749]), .C(n198), .D(regs[685]), .Q(n573) );
  AOI220 U646 ( .A(n201), .B(regs[238]), .C(n198), .D(regs[174]), .Q(n599) );
  AOI220 U647 ( .A(regs[236]), .B(n245), .C(regs[172]), .D(n199), .Q(n1189) );
  AOI220 U648 ( .A(n201), .B(regs[1010]), .C(n198), .D(regs[946]), .Q(n673) );
  AOI220 U649 ( .A(regs[1009]), .B(n245), .C(regs[945]), .D(n199), .Q(n1263)
         );
  AOI220 U650 ( .A(regs[1007]), .B(n245), .C(regs[943]), .D(n199), .Q(n1219)
         );
  AOI220 U651 ( .A(n975), .B(regs[223]), .C(n202), .D(regs[159]), .Q(n982) );
  NAND22 U652 ( .A(n1581), .B(i_addr_Rd[3]), .Q(n1592) );
  NAND31 U653 ( .A(i_addr_Rd[0]), .B(n240), .C(n1586), .Q(n1591) );
  NOR21 U654 ( .A(i_addr_Rd[4]), .B(n1580), .Q(n1581) );
  NAND31 U655 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n240), .Q(n1589) );
  NAND31 U656 ( .A(n240), .B(n1587), .C(n1586), .Q(n1585) );
  NOR22 U657 ( .A(i_addr_Rs[4]), .B(n994), .Q(n1555) );
  NOR32 U658 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .C(n268), .Q(n974) );
  NOR22 U659 ( .A(i_addr_Rt_3_), .B(n283), .Q(n987) );
  NAND31 U660 ( .A(i_addr_Rd[1]), .B(n240), .C(n1587), .Q(n1590) );
  NOR22 U661 ( .A(i_addr_Rs[3]), .B(n995), .Q(n1577) );
  NOR32 U662 ( .A(i_addr_Rt_0_), .B(n271), .C(n268), .Q(n975) );
  INV2 U663 ( .A(i_addr_Rs[0]), .Q(n992) );
  INV3 U664 ( .A(i_addr_Rs[3]), .Q(n994) );
  INV2 U665 ( .A(i_addr_Rs[1]), .Q(n993) );
  NOR33 U666 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[1]), .C(i_addr_Rs[2]), .Q(n1568)
         );
  INV3 U667 ( .A(i_addr_Rs[4]), .Q(n995) );
  NAND21 U668 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[1]), .Q(n991) );
  INV2 U669 ( .A(i_con_RegWr), .Q(n1580) );
  INV3 U670 ( .A(i_addr_Rt_1_), .Q(n271) );
  INV3 U671 ( .A(i_addr_Rt_0_), .Q(n270) );
  NAND22 U672 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .Q(n269) );
  INV3 U673 ( .A(i_addr_Rt_4_), .Q(n283) );
  NAND31 U674 ( .A(i_con_RegWr), .B(i_addr_Rd[4]), .C(n1584), .Q(n1588) );
  INV3 U675 ( .A(i_addr_Rd[3]), .Q(n1584) );
  NAND31 U676 ( .A(i_addr_Rd[4]), .B(i_con_RegWr), .C(i_addr_Rd[3]), .Q(n1583)
         );
  INV3 U677 ( .A(i_addr_Rd[0]), .Q(n1587) );
  INV3 U678 ( .A(i_addr_Rd[1]), .Q(n1586) );
  INV3 U679 ( .A(i_addr_Rt_3_), .Q(n276) );
  NOR31 U680 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_1_), .C(i_addr_Rt_2_), .Q(n978)
         );
  NAND22 U681 ( .A(n1581), .B(n1584), .Q(n1582) );
  AOI220 U682 ( .A(n243), .B(regs[358]), .C(n206), .D(regs[294]), .Q(n411) );
  AOI220 U683 ( .A(n243), .B(regs[870]), .C(n206), .D(regs[806]), .Q(n407) );
  AOI220 U684 ( .A(n243), .B(regs[101]), .C(n206), .D(regs[37]), .Q(n399) );
  AOI220 U685 ( .A(n243), .B(regs[613]), .C(n206), .D(regs[549]), .Q(n395) );
  AOI220 U686 ( .A(n243), .B(regs[357]), .C(n206), .D(regs[293]), .Q(n389) );
  AOI220 U687 ( .A(n243), .B(regs[869]), .C(n206), .D(regs[805]), .Q(n385) );
  AOI220 U688 ( .A(n201), .B(regs[245]), .C(n972), .D(regs[181]), .Q(n753) );
  AOI220 U689 ( .A(n243), .B(regs[629]), .C(n206), .D(regs[565]), .Q(n747) );
  AOI220 U690 ( .A(n201), .B(regs[501]), .C(n972), .D(regs[437]), .Q(n743) );
  AOI220 U691 ( .A(n243), .B(regs[885]), .C(n206), .D(regs[821]), .Q(n737) );
  AOI220 U692 ( .A(n243), .B(regs[871]), .C(n206), .D(regs[807]), .Q(n429) );
  AOI220 U693 ( .A(n243), .B(regs[124]), .C(n206), .D(regs[60]), .Q(n905) );
  AOI220 U694 ( .A(n243), .B(regs[636]), .C(n206), .D(regs[572]), .Q(n901) );
  AOI220 U695 ( .A(n243), .B(regs[380]), .C(n206), .D(regs[316]), .Q(n895) );
  AOI220 U696 ( .A(n975), .B(regs[988]), .C(n202), .D(regs[924]), .Q(n892) );
  AOI220 U697 ( .A(n243), .B(regs[108]), .C(n206), .D(regs[44]), .Q(n553) );
  AOI220 U698 ( .A(n243), .B(regs[620]), .C(n206), .D(regs[556]), .Q(n549) );
  AOI220 U699 ( .A(n975), .B(regs[218]), .C(n974), .D(regs[154]), .Q(n862) );
  AOI220 U700 ( .A(n243), .B(regs[887]), .C(n206), .D(regs[823]), .Q(n781) );
  AOI220 U701 ( .A(n243), .B(regs[123]), .C(n206), .D(regs[59]), .Q(n883) );
  AOI220 U702 ( .A(n975), .B(regs[731]), .C(n202), .D(regs[667]), .Q(n880) );
  AOI220 U703 ( .A(n243), .B(regs[379]), .C(n206), .D(regs[315]), .Q(n873) );
  AOI220 U704 ( .A(n975), .B(regs[987]), .C(n202), .D(regs[923]), .Q(n870) );
  AOI220 U705 ( .A(n243), .B(regs[118]), .C(n206), .D(regs[54]), .Q(n773) );
  AOI220 U706 ( .A(n243), .B(regs[630]), .C(n206), .D(regs[566]), .Q(n769) );
  AOI220 U707 ( .A(n243), .B(regs[886]), .C(n206), .D(regs[822]), .Q(n759) );
  AOI220 U708 ( .A(n975), .B(regs[208]), .C(n202), .D(regs[144]), .Q(n642) );
  AOI220 U709 ( .A(n975), .B(regs[720]), .C(n202), .D(regs[656]), .Q(n638) );
  AOI220 U710 ( .A(n975), .B(regs[976]), .C(n202), .D(regs[912]), .Q(n628) );
  AOI220 U711 ( .A(n975), .B(regs[192]), .C(n202), .D(regs[128]), .Q(n290) );
  AOI220 U712 ( .A(n975), .B(regs[448]), .C(n202), .D(regs[384]), .Q(n279) );
  AOI220 U713 ( .A(n975), .B(regs[193]), .C(n202), .D(regs[129]), .Q(n312) );
  AOI220 U714 ( .A(n975), .B(regs[705]), .C(n202), .D(regs[641]), .Q(n308) );
  AOI220 U715 ( .A(n975), .B(regs[449]), .C(n202), .D(regs[385]), .Q(n302) );
  AOI220 U716 ( .A(n975), .B(regs[961]), .C(n202), .D(regs[897]), .Q(n298) );
  AOI220 U717 ( .A(n975), .B(regs[719]), .C(n202), .D(regs[655]), .Q(n616) );
  AOI220 U718 ( .A(n975), .B(regs[463]), .C(n202), .D(regs[399]), .Q(n610) );
  AOI220 U719 ( .A(n243), .B(regs[109]), .C(n206), .D(regs[45]), .Q(n575) );
  AOI220 U720 ( .A(n243), .B(regs[877]), .C(n206), .D(regs[813]), .Q(n561) );
  AOI220 U721 ( .A(n975), .B(regs[209]), .C(n202), .D(regs[145]), .Q(n664) );
  AOI220 U722 ( .A(n975), .B(regs[721]), .C(n202), .D(regs[657]), .Q(n660) );
  AOI220 U723 ( .A(n975), .B(regs[450]), .C(n202), .D(regs[386]), .Q(n324) );
  AOI220 U724 ( .A(n975), .B(regs[962]), .C(n974), .D(regs[898]), .Q(n320) );
  AOI220 U725 ( .A(n243), .B(regs[619]), .C(n206), .D(regs[555]), .Q(n527) );
  AOI220 U726 ( .A(n243), .B(regs[875]), .C(n206), .D(regs[811]), .Q(n517) );
  AOI220 U727 ( .A(n975), .B(regs[206]), .C(n202), .D(regs[142]), .Q(n598) );
  AOI220 U728 ( .A(n975), .B(regs[718]), .C(n974), .D(regs[654]), .Q(n594) );
  AOI220 U729 ( .A(n243), .B(regs[116]), .C(n206), .D(regs[52]), .Q(n729) );
  AOI220 U730 ( .A(n201), .B(regs[244]), .C(n972), .D(regs[180]), .Q(n731) );
  AOI220 U731 ( .A(n201), .B(regs[500]), .C(n972), .D(regs[436]), .Q(n721) );
  NOR31 U732 ( .A(i_addr_Rt_0_), .B(i_addr_Rt_2_), .C(n271), .Q(n979) );
  NOR31 U733 ( .A(i_addr_Rt_1_), .B(i_addr_Rt_2_), .C(n270), .Q(n976) );
  INV3 U734 ( .A(i_addr_Rt_2_), .Q(n268) );
  AOI220 U735 ( .A(regs[201]), .B(n246), .C(regs[137]), .D(n200), .Q(n1144) );
  AOI220 U736 ( .A(regs[233]), .B(n245), .C(regs[169]), .D(n199), .Q(n1145) );
  AOI220 U737 ( .A(regs[713]), .B(n246), .C(regs[649]), .D(n200), .Q(n1140) );
  AOI220 U738 ( .A(regs[745]), .B(n245), .C(regs[681]), .D(n199), .Q(n1141) );
  AOI220 U739 ( .A(regs[457]), .B(n246), .C(regs[393]), .D(n200), .Q(n1134) );
  AOI220 U740 ( .A(regs[969]), .B(n246), .C(regs[905]), .D(n200), .Q(n1130) );
  AOI220 U741 ( .A(regs[1001]), .B(n245), .C(regs[937]), .D(n199), .Q(n1131)
         );
  AOI220 U742 ( .A(regs[122]), .B(n247), .C(regs[58]), .D(n205), .Q(n1451) );
  AOI220 U743 ( .A(regs[218]), .B(n246), .C(regs[154]), .D(n200), .Q(n1452) );
  AOI220 U744 ( .A(regs[250]), .B(n245), .C(regs[186]), .D(n199), .Q(n1453) );
  AOI220 U745 ( .A(regs[634]), .B(n247), .C(regs[570]), .D(n205), .Q(n1447) );
  AOI220 U746 ( .A(regs[378]), .B(n247), .C(regs[314]), .D(n205), .Q(n1441) );
  AOI220 U747 ( .A(regs[474]), .B(n246), .C(regs[410]), .D(n200), .Q(n1442) );
  AOI220 U748 ( .A(regs[506]), .B(n245), .C(regs[442]), .D(n199), .Q(n1443) );
  AOI220 U749 ( .A(regs[986]), .B(n246), .C(regs[922]), .D(n200), .Q(n1438) );
  AOI220 U750 ( .A(regs[108]), .B(n247), .C(regs[44]), .D(n205), .Q(n1187) );
  AOI220 U751 ( .A(regs[204]), .B(n246), .C(regs[140]), .D(n200), .Q(n1188) );
  AOI220 U752 ( .A(regs[620]), .B(n247), .C(regs[556]), .D(n205), .Q(n1183) );
  AOI220 U753 ( .A(regs[716]), .B(n246), .C(regs[652]), .D(n200), .Q(n1184) );
  AOI220 U754 ( .A(regs[972]), .B(n246), .C(regs[908]), .D(n200), .Q(n1174) );
  AOI220 U755 ( .A(regs[1004]), .B(n245), .C(regs[940]), .D(n199), .Q(n1175)
         );
  AOI220 U756 ( .A(regs[125]), .B(n247), .C(regs[61]), .D(n205), .Q(n1517) );
  AOI220 U757 ( .A(regs[637]), .B(n247), .C(regs[573]), .D(n205), .Q(n1513) );
  AOI220 U758 ( .A(regs[893]), .B(n247), .C(regs[829]), .D(n205), .Q(n1503) );
  AOI220 U759 ( .A(regs[214]), .B(n246), .C(regs[150]), .D(n200), .Q(n1364) );
  AOI220 U760 ( .A(regs[246]), .B(n245), .C(regs[182]), .D(n199), .Q(n1365) );
  AOI220 U761 ( .A(regs[630]), .B(n247), .C(regs[566]), .D(n205), .Q(n1359) );
  AOI220 U762 ( .A(regs[726]), .B(n246), .C(regs[662]), .D(n200), .Q(n1360) );
  AOI220 U763 ( .A(regs[758]), .B(n245), .C(regs[694]), .D(n199), .Q(n1361) );
  AOI220 U764 ( .A(regs[470]), .B(n246), .C(regs[406]), .D(n200), .Q(n1354) );
  AOI220 U765 ( .A(regs[502]), .B(n245), .C(regs[438]), .D(n199), .Q(n1355) );
  AOI220 U766 ( .A(regs[886]), .B(n247), .C(regs[822]), .D(n205), .Q(n1349) );
  AOI220 U767 ( .A(regs[1014]), .B(n245), .C(regs[950]), .D(n199), .Q(n1351)
         );
  AOI220 U768 ( .A(regs[109]), .B(n247), .C(regs[45]), .D(n205), .Q(n1209) );
  AOI220 U769 ( .A(regs[205]), .B(n246), .C(regs[141]), .D(n200), .Q(n1210) );
  AOI220 U770 ( .A(regs[621]), .B(n247), .C(regs[557]), .D(n205), .Q(n1205) );
  AOI220 U771 ( .A(regs[717]), .B(n246), .C(regs[653]), .D(n200), .Q(n1206) );
  AOI220 U772 ( .A(regs[365]), .B(n247), .C(regs[301]), .D(n205), .Q(n1199) );
  AOI220 U773 ( .A(regs[461]), .B(n246), .C(regs[397]), .D(n200), .Q(n1200) );
  AOI220 U774 ( .A(regs[877]), .B(n247), .C(regs[813]), .D(n205), .Q(n1195) );
  AOI220 U775 ( .A(regs[973]), .B(n246), .C(regs[909]), .D(n200), .Q(n1196) );
  AOI220 U776 ( .A(regs[123]), .B(n247), .C(regs[59]), .D(n205), .Q(n1473) );
  AOI220 U777 ( .A(regs[219]), .B(n246), .C(regs[155]), .D(n200), .Q(n1474) );
  AOI220 U778 ( .A(regs[635]), .B(n247), .C(regs[571]), .D(n205), .Q(n1469) );
  AOI220 U779 ( .A(regs[379]), .B(n247), .C(regs[315]), .D(n205), .Q(n1463) );
  AOI220 U780 ( .A(regs[891]), .B(n247), .C(regs[827]), .D(n205), .Q(n1459) );
  AOI220 U781 ( .A(regs[1019]), .B(n245), .C(regs[955]), .D(n199), .Q(n1461)
         );
  AOI220 U782 ( .A(regs[723]), .B(n246), .C(regs[659]), .D(n200), .Q(n1316) );
  AOI220 U783 ( .A(regs[755]), .B(n245), .C(regs[691]), .D(n199), .Q(n1317) );
  AOI220 U784 ( .A(regs[979]), .B(n246), .C(regs[915]), .D(n200), .Q(n1306) );
  AOI220 U785 ( .A(regs[1011]), .B(n245), .C(regs[947]), .D(n199), .Q(n1307)
         );
  AOI220 U786 ( .A(regs[124]), .B(n247), .C(regs[60]), .D(n205), .Q(n1495) );
  AOI220 U787 ( .A(regs[636]), .B(n247), .C(regs[572]), .D(n205), .Q(n1491) );
  AOI220 U788 ( .A(regs[476]), .B(n246), .C(regs[412]), .D(n200), .Q(n1486) );
  AOI220 U789 ( .A(regs[892]), .B(n247), .C(regs[828]), .D(n205), .Q(n1481) );
  AOI220 U790 ( .A(regs[988]), .B(n246), .C(regs[924]), .D(n200), .Q(n1482) );
  AOI220 U791 ( .A(regs[626]), .B(n247), .C(regs[562]), .D(n205), .Q(n1293) );
  AOI220 U792 ( .A(regs[722]), .B(n246), .C(regs[658]), .D(n200), .Q(n1294) );
  AOI220 U793 ( .A(regs[754]), .B(n245), .C(regs[690]), .D(n199), .Q(n1295) );
  AOI220 U794 ( .A(regs[466]), .B(n246), .C(regs[402]), .D(n200), .Q(n1288) );
  AOI220 U795 ( .A(regs[498]), .B(n245), .C(regs[434]), .D(n199), .Q(n1289) );
  AOI220 U796 ( .A(regs[882]), .B(n247), .C(regs[818]), .D(n205), .Q(n1283) );
  AOI220 U797 ( .A(regs[978]), .B(n246), .C(regs[914]), .D(n200), .Q(n1284) );
  AOI220 U798 ( .A(regs[1010]), .B(n245), .C(regs[946]), .D(n199), .Q(n1285)
         );
  AOI220 U799 ( .A(regs[625]), .B(n247), .C(regs[561]), .D(n205), .Q(n1271) );
  AOI220 U800 ( .A(regs[721]), .B(n246), .C(regs[657]), .D(n200), .Q(n1272) );
  AOI220 U801 ( .A(regs[753]), .B(n245), .C(regs[689]), .D(n199), .Q(n1273) );
  AOI220 U802 ( .A(regs[881]), .B(n247), .C(regs[817]), .D(n205), .Q(n1261) );
  AOI220 U803 ( .A(regs[977]), .B(n246), .C(regs[913]), .D(n200), .Q(n1262) );
  AOI220 U804 ( .A(regs[216]), .B(n246), .C(regs[152]), .D(n200), .Q(n1408) );
  AOI220 U805 ( .A(regs[248]), .B(n245), .C(regs[184]), .D(n199), .Q(n1409) );
  AOI220 U806 ( .A(regs[472]), .B(n246), .C(regs[408]), .D(n200), .Q(n1398) );
  AOI220 U807 ( .A(regs[504]), .B(n245), .C(regs[440]), .D(n199), .Q(n1399) );
  AOI220 U808 ( .A(regs[984]), .B(n246), .C(regs[920]), .D(n200), .Q(n1394) );
  AOI220 U809 ( .A(regs[215]), .B(n246), .C(regs[151]), .D(n200), .Q(n1386) );
  AOI220 U810 ( .A(regs[247]), .B(n245), .C(regs[183]), .D(n199), .Q(n1387) );
  AOI220 U811 ( .A(regs[727]), .B(n246), .C(regs[663]), .D(n200), .Q(n1382) );
  AOI220 U812 ( .A(regs[759]), .B(n245), .C(regs[695]), .D(n199), .Q(n1383) );
  AOI220 U813 ( .A(regs[471]), .B(n246), .C(regs[407]), .D(n200), .Q(n1376) );
  AOI220 U814 ( .A(regs[503]), .B(n245), .C(regs[439]), .D(n199), .Q(n1377) );
  AOI220 U815 ( .A(regs[1015]), .B(n245), .C(regs[951]), .D(n199), .Q(n1373)
         );
  AOI220 U816 ( .A(regs[715]), .B(n246), .C(regs[651]), .D(n200), .Q(n1162) );
  AOI220 U817 ( .A(regs[747]), .B(n245), .C(regs[683]), .D(n199), .Q(n1163) );
  AOI220 U818 ( .A(regs[459]), .B(n246), .C(regs[395]), .D(n200), .Q(n1156) );
  AOI220 U819 ( .A(regs[491]), .B(n245), .C(regs[427]), .D(n199), .Q(n1157) );
  AOI220 U820 ( .A(regs[194]), .B(n246), .C(regs[130]), .D(n200), .Q(n1012) );
  AOI220 U821 ( .A(regs[226]), .B(n245), .C(regs[162]), .D(n199), .Q(n1013) );
  AOI220 U822 ( .A(regs[706]), .B(n246), .C(regs[642]), .D(n200), .Q(n1008) );
  AOI220 U823 ( .A(regs[738]), .B(n245), .C(regs[674]), .D(n199), .Q(n1009) );
  AOI220 U824 ( .A(regs[450]), .B(n246), .C(regs[386]), .D(n200), .Q(n1002) );
  AOI220 U825 ( .A(regs[482]), .B(n245), .C(regs[418]), .D(n199), .Q(n1003) );
  AOI220 U826 ( .A(regs[962]), .B(n246), .C(regs[898]), .D(n200), .Q(n998) );
  AOI220 U827 ( .A(regs[994]), .B(n245), .C(regs[930]), .D(n199), .Q(n999) );
  AOI220 U828 ( .A(regs[197]), .B(n246), .C(regs[133]), .D(n200), .Q(n1056) );
  AOI220 U829 ( .A(regs[709]), .B(n246), .C(regs[645]), .D(n200), .Q(n1052) );
  AOI220 U830 ( .A(regs[112]), .B(n247), .C(regs[48]), .D(n205), .Q(n1253) );
  AOI220 U831 ( .A(regs[624]), .B(n247), .C(regs[560]), .D(n205), .Q(n1249) );
  AOI220 U832 ( .A(regs[720]), .B(n246), .C(regs[656]), .D(n200), .Q(n1250) );
  AOI220 U833 ( .A(regs[464]), .B(n246), .C(regs[400]), .D(n200), .Q(n1244) );
  AOI220 U834 ( .A(regs[880]), .B(n247), .C(regs[816]), .D(n205), .Q(n1239) );
  AOI220 U835 ( .A(regs[111]), .B(n247), .C(regs[47]), .D(n205), .Q(n1231) );
  AOI220 U836 ( .A(regs[623]), .B(n247), .C(regs[559]), .D(n205), .Q(n1227) );
  AOI220 U837 ( .A(regs[719]), .B(n246), .C(regs[655]), .D(n200), .Q(n1228) );
  AOI220 U838 ( .A(regs[367]), .B(n247), .C(regs[303]), .D(n205), .Q(n1221) );
  AOI220 U839 ( .A(regs[463]), .B(n246), .C(regs[399]), .D(n200), .Q(n1222) );
  AOI220 U840 ( .A(regs[879]), .B(n247), .C(regs[815]), .D(n205), .Q(n1217) );
  AOI220 U841 ( .A(regs[975]), .B(n246), .C(regs[911]), .D(n200), .Q(n1218) );
  AOI220 U842 ( .A(regs[212]), .B(n246), .C(regs[148]), .D(n200), .Q(n1342) );
  AOI220 U843 ( .A(regs[244]), .B(n245), .C(regs[180]), .D(n199), .Q(n1343) );
  AOI220 U844 ( .A(regs[628]), .B(n247), .C(regs[564]), .D(n205), .Q(n1337) );
  AOI220 U845 ( .A(regs[724]), .B(n246), .C(regs[660]), .D(n200), .Q(n1338) );
  AOI220 U846 ( .A(regs[756]), .B(n245), .C(regs[692]), .D(n199), .Q(n1339) );
  AOI220 U847 ( .A(regs[884]), .B(n247), .C(regs[820]), .D(n205), .Q(n1327) );
  AOI220 U848 ( .A(regs[980]), .B(n246), .C(regs[916]), .D(n200), .Q(n1328) );
  AOI220 U849 ( .A(regs[1012]), .B(n245), .C(regs[948]), .D(n199), .Q(n1329)
         );
  AOI220 U850 ( .A(regs[217]), .B(n246), .C(regs[153]), .D(n200), .Q(n1430) );
  AOI220 U851 ( .A(regs[249]), .B(n245), .C(regs[185]), .D(n199), .Q(n1431) );
  AOI220 U852 ( .A(regs[729]), .B(n246), .C(regs[665]), .D(n200), .Q(n1426) );
  AOI220 U853 ( .A(regs[761]), .B(n245), .C(regs[697]), .D(n199), .Q(n1427) );
  AOI220 U854 ( .A(regs[473]), .B(n246), .C(regs[409]), .D(n200), .Q(n1420) );
  AOI220 U855 ( .A(regs[505]), .B(n245), .C(regs[441]), .D(n199), .Q(n1421) );
  AOI220 U856 ( .A(regs[985]), .B(n246), .C(regs[921]), .D(n200), .Q(n1416) );
  AOI220 U857 ( .A(regs[1017]), .B(n245), .C(regs[953]), .D(n199), .Q(n1417)
         );
  AOI220 U858 ( .A(regs[200]), .B(n246), .C(regs[136]), .D(n200), .Q(n1122) );
  AOI220 U859 ( .A(regs[232]), .B(n245), .C(regs[168]), .D(n199), .Q(n1123) );
  AOI220 U860 ( .A(regs[198]), .B(n246), .C(regs[134]), .D(n200), .Q(n1078) );
  AOI220 U861 ( .A(regs[230]), .B(n245), .C(regs[166]), .D(n199), .Q(n1079) );
  AOI220 U862 ( .A(regs[966]), .B(n246), .C(regs[902]), .D(n200), .Q(n1064) );
  AOI220 U863 ( .A(regs[126]), .B(n247), .C(regs[62]), .D(n205), .Q(n1539) );
  AOI220 U864 ( .A(regs[222]), .B(n246), .C(regs[158]), .D(n200), .Q(n1540) );
  AOI220 U865 ( .A(regs[638]), .B(n247), .C(regs[574]), .D(n205), .Q(n1535) );
  AOI220 U866 ( .A(regs[734]), .B(n246), .C(regs[670]), .D(n200), .Q(n1536) );
  AOI220 U867 ( .A(regs[478]), .B(n246), .C(regs[414]), .D(n200), .Q(n1530) );
  AOI220 U868 ( .A(regs[894]), .B(n247), .C(regs[830]), .D(n205), .Q(n1525) );
  AOI220 U869 ( .A(regs[639]), .B(n247), .C(regs[575]), .D(n205), .Q(n1559) );
  AOI220 U870 ( .A(regs[479]), .B(n246), .C(regs[415]), .D(n200), .Q(n1552) );
  AOI220 U871 ( .A(regs[511]), .B(n245), .C(regs[447]), .D(n199), .Q(n1553) );
  AOI220 U872 ( .A(regs[895]), .B(n247), .C(regs[831]), .D(n205), .Q(n1547) );
  AOI220 U873 ( .A(regs[991]), .B(n246), .C(regs[927]), .D(n200), .Q(n1548) );
  AOI220 U874 ( .A(regs[1023]), .B(n245), .C(regs[959]), .D(n199), .Q(n1549)
         );
  NOR31 U875 ( .A(i_addr_Rs[1]), .B(n992), .C(n990), .Q(n1562) );
  INV3 U876 ( .A(i_addr_Rs[2]), .Q(n990) );
  AOI221 U877 ( .A(n244), .B(regs[860]), .C(n232), .D(regs[796]), .Q(n890) );
  AOI221 U878 ( .A(n244), .B(regs[588]), .C(n232), .D(regs[524]), .Q(n548) );
  AOI221 U879 ( .A(n244), .B(regs[602]), .C(n232), .D(regs[538]), .Q(n856) );
  AOI221 U880 ( .A(n244), .B(regs[603]), .C(n232), .D(regs[539]), .Q(n878) );
  AOI221 U881 ( .A(n244), .B(regs[856]), .C(n232), .D(regs[792]), .Q(n802) );
  AOI221 U882 ( .A(n244), .B(regs[77]), .C(n232), .D(regs[13]), .Q(n574) );
  AOI221 U883 ( .A(n244), .B(regs[589]), .C(n232), .D(regs[525]), .Q(n570) );
  AOI220 U884 ( .A(regs[858]), .B(n203), .C(regs[794]), .D(n204), .Q(n1436) );
  AOI220 U885 ( .A(regs[844]), .B(n203), .C(regs[780]), .D(n204), .Q(n1172) );
  AOI220 U886 ( .A(regs[861]), .B(n203), .C(regs[797]), .D(n204), .Q(n1502) );
  AOI220 U887 ( .A(regs[83]), .B(n203), .C(regs[19]), .D(n204), .Q(n1318) );
  AOI220 U888 ( .A(regs[75]), .B(n203), .C(regs[11]), .D(n204), .Q(n1164) );
  AOI220 U889 ( .A(regs[834]), .B(n203), .C(regs[770]), .D(n204), .Q(n996) );
  AOI220 U890 ( .A(regs[581]), .B(n203), .C(regs[517]), .D(n204), .Q(n1050) );
  AOI220 U891 ( .A(regs[606]), .B(n203), .C(regs[542]), .D(n204), .Q(n1534) );
  AOI220 U892 ( .A(regs[350]), .B(n203), .C(regs[286]), .D(n204), .Q(n1528) );
  AOI220 U893 ( .A(regs[862]), .B(n203), .C(regs[798]), .D(n204), .Q(n1524) );
  AOI220 U894 ( .A(regs[607]), .B(n203), .C(regs[543]), .D(n204), .Q(n1558) );
  AOI220 U895 ( .A(regs[863]), .B(n203), .C(regs[799]), .D(n204), .Q(n1546) );
  AOI221 U896 ( .A(n201), .B(regs[743]), .C(n198), .D(regs[679]), .Q(n441) );
  AOI221 U897 ( .A(n201), .B(regs[1008]), .C(n198), .D(regs[944]), .Q(n629) );
  AOI221 U898 ( .A(n201), .B(regs[1007]), .C(n198), .D(regs[943]), .Q(n607) );
  AOI221 U899 ( .A(n201), .B(regs[241]), .C(n198), .D(regs[177]), .Q(n665) );
  AOI221 U900 ( .A(n201), .B(regs[1006]), .C(n198), .D(regs[942]), .Q(n585) );
  AOI220 U901 ( .A(regs[598]), .B(n203), .C(regs[534]), .D(n204), .Q(n1358) );
  AOI220 U902 ( .A(regs[351]), .B(n203), .C(regs[287]), .D(n204), .Q(n1550) );
  AOI221 U903 ( .A(n967), .B(n349), .C(n965), .D(n348), .Q(n361) );
  AOI220 U904 ( .A(n243), .B(regs[873]), .C(n206), .D(regs[809]), .Q(n473) );
  AOI220 U905 ( .A(n243), .B(regs[616]), .C(n206), .D(regs[552]), .Q(n461) );
  AOI221 U906 ( .A(n967), .B(n282), .C(n965), .D(n281), .Q(n295) );
  AOI221 U907 ( .A(n967), .B(n305), .C(n965), .D(n304), .Q(n317) );
  AOI221 U908 ( .A(n967), .B(n613), .C(n965), .D(n612), .Q(n625) );
  AOI221 U909 ( .A(n244), .B(regs[82]), .C(n232), .D(regs[18]), .Q(n684) );
  AOI220 U910 ( .A(regs[595]), .B(n203), .C(regs[531]), .D(n204), .Q(n1314) );
  AOI220 U911 ( .A(regs[339]), .B(n203), .C(regs[275]), .D(n204), .Q(n1308) );
  AOI220 U912 ( .A(regs[82]), .B(n203), .C(regs[18]), .D(n204), .Q(n1296) );
  AOI220 U913 ( .A(regs[594]), .B(n203), .C(regs[530]), .D(n204), .Q(n1292) );
  AOI220 U914 ( .A(regs[338]), .B(n203), .C(regs[274]), .D(n204), .Q(n1286) );
  AOI220 U915 ( .A(regs[850]), .B(n203), .C(regs[786]), .D(n204), .Q(n1282) );
  AOI220 U916 ( .A(regs[836]), .B(n203), .C(regs[772]), .D(n204), .Q(n1018) );
  AOI220 U917 ( .A(regs[81]), .B(n203), .C(regs[17]), .D(n204), .Q(n1274) );
  AOI220 U918 ( .A(regs[88]), .B(n203), .C(regs[24]), .D(n204), .Q(n1406) );
  AOI220 U919 ( .A(regs[344]), .B(n203), .C(regs[280]), .D(n204), .Q(n1396) );
  AOI220 U920 ( .A(regs[856]), .B(n203), .C(regs[792]), .D(n204), .Q(n1392) );
  AOI220 U921 ( .A(regs[87]), .B(n203), .C(regs[23]), .D(n204), .Q(n1384) );
  AOI220 U922 ( .A(regs[599]), .B(n203), .C(regs[535]), .D(n204), .Q(n1380) );
  AOI220 U923 ( .A(regs[855]), .B(n203), .C(regs[791]), .D(n204), .Q(n1370) );
  AOI220 U924 ( .A(regs[587]), .B(n203), .C(regs[523]), .D(n204), .Q(n1160) );
  AOI220 U925 ( .A(regs[331]), .B(n203), .C(regs[267]), .D(n204), .Q(n1154) );
  AOI220 U926 ( .A(regs[325]), .B(n203), .C(regs[261]), .D(n204), .Q(n1044) );
  AOI220 U927 ( .A(regs[591]), .B(n203), .C(regs[527]), .D(n204), .Q(n1226) );
  AOI220 U928 ( .A(regs[84]), .B(n203), .C(regs[20]), .D(n204), .Q(n1340) );
  AOI220 U929 ( .A(regs[596]), .B(n203), .C(regs[532]), .D(n204), .Q(n1336) );
  AOI220 U930 ( .A(regs[852]), .B(n203), .C(regs[788]), .D(n204), .Q(n1326) );
  AOI220 U931 ( .A(regs[89]), .B(n203), .C(regs[25]), .D(n204), .Q(n1428) );
  AOI220 U932 ( .A(regs[601]), .B(n203), .C(regs[537]), .D(n204), .Q(n1424) );
  AOI220 U933 ( .A(regs[857]), .B(n203), .C(regs[793]), .D(n204), .Q(n1414) );
  AOI220 U934 ( .A(regs[584]), .B(n203), .C(regs[520]), .D(n204), .Q(n1116) );
  AOI220 U935 ( .A(regs[840]), .B(n203), .C(regs[776]), .D(n204), .Q(n1106) );
  AOI221 U936 ( .A(n201), .B(regs[509]), .C(n198), .D(regs[445]), .Q(n919) );
  AOI221 U937 ( .A(n201), .B(regs[1021]), .C(n198), .D(regs[957]), .Q(n915) );
  AOI221 U938 ( .A(n201), .B(regs[486]), .C(n198), .D(regs[422]), .Q(n413) );
  AOI221 U939 ( .A(n201), .B(regs[998]), .C(n198), .D(regs[934]), .Q(n409) );
  AOI221 U940 ( .A(n201), .B(regs[229]), .C(n198), .D(regs[165]), .Q(n401) );
  AOI221 U941 ( .A(n201), .B(regs[741]), .C(n198), .D(regs[677]), .Q(n397) );
  AOI221 U942 ( .A(n201), .B(regs[485]), .C(n198), .D(regs[421]), .Q(n391) );
  AOI221 U943 ( .A(n201), .B(regs[997]), .C(n198), .D(regs[933]), .Q(n387) );
  AOI221 U944 ( .A(n201), .B(regs[255]), .C(n198), .D(regs[191]), .Q(n983) );
  AOI221 U945 ( .A(n201), .B(regs[510]), .C(n198), .D(regs[446]), .Q(n941) );
  AOI221 U946 ( .A(n201), .B(regs[252]), .C(n198), .D(regs[188]), .Q(n907) );
  AOI221 U947 ( .A(n201), .B(regs[764]), .C(n198), .D(regs[700]), .Q(n903) );
  AOI221 U948 ( .A(n201), .B(regs[236]), .C(n198), .D(regs[172]), .Q(n555) );
  AOI221 U949 ( .A(n201), .B(regs[763]), .C(n198), .D(regs[699]), .Q(n881) );
  AOI221 U950 ( .A(n201), .B(regs[1019]), .C(n198), .D(regs[955]), .Q(n871) );
  AOI221 U951 ( .A(regs[736]), .B(n201), .C(regs[672]), .D(n198), .Q(n287) );
  AOI221 U952 ( .A(n201), .B(regs[228]), .C(n198), .D(regs[164]), .Q(n379) );
  AOI221 U953 ( .A(n201), .B(regs[740]), .C(n198), .D(regs[676]), .Q(n375) );
  AOI221 U954 ( .A(n201), .B(regs[1009]), .C(n198), .D(regs[945]), .Q(n651) );
  AOI221 U955 ( .A(n967), .B(n591), .C(n965), .D(n590), .Q(n603) );
  AOI221 U956 ( .A(n201), .B(regs[242]), .C(n198), .D(regs[178]), .Q(n687) );
  AOI221 U957 ( .A(n967), .B(n701), .C(n965), .D(n700), .Q(n713) );
  NOR21 U958 ( .A(i_addr_Rt_2_), .B(n269), .Q(n977) );
  NOR31 U959 ( .A(i_addr_Rt_1_), .B(n270), .C(n268), .Q(n972) );
  NOR21 U960 ( .A(n269), .B(n268), .Q(n973) );
  AOI220 U961 ( .A(regs[86]), .B(n203), .C(regs[22]), .D(n204), .Q(n1362) );
  AOI220 U962 ( .A(regs[92]), .B(n203), .C(regs[28]), .D(n204), .Q(n1494) );
  AOI220 U963 ( .A(regs[604]), .B(n203), .C(regs[540]), .D(n204), .Q(n1490) );
  AOI220 U964 ( .A(regs[348]), .B(n203), .C(regs[284]), .D(n204), .Q(n1484) );
  AOI220 U965 ( .A(regs[860]), .B(n203), .C(regs[796]), .D(n204), .Q(n1480) );
  AOI220 U966 ( .A(regs[849]), .B(n203), .C(regs[785]), .D(n204), .Q(n1260) );
  AOI220 U967 ( .A(regs[837]), .B(n203), .C(regs[773]), .D(n204), .Q(n1040) );
  AOI220 U968 ( .A(regs[592]), .B(n203), .C(regs[528]), .D(n204), .Q(n1248) );
  AOI220 U969 ( .A(regs[345]), .B(n203), .C(regs[281]), .D(n204), .Q(n1418) );
  AOI220 U970 ( .A(regs[838]), .B(n203), .C(regs[774]), .D(n204), .Q(n1062) );
  AOI220 U971 ( .A(regs[95]), .B(n203), .C(regs[31]), .D(n204), .Q(n1570) );
  NOR21 U972 ( .A(n991), .B(n990), .Q(n1563) );
  BUF2 U973 ( .A(n22), .Q(n260) );
  BUF2 U974 ( .A(n21), .Q(n261) );
  BUF2 U975 ( .A(n20), .Q(n262) );
  BUF2 U976 ( .A(n18), .Q(n263) );
  BUF2 U977 ( .A(n25), .Q(n258) );
  BUF2 U978 ( .A(n26), .Q(n257) );
  BUF2 U979 ( .A(n23), .Q(n259) );
  BUF2 U980 ( .A(n15), .Q(n266) );
  BUF2 U981 ( .A(n16), .Q(n265) );
  BUF2 U982 ( .A(n13), .Q(n267) );
  BUF2 U983 ( .A(n42), .Q(n250) );
  BUF2 U984 ( .A(n41), .Q(n251) );
  BUF2 U985 ( .A(n43), .Q(n249) );
  BUF2 U986 ( .A(n32), .Q(n255) );
  BUF2 U987 ( .A(n35), .Q(n253) );
  BUF2 U988 ( .A(n34), .Q(n254) );
  BUF2 U989 ( .A(i_addr_Rd[2]), .Q(n240) );
  AOI221 U990 ( .A(n987), .B(n403), .C(n985), .D(n402), .Q(n404) );
  AOI221 U991 ( .A(n201), .B(regs[767]), .C(n198), .D(regs[703]), .Q(n971) );
  AOI221 U992 ( .A(n201), .B(regs[511]), .C(n198), .D(regs[447]), .Q(n963) );
  AOI221 U993 ( .A(n201), .B(regs[1023]), .C(n198), .D(regs[959]), .Q(n959) );
  AOI221 U994 ( .A(n242), .B(regs[201]), .C(n202), .D(regs[137]), .Q(n488) );
  AOI221 U995 ( .A(n201), .B(regs[254]), .C(n198), .D(regs[190]), .Q(n951) );
  AOI221 U996 ( .A(n201), .B(regs[766]), .C(n198), .D(regs[702]), .Q(n947) );
  AOI221 U997 ( .A(n201), .B(regs[992]), .C(n198), .D(regs[928]), .Q(n275) );
  AOI221 U998 ( .A(n987), .B(n667), .C(n985), .D(n666), .Q(n668) );
  AOI220 U999 ( .A(regs[883]), .B(n247), .C(regs[819]), .D(n205), .Q(n1305) );
  AOI220 U1000 ( .A(regs[370]), .B(n247), .C(regs[306]), .D(n205), .Q(n1287)
         );
  NOR31 U1001 ( .A(i_addr_Rs[0]), .B(i_addr_Rs[2]), .C(n993), .Q(n1569) );
  NOR21 U1002 ( .A(i_addr_Rs[2]), .B(n991), .Q(n1567) );
  BUF2 U1003 ( .A(n27), .Q(n256) );
  BUF2 U1004 ( .A(n17), .Q(n264) );
  BUF2 U1005 ( .A(n44), .Q(n248) );
  NOR40 U1006 ( .A(n240), .B(n1587), .C(n1592), .D(n1586), .Q(n44) );
  AOI221 U1007 ( .A(n987), .B(n425), .C(n985), .D(n424), .Q(n426) );
  AOI221 U1008 ( .A(n987), .B(n491), .C(n985), .D(n490), .Q(n492) );
  AOI221 U1009 ( .A(n987), .B(n447), .C(n985), .D(n446), .Q(n448) );
  AOI220 U1010 ( .A(n243), .B(regs[382]), .C(n206), .D(regs[318]), .Q(n939) );
  AOI220 U1011 ( .A(n243), .B(regs[122]), .C(n206), .D(regs[58]), .Q(n861) );
  AOI221 U1012 ( .A(n987), .B(n645), .C(n985), .D(n644), .Q(n646) );
  AOI221 U1013 ( .A(n987), .B(n293), .C(n985), .D(n292), .Q(n294) );
  AOI220 U1014 ( .A(regs[576]), .B(n244), .C(regs[512]), .D(n232), .Q(n284) );
  AOI221 U1015 ( .A(n987), .B(n623), .C(n985), .D(n622), .Q(n624) );
  AOI221 U1016 ( .A(n987), .B(n337), .C(n985), .D(n336), .Q(n338) );
  AOI221 U1017 ( .A(n1577), .B(n1147), .C(n1575), .D(n1146), .Q(n1148) );
  AOI220 U1018 ( .A(regs[114]), .B(n247), .C(regs[50]), .D(n205), .Q(n1297) );
  AOI221 U1019 ( .A(n1577), .B(n1037), .C(n1575), .D(n1036), .Q(n1038) );
  AOI220 U1020 ( .A(regs[113]), .B(n247), .C(regs[49]), .D(n205), .Q(n1275) );
  AOI220 U1021 ( .A(regs[600]), .B(n203), .C(regs[536]), .D(n204), .Q(n1402)
         );
  AOI221 U1022 ( .A(n1577), .B(n1015), .C(n1575), .D(n1014), .Q(n1016) );
  AOI221 U1023 ( .A(n1577), .B(n1059), .C(n1575), .D(n1058), .Q(n1060) );
  AOI221 U1024 ( .A(n1577), .B(n1257), .C(n1575), .D(n1256), .Q(n1258) );
  AOI221 U1025 ( .A(n1577), .B(n1235), .C(n1575), .D(n1234), .Q(n1236) );
  AOI220 U1026 ( .A(regs[116]), .B(n247), .C(regs[52]), .D(n205), .Q(n1341) );
  AOI221 U1027 ( .A(n1577), .B(n1125), .C(n1575), .D(n1124), .Q(n1126) );
  AOI221 U1028 ( .A(n1577), .B(n1081), .C(n1575), .D(n1080), .Q(n1082) );
  NOR31 U1029 ( .A(i_addr_Rs[0]), .B(n993), .C(n990), .Q(n1565) );
  NOR40 U1030 ( .A(n240), .B(n1586), .C(n1587), .D(n1583), .Q(n27) );
  NOR40 U1031 ( .A(n240), .B(i_addr_Rd[1]), .C(n1587), .D(n1583), .Q(n25) );
  NOR40 U1032 ( .A(n240), .B(n1586), .C(n1587), .D(n1588), .Q(n17) );
  NOR40 U1033 ( .A(n240), .B(i_addr_Rd[1]), .C(n1587), .D(n1588), .Q(n15) );
  NOR40 U1034 ( .A(i_addr_Rd[1]), .B(n240), .C(n1587), .D(n1592), .Q(n42) );
  NOR40 U1035 ( .A(i_addr_Rd[0]), .B(n240), .C(n1592), .D(n1586), .Q(n43) );
  NOR40 U1036 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n240), .D(n1582), .Q(
        n32) );
  NOR40 U1037 ( .A(i_addr_Rd[0]), .B(n240), .C(n1586), .D(n1582), .Q(n35) );
  NOR40 U1038 ( .A(n240), .B(i_addr_Rd[1]), .C(n1587), .D(n1582), .Q(n34) );
  BUF2 U1039 ( .A(n36), .Q(n252) );
  NOR40 U1040 ( .A(n240), .B(n1586), .C(n1587), .D(n1582), .Q(n36) );
  AOI220 U1041 ( .A(n244), .B(regs[838]), .C(n232), .D(regs[774]), .Q(n406) );
  AOI220 U1042 ( .A(n244), .B(regs[69]), .C(n232), .D(regs[5]), .Q(n398) );
  AOI220 U1043 ( .A(n244), .B(regs[581]), .C(n232), .D(regs[517]), .Q(n394) );
  AOI220 U1044 ( .A(n244), .B(regs[837]), .C(n232), .D(regs[773]), .Q(n384) );
  AOI220 U1045 ( .A(n244), .B(regs[95]), .C(n232), .D(regs[31]), .Q(n980) );
  AOI220 U1046 ( .A(n243), .B(regs[383]), .C(n206), .D(regs[319]), .Q(n961) );
  AOI220 U1047 ( .A(n243), .B(regs[361]), .C(n206), .D(regs[297]), .Q(n477) );
  AOI220 U1048 ( .A(n244), .B(regs[336]), .C(n232), .D(regs[272]), .Q(n630) );
  AOI220 U1049 ( .A(n244), .B(regs[580]), .C(n232), .D(regs[516]), .Q(n372) );
  AOI220 U1050 ( .A(n243), .B(regs[98]), .C(n206), .D(regs[34]), .Q(n333) );
  AOI220 U1051 ( .A(n243), .B(regs[610]), .C(n206), .D(regs[546]), .Q(n329) );
  AOI220 U1052 ( .A(regs[876]), .B(n247), .C(regs[812]), .D(n205), .Q(n1173)
         );
  AOI220 U1053 ( .A(regs[359]), .B(n247), .C(regs[295]), .D(n205), .Q(n1089)
         );
  AOI220 U1054 ( .A(regs[100]), .B(n247), .C(regs[36]), .D(n205), .Q(n1033) );
  AOI220 U1055 ( .A(regs[107]), .B(n247), .C(regs[43]), .D(n205), .Q(n1165) );
  AOI220 U1056 ( .A(regs[619]), .B(n247), .C(regs[555]), .D(n205), .Q(n1161)
         );
  AOI220 U1057 ( .A(regs[363]), .B(n247), .C(regs[299]), .D(n205), .Q(n1155)
         );
  AOI220 U1058 ( .A(regs[875]), .B(n247), .C(regs[811]), .D(n205), .Q(n1151)
         );
  AOI220 U1059 ( .A(regs[98]), .B(n247), .C(regs[34]), .D(n205), .Q(n1011) );
  AOI220 U1060 ( .A(regs[354]), .B(n247), .C(regs[290]), .D(n205), .Q(n1001)
         );
  AOI220 U1061 ( .A(regs[866]), .B(n247), .C(regs[802]), .D(n205), .Q(n997) );
  AOI220 U1062 ( .A(regs[101]), .B(n247), .C(regs[37]), .D(n205), .Q(n1055) );
  AOI220 U1063 ( .A(regs[613]), .B(n247), .C(regs[549]), .D(n205), .Q(n1051)
         );
  AOI220 U1064 ( .A(regs[357]), .B(n247), .C(regs[293]), .D(n205), .Q(n1045)
         );
  AOI220 U1065 ( .A(regs[869]), .B(n247), .C(regs[805]), .D(n205), .Q(n1041)
         );
  AOI220 U1066 ( .A(regs[102]), .B(n247), .C(regs[38]), .D(n205), .Q(n1077) );
  AOI220 U1067 ( .A(regs[870]), .B(n247), .C(regs[806]), .D(n205), .Q(n1063)
         );
  NOR40 U1068 ( .A(i_addr_Rd[0]), .B(n240), .C(n1586), .D(n1583), .Q(n26) );
  NOR40 U1069 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n240), .D(n1583), .Q(
        n23) );
  NOR40 U1070 ( .A(i_addr_Rd[0]), .B(n240), .C(n1586), .D(n1588), .Q(n16) );
  NOR40 U1071 ( .A(i_addr_Rd[0]), .B(i_addr_Rd[1]), .C(n240), .D(n1588), .Q(
        n13) );
  NOR40 U1072 ( .A(i_addr_Rd[1]), .B(i_addr_Rd[0]), .C(n240), .D(n1592), .Q(
        n41) );
  NAND22 U1073 ( .A(n933), .B(n932), .Q(o_data_Rt[29]) );
  AOI221 U1074 ( .A(n987), .B(n931), .C(n985), .D(n930), .Q(n932) );
  NAND41 U1075 ( .A(n929), .B(n928), .C(n927), .D(n926), .Q(n930) );
  NAND41 U1076 ( .A(n925), .B(n924), .C(n923), .D(n922), .Q(n931) );
  NAND41 U1077 ( .A(n919), .B(n918), .C(n917), .D(n916), .Q(n920) );
  NAND41 U1078 ( .A(n915), .B(n914), .C(n913), .D(n912), .Q(n921) );
  NAND22 U1079 ( .A(n427), .B(n426), .Q(o_data_Rt[6]) );
  NAND41 U1080 ( .A(n423), .B(n422), .C(n421), .D(n420), .Q(n424) );
  NAND41 U1081 ( .A(n419), .B(n418), .C(n417), .D(n416), .Q(n425) );
  NAND41 U1082 ( .A(n413), .B(n412), .C(n411), .D(n410), .Q(n414) );
  NAND41 U1083 ( .A(n409), .B(n408), .C(n407), .D(n406), .Q(n415) );
  NAND22 U1084 ( .A(n405), .B(n404), .Q(o_data_Rt[5]) );
  NAND41 U1085 ( .A(n401), .B(n400), .C(n399), .D(n398), .Q(n402) );
  NAND41 U1086 ( .A(n397), .B(n396), .C(n395), .D(n394), .Q(n403) );
  NAND41 U1087 ( .A(n391), .B(n390), .C(n389), .D(n388), .Q(n392) );
  NAND41 U1088 ( .A(n387), .B(n386), .C(n385), .D(n384), .Q(n393) );
  NAND41 U1089 ( .A(n983), .B(n982), .C(n981), .D(n980), .Q(n984) );
  NAND41 U1090 ( .A(n971), .B(n970), .C(n969), .D(n968), .Q(n986) );
  NAND41 U1091 ( .A(n963), .B(n962), .C(n961), .D(n960), .Q(n964) );
  NAND41 U1092 ( .A(n959), .B(n958), .C(n957), .D(n956), .Q(n966) );
  NAND22 U1093 ( .A(n845), .B(n844), .Q(o_data_Rt[25]) );
  AOI221 U1094 ( .A(n987), .B(n843), .C(n985), .D(n842), .Q(n844) );
  NAND41 U1095 ( .A(n841), .B(n840), .C(n839), .D(n838), .Q(n842) );
  NAND41 U1096 ( .A(n837), .B(n836), .C(n835), .D(n834), .Q(n843) );
  AOI221 U1097 ( .A(n967), .B(n833), .C(n965), .D(n832), .Q(n845) );
  NAND41 U1098 ( .A(n831), .B(n830), .C(n829), .D(n828), .Q(n832) );
  NAND41 U1099 ( .A(n827), .B(n826), .C(n825), .D(n824), .Q(n833) );
  NAND22 U1100 ( .A(n757), .B(n756), .Q(o_data_Rt[21]) );
  AOI221 U1101 ( .A(n987), .B(n755), .C(n985), .D(n754), .Q(n756) );
  NAND41 U1102 ( .A(n753), .B(n752), .C(n751), .D(n750), .Q(n754) );
  NAND41 U1103 ( .A(n749), .B(n748), .C(n747), .D(n746), .Q(n755) );
  NAND41 U1104 ( .A(n743), .B(n742), .C(n741), .D(n740), .Q(n744) );
  NAND41 U1105 ( .A(n739), .B(n738), .C(n737), .D(n736), .Q(n745) );
  NAND22 U1106 ( .A(n361), .B(n360), .Q(o_data_Rt[3]) );
  AOI221 U1107 ( .A(n987), .B(n359), .C(n985), .D(n358), .Q(n360) );
  NAND41 U1108 ( .A(n357), .B(n356), .C(n355), .D(n354), .Q(n358) );
  NAND41 U1109 ( .A(n353), .B(n352), .C(n351), .D(n350), .Q(n359) );
  NAND41 U1110 ( .A(n347), .B(n346), .C(n345), .D(n344), .Q(n348) );
  NAND41 U1111 ( .A(n343), .B(n342), .C(n341), .D(n340), .Q(n349) );
  NAND22 U1112 ( .A(n493), .B(n492), .Q(o_data_Rt[9]) );
  NAND41 U1113 ( .A(n489), .B(n488), .C(n487), .D(n486), .Q(n490) );
  NAND41 U1114 ( .A(n485), .B(n484), .C(n483), .D(n482), .Q(n491) );
  AOI221 U1115 ( .A(n241), .B(regs[713]), .C(n202), .D(regs[649]), .Q(n484) );
  NAND41 U1116 ( .A(n479), .B(n478), .C(n477), .D(n476), .Q(n480) );
  NAND41 U1117 ( .A(n475), .B(n474), .C(n473), .D(n472), .Q(n481) );
  NAND22 U1118 ( .A(n449), .B(n448), .Q(o_data_Rt[7]) );
  NAND41 U1119 ( .A(n445), .B(n444), .C(n443), .D(n442), .Q(n446) );
  NAND41 U1120 ( .A(n441), .B(n440), .C(n439), .D(n438), .Q(n447) );
  NAND41 U1121 ( .A(n435), .B(n434), .C(n433), .D(n432), .Q(n436) );
  NAND41 U1122 ( .A(n431), .B(n430), .C(n429), .D(n428), .Q(n437) );
  NAND22 U1123 ( .A(n471), .B(n470), .Q(o_data_Rt[8]) );
  NAND41 U1124 ( .A(n467), .B(n466), .C(n465), .D(n464), .Q(n468) );
  NAND41 U1125 ( .A(n463), .B(n462), .C(n461), .D(n460), .Q(n469) );
  NAND41 U1126 ( .A(n457), .B(n456), .C(n455), .D(n454), .Q(n458) );
  NAND41 U1127 ( .A(n453), .B(n452), .C(n451), .D(n450), .Q(n459) );
  NAND22 U1128 ( .A(n515), .B(n514), .Q(o_data_Rt[10]) );
  AOI221 U1129 ( .A(n987), .B(n513), .C(n985), .D(n512), .Q(n514) );
  NAND41 U1130 ( .A(n511), .B(n510), .C(n509), .D(n508), .Q(n512) );
  NAND41 U1131 ( .A(n507), .B(n506), .C(n505), .D(n504), .Q(n513) );
  NAND41 U1132 ( .A(n501), .B(n500), .C(n499), .D(n498), .Q(n502) );
  NAND41 U1133 ( .A(n497), .B(n496), .C(n495), .D(n494), .Q(n503) );
  NAND22 U1134 ( .A(n955), .B(n954), .Q(o_data_Rt[30]) );
  AOI221 U1135 ( .A(n987), .B(n953), .C(n985), .D(n952), .Q(n954) );
  NAND41 U1136 ( .A(n951), .B(n950), .C(n949), .D(n948), .Q(n952) );
  NAND41 U1137 ( .A(n947), .B(n946), .C(n945), .D(n944), .Q(n953) );
  NAND41 U1138 ( .A(n941), .B(n940), .C(n939), .D(n938), .Q(n942) );
  NAND41 U1139 ( .A(n937), .B(n936), .C(n935), .D(n934), .Q(n943) );
  NAND22 U1140 ( .A(n911), .B(n910), .Q(o_data_Rt[28]) );
  NAND41 U1141 ( .A(n907), .B(n906), .C(n905), .D(n904), .Q(n908) );
  NAND41 U1142 ( .A(n903), .B(n902), .C(n901), .D(n900), .Q(n909) );
  NAND41 U1143 ( .A(n897), .B(n896), .C(n895), .D(n894), .Q(n898) );
  NAND41 U1144 ( .A(n893), .B(n892), .C(n891), .D(n890), .Q(n899) );
  AOI221 U1145 ( .A(n201), .B(regs[1020]), .C(n198), .D(regs[956]), .Q(n893)
         );
  NAND22 U1146 ( .A(n559), .B(n558), .Q(o_data_Rt[12]) );
  AOI221 U1147 ( .A(n987), .B(n557), .C(n985), .D(n556), .Q(n558) );
  NAND41 U1148 ( .A(n555), .B(n554), .C(n553), .D(n552), .Q(n556) );
  NAND41 U1149 ( .A(n551), .B(n550), .C(n549), .D(n548), .Q(n557) );
  NAND41 U1150 ( .A(n545), .B(n544), .C(n543), .D(n542), .Q(n546) );
  NAND41 U1151 ( .A(n541), .B(n540), .C(n539), .D(n538), .Q(n547) );
  NAND22 U1152 ( .A(n867), .B(n866), .Q(o_data_Rt[26]) );
  AOI221 U1153 ( .A(n987), .B(n865), .C(n985), .D(n864), .Q(n866) );
  NAND41 U1154 ( .A(n863), .B(n862), .C(n861), .D(n860), .Q(n864) );
  NAND41 U1155 ( .A(n859), .B(n858), .C(n857), .D(n856), .Q(n865) );
  AOI221 U1156 ( .A(n201), .B(regs[762]), .C(n198), .D(regs[698]), .Q(n859) );
  AOI221 U1157 ( .A(n967), .B(n855), .C(n965), .D(n854), .Q(n867) );
  NAND41 U1158 ( .A(n853), .B(n852), .C(n851), .D(n850), .Q(n854) );
  NAND41 U1159 ( .A(n849), .B(n848), .C(n847), .D(n846), .Q(n855) );
  NAND22 U1160 ( .A(n801), .B(n800), .Q(o_data_Rt[23]) );
  AOI221 U1161 ( .A(n987), .B(n799), .C(n985), .D(n798), .Q(n800) );
  NAND41 U1162 ( .A(n797), .B(n796), .C(n795), .D(n794), .Q(n798) );
  NAND41 U1163 ( .A(n793), .B(n792), .C(n791), .D(n790), .Q(n799) );
  NAND41 U1164 ( .A(n787), .B(n786), .C(n785), .D(n784), .Q(n788) );
  NAND41 U1165 ( .A(n783), .B(n782), .C(n781), .D(n780), .Q(n789) );
  NAND22 U1166 ( .A(n889), .B(n888), .Q(o_data_Rt[27]) );
  AOI221 U1167 ( .A(n987), .B(n887), .C(n985), .D(n886), .Q(n888) );
  NAND41 U1168 ( .A(n885), .B(n884), .C(n883), .D(n882), .Q(n886) );
  AOI221 U1169 ( .A(n201), .B(regs[251]), .C(n198), .D(regs[187]), .Q(n885) );
  NAND41 U1170 ( .A(n881), .B(n880), .C(n879), .D(n878), .Q(n887) );
  AOI221 U1171 ( .A(n967), .B(n877), .C(n965), .D(n876), .Q(n889) );
  NAND41 U1172 ( .A(n875), .B(n874), .C(n873), .D(n872), .Q(n876) );
  AOI221 U1173 ( .A(n201), .B(regs[507]), .C(n198), .D(regs[443]), .Q(n875) );
  NAND41 U1174 ( .A(n871), .B(n870), .C(n869), .D(n868), .Q(n877) );
  NAND22 U1175 ( .A(n823), .B(n822), .Q(o_data_Rt[24]) );
  AOI221 U1176 ( .A(n987), .B(n821), .C(n985), .D(n820), .Q(n822) );
  NAND41 U1177 ( .A(n819), .B(n818), .C(n817), .D(n816), .Q(n820) );
  NAND41 U1178 ( .A(n815), .B(n814), .C(n813), .D(n812), .Q(n821) );
  NAND41 U1179 ( .A(n809), .B(n808), .C(n807), .D(n806), .Q(n810) );
  NAND41 U1180 ( .A(n805), .B(n804), .C(n803), .D(n802), .Q(n811) );
  NAND22 U1181 ( .A(n779), .B(n778), .Q(o_data_Rt[22]) );
  AOI221 U1182 ( .A(n987), .B(n777), .C(n985), .D(n776), .Q(n778) );
  NAND41 U1183 ( .A(n775), .B(n774), .C(n773), .D(n772), .Q(n776) );
  NAND41 U1184 ( .A(n771), .B(n770), .C(n769), .D(n768), .Q(n777) );
  NAND41 U1185 ( .A(n765), .B(n764), .C(n763), .D(n762), .Q(n766) );
  AOI221 U1186 ( .A(n201), .B(regs[502]), .C(n198), .D(regs[438]), .Q(n765) );
  NAND41 U1187 ( .A(n761), .B(n760), .C(n759), .D(n758), .Q(n767) );
  NAND22 U1188 ( .A(n647), .B(n646), .Q(o_data_Rt[16]) );
  NAND41 U1189 ( .A(n643), .B(n642), .C(n641), .D(n640), .Q(n644) );
  NAND41 U1190 ( .A(n639), .B(n638), .C(n637), .D(n636), .Q(n645) );
  AOI221 U1191 ( .A(n967), .B(n635), .C(n965), .D(n634), .Q(n647) );
  NAND41 U1192 ( .A(n633), .B(n632), .C(n631), .D(n630), .Q(n634) );
  NAND41 U1193 ( .A(n629), .B(n628), .C(n627), .D(n626), .Q(n635) );
  NAND22 U1194 ( .A(n295), .B(n294), .Q(o_data_Rt[0]) );
  NAND41 U1195 ( .A(n291), .B(n290), .C(n289), .D(n288), .Q(n292) );
  NAND41 U1196 ( .A(n287), .B(n286), .C(n285), .D(n284), .Q(n293) );
  NAND41 U1197 ( .A(n280), .B(n279), .C(n278), .D(n277), .Q(n281) );
  NAND41 U1198 ( .A(n275), .B(n274), .C(n273), .D(n272), .Q(n282) );
  NAND22 U1199 ( .A(n317), .B(n316), .Q(o_data_Rt[1]) );
  AOI221 U1200 ( .A(n987), .B(n315), .C(n985), .D(n314), .Q(n316) );
  NAND41 U1201 ( .A(n313), .B(n312), .C(n311), .D(n310), .Q(n314) );
  NAND41 U1202 ( .A(n309), .B(n308), .C(n307), .D(n306), .Q(n315) );
  NAND41 U1203 ( .A(n303), .B(n302), .C(n301), .D(n300), .Q(n304) );
  NAND41 U1204 ( .A(n299), .B(n298), .C(n297), .D(n296), .Q(n305) );
  NAND22 U1205 ( .A(n625), .B(n624), .Q(o_data_Rt[15]) );
  NAND41 U1206 ( .A(n621), .B(n620), .C(n619), .D(n618), .Q(n622) );
  NAND41 U1207 ( .A(n617), .B(n616), .C(n615), .D(n614), .Q(n623) );
  NAND41 U1208 ( .A(n611), .B(n610), .C(n609), .D(n608), .Q(n612) );
  NAND41 U1209 ( .A(n607), .B(n606), .C(n605), .D(n604), .Q(n613) );
  NAND22 U1210 ( .A(n581), .B(n580), .Q(o_data_Rt[13]) );
  AOI221 U1211 ( .A(n987), .B(n579), .C(n985), .D(n578), .Q(n580) );
  NAND41 U1212 ( .A(n577), .B(n576), .C(n575), .D(n574), .Q(n578) );
  NAND41 U1213 ( .A(n573), .B(n572), .C(n571), .D(n570), .Q(n579) );
  NAND41 U1214 ( .A(n567), .B(n566), .C(n565), .D(n564), .Q(n568) );
  NAND41 U1215 ( .A(n563), .B(n562), .C(n561), .D(n560), .Q(n569) );
  NAND22 U1216 ( .A(n383), .B(n382), .Q(o_data_Rt[4]) );
  AOI221 U1217 ( .A(n987), .B(n381), .C(n985), .D(n380), .Q(n382) );
  NAND41 U1218 ( .A(n379), .B(n378), .C(n377), .D(n376), .Q(n380) );
  NAND41 U1219 ( .A(n375), .B(n374), .C(n373), .D(n372), .Q(n381) );
  NAND41 U1220 ( .A(n369), .B(n368), .C(n367), .D(n366), .Q(n370) );
  NAND41 U1221 ( .A(n365), .B(n364), .C(n363), .D(n362), .Q(n371) );
  NAND22 U1222 ( .A(n669), .B(n668), .Q(o_data_Rt[17]) );
  NAND41 U1223 ( .A(n665), .B(n664), .C(n663), .D(n662), .Q(n666) );
  NAND41 U1224 ( .A(n661), .B(n660), .C(n659), .D(n658), .Q(n667) );
  AOI221 U1225 ( .A(n967), .B(n657), .C(n965), .D(n656), .Q(n669) );
  NAND41 U1226 ( .A(n655), .B(n654), .C(n653), .D(n652), .Q(n656) );
  NAND41 U1227 ( .A(n651), .B(n650), .C(n649), .D(n648), .Q(n657) );
  NAND22 U1228 ( .A(n339), .B(n338), .Q(o_data_Rt[2]) );
  NAND41 U1229 ( .A(n335), .B(n334), .C(n333), .D(n332), .Q(n336) );
  NAND41 U1230 ( .A(n331), .B(n330), .C(n329), .D(n328), .Q(n337) );
  NAND41 U1231 ( .A(n325), .B(n324), .C(n323), .D(n322), .Q(n326) );
  NAND41 U1232 ( .A(n321), .B(n320), .C(n319), .D(n318), .Q(n327) );
  NAND22 U1233 ( .A(n537), .B(n536), .Q(o_data_Rt[11]) );
  AOI221 U1234 ( .A(n987), .B(n535), .C(n985), .D(n534), .Q(n536) );
  NAND41 U1235 ( .A(n533), .B(n532), .C(n531), .D(n530), .Q(n534) );
  NAND41 U1236 ( .A(n529), .B(n528), .C(n527), .D(n526), .Q(n535) );
  NAND41 U1237 ( .A(n523), .B(n522), .C(n521), .D(n520), .Q(n524) );
  NAND41 U1238 ( .A(n519), .B(n518), .C(n517), .D(n516), .Q(n525) );
  NAND22 U1239 ( .A(n603), .B(n602), .Q(o_data_Rt[14]) );
  AOI221 U1240 ( .A(n987), .B(n601), .C(n985), .D(n600), .Q(n602) );
  NAND41 U1241 ( .A(n599), .B(n598), .C(n597), .D(n596), .Q(n600) );
  NAND41 U1242 ( .A(n595), .B(n594), .C(n593), .D(n592), .Q(n601) );
  NAND41 U1243 ( .A(n589), .B(n588), .C(n587), .D(n586), .Q(n590) );
  AOI221 U1244 ( .A(n244), .B(regs[334]), .C(n232), .D(regs[270]), .Q(n586) );
  NAND41 U1245 ( .A(n585), .B(n584), .C(n583), .D(n582), .Q(n591) );
  NAND22 U1246 ( .A(n691), .B(n690), .Q(o_data_Rt[18]) );
  AOI221 U1247 ( .A(n987), .B(n689), .C(n985), .D(n688), .Q(n690) );
  NAND41 U1248 ( .A(n687), .B(n686), .C(n685), .D(n684), .Q(n688) );
  NAND41 U1249 ( .A(n683), .B(n682), .C(n681), .D(n680), .Q(n689) );
  NAND41 U1250 ( .A(n677), .B(n676), .C(n675), .D(n674), .Q(n678) );
  AOI221 U1251 ( .A(n244), .B(regs[338]), .C(n232), .D(regs[274]), .Q(n674) );
  NAND41 U1252 ( .A(n673), .B(n672), .C(n671), .D(n670), .Q(n679) );
  NAND22 U1253 ( .A(n713), .B(n712), .Q(o_data_Rt[19]) );
  AOI221 U1254 ( .A(n987), .B(n711), .C(n985), .D(n710), .Q(n712) );
  NAND41 U1255 ( .A(n709), .B(n708), .C(n707), .D(n706), .Q(n710) );
  NAND41 U1256 ( .A(n705), .B(n704), .C(n703), .D(n702), .Q(n711) );
  AOI221 U1257 ( .A(n244), .B(regs[595]), .C(n232), .D(regs[531]), .Q(n702) );
  NAND41 U1258 ( .A(n699), .B(n698), .C(n697), .D(n696), .Q(n700) );
  NAND41 U1259 ( .A(n695), .B(n694), .C(n693), .D(n692), .Q(n701) );
  AOI221 U1260 ( .A(n244), .B(regs[851]), .C(n232), .D(regs[787]), .Q(n692) );
  NAND22 U1261 ( .A(n735), .B(n734), .Q(o_data_Rt[20]) );
  AOI221 U1262 ( .A(n987), .B(n733), .C(n985), .D(n732), .Q(n734) );
  NAND41 U1263 ( .A(n731), .B(n730), .C(n729), .D(n728), .Q(n732) );
  NAND41 U1264 ( .A(n727), .B(n726), .C(n725), .D(n724), .Q(n733) );
  AOI221 U1265 ( .A(n967), .B(n723), .C(n965), .D(n722), .Q(n735) );
  NAND41 U1266 ( .A(n721), .B(n720), .C(n719), .D(n718), .Q(n722) );
  NAND41 U1267 ( .A(n717), .B(n716), .C(n715), .D(n714), .Q(n723) );
  NAND22 U1268 ( .A(n1149), .B(n1148), .Q(o_data_Rs[9]) );
  NAND41 U1269 ( .A(n1145), .B(n1144), .C(n1143), .D(n1142), .Q(n1146) );
  NAND41 U1270 ( .A(n1141), .B(n1140), .C(n1139), .D(n1138), .Q(n1147) );
  AOI221 U1271 ( .A(n1557), .B(n1137), .C(n1555), .D(n1136), .Q(n1149) );
  NAND41 U1272 ( .A(n1135), .B(n1134), .C(n1133), .D(n1132), .Q(n1136) );
  NAND41 U1273 ( .A(n1131), .B(n1130), .C(n1129), .D(n1128), .Q(n1137) );
  NAND22 U1274 ( .A(n1457), .B(n1456), .Q(o_data_Rs[26]) );
  AOI221 U1275 ( .A(n1577), .B(n1455), .C(n1575), .D(n1454), .Q(n1456) );
  NAND41 U1276 ( .A(n1453), .B(n1452), .C(n1451), .D(n1450), .Q(n1454) );
  NAND41 U1277 ( .A(n1449), .B(n1448), .C(n1447), .D(n1446), .Q(n1455) );
  AOI221 U1278 ( .A(n1557), .B(n1445), .C(n1555), .D(n1444), .Q(n1457) );
  NAND41 U1279 ( .A(n1443), .B(n1442), .C(n1441), .D(n1440), .Q(n1444) );
  NAND41 U1280 ( .A(n1439), .B(n1438), .C(n1437), .D(n1436), .Q(n1445) );
  NAND22 U1281 ( .A(n1193), .B(n1192), .Q(o_data_Rs[12]) );
  AOI221 U1282 ( .A(n1577), .B(n1191), .C(n1575), .D(n1190), .Q(n1192) );
  NAND41 U1283 ( .A(n1189), .B(n1188), .C(n1187), .D(n1186), .Q(n1190) );
  NAND41 U1284 ( .A(n1185), .B(n1184), .C(n1183), .D(n1182), .Q(n1191) );
  AOI221 U1285 ( .A(n1557), .B(n1181), .C(n1555), .D(n1180), .Q(n1193) );
  NAND41 U1286 ( .A(n1179), .B(n1178), .C(n1177), .D(n1176), .Q(n1180) );
  NAND41 U1287 ( .A(n1175), .B(n1174), .C(n1173), .D(n1172), .Q(n1181) );
  NAND22 U1288 ( .A(n1523), .B(n1522), .Q(o_data_Rs[29]) );
  AOI221 U1289 ( .A(n1577), .B(n1521), .C(n1575), .D(n1520), .Q(n1522) );
  NAND41 U1290 ( .A(n1519), .B(n1518), .C(n1517), .D(n1516), .Q(n1520) );
  NAND41 U1291 ( .A(n1515), .B(n1514), .C(n1513), .D(n1512), .Q(n1521) );
  AOI221 U1292 ( .A(n1557), .B(n1511), .C(n1555), .D(n1510), .Q(n1523) );
  NAND41 U1293 ( .A(n1509), .B(n1508), .C(n1507), .D(n1506), .Q(n1510) );
  NAND41 U1294 ( .A(n1505), .B(n1504), .C(n1503), .D(n1502), .Q(n1511) );
  NAND22 U1295 ( .A(n1105), .B(n1104), .Q(o_data_Rs[7]) );
  AOI221 U1296 ( .A(n1577), .B(n1103), .C(n1575), .D(n1102), .Q(n1104) );
  NAND41 U1297 ( .A(n1101), .B(n1100), .C(n1099), .D(n1098), .Q(n1102) );
  NAND41 U1298 ( .A(n1097), .B(n1096), .C(n1095), .D(n1094), .Q(n1103) );
  AOI221 U1299 ( .A(n1557), .B(n1093), .C(n1555), .D(n1092), .Q(n1105) );
  NAND41 U1300 ( .A(n1091), .B(n1090), .C(n1089), .D(n1088), .Q(n1092) );
  NAND41 U1301 ( .A(n1087), .B(n1086), .C(n1085), .D(n1084), .Q(n1093) );
  NAND22 U1302 ( .A(n1369), .B(n1368), .Q(o_data_Rs[22]) );
  AOI221 U1303 ( .A(n1577), .B(n1367), .C(n1575), .D(n1366), .Q(n1368) );
  NAND41 U1304 ( .A(n1365), .B(n1364), .C(n1363), .D(n1362), .Q(n1366) );
  NAND41 U1305 ( .A(n1361), .B(n1360), .C(n1359), .D(n1358), .Q(n1367) );
  AOI221 U1306 ( .A(n1557), .B(n1357), .C(n1555), .D(n1356), .Q(n1369) );
  NAND41 U1307 ( .A(n1355), .B(n1354), .C(n1353), .D(n1352), .Q(n1356) );
  NAND41 U1308 ( .A(n1351), .B(n1350), .C(n1349), .D(n1348), .Q(n1357) );
  NAND22 U1309 ( .A(n1215), .B(n1214), .Q(o_data_Rs[13]) );
  AOI221 U1310 ( .A(n1577), .B(n1213), .C(n1575), .D(n1212), .Q(n1214) );
  NAND41 U1311 ( .A(n1211), .B(n1210), .C(n1209), .D(n1208), .Q(n1212) );
  NAND41 U1312 ( .A(n1207), .B(n1206), .C(n1205), .D(n1204), .Q(n1213) );
  NAND41 U1313 ( .A(n1201), .B(n1200), .C(n1199), .D(n1198), .Q(n1202) );
  NAND41 U1314 ( .A(n1197), .B(n1196), .C(n1195), .D(n1194), .Q(n1203) );
  NAND22 U1315 ( .A(n1479), .B(n1478), .Q(o_data_Rs[27]) );
  AOI221 U1316 ( .A(n1577), .B(n1477), .C(n1575), .D(n1476), .Q(n1478) );
  NAND41 U1317 ( .A(n1475), .B(n1474), .C(n1473), .D(n1472), .Q(n1476) );
  NAND41 U1318 ( .A(n1471), .B(n1470), .C(n1469), .D(n1468), .Q(n1477) );
  AOI221 U1319 ( .A(n1557), .B(n1467), .C(n1555), .D(n1466), .Q(n1479) );
  NAND41 U1320 ( .A(n1465), .B(n1464), .C(n1463), .D(n1462), .Q(n1466) );
  NAND41 U1321 ( .A(n1461), .B(n1460), .C(n1459), .D(n1458), .Q(n1467) );
  NAND22 U1322 ( .A(n1325), .B(n1324), .Q(o_data_Rs[19]) );
  AOI221 U1323 ( .A(n1577), .B(n1323), .C(n1575), .D(n1322), .Q(n1324) );
  NAND41 U1324 ( .A(n1321), .B(n1320), .C(n1319), .D(n1318), .Q(n1322) );
  NAND41 U1325 ( .A(n1317), .B(n1316), .C(n1315), .D(n1314), .Q(n1323) );
  AOI221 U1326 ( .A(n1557), .B(n1313), .C(n1555), .D(n1312), .Q(n1325) );
  NAND41 U1327 ( .A(n1311), .B(n1310), .C(n1309), .D(n1308), .Q(n1312) );
  NAND41 U1328 ( .A(n1307), .B(n1306), .C(n1305), .D(n1304), .Q(n1313) );
  NAND22 U1329 ( .A(n1501), .B(n1500), .Q(o_data_Rs[28]) );
  AOI221 U1330 ( .A(n1577), .B(n1499), .C(n1575), .D(n1498), .Q(n1500) );
  NAND41 U1331 ( .A(n1497), .B(n1496), .C(n1495), .D(n1494), .Q(n1498) );
  NAND41 U1332 ( .A(n1493), .B(n1492), .C(n1491), .D(n1490), .Q(n1499) );
  AOI221 U1333 ( .A(n1557), .B(n1489), .C(n1555), .D(n1488), .Q(n1501) );
  NAND41 U1334 ( .A(n1487), .B(n1486), .C(n1485), .D(n1484), .Q(n1488) );
  NAND41 U1335 ( .A(n1483), .B(n1482), .C(n1481), .D(n1480), .Q(n1489) );
  NAND22 U1336 ( .A(n1303), .B(n1302), .Q(o_data_Rs[18]) );
  AOI221 U1337 ( .A(n1577), .B(n1301), .C(n1575), .D(n1300), .Q(n1302) );
  NAND41 U1338 ( .A(n1299), .B(n1298), .C(n1297), .D(n1296), .Q(n1300) );
  NAND41 U1339 ( .A(n1295), .B(n1294), .C(n1293), .D(n1292), .Q(n1301) );
  AOI221 U1340 ( .A(n1557), .B(n1291), .C(n1555), .D(n1290), .Q(n1303) );
  NAND41 U1341 ( .A(n1289), .B(n1288), .C(n1287), .D(n1286), .Q(n1290) );
  NAND41 U1342 ( .A(n1285), .B(n1284), .C(n1283), .D(n1282), .Q(n1291) );
  NAND22 U1343 ( .A(n1039), .B(n1038), .Q(o_data_Rs[4]) );
  NAND41 U1344 ( .A(n1035), .B(n1034), .C(n1033), .D(n1032), .Q(n1036) );
  NAND41 U1345 ( .A(n1031), .B(n1030), .C(n1029), .D(n1028), .Q(n1037) );
  AOI221 U1346 ( .A(n1557), .B(n1027), .C(n1555), .D(n1026), .Q(n1039) );
  NAND41 U1347 ( .A(n1025), .B(n1024), .C(n1023), .D(n1022), .Q(n1026) );
  NAND41 U1348 ( .A(n1021), .B(n1020), .C(n1019), .D(n1018), .Q(n1027) );
  NAND22 U1349 ( .A(n1281), .B(n1280), .Q(o_data_Rs[17]) );
  AOI221 U1350 ( .A(n1577), .B(n1279), .C(n1575), .D(n1278), .Q(n1280) );
  NAND41 U1351 ( .A(n1277), .B(n1276), .C(n1275), .D(n1274), .Q(n1278) );
  NAND41 U1352 ( .A(n1273), .B(n1272), .C(n1271), .D(n1270), .Q(n1279) );
  AOI221 U1353 ( .A(n1557), .B(n1269), .C(n1555), .D(n1268), .Q(n1281) );
  NAND41 U1354 ( .A(n1267), .B(n1266), .C(n1265), .D(n1264), .Q(n1268) );
  NAND41 U1355 ( .A(n1263), .B(n1262), .C(n1261), .D(n1260), .Q(n1269) );
  NAND22 U1356 ( .A(n1413), .B(n1412), .Q(o_data_Rs[24]) );
  AOI221 U1357 ( .A(n1577), .B(n1411), .C(n1575), .D(n1410), .Q(n1412) );
  NAND41 U1358 ( .A(n1409), .B(n1408), .C(n1407), .D(n1406), .Q(n1410) );
  NAND41 U1359 ( .A(n1405), .B(n1404), .C(n1403), .D(n1402), .Q(n1411) );
  AOI221 U1360 ( .A(n1557), .B(n1401), .C(n1555), .D(n1400), .Q(n1413) );
  NAND41 U1361 ( .A(n1399), .B(n1398), .C(n1397), .D(n1396), .Q(n1400) );
  NAND41 U1362 ( .A(n1395), .B(n1394), .C(n1393), .D(n1392), .Q(n1401) );
  NAND22 U1363 ( .A(n1391), .B(n1390), .Q(o_data_Rs[23]) );
  AOI221 U1364 ( .A(n1577), .B(n1389), .C(n1575), .D(n1388), .Q(n1390) );
  NAND41 U1365 ( .A(n1387), .B(n1386), .C(n1385), .D(n1384), .Q(n1388) );
  NAND41 U1366 ( .A(n1383), .B(n1382), .C(n1381), .D(n1380), .Q(n1389) );
  AOI221 U1367 ( .A(n1557), .B(n1379), .C(n1555), .D(n1378), .Q(n1391) );
  NAND41 U1368 ( .A(n1377), .B(n1376), .C(n1375), .D(n1374), .Q(n1378) );
  NAND41 U1369 ( .A(n1373), .B(n1372), .C(n1371), .D(n1370), .Q(n1379) );
  NAND22 U1370 ( .A(n1171), .B(n1170), .Q(o_data_Rs[11]) );
  AOI221 U1371 ( .A(n1577), .B(n1169), .C(n1575), .D(n1168), .Q(n1170) );
  NAND41 U1372 ( .A(n1167), .B(n1166), .C(n1165), .D(n1164), .Q(n1168) );
  NAND41 U1373 ( .A(n1163), .B(n1162), .C(n1161), .D(n1160), .Q(n1169) );
  AOI221 U1374 ( .A(n1557), .B(n1159), .C(n1555), .D(n1158), .Q(n1171) );
  NAND41 U1375 ( .A(n1157), .B(n1156), .C(n1155), .D(n1154), .Q(n1158) );
  NAND41 U1376 ( .A(n1153), .B(n1152), .C(n1151), .D(n1150), .Q(n1159) );
  NAND22 U1377 ( .A(n1017), .B(n1016), .Q(o_data_Rs[2]) );
  NAND41 U1378 ( .A(n1013), .B(n1012), .C(n1011), .D(n1010), .Q(n1014) );
  NAND41 U1379 ( .A(n1009), .B(n1008), .C(n1007), .D(n1006), .Q(n1015) );
  AOI221 U1380 ( .A(n1557), .B(n1005), .C(n1555), .D(n1004), .Q(n1017) );
  NAND41 U1381 ( .A(n1003), .B(n1002), .C(n1001), .D(n1000), .Q(n1004) );
  NAND41 U1382 ( .A(n999), .B(n998), .C(n997), .D(n996), .Q(n1005) );
  NAND22 U1383 ( .A(n1061), .B(n1060), .Q(o_data_Rs[5]) );
  NAND41 U1384 ( .A(n1057), .B(n1056), .C(n1055), .D(n1054), .Q(n1058) );
  NAND41 U1385 ( .A(n1053), .B(n1052), .C(n1051), .D(n1050), .Q(n1059) );
  AOI221 U1386 ( .A(n1557), .B(n1049), .C(n1555), .D(n1048), .Q(n1061) );
  NAND41 U1387 ( .A(n1047), .B(n1046), .C(n1045), .D(n1044), .Q(n1048) );
  NAND41 U1388 ( .A(n1043), .B(n1042), .C(n1041), .D(n1040), .Q(n1049) );
  NAND22 U1389 ( .A(n1259), .B(n1258), .Q(o_data_Rs[16]) );
  NAND41 U1390 ( .A(n1255), .B(n1254), .C(n1253), .D(n1252), .Q(n1256) );
  NAND41 U1391 ( .A(n1251), .B(n1250), .C(n1249), .D(n1248), .Q(n1257) );
  AOI221 U1392 ( .A(n1557), .B(n1247), .C(n1555), .D(n1246), .Q(n1259) );
  NAND41 U1393 ( .A(n1245), .B(n1244), .C(n1243), .D(n1242), .Q(n1246) );
  NAND41 U1394 ( .A(n1241), .B(n1240), .C(n1239), .D(n1238), .Q(n1247) );
  NAND22 U1395 ( .A(n1237), .B(n1236), .Q(o_data_Rs[15]) );
  NAND41 U1396 ( .A(n1233), .B(n1232), .C(n1231), .D(n1230), .Q(n1234) );
  NAND41 U1397 ( .A(n1229), .B(n1228), .C(n1227), .D(n1226), .Q(n1235) );
  AOI221 U1398 ( .A(n1557), .B(n1225), .C(n1555), .D(n1224), .Q(n1237) );
  NAND41 U1399 ( .A(n1223), .B(n1222), .C(n1221), .D(n1220), .Q(n1224) );
  NAND41 U1400 ( .A(n1219), .B(n1218), .C(n1217), .D(n1216), .Q(n1225) );
  NAND22 U1401 ( .A(n1347), .B(n1346), .Q(o_data_Rs[20]) );
  AOI221 U1402 ( .A(n1577), .B(n1345), .C(n1575), .D(n1344), .Q(n1346) );
  NAND41 U1403 ( .A(n1343), .B(n1342), .C(n1341), .D(n1340), .Q(n1344) );
  NAND41 U1404 ( .A(n1339), .B(n1338), .C(n1337), .D(n1336), .Q(n1345) );
  AOI221 U1405 ( .A(n1557), .B(n1335), .C(n1555), .D(n1334), .Q(n1347) );
  NAND41 U1406 ( .A(n1333), .B(n1332), .C(n1331), .D(n1330), .Q(n1334) );
  NAND41 U1407 ( .A(n1329), .B(n1328), .C(n1327), .D(n1326), .Q(n1335) );
  NAND22 U1408 ( .A(n1435), .B(n1434), .Q(o_data_Rs[25]) );
  AOI221 U1409 ( .A(n1577), .B(n1433), .C(n1575), .D(n1432), .Q(n1434) );
  NAND41 U1410 ( .A(n1431), .B(n1430), .C(n1429), .D(n1428), .Q(n1432) );
  NAND41 U1411 ( .A(n1427), .B(n1426), .C(n1425), .D(n1424), .Q(n1433) );
  AOI221 U1412 ( .A(n1557), .B(n1423), .C(n1555), .D(n1422), .Q(n1435) );
  NAND41 U1413 ( .A(n1421), .B(n1420), .C(n1419), .D(n1418), .Q(n1422) );
  NAND41 U1414 ( .A(n1417), .B(n1416), .C(n1415), .D(n1414), .Q(n1423) );
  NAND22 U1415 ( .A(n1127), .B(n1126), .Q(o_data_Rs[8]) );
  NAND41 U1416 ( .A(n1123), .B(n1122), .C(n1121), .D(n1120), .Q(n1124) );
  NAND41 U1417 ( .A(n1119), .B(n1118), .C(n1117), .D(n1116), .Q(n1125) );
  AOI221 U1418 ( .A(n1557), .B(n1115), .C(n1555), .D(n1114), .Q(n1127) );
  NAND41 U1419 ( .A(n1113), .B(n1112), .C(n1111), .D(n1110), .Q(n1114) );
  NAND41 U1420 ( .A(n1109), .B(n1108), .C(n1107), .D(n1106), .Q(n1115) );
  NAND22 U1421 ( .A(n1083), .B(n1082), .Q(o_data_Rs[6]) );
  NAND41 U1422 ( .A(n1079), .B(n1078), .C(n1077), .D(n1076), .Q(n1080) );
  NAND41 U1423 ( .A(n1075), .B(n1074), .C(n1073), .D(n1072), .Q(n1081) );
  AOI221 U1424 ( .A(n1557), .B(n1071), .C(n1555), .D(n1070), .Q(n1083) );
  NAND41 U1425 ( .A(n1069), .B(n1068), .C(n1067), .D(n1066), .Q(n1070) );
  NAND41 U1426 ( .A(n1065), .B(n1064), .C(n1063), .D(n1062), .Q(n1071) );
  NAND22 U1427 ( .A(n1545), .B(n1544), .Q(o_data_Rs[30]) );
  AOI221 U1428 ( .A(n1577), .B(n1543), .C(n1575), .D(n1542), .Q(n1544) );
  NAND41 U1429 ( .A(n1541), .B(n1540), .C(n1539), .D(n1538), .Q(n1542) );
  NAND41 U1430 ( .A(n1537), .B(n1536), .C(n1535), .D(n1534), .Q(n1543) );
  AOI221 U1431 ( .A(n1557), .B(n1533), .C(n1555), .D(n1532), .Q(n1545) );
  NAND41 U1432 ( .A(n1531), .B(n1530), .C(n1529), .D(n1528), .Q(n1532) );
  NAND41 U1433 ( .A(n1527), .B(n1526), .C(n1525), .D(n1524), .Q(n1533) );
  NAND22 U1434 ( .A(n1579), .B(n1578), .Q(o_data_Rs[31]) );
  AOI221 U1435 ( .A(n1577), .B(n1576), .C(n1575), .D(n1574), .Q(n1578) );
  NAND41 U1436 ( .A(n1573), .B(n1572), .C(n1571), .D(n1570), .Q(n1574) );
  NAND41 U1437 ( .A(n1561), .B(n1560), .C(n1559), .D(n1558), .Q(n1576) );
  AOI221 U1438 ( .A(n1557), .B(n1556), .C(n1555), .D(n1554), .Q(n1579) );
  NAND41 U1439 ( .A(n1553), .B(n1552), .C(n1551), .D(n1550), .Q(n1554) );
  NAND41 U1440 ( .A(n1549), .B(n1548), .C(n1547), .D(n1546), .Q(n1556) );
  NOR21 U1441 ( .A(n1589), .B(n1588), .Q(n22) );
  NOR21 U1442 ( .A(n1590), .B(n1588), .Q(n21) );
  NOR21 U1443 ( .A(n1591), .B(n1588), .Q(n20) );
  NOR21 U1444 ( .A(n1585), .B(n1588), .Q(n18) );
  BUF2 U1445 ( .A(n975), .Q(n242) );
  BUF2 U1446 ( .A(n975), .Q(n241) );
  AOI220 U1447 ( .A(n201), .B(regs[480]), .C(n972), .D(regs[416]), .Q(n280) );
  AOI220 U1448 ( .A(regs[608]), .B(n243), .C(regs[544]), .D(n206), .Q(n285) );
  AOI220 U1449 ( .A(n973), .B(regs[224]), .C(n972), .D(regs[160]), .Q(n291) );
  AOI220 U1450 ( .A(n973), .B(regs[993]), .C(n972), .D(regs[929]), .Q(n299) );
  AOI220 U1451 ( .A(n201), .B(regs[481]), .C(n972), .D(regs[417]), .Q(n303) );
  AOI220 U1452 ( .A(n201), .B(regs[737]), .C(n972), .D(regs[673]), .Q(n309) );
  AOI220 U1453 ( .A(n201), .B(regs[225]), .C(n972), .D(regs[161]), .Q(n313) );
  AOI220 U1454 ( .A(n201), .B(regs[994]), .C(n972), .D(regs[930]), .Q(n321) );
  AOI220 U1455 ( .A(n201), .B(regs[482]), .C(n972), .D(regs[418]), .Q(n325) );
  AOI220 U1456 ( .A(n243), .B(regs[867]), .C(n206), .D(regs[803]), .Q(n341) );
  AOI220 U1457 ( .A(n243), .B(regs[355]), .C(n206), .D(regs[291]), .Q(n345) );
  AOI220 U1458 ( .A(n242), .B(regs[707]), .C(n974), .D(regs[643]), .Q(n352) );
  AOI220 U1459 ( .A(n243), .B(regs[611]), .C(n206), .D(regs[547]), .Q(n351) );
  AOI220 U1460 ( .A(n243), .B(regs[99]), .C(n206), .D(regs[35]), .Q(n355) );
  AOI220 U1461 ( .A(n243), .B(regs[868]), .C(n206), .D(regs[804]), .Q(n363) );
  AOI220 U1462 ( .A(n241), .B(regs[452]), .C(n974), .D(regs[388]), .Q(n368) );
  AOI220 U1463 ( .A(n977), .B(regs[612]), .C(n206), .D(regs[548]), .Q(n373) );
  AOI220 U1464 ( .A(n242), .B(regs[196]), .C(n974), .D(regs[132]), .Q(n378) );
  AOI220 U1465 ( .A(n242), .B(regs[453]), .C(n974), .D(regs[389]), .Q(n390) );
  AOI220 U1466 ( .A(n979), .B(regs[582]), .C(n232), .D(regs[518]), .Q(n416) );
  AOI220 U1467 ( .A(n973), .B(regs[230]), .C(n198), .D(regs[166]), .Q(n423) );
  AOI220 U1468 ( .A(n977), .B(regs[102]), .C(n206), .D(regs[38]), .Q(n421) );
  AOI220 U1469 ( .A(n979), .B(regs[70]), .C(n232), .D(regs[6]), .Q(n420) );
  AOI220 U1470 ( .A(n973), .B(regs[999]), .C(n198), .D(regs[935]), .Q(n431) );
  AOI220 U1471 ( .A(n979), .B(regs[839]), .C(n232), .D(regs[775]), .Q(n428) );
  AOI220 U1472 ( .A(n977), .B(regs[359]), .C(n206), .D(regs[295]), .Q(n433) );
  AOI220 U1473 ( .A(n979), .B(regs[327]), .C(n232), .D(regs[263]), .Q(n432) );
  AOI220 U1474 ( .A(n979), .B(regs[583]), .C(n232), .D(regs[519]), .Q(n438) );
  AOI220 U1475 ( .A(n973), .B(regs[231]), .C(n198), .D(regs[167]), .Q(n445) );
  AOI220 U1476 ( .A(n977), .B(regs[103]), .C(n206), .D(regs[39]), .Q(n443) );
  AOI220 U1477 ( .A(n979), .B(regs[71]), .C(n232), .D(regs[7]), .Q(n442) );
  AOI220 U1478 ( .A(n979), .B(regs[840]), .C(n232), .D(regs[776]), .Q(n450) );
  AOI220 U1479 ( .A(n977), .B(regs[360]), .C(n206), .D(regs[296]), .Q(n455) );
  AOI220 U1480 ( .A(n979), .B(regs[328]), .C(n232), .D(regs[264]), .Q(n454) );
  AOI220 U1481 ( .A(n243), .B(regs[362]), .C(n206), .D(regs[298]), .Q(n499) );
  AOI220 U1482 ( .A(n243), .B(regs[363]), .C(n206), .D(regs[299]), .Q(n521) );
  AOI220 U1483 ( .A(n243), .B(regs[876]), .C(n976), .D(regs[812]), .Q(n539) );
  AOI220 U1484 ( .A(n973), .B(regs[492]), .C(n198), .D(regs[428]), .Q(n545) );
  AOI220 U1485 ( .A(n973), .B(regs[1005]), .C(n198), .D(regs[941]), .Q(n563)
         );
  AOI220 U1486 ( .A(n244), .B(regs[845]), .C(n978), .D(regs[781]), .Q(n560) );
  AOI220 U1487 ( .A(n977), .B(regs[878]), .C(n206), .D(regs[814]), .Q(n583) );
  AOI220 U1488 ( .A(n979), .B(regs[846]), .C(n232), .D(regs[782]), .Q(n582) );
  AOI220 U1489 ( .A(n977), .B(regs[110]), .C(n206), .D(regs[46]), .Q(n597) );
  AOI220 U1490 ( .A(n243), .B(regs[879]), .C(n976), .D(regs[815]), .Q(n605) );
  AOI220 U1491 ( .A(n977), .B(regs[367]), .C(n206), .D(regs[303]), .Q(n609) );
  AOI220 U1492 ( .A(n243), .B(regs[111]), .C(n206), .D(regs[47]), .Q(n619) );
  AOI220 U1493 ( .A(n973), .B(regs[496]), .C(n198), .D(regs[432]), .Q(n633) );
  AOI220 U1494 ( .A(n243), .B(regs[112]), .C(n976), .D(regs[48]), .Q(n641) );
  AOI220 U1495 ( .A(n975), .B(regs[977]), .C(n202), .D(regs[913]), .Q(n650) );
  AOI220 U1496 ( .A(n243), .B(regs[625]), .C(n976), .D(regs[561]), .Q(n659) );
  AOI220 U1497 ( .A(n243), .B(regs[113]), .C(n976), .D(regs[49]), .Q(n663) );
  AOI220 U1498 ( .A(n975), .B(regs[978]), .C(n202), .D(regs[914]), .Q(n672) );
  AOI220 U1499 ( .A(n244), .B(regs[852]), .C(n978), .D(regs[788]), .Q(n714) );
  AOI220 U1500 ( .A(n975), .B(regs[468]), .C(n202), .D(regs[404]), .Q(n720) );
  AOI220 U1501 ( .A(n243), .B(regs[372]), .C(n976), .D(regs[308]), .Q(n719) );
  AOI220 U1502 ( .A(n244), .B(regs[340]), .C(n978), .D(regs[276]), .Q(n718) );
  AOI220 U1503 ( .A(n243), .B(regs[628]), .C(n206), .D(regs[564]), .Q(n725) );
  AOI220 U1504 ( .A(n244), .B(regs[84]), .C(n978), .D(regs[20]), .Q(n728) );
  AOI220 U1505 ( .A(n244), .B(regs[853]), .C(n978), .D(regs[789]), .Q(n736) );
  AOI220 U1506 ( .A(n975), .B(regs[469]), .C(n974), .D(regs[405]), .Q(n742) );
  AOI220 U1507 ( .A(n243), .B(regs[373]), .C(n976), .D(regs[309]), .Q(n741) );
  AOI220 U1508 ( .A(n244), .B(regs[341]), .C(n978), .D(regs[277]), .Q(n740) );
  AOI220 U1509 ( .A(n975), .B(regs[213]), .C(n974), .D(regs[149]), .Q(n752) );
  AOI220 U1510 ( .A(n243), .B(regs[117]), .C(n976), .D(regs[53]), .Q(n751) );
  AOI220 U1511 ( .A(n244), .B(regs[85]), .C(n978), .D(regs[21]), .Q(n750) );
  AOI220 U1512 ( .A(n244), .B(regs[854]), .C(n978), .D(regs[790]), .Q(n758) );
  AOI220 U1513 ( .A(n243), .B(regs[375]), .C(n206), .D(regs[311]), .Q(n785) );
  AOI220 U1514 ( .A(n243), .B(regs[631]), .C(n206), .D(regs[567]), .Q(n791) );
  AOI220 U1515 ( .A(n243), .B(regs[119]), .C(n206), .D(regs[55]), .Q(n795) );
  AOI220 U1516 ( .A(n244), .B(regs[87]), .C(n978), .D(regs[23]), .Q(n794) );
  AOI220 U1517 ( .A(n243), .B(regs[888]), .C(n206), .D(regs[824]), .Q(n803) );
  AOI220 U1518 ( .A(n243), .B(regs[376]), .C(n206), .D(regs[312]), .Q(n807) );
  AOI220 U1519 ( .A(n243), .B(regs[377]), .C(n206), .D(regs[313]), .Q(n829) );
  AOI220 U1520 ( .A(n975), .B(regs[729]), .C(n974), .D(regs[665]), .Q(n836) );
  AOI220 U1521 ( .A(n243), .B(regs[121]), .C(n206), .D(regs[57]), .Q(n839) );
  AOI220 U1522 ( .A(n243), .B(regs[890]), .C(n206), .D(regs[826]), .Q(n847) );
  AOI220 U1523 ( .A(n975), .B(regs[475]), .C(n974), .D(regs[411]), .Q(n874) );
  AOI220 U1524 ( .A(n975), .B(regs[219]), .C(n974), .D(regs[155]), .Q(n884) );
  AOI220 U1525 ( .A(n975), .B(regs[732]), .C(n974), .D(regs[668]), .Q(n902) );
  AOI220 U1526 ( .A(n977), .B(regs[893]), .C(n206), .D(regs[829]), .Q(n913) );
  AOI220 U1527 ( .A(n979), .B(regs[605]), .C(n232), .D(regs[541]), .Q(n922) );
  AOI220 U1528 ( .A(n243), .B(regs[638]), .C(n976), .D(regs[574]), .Q(n945) );
  AOI220 U1529 ( .A(n243), .B(regs[126]), .C(n206), .D(regs[62]), .Q(n949) );
  AOI220 U1530 ( .A(n243), .B(regs[895]), .C(n206), .D(regs[831]), .Q(n957) );
  AOI220 U1531 ( .A(n243), .B(regs[639]), .C(n206), .D(regs[575]), .Q(n969) );
  AOI220 U1532 ( .A(n977), .B(regs[127]), .C(n206), .D(regs[63]), .Q(n981) );
  AOI220 U1533 ( .A(regs[322]), .B(n203), .C(regs[258]), .D(n1568), .Q(n1000)
         );
  AOI220 U1534 ( .A(regs[578]), .B(n203), .C(regs[514]), .D(n1568), .Q(n1006)
         );
  AOI220 U1535 ( .A(regs[66]), .B(n203), .C(regs[2]), .D(n1568), .Q(n1010) );
  AOI220 U1536 ( .A(regs[868]), .B(n247), .C(regs[804]), .D(n205), .Q(n1019)
         );
  AOI220 U1537 ( .A(regs[356]), .B(n247), .C(regs[292]), .D(n205), .Q(n1023)
         );
  AOI220 U1538 ( .A(regs[324]), .B(n1569), .C(regs[260]), .D(n204), .Q(n1022)
         );
  AOI220 U1539 ( .A(regs[580]), .B(n203), .C(regs[516]), .D(n1568), .Q(n1028)
         );
  AOI220 U1540 ( .A(regs[68]), .B(n203), .C(regs[4]), .D(n1568), .Q(n1032) );
  AOI220 U1541 ( .A(regs[485]), .B(n1563), .C(regs[421]), .D(n199), .Q(n1047)
         );
  AOI220 U1542 ( .A(regs[453]), .B(n1565), .C(regs[389]), .D(n200), .Q(n1046)
         );
  AOI220 U1543 ( .A(regs[229]), .B(n1563), .C(regs[165]), .D(n199), .Q(n1057)
         );
  AOI220 U1544 ( .A(regs[69]), .B(n203), .C(regs[5]), .D(n1568), .Q(n1054) );
  AOI220 U1545 ( .A(regs[486]), .B(n1563), .C(regs[422]), .D(n199), .Q(n1069)
         );
  AOI220 U1546 ( .A(regs[454]), .B(n1565), .C(regs[390]), .D(n200), .Q(n1068)
         );
  AOI220 U1547 ( .A(regs[358]), .B(n1567), .C(regs[294]), .D(n205), .Q(n1067)
         );
  AOI220 U1548 ( .A(regs[326]), .B(n203), .C(regs[262]), .D(n1568), .Q(n1066)
         );
  AOI220 U1549 ( .A(regs[614]), .B(n1567), .C(regs[550]), .D(n205), .Q(n1073)
         );
  AOI220 U1550 ( .A(regs[582]), .B(n203), .C(regs[518]), .D(n1568), .Q(n1072)
         );
  AOI220 U1551 ( .A(regs[70]), .B(n203), .C(regs[6]), .D(n1568), .Q(n1076) );
  AOI220 U1552 ( .A(regs[839]), .B(n1569), .C(regs[775]), .D(n1568), .Q(n1084)
         );
  AOI220 U1553 ( .A(regs[327]), .B(n1569), .C(regs[263]), .D(n1568), .Q(n1088)
         );
  AOI220 U1554 ( .A(regs[583]), .B(n203), .C(regs[519]), .D(n1568), .Q(n1094)
         );
  AOI220 U1555 ( .A(regs[71]), .B(n1569), .C(regs[7]), .D(n1568), .Q(n1098) );
  AOI220 U1556 ( .A(regs[328]), .B(n1569), .C(regs[264]), .D(n204), .Q(n1110)
         );
  AOI220 U1557 ( .A(regs[72]), .B(n203), .C(regs[8]), .D(n1568), .Q(n1120) );
  AOI220 U1558 ( .A(regs[841]), .B(n203), .C(regs[777]), .D(n1568), .Q(n1128)
         );
  AOI220 U1559 ( .A(regs[329]), .B(n1569), .C(regs[265]), .D(n204), .Q(n1132)
         );
  AOI220 U1560 ( .A(regs[585]), .B(n203), .C(regs[521]), .D(n1568), .Q(n1138)
         );
  AOI220 U1561 ( .A(regs[73]), .B(n1569), .C(regs[9]), .D(n204), .Q(n1142) );
  AOI220 U1562 ( .A(regs[843]), .B(n203), .C(regs[779]), .D(n1568), .Q(n1150)
         );
  AOI220 U1563 ( .A(regs[235]), .B(n1563), .C(regs[171]), .D(n199), .Q(n1167)
         );
  AOI220 U1564 ( .A(regs[203]), .B(n1565), .C(regs[139]), .D(n200), .Q(n1166)
         );
  AOI220 U1565 ( .A(regs[492]), .B(n245), .C(regs[428]), .D(n1562), .Q(n1179)
         );
  AOI220 U1566 ( .A(regs[460]), .B(n246), .C(regs[396]), .D(n1564), .Q(n1178)
         );
  AOI220 U1567 ( .A(regs[364]), .B(n247), .C(regs[300]), .D(n1566), .Q(n1177)
         );
  AOI220 U1568 ( .A(regs[332]), .B(n1569), .C(regs[268]), .D(n1568), .Q(n1176)
         );
  AOI220 U1569 ( .A(regs[588]), .B(n203), .C(regs[524]), .D(n1568), .Q(n1182)
         );
  AOI220 U1570 ( .A(regs[76]), .B(n203), .C(regs[12]), .D(n1568), .Q(n1186) );
  AOI220 U1571 ( .A(regs[845]), .B(n203), .C(regs[781]), .D(n1568), .Q(n1194)
         );
  AOI220 U1572 ( .A(regs[493]), .B(n245), .C(regs[429]), .D(n1562), .Q(n1201)
         );
  AOI220 U1573 ( .A(regs[333]), .B(n203), .C(regs[269]), .D(n1568), .Q(n1198)
         );
  AOI220 U1574 ( .A(regs[589]), .B(n203), .C(regs[525]), .D(n1568), .Q(n1204)
         );
  AOI220 U1575 ( .A(regs[77]), .B(n203), .C(regs[13]), .D(n1568), .Q(n1208) );
  AOI220 U1576 ( .A(regs[847]), .B(n203), .C(regs[783]), .D(n1568), .Q(n1216)
         );
  AOI220 U1577 ( .A(regs[335]), .B(n203), .C(regs[271]), .D(n1568), .Q(n1220)
         );
  AOI220 U1578 ( .A(regs[239]), .B(n1563), .C(regs[175]), .D(n199), .Q(n1233)
         );
  AOI220 U1579 ( .A(regs[207]), .B(n1565), .C(regs[143]), .D(n200), .Q(n1232)
         );
  AOI220 U1580 ( .A(regs[79]), .B(n203), .C(regs[15]), .D(n1568), .Q(n1230) );
  AOI220 U1581 ( .A(regs[848]), .B(n203), .C(regs[784]), .D(n1568), .Q(n1238)
         );
  AOI220 U1582 ( .A(regs[368]), .B(n1567), .C(regs[304]), .D(n205), .Q(n1243)
         );
  AOI220 U1583 ( .A(regs[336]), .B(n203), .C(regs[272]), .D(n1568), .Q(n1242)
         );
  AOI220 U1584 ( .A(regs[80]), .B(n203), .C(regs[16]), .D(n1568), .Q(n1252) );
  AOI220 U1585 ( .A(regs[465]), .B(n246), .C(regs[401]), .D(n1564), .Q(n1266)
         );
  AOI220 U1586 ( .A(regs[369]), .B(n247), .C(regs[305]), .D(n1566), .Q(n1265)
         );
  AOI220 U1587 ( .A(regs[337]), .B(n203), .C(regs[273]), .D(n1568), .Q(n1264)
         );
  AOI220 U1588 ( .A(regs[593]), .B(n203), .C(regs[529]), .D(n1568), .Q(n1270)
         );
  AOI220 U1589 ( .A(regs[851]), .B(n203), .C(regs[787]), .D(n1568), .Q(n1304)
         );
  AOI220 U1590 ( .A(regs[499]), .B(n245), .C(regs[435]), .D(n1562), .Q(n1311)
         );
  AOI220 U1591 ( .A(regs[467]), .B(n246), .C(regs[403]), .D(n1564), .Q(n1310)
         );
  AOI220 U1592 ( .A(regs[371]), .B(n247), .C(regs[307]), .D(n1566), .Q(n1309)
         );
  AOI220 U1593 ( .A(regs[243]), .B(n1563), .C(regs[179]), .D(n1562), .Q(n1321)
         );
  AOI220 U1594 ( .A(regs[211]), .B(n1565), .C(regs[147]), .D(n1564), .Q(n1320)
         );
  AOI220 U1595 ( .A(regs[115]), .B(n247), .C(regs[51]), .D(n1566), .Q(n1319)
         );
  AOI220 U1596 ( .A(regs[500]), .B(n245), .C(regs[436]), .D(n1562), .Q(n1333)
         );
  AOI220 U1597 ( .A(regs[468]), .B(n246), .C(regs[404]), .D(n1564), .Q(n1332)
         );
  AOI220 U1598 ( .A(regs[372]), .B(n247), .C(regs[308]), .D(n1566), .Q(n1331)
         );
  AOI220 U1599 ( .A(regs[340]), .B(n203), .C(regs[276]), .D(n1568), .Q(n1330)
         );
  AOI220 U1600 ( .A(regs[854]), .B(n203), .C(regs[790]), .D(n1568), .Q(n1348)
         );
  AOI220 U1601 ( .A(regs[374]), .B(n1567), .C(regs[310]), .D(n205), .Q(n1353)
         );
  AOI220 U1602 ( .A(regs[342]), .B(n203), .C(regs[278]), .D(n1568), .Q(n1352)
         );
  AOI220 U1603 ( .A(regs[983]), .B(n246), .C(regs[919]), .D(n1564), .Q(n1372)
         );
  AOI220 U1604 ( .A(regs[343]), .B(n1569), .C(regs[279]), .D(n204), .Q(n1374)
         );
  AOI220 U1605 ( .A(regs[1018]), .B(n245), .C(regs[954]), .D(n1562), .Q(n1439)
         );
  AOI220 U1606 ( .A(regs[346]), .B(n203), .C(regs[282]), .D(n1568), .Q(n1440)
         );
  AOI220 U1607 ( .A(regs[602]), .B(n1569), .C(regs[538]), .D(n1568), .Q(n1446)
         );
  AOI220 U1608 ( .A(regs[90]), .B(n203), .C(regs[26]), .D(n1568), .Q(n1450) );
  AOI220 U1609 ( .A(regs[859]), .B(n203), .C(regs[795]), .D(n1568), .Q(n1458)
         );
  AOI220 U1610 ( .A(regs[347]), .B(n1569), .C(regs[283]), .D(n1568), .Q(n1462)
         );
  AOI220 U1611 ( .A(regs[603]), .B(n1569), .C(regs[539]), .D(n1568), .Q(n1468)
         );
  AOI220 U1612 ( .A(regs[91]), .B(n203), .C(regs[27]), .D(n1568), .Q(n1472) );
  AOI220 U1613 ( .A(regs[380]), .B(n1567), .C(regs[316]), .D(n205), .Q(n1485)
         );
  AOI220 U1614 ( .A(regs[381]), .B(n1567), .C(regs[317]), .D(n205), .Q(n1507)
         );
  AOI220 U1615 ( .A(regs[349]), .B(n203), .C(regs[285]), .D(n1568), .Q(n1506)
         );
  AOI220 U1616 ( .A(regs[605]), .B(n203), .C(regs[541]), .D(n1568), .Q(n1512)
         );
  AOI220 U1617 ( .A(regs[253]), .B(n1563), .C(regs[189]), .D(n199), .Q(n1519)
         );
  AOI220 U1618 ( .A(regs[221]), .B(n1565), .C(regs[157]), .D(n200), .Q(n1518)
         );
  AOI220 U1619 ( .A(regs[93]), .B(n203), .C(regs[29]), .D(n1568), .Q(n1516) );
  AOI220 U1620 ( .A(regs[382]), .B(n1567), .C(regs[318]), .D(n1566), .Q(n1529)
         );
  AOI220 U1621 ( .A(regs[94]), .B(n203), .C(regs[30]), .D(n1568), .Q(n1538) );
  AOI220 U1622 ( .A(regs[767]), .B(n1563), .C(regs[703]), .D(n199), .Q(n1561)
         );
  AOI220 U1623 ( .A(regs[735]), .B(n1565), .C(regs[671]), .D(n200), .Q(n1560)
         );
  AOI220 U1624 ( .A(regs[127]), .B(n1567), .C(regs[63]), .D(n205), .Q(n1571)
         );
endmodule


module core ( clk, rst_n, read_instruction, read_data, instruction_address, 
        data_address, write_data, mem_write, mem_read );
  input [31:0] read_instruction;
  input [31:0] read_data;
  output [31:0] instruction_address;
  output [31:0] data_address;
  output [31:0] write_data;
  input clk, rst_n;
  output mem_write, mem_read;
  wire   if_con_b, if_con_ifstall, id_con_Wregwrite, ex_con_Wregwrite,
         mem_con_Wregwrite, for_FWmemread, ex_con_Ealusrc, ex_con_Eregdst,
         ex_con_Mmemread, ex_con_Mmemwrite, ex_con_Malupc8, ex_con_Wmemtoreg,
         mem_con_Malupc8, mem_con_Wmemtoreg, wb_con_Wmemtoreg,
         u_fetch_jmux_i_addr_pc4_2_, u_fetch_jmux_i_addr_pc4_3_,
         u_fetch_jmux_i_addr_pc4_4_, u_fetch_jmux_i_addr_pc4_5_,
         u_fetch_jmux_i_addr_pc4_6_, u_fetch_jmux_i_addr_pc4_7_,
         u_fetch_jmux_i_addr_pc4_8_, u_fetch_jmux_i_addr_pc4_9_,
         u_fetch_jmux_i_addr_pc4_10_, u_fetch_jmux_i_addr_pc4_11_,
         u_fetch_jmux_i_addr_pc4_12_, u_fetch_jmux_i_addr_pc4_13_,
         u_fetch_jmux_i_addr_pc4_14_, u_fetch_jmux_i_addr_pc4_15_,
         u_fetch_jmux_i_addr_pc4_16_, u_fetch_jmux_i_addr_pc4_17_,
         u_fetch_jmux_i_addr_pc4_18_, u_fetch_jmux_i_addr_pc4_19_,
         u_fetch_jmux_i_addr_pc4_20_, u_fetch_jmux_i_addr_pc4_21_,
         u_fetch_jmux_i_addr_pc4_22_, u_fetch_jmux_i_addr_pc4_23_,
         u_fetch_jmux_i_addr_pc4_24_, u_fetch_jmux_i_addr_pc4_25_,
         u_fetch_jmux_i_addr_pc4_26_, u_fetch_jmux_i_addr_pc4_27_,
         u_fetch_jmux_i_addr_pc4_28_, u_fetch_jmux_i_addr_pc4_29_,
         u_fetch_jmux_i_addr_pc4_30_, u_fetch_jmux_i_addr_pc4_31_, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, u_decode_n6,
         u_decode_n1, u_decode_for_o_con_fa_0_, u_decode_for_o_con_fa_1_,
         u_decode_for_o_con_fa_2_, u_decode_control_o_con_regwrite,
         u_decode_control_o_con_memtoreg, u_decode_control_o_con_memwrite,
         u_decode_control_o_con_memread, u_decode_jbcon_o_con_aluPC4,
         u_decode_control_o_con_regdst, u_decode_control_o_con_alusrc,
         u_decode_control_o_con_aluop_0_, u_decode_control_o_con_aluop_1_,
         u_decode_control_o_con_aluop_2_, u_decode_control_o_con_aluop_3_,
         u_decode_control_o_con_aluop_4_, u_decode_control_o_con_aluop_5_,
         u_decode_add_x_16_n135, u_decode_add_x_16_n131,
         u_decode_add_x_16_n129, u_decode_add_x_16_n117,
         u_decode_add_x_16_n115, u_decode_add_x_16_n114,
         u_decode_add_x_16_n113, u_decode_add_x_16_n112,
         u_decode_add_x_16_n111, u_decode_add_x_16_n110,
         u_decode_add_x_16_n109, u_decode_add_x_16_n108,
         u_decode_add_x_16_n107, u_decode_add_x_16_n106,
         u_decode_add_x_16_n105, u_decode_add_x_16_n104,
         u_decode_add_x_16_n103, u_decode_add_x_16_n102,
         u_decode_add_x_16_n101, u_decode_add_x_16_n99, u_decode_add_x_16_n97,
         u_decode_add_x_16_n96, u_decode_add_x_16_n95, u_decode_add_x_16_n94,
         u_decode_add_x_16_n93, u_decode_add_x_16_n92, u_decode_add_x_16_n91,
         u_decode_add_x_16_n90, u_decode_add_x_16_n89, u_decode_add_x_16_n88,
         u_decode_add_x_16_n87, u_decode_add_x_16_n86, u_decode_add_x_16_n85,
         u_decode_add_x_16_n84, u_decode_add_x_16_n83, u_decode_add_x_16_n82,
         u_decode_add_x_16_n81, u_decode_add_x_16_n80, u_decode_add_x_16_n79,
         u_decode_add_x_16_n78, u_decode_add_x_16_n77, u_decode_add_x_16_n76,
         u_decode_add_x_16_n75, u_decode_add_x_16_n74, u_decode_add_x_16_n73,
         u_decode_add_x_16_n72, u_decode_add_x_16_n71, u_decode_add_x_16_n70,
         u_decode_add_x_16_n69, u_decode_add_x_16_n68, u_decode_add_x_16_n67,
         u_decode_add_x_16_n66, u_decode_add_x_16_n65, u_decode_add_x_16_n64,
         u_decode_add_x_16_n63, u_decode_add_x_16_n62, u_decode_add_x_16_n61,
         u_decode_add_x_16_n60, u_decode_add_x_16_n59, u_decode_add_x_16_n58,
         u_decode_add_x_16_n57, u_decode_add_x_16_n56, u_decode_add_x_16_n55,
         u_decode_add_x_16_n54, u_decode_add_x_16_n53, u_decode_add_x_16_n52,
         u_decode_add_x_16_n51, u_decode_add_x_16_n50, u_decode_add_x_16_n49,
         u_decode_add_x_16_n48, u_decode_add_x_16_n47, u_decode_add_x_16_n46,
         u_decode_add_x_16_n45, u_decode_add_x_16_n44, u_decode_add_x_16_n43,
         u_decode_add_x_16_n42, u_decode_add_x_16_n41, u_decode_add_x_16_n40,
         u_decode_add_x_16_n39, u_decode_add_x_16_n38, u_decode_add_x_16_n37,
         u_decode_add_x_16_n36, u_decode_add_x_16_n35, u_decode_add_x_16_n34,
         u_decode_add_x_16_n33, u_decode_add_x_16_n32, u_decode_add_x_16_n31,
         u_decode_add_x_16_n30, u_decode_add_x_16_n29, u_decode_add_x_16_n28,
         u_decode_add_x_16_n27, u_decode_add_x_16_n26, u_decode_add_x_16_n25,
         u_decode_add_x_16_n24, u_decode_add_x_16_n23, u_decode_add_x_16_n19,
         u_decode_add_x_16_n18, u_decode_add_x_16_n15, u_decode_add_x_16_n13,
         u_decode_add_x_16_n11, u_decode_add_x_16_n9, u_decode_add_x_16_n7,
         u_decode_add_x_16_n5, u_decode_add_x_16_n3, add_x_4_n28, add_x_4_n27,
         add_x_4_n26, add_x_4_n25, add_x_4_n24, add_x_4_n23, add_x_4_n22,
         add_x_4_n21, add_x_4_n20, add_x_4_n19, add_x_4_n18, add_x_4_n17,
         add_x_4_n16, add_x_4_n15, add_x_4_n12, add_x_4_n11, add_x_4_n10,
         add_x_4_n9, add_x_4_n8, add_x_4_n7, add_x_4_n6, add_x_4_n5,
         add_x_4_n4, add_x_4_n3, add_x_4_n2, add_x_4_n1, add_x_1_n28,
         add_x_1_n27, add_x_1_n26, add_x_1_n25, add_x_1_n24, add_x_1_n23,
         add_x_1_n22, add_x_1_n21, add_x_1_n20, add_x_1_n17, add_x_1_n16,
         add_x_1_n15, add_x_1_n14, add_x_1_n13, add_x_1_n12, add_x_1_n11,
         add_x_1_n10, add_x_1_n9, add_x_1_n8, add_x_1_n7, add_x_1_n6,
         add_x_1_n5, add_x_1_n4, add_x_1_n3, add_x_1_n2, add_x_1_n1, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405;
  wire   [31:2] if_addr_b;
  wire   [31:2] if_addr_j;
  wire   [31:0] id_data_jr;
  wire   [1:0] if_con_j;
  wire   [27:2] id_addr_pc4;
  wire   [31:26] id_data_instr;
  wire   [31:0] id_data_Wregwrite;
  wire   [4:0] id_addr_Wregwrite;
  wire   [4:0] for_o_addr_Erd;
  wire   [4:0] mem_addr_regdst;
  wire   [4:0] for_addr_rtM;
  wire   [4:0] for_addr_rtW;
  wire   [31:0] wb_data_memout;
  wire   [31:0] id_data_rs;
  wire   [31:0] ex_data_rt;
  wire   [4:0] ex_addr_rd;
  wire   [4:0] ex_addr_rt;
  wire   [31:0] ex_data_pc4;
  wire   [5:0] ex_con_Ealuop;
  wire   [2:0] ex_con_bop;
  wire   [31:0] ex_data_immext;
  wire   [2:0] for_o_con_Efamux;
  wire   [2:0] for_o_con_Efbmux;
  wire   [31:0] for_memout;
  wire   [31:0] mem_data_alures;
  wire   [31:2] mem_data_pc4;
  wire   [31:0] u_mem_resmux_o_data_alu;
  wire   [31:0] u_mem_pc8;
  wire   [1:0] u_decode_jbcon_o_con_bop;
  wire   [31:0] u_decode_pcadd_o_addr_pcbranchE;
  wire   [2:0] u_decode_for_o_con_fb;
  wire   [31:0] u_decode_regbank_o_data_Rt;

  execute u_execute ( .i_clk(clk), .i_nrst(rst_n), .i_data_pc4(ex_data_pc4), 
        .i_data_rs(id_data_rs), .i_data_rt(ex_data_rt), .i_data_immext({n204, 
        n204, n204, n204, n204, n204, n204, n204, n204, n204, n204, n204, n204, 
        n204, n204, ex_data_immext[31], ex_addr_rd, ex_data_immext[10:9], n207, 
        ex_data_immext[7], n206, ex_data_immext[5:0]}), .i_addr_rt(ex_addr_rt), 
        .i_addr_rd({n204, n204, n204, n204, n204}), .i_data_FEalures(
        data_address), .i_data_FMalures(mem_data_alures), .i_data_FMmemout(
        wb_data_memout), .i_data_FWmemout(for_memout), .i_con_Efamux(
        for_o_con_Efamux), .i_con_Efbmux(for_o_con_Efbmux), .i_con_Ealuop(
        ex_con_Ealuop), .i_con_Ealusrc(ex_con_Ealusrc), .i_con_Eregdst(
        ex_con_Eregdst), .i_con_Mmemread(ex_con_Mmemread), .i_con_Mmemwrite(
        ex_con_Mmemwrite), .i_con_Malupc8(ex_con_Malupc8), .i_con_Wmemtoreg(
        ex_con_Wmemtoreg), .i_con_Wregwrite(ex_con_Wregwrite), .i_con_bop(
        ex_con_bop), .o_data_pc4({mem_data_pc4, u_mem_pc8[1:0]}), 
        .o_data_alures(data_address), .o_data_rt(write_data), .o_addr_regdst(
        mem_addr_regdst), .o_con_Mmemread(mem_read), .o_con_Mmemwrite(
        mem_write), .o_con_Malupc8(mem_con_Malupc8), .o_con_Wmemtoreg(
        mem_con_Wmemtoreg), .o_con_Wregwrite(mem_con_Wregwrite), .o_addr_Erd(
        for_o_addr_Erd), .o_addr_Mrt(for_addr_rtM), .o_con_ifbranch(if_con_b)
         );
  DFC1 u_fetch_pipe_pc4_reg_0_ ( .D(instruction_address[0]), .C(clk), .RN(
        rst_n), .Q(u_decode_pcadd_o_addr_pcbranchE[0]) );
  DFC1 u_fetch_pipe_pc4_reg_1_ ( .D(instruction_address[1]), .C(clk), .RN(
        rst_n), .Q(u_decode_pcadd_o_addr_pcbranchE[1]) );
  DFC1 u_fetch_pipe_pc4_reg_2_ ( .D(u_fetch_jmux_i_addr_pc4_2_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[2]) );
  DFC1 u_fetch_pipe_pc4_reg_3_ ( .D(u_fetch_jmux_i_addr_pc4_3_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[3]) );
  DFC1 u_fetch_pipe_pc4_reg_4_ ( .D(u_fetch_jmux_i_addr_pc4_4_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[4]) );
  DFC1 u_fetch_pipe_pc4_reg_5_ ( .D(u_fetch_jmux_i_addr_pc4_5_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[5]) );
  DFC1 u_fetch_pipe_pc4_reg_6_ ( .D(u_fetch_jmux_i_addr_pc4_6_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[6]) );
  DFC1 u_fetch_pipe_pc4_reg_7_ ( .D(u_fetch_jmux_i_addr_pc4_7_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[7]) );
  DFC1 u_fetch_pipe_pc4_reg_8_ ( .D(u_fetch_jmux_i_addr_pc4_8_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[8]) );
  DFC1 u_fetch_pipe_pc4_reg_9_ ( .D(u_fetch_jmux_i_addr_pc4_9_), .C(clk), .RN(
        rst_n), .Q(id_addr_pc4[9]) );
  DFC1 u_fetch_pipe_pc4_reg_10_ ( .D(u_fetch_jmux_i_addr_pc4_10_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[10]) );
  DFC1 u_fetch_pipe_pc4_reg_11_ ( .D(u_fetch_jmux_i_addr_pc4_11_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[11]) );
  DFC1 u_fetch_pipe_pc4_reg_12_ ( .D(u_fetch_jmux_i_addr_pc4_12_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[12]) );
  DFC1 u_fetch_pipe_pc4_reg_13_ ( .D(u_fetch_jmux_i_addr_pc4_13_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[13]) );
  DFC1 u_fetch_pipe_pc4_reg_14_ ( .D(u_fetch_jmux_i_addr_pc4_14_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[14]) );
  DFC1 u_fetch_pipe_pc4_reg_15_ ( .D(u_fetch_jmux_i_addr_pc4_15_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[15]) );
  DFC1 u_fetch_pipe_pc4_reg_16_ ( .D(u_fetch_jmux_i_addr_pc4_16_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[16]) );
  DFC1 u_fetch_pipe_pc4_reg_17_ ( .D(u_fetch_jmux_i_addr_pc4_17_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[17]) );
  DFC1 u_fetch_pipe_pc4_reg_18_ ( .D(u_fetch_jmux_i_addr_pc4_18_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[18]) );
  DFC1 u_fetch_pipe_pc4_reg_19_ ( .D(u_fetch_jmux_i_addr_pc4_19_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[19]) );
  DFC1 u_fetch_pipe_pc4_reg_20_ ( .D(u_fetch_jmux_i_addr_pc4_20_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[20]) );
  DFC1 u_fetch_pipe_pc4_reg_21_ ( .D(u_fetch_jmux_i_addr_pc4_21_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[21]) );
  DFC1 u_fetch_pipe_pc4_reg_22_ ( .D(u_fetch_jmux_i_addr_pc4_22_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[22]) );
  DFC1 u_fetch_pipe_pc4_reg_23_ ( .D(u_fetch_jmux_i_addr_pc4_23_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[23]) );
  DFC1 u_fetch_pipe_pc4_reg_24_ ( .D(u_fetch_jmux_i_addr_pc4_24_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[24]) );
  DFC1 u_fetch_pipe_pc4_reg_25_ ( .D(u_fetch_jmux_i_addr_pc4_25_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[25]) );
  DFC1 u_fetch_pipe_pc4_reg_26_ ( .D(u_fetch_jmux_i_addr_pc4_26_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[26]) );
  DFC1 u_fetch_pipe_pc4_reg_27_ ( .D(u_fetch_jmux_i_addr_pc4_27_), .C(clk), 
        .RN(rst_n), .Q(id_addr_pc4[27]) );
  DFC1 u_fetch_pipe_pc4_reg_28_ ( .D(u_fetch_jmux_i_addr_pc4_28_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[28]) );
  DFC1 u_fetch_pipe_pc4_reg_29_ ( .D(u_fetch_jmux_i_addr_pc4_29_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[29]) );
  DFC1 u_fetch_pipe_pc4_reg_30_ ( .D(u_fetch_jmux_i_addr_pc4_30_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[30]) );
  DFC1 u_fetch_pipe_pc4_reg_31_ ( .D(u_fetch_jmux_i_addr_pc4_31_), .C(clk), 
        .RN(rst_n), .Q(if_addr_j[31]) );
  DFC1 u_fetch_pipe_instr_reg_0_ ( .D(read_instruction[0]), .C(clk), .RN(rst_n), .Q(if_addr_j[2]) );
  DFC1 u_fetch_pipe_instr_reg_1_ ( .D(read_instruction[1]), .C(clk), .RN(rst_n), .Q(if_addr_j[3]) );
  DFC1 u_fetch_pipe_instr_reg_2_ ( .D(read_instruction[2]), .C(clk), .RN(rst_n), .Q(if_addr_j[4]) );
  DFC1 u_fetch_pipe_instr_reg_3_ ( .D(read_instruction[3]), .C(clk), .RN(rst_n), .Q(if_addr_j[5]) );
  DFC1 u_fetch_pipe_instr_reg_4_ ( .D(read_instruction[4]), .C(clk), .RN(rst_n), .Q(if_addr_j[6]) );
  DFC1 u_fetch_pipe_instr_reg_5_ ( .D(read_instruction[5]), .C(clk), .RN(rst_n), .Q(if_addr_j[7]), .QN(n196) );
  DFC1 u_fetch_pipe_instr_reg_6_ ( .D(read_instruction[6]), .C(clk), .RN(rst_n), .Q(if_addr_j[8]) );
  DFC1 u_fetch_pipe_instr_reg_7_ ( .D(read_instruction[7]), .C(clk), .RN(rst_n), .Q(if_addr_j[9]) );
  DFC1 u_fetch_pipe_instr_reg_8_ ( .D(read_instruction[8]), .C(clk), .RN(rst_n), .Q(if_addr_j[10]) );
  DFC1 u_fetch_pipe_instr_reg_9_ ( .D(read_instruction[9]), .C(clk), .RN(rst_n), .Q(if_addr_j[11]) );
  DFC1 u_fetch_pipe_instr_reg_10_ ( .D(read_instruction[10]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[12]) );
  DFC1 u_fetch_pipe_instr_reg_11_ ( .D(read_instruction[11]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[13]) );
  DFC1 u_fetch_pipe_instr_reg_12_ ( .D(read_instruction[12]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[14]) );
  DFC1 u_fetch_pipe_instr_reg_13_ ( .D(read_instruction[13]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[15]) );
  DFC1 u_fetch_pipe_instr_reg_14_ ( .D(read_instruction[14]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[16]) );
  DFC1 u_fetch_pipe_instr_reg_21_ ( .D(read_instruction[21]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[23]), .QN(n193) );
  DFC1 u_fetch_pipe_instr_reg_22_ ( .D(read_instruction[22]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[24]), .QN(n191) );
  DFC1 u_fetch_pipe_instr_reg_23_ ( .D(read_instruction[23]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[25]), .QN(n190) );
  DFC1 u_fetch_pipe_instr_reg_24_ ( .D(read_instruction[24]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[26]), .QN(n195) );
  DFC1 u_fetch_pipe_instr_reg_25_ ( .D(read_instruction[25]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[27]), .QN(n194) );
  DFC1 u_fetch_pipe_instr_reg_26_ ( .D(read_instruction[26]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[26]), .QN(n185) );
  DFC1 u_fetch_pipe_instr_reg_27_ ( .D(read_instruction[27]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[27]), .QN(n192) );
  DFC1 u_fetch_pipe_instr_reg_28_ ( .D(read_instruction[28]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[28]), .QN(n189) );
  DFC1 u_fetch_pipe_instr_reg_29_ ( .D(read_instruction[29]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[29]), .QN(n186) );
  DFC1 u_fetch_pipe_instr_reg_30_ ( .D(read_instruction[30]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[30]) );
  DFC1 u_fetch_pipe_instr_reg_31_ ( .D(read_instruction[31]), .C(clk), .RN(
        rst_n), .Q(id_data_instr[31]), .QN(n200) );
  DFC1 u_mem_pipe_data_memout_reg_0_ ( .D(read_data[0]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[0]) );
  DFC1 u_mem_pipe_data_memout_reg_1_ ( .D(read_data[1]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[1]) );
  DFC1 u_mem_pipe_data_memout_reg_2_ ( .D(read_data[2]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[2]) );
  DFC1 u_mem_pipe_data_memout_reg_3_ ( .D(read_data[3]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[3]) );
  DFC1 u_mem_pipe_data_memout_reg_4_ ( .D(read_data[4]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[4]) );
  DFC1 u_mem_pipe_data_memout_reg_5_ ( .D(read_data[5]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[5]) );
  DFC1 u_mem_pipe_data_memout_reg_6_ ( .D(read_data[6]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[6]) );
  DFC1 u_mem_pipe_data_memout_reg_7_ ( .D(read_data[7]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[7]) );
  DFC1 u_mem_pipe_data_memout_reg_8_ ( .D(read_data[8]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[8]) );
  DFC1 u_mem_pipe_data_memout_reg_9_ ( .D(read_data[9]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[9]) );
  DFC1 u_mem_pipe_data_memout_reg_10_ ( .D(read_data[10]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[10]) );
  DFC1 u_mem_pipe_data_memout_reg_11_ ( .D(read_data[11]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[11]) );
  DFC1 u_mem_pipe_data_memout_reg_12_ ( .D(read_data[12]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[12]) );
  DFC1 u_mem_pipe_data_memout_reg_13_ ( .D(read_data[13]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[13]) );
  DFC1 u_mem_pipe_data_memout_reg_14_ ( .D(read_data[14]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[14]) );
  DFC1 u_mem_pipe_data_memout_reg_15_ ( .D(read_data[15]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[15]) );
  DFC1 u_mem_pipe_data_memout_reg_16_ ( .D(read_data[16]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[16]) );
  DFC1 u_mem_pipe_data_memout_reg_17_ ( .D(read_data[17]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[17]) );
  DFC1 u_mem_pipe_data_memout_reg_18_ ( .D(read_data[18]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[18]) );
  DFC1 u_mem_pipe_data_memout_reg_19_ ( .D(read_data[19]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[19]) );
  DFC1 u_mem_pipe_data_memout_reg_20_ ( .D(read_data[20]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[20]) );
  DFC1 u_mem_pipe_data_memout_reg_21_ ( .D(read_data[21]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[21]) );
  DFC1 u_mem_pipe_data_memout_reg_22_ ( .D(read_data[22]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[22]) );
  DFC1 u_mem_pipe_data_memout_reg_23_ ( .D(read_data[23]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[23]) );
  DFC1 u_mem_pipe_data_memout_reg_24_ ( .D(read_data[24]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[24]) );
  DFC1 u_mem_pipe_data_memout_reg_25_ ( .D(read_data[25]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[25]) );
  DFC1 u_mem_pipe_data_memout_reg_26_ ( .D(read_data[26]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[26]) );
  DFC1 u_mem_pipe_data_memout_reg_27_ ( .D(read_data[27]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[27]) );
  DFC1 u_mem_pipe_data_memout_reg_28_ ( .D(read_data[28]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[28]) );
  DFC1 u_mem_pipe_data_memout_reg_29_ ( .D(read_data[29]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[29]) );
  DFC1 u_mem_pipe_data_memout_reg_30_ ( .D(read_data[30]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[30]) );
  DFC1 u_mem_pipe_data_memout_reg_31_ ( .D(read_data[31]), .C(clk), .RN(rst_n), 
        .Q(wb_data_memout[31]) );
  DFC1 u_mem_pipe_rt_reg_4_ ( .D(for_addr_rtM[4]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[4]) );
  DFC1 u_mem_pipe_con_FWmemread_reg ( .D(ex_con_Mmemread), .C(clk), .RN(rst_n), 
        .Q(for_FWmemread) );
  DFC1 u_mem_pipe_rt_reg_0_ ( .D(for_addr_rtM[0]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[0]) );
  DFC1 u_mem_pipe_rt_reg_1_ ( .D(for_addr_rtM[1]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[1]) );
  DFC1 u_mem_pipe_rt_reg_2_ ( .D(for_addr_rtM[2]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[2]) );
  DFC1 u_mem_pipe_rt_reg_3_ ( .D(for_addr_rtM[3]), .C(clk), .RN(rst_n), .Q(
        for_addr_rtW[3]) );
  DFC1 u_mem_pipe_con_Wregwrite_reg ( .D(mem_con_Wregwrite), .C(clk), .RN(
        rst_n), .Q(id_con_Wregwrite) );
  DFC1 u_mem_pipe_addr_regdst_reg_1_ ( .D(mem_addr_regdst[1]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[1]) );
  DFC1 u_mem_pipe_addr_regdst_reg_2_ ( .D(mem_addr_regdst[2]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[2]) );
  DFC1 u_mem_pipe_addr_regdst_reg_4_ ( .D(mem_addr_regdst[4]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[4]) );
  DFC1 u_mem_pipe_data_alures_reg_0_ ( .D(u_mem_resmux_o_data_alu[0]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[0]) );
  DFC1 u_mem_pipe_data_alures_reg_1_ ( .D(u_mem_resmux_o_data_alu[1]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[1]) );
  DFC1 u_mem_pipe_data_alures_reg_2_ ( .D(u_mem_resmux_o_data_alu[2]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[2]) );
  DFC1 u_mem_pipe_data_alures_reg_3_ ( .D(u_mem_resmux_o_data_alu[3]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[3]) );
  DFC1 u_mem_pipe_data_alures_reg_4_ ( .D(u_mem_resmux_o_data_alu[4]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[4]) );
  DFC1 u_mem_pipe_data_alures_reg_5_ ( .D(u_mem_resmux_o_data_alu[5]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[5]) );
  DFC1 u_mem_pipe_data_alures_reg_6_ ( .D(u_mem_resmux_o_data_alu[6]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[6]) );
  DFC1 u_mem_pipe_data_alures_reg_7_ ( .D(u_mem_resmux_o_data_alu[7]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[7]) );
  DFC1 u_mem_pipe_data_alures_reg_8_ ( .D(u_mem_resmux_o_data_alu[8]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[8]) );
  DFC1 u_mem_pipe_data_alures_reg_9_ ( .D(u_mem_resmux_o_data_alu[9]), .C(clk), 
        .RN(rst_n), .Q(mem_data_alures[9]) );
  DFC1 u_mem_pipe_data_alures_reg_10_ ( .D(u_mem_resmux_o_data_alu[10]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[10]) );
  DFC1 u_mem_pipe_data_alures_reg_11_ ( .D(u_mem_resmux_o_data_alu[11]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[11]) );
  DFC1 u_mem_pipe_data_alures_reg_12_ ( .D(u_mem_resmux_o_data_alu[12]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[12]) );
  DFC1 u_mem_pipe_data_alures_reg_13_ ( .D(u_mem_resmux_o_data_alu[13]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[13]) );
  DFC1 u_mem_pipe_data_alures_reg_14_ ( .D(u_mem_resmux_o_data_alu[14]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[14]) );
  DFC1 u_mem_pipe_data_alures_reg_15_ ( .D(u_mem_resmux_o_data_alu[15]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[15]) );
  DFC1 u_mem_pipe_data_alures_reg_16_ ( .D(u_mem_resmux_o_data_alu[16]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[16]) );
  DFC1 u_mem_pipe_data_alures_reg_17_ ( .D(u_mem_resmux_o_data_alu[17]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[17]) );
  DFC1 u_mem_pipe_data_alures_reg_18_ ( .D(u_mem_resmux_o_data_alu[18]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[18]) );
  DFC1 u_mem_pipe_data_alures_reg_19_ ( .D(u_mem_resmux_o_data_alu[19]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[19]) );
  DFC1 u_mem_pipe_data_alures_reg_20_ ( .D(u_mem_resmux_o_data_alu[20]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[20]) );
  DFC1 u_mem_pipe_data_alures_reg_21_ ( .D(u_mem_resmux_o_data_alu[21]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[21]) );
  DFC1 u_mem_pipe_data_alures_reg_22_ ( .D(u_mem_resmux_o_data_alu[22]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[22]) );
  DFC1 u_mem_pipe_data_alures_reg_23_ ( .D(u_mem_resmux_o_data_alu[23]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[23]) );
  DFC1 u_mem_pipe_data_alures_reg_24_ ( .D(u_mem_resmux_o_data_alu[24]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[24]) );
  DFC1 u_mem_pipe_data_alures_reg_25_ ( .D(u_mem_resmux_o_data_alu[25]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[25]) );
  DFC1 u_mem_pipe_data_alures_reg_26_ ( .D(u_mem_resmux_o_data_alu[26]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[26]) );
  DFC1 u_mem_pipe_data_alures_reg_27_ ( .D(u_mem_resmux_o_data_alu[27]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[27]) );
  DFC1 u_mem_pipe_data_alures_reg_28_ ( .D(u_mem_resmux_o_data_alu[28]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[28]) );
  DFC1 u_mem_pipe_data_alures_reg_29_ ( .D(u_mem_resmux_o_data_alu[29]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[29]) );
  DFC1 u_mem_pipe_data_alures_reg_30_ ( .D(u_mem_resmux_o_data_alu[30]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[30]) );
  DFC1 u_mem_pipe_data_alures_reg_31_ ( .D(u_mem_resmux_o_data_alu[31]), .C(
        clk), .RN(rst_n), .Q(mem_data_alures[31]) );
  DFC1 u_fetch_u_pc_program_counter_reg_0_ ( .D(n137), .C(clk), .RN(rst_n), 
        .Q(instruction_address[0]), .QN(n202) );
  DFC1 u_fetch_u_pc_program_counter_reg_1_ ( .D(n136), .C(clk), .RN(rst_n), 
        .Q(instruction_address[1]), .QN(n203) );
  DFC1 u_fetch_u_pc_program_counter_reg_4_ ( .D(n133), .C(clk), .RN(rst_n), 
        .Q(instruction_address[4]) );
  DFC1 u_fetch_u_pc_program_counter_reg_5_ ( .D(n132), .C(clk), .RN(rst_n), 
        .Q(instruction_address[5]) );
  DFC1 u_fetch_u_pc_program_counter_reg_6_ ( .D(n131), .C(clk), .RN(rst_n), 
        .Q(instruction_address[6]) );
  DFC1 u_fetch_u_pc_program_counter_reg_7_ ( .D(n130), .C(clk), .RN(rst_n), 
        .Q(instruction_address[7]) );
  DFC1 u_fetch_u_pc_program_counter_reg_8_ ( .D(n129), .C(clk), .RN(rst_n), 
        .Q(instruction_address[8]) );
  DFC1 u_fetch_u_pc_program_counter_reg_9_ ( .D(n128), .C(clk), .RN(rst_n), 
        .Q(instruction_address[9]) );
  DFC1 u_fetch_u_pc_program_counter_reg_10_ ( .D(n127), .C(clk), .RN(rst_n), 
        .Q(instruction_address[10]) );
  DFC1 u_fetch_u_pc_program_counter_reg_11_ ( .D(n126), .C(clk), .RN(rst_n), 
        .Q(instruction_address[11]) );
  DFC1 u_fetch_u_pc_program_counter_reg_12_ ( .D(n125), .C(clk), .RN(rst_n), 
        .Q(instruction_address[12]) );
  DFC1 u_fetch_u_pc_program_counter_reg_13_ ( .D(n124), .C(clk), .RN(rst_n), 
        .Q(instruction_address[13]) );
  DFC1 u_fetch_u_pc_program_counter_reg_14_ ( .D(n123), .C(clk), .RN(rst_n), 
        .Q(instruction_address[14]) );
  DFC1 u_fetch_u_pc_program_counter_reg_15_ ( .D(n122), .C(clk), .RN(rst_n), 
        .Q(instruction_address[15]) );
  DFC1 u_fetch_u_pc_program_counter_reg_16_ ( .D(n121), .C(clk), .RN(rst_n), 
        .Q(instruction_address[16]) );
  DFC1 u_fetch_u_pc_program_counter_reg_17_ ( .D(n120), .C(clk), .RN(rst_n), 
        .Q(instruction_address[17]) );
  DFC1 u_fetch_u_pc_program_counter_reg_18_ ( .D(n119), .C(clk), .RN(rst_n), 
        .Q(instruction_address[18]), .QN(n168) );
  DFC1 u_fetch_u_pc_program_counter_reg_19_ ( .D(n118), .C(clk), .RN(rst_n), 
        .Q(instruction_address[19]) );
  DFC1 u_fetch_u_pc_program_counter_reg_20_ ( .D(n117), .C(clk), .RN(rst_n), 
        .Q(instruction_address[20]) );
  DFC1 u_fetch_u_pc_program_counter_reg_21_ ( .D(n116), .C(clk), .RN(rst_n), 
        .Q(instruction_address[21]) );
  DFC1 u_fetch_u_pc_program_counter_reg_22_ ( .D(n115), .C(clk), .RN(rst_n), 
        .Q(instruction_address[22]) );
  DFC1 u_fetch_u_pc_program_counter_reg_23_ ( .D(n114), .C(clk), .RN(rst_n), 
        .Q(instruction_address[23]) );
  DFC1 u_fetch_u_pc_program_counter_reg_24_ ( .D(n113), .C(clk), .RN(rst_n), 
        .Q(instruction_address[24]) );
  DFC1 u_fetch_u_pc_program_counter_reg_25_ ( .D(n112), .C(clk), .RN(rst_n), 
        .Q(instruction_address[25]) );
  DFC1 u_fetch_u_pc_program_counter_reg_26_ ( .D(n111), .C(clk), .RN(rst_n), 
        .Q(instruction_address[26]) );
  DFC1 u_fetch_u_pc_program_counter_reg_27_ ( .D(n110), .C(clk), .RN(rst_n), 
        .Q(instruction_address[27]) );
  DFC1 u_fetch_u_pc_program_counter_reg_28_ ( .D(n109), .C(clk), .RN(rst_n), 
        .Q(instruction_address[28]) );
  DFC1 u_fetch_u_pc_program_counter_reg_29_ ( .D(n108), .C(clk), .RN(rst_n), 
        .Q(instruction_address[29]) );
  DFC1 u_fetch_u_pc_program_counter_reg_30_ ( .D(n107), .C(clk), .RN(rst_n), 
        .Q(instruction_address[30]) );
  DFC1 u_fetch_u_pc_program_counter_reg_31_ ( .D(n138), .C(clk), .RN(rst_n), 
        .Q(instruction_address[31]), .QN(n179) );
  DFC1 u_decode_pipe_addr_branch_reg_0_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[0]), .C(clk), .RN(rst_n), .Q(
        ex_data_pc4[0]) );
  DFC1 u_decode_pipe_addr_branch_reg_1_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[1]), .C(clk), .RN(rst_n), .Q(
        ex_data_pc4[1]) );
  DFC1 u_decode_pipe_addr_branch_reg_2_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[2]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[2]) );
  DFC1 u_decode_pipe_addr_branch_reg_3_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[3]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[3]) );
  DFC1 u_decode_pipe_addr_branch_reg_4_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[4]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[4]) );
  DFC1 u_decode_pipe_addr_branch_reg_5_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[5]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[5]) );
  DFC1 u_decode_pipe_addr_branch_reg_6_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[6]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[6]) );
  DFC1 u_decode_pipe_addr_branch_reg_7_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[7]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[7]) );
  DFC1 u_decode_pipe_addr_branch_reg_8_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[8]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[8]) );
  DFC1 u_decode_pipe_addr_branch_reg_9_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[9]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[9]) );
  DFC1 u_decode_pipe_addr_branch_reg_10_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[10]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[10]) );
  DFC1 u_decode_pipe_addr_branch_reg_11_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[11]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[11]) );
  DFC1 u_decode_pipe_addr_branch_reg_12_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[12]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[12]) );
  DFC1 u_decode_pipe_addr_branch_reg_13_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[13]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[13]) );
  DFC1 u_decode_pipe_addr_branch_reg_14_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[14]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[14]) );
  DFC1 u_decode_pipe_addr_branch_reg_15_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[15]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[15]) );
  DFC1 u_decode_pipe_addr_branch_reg_16_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[16]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[16]) );
  DFC1 u_decode_pipe_addr_branch_reg_17_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[17]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[17]) );
  DFC1 u_decode_pipe_addr_branch_reg_18_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[18]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[18]) );
  DFC1 u_decode_pipe_addr_branch_reg_19_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[19]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[19]) );
  DFC1 u_decode_pipe_addr_branch_reg_20_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[20]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[20]) );
  DFC1 u_decode_pipe_addr_branch_reg_21_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[21]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[21]) );
  DFC1 u_decode_pipe_addr_branch_reg_22_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[22]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[22]) );
  DFC1 u_decode_pipe_addr_branch_reg_23_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[23]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[23]) );
  DFC1 u_decode_pipe_addr_branch_reg_24_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[24]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[24]) );
  DFC1 u_decode_pipe_addr_branch_reg_25_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[25]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[25]) );
  DFC1 u_decode_pipe_addr_branch_reg_26_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[26]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[26]) );
  DFC1 u_decode_pipe_addr_branch_reg_27_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[27]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[27]) );
  DFC1 u_decode_pipe_addr_branch_reg_28_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[28]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[28]) );
  DFC1 u_decode_pipe_addr_branch_reg_29_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[29]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[29]) );
  DFC1 u_decode_pipe_addr_branch_reg_30_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[30]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[30]) );
  DFC1 u_decode_pipe_addr_branch_reg_31_ ( .D(
        u_decode_pcadd_o_addr_pcbranchE[31]), .C(clk), .RN(rst_n), .Q(
        if_addr_b[31]) );
  DFC1 u_decode_pipe_FWmemout_reg_0_ ( .D(wb_data_memout[0]), .C(clk), .RN(
        rst_n), .Q(for_memout[0]) );
  DFC1 u_decode_pipe_FWmemout_reg_1_ ( .D(wb_data_memout[1]), .C(clk), .RN(
        rst_n), .Q(for_memout[1]) );
  DFC1 u_decode_pipe_FWmemout_reg_2_ ( .D(wb_data_memout[2]), .C(clk), .RN(
        rst_n), .Q(for_memout[2]) );
  DFC1 u_decode_pipe_FWmemout_reg_3_ ( .D(wb_data_memout[3]), .C(clk), .RN(
        rst_n), .Q(for_memout[3]) );
  DFC1 u_decode_pipe_FWmemout_reg_4_ ( .D(wb_data_memout[4]), .C(clk), .RN(
        rst_n), .Q(for_memout[4]) );
  DFC1 u_decode_pipe_FWmemout_reg_5_ ( .D(wb_data_memout[5]), .C(clk), .RN(
        rst_n), .Q(for_memout[5]) );
  DFC1 u_decode_pipe_FWmemout_reg_6_ ( .D(wb_data_memout[6]), .C(clk), .RN(
        rst_n), .Q(for_memout[6]) );
  DFC1 u_decode_pipe_FWmemout_reg_7_ ( .D(wb_data_memout[7]), .C(clk), .RN(
        rst_n), .Q(for_memout[7]) );
  DFC1 u_decode_pipe_FWmemout_reg_8_ ( .D(wb_data_memout[8]), .C(clk), .RN(
        rst_n), .Q(for_memout[8]) );
  DFC1 u_decode_pipe_FWmemout_reg_9_ ( .D(wb_data_memout[9]), .C(clk), .RN(
        rst_n), .Q(for_memout[9]) );
  DFC1 u_decode_pipe_FWmemout_reg_10_ ( .D(wb_data_memout[10]), .C(clk), .RN(
        rst_n), .Q(for_memout[10]) );
  DFC1 u_decode_pipe_FWmemout_reg_11_ ( .D(wb_data_memout[11]), .C(clk), .RN(
        rst_n), .Q(for_memout[11]) );
  DFC1 u_decode_pipe_FWmemout_reg_12_ ( .D(wb_data_memout[12]), .C(clk), .RN(
        rst_n), .Q(for_memout[12]) );
  DFC1 u_decode_pipe_FWmemout_reg_13_ ( .D(wb_data_memout[13]), .C(clk), .RN(
        rst_n), .Q(for_memout[13]) );
  DFC1 u_decode_pipe_FWmemout_reg_14_ ( .D(wb_data_memout[14]), .C(clk), .RN(
        rst_n), .Q(for_memout[14]) );
  DFC1 u_decode_pipe_FWmemout_reg_15_ ( .D(wb_data_memout[15]), .C(clk), .RN(
        rst_n), .Q(for_memout[15]) );
  DFC1 u_decode_pipe_FWmemout_reg_16_ ( .D(wb_data_memout[16]), .C(clk), .RN(
        rst_n), .Q(for_memout[16]) );
  DFC1 u_decode_pipe_FWmemout_reg_17_ ( .D(wb_data_memout[17]), .C(clk), .RN(
        rst_n), .Q(for_memout[17]) );
  DFC1 u_decode_pipe_FWmemout_reg_18_ ( .D(wb_data_memout[18]), .C(clk), .RN(
        rst_n), .Q(for_memout[18]) );
  DFC1 u_decode_pipe_FWmemout_reg_19_ ( .D(wb_data_memout[19]), .C(clk), .RN(
        rst_n), .Q(for_memout[19]) );
  DFC1 u_decode_pipe_FWmemout_reg_20_ ( .D(wb_data_memout[20]), .C(clk), .RN(
        rst_n), .Q(for_memout[20]) );
  DFC1 u_decode_pipe_FWmemout_reg_21_ ( .D(wb_data_memout[21]), .C(clk), .RN(
        rst_n), .Q(for_memout[21]) );
  DFC1 u_decode_pipe_FWmemout_reg_22_ ( .D(wb_data_memout[22]), .C(clk), .RN(
        rst_n), .Q(for_memout[22]) );
  DFC1 u_decode_pipe_FWmemout_reg_23_ ( .D(wb_data_memout[23]), .C(clk), .RN(
        rst_n), .Q(for_memout[23]) );
  DFC1 u_decode_pipe_FWmemout_reg_24_ ( .D(wb_data_memout[24]), .C(clk), .RN(
        rst_n), .Q(for_memout[24]) );
  DFC1 u_decode_pipe_FWmemout_reg_25_ ( .D(wb_data_memout[25]), .C(clk), .RN(
        rst_n), .Q(for_memout[25]) );
  DFC1 u_decode_pipe_FWmemout_reg_26_ ( .D(wb_data_memout[26]), .C(clk), .RN(
        rst_n), .Q(for_memout[26]) );
  DFC1 u_decode_pipe_FWmemout_reg_27_ ( .D(wb_data_memout[27]), .C(clk), .RN(
        rst_n), .Q(for_memout[27]) );
  DFC1 u_decode_pipe_FWmemout_reg_28_ ( .D(wb_data_memout[28]), .C(clk), .RN(
        rst_n), .Q(for_memout[28]) );
  DFC1 u_decode_pipe_FWmemout_reg_29_ ( .D(wb_data_memout[29]), .C(clk), .RN(
        rst_n), .Q(for_memout[29]) );
  DFC1 u_decode_pipe_FWmemout_reg_30_ ( .D(wb_data_memout[30]), .C(clk), .RN(
        rst_n), .Q(for_memout[30]) );
  DFC1 u_decode_pipe_FWmemout_reg_31_ ( .D(wb_data_memout[31]), .C(clk), .RN(
        rst_n), .Q(for_memout[31]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_0_ ( .D(if_addr_j[2]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[0]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_2_ ( .D(if_addr_j[4]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[2]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_3_ ( .D(if_addr_j[5]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[3]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_4_ ( .D(if_addr_j[6]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[4]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_5_ ( .D(if_addr_j[7]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[5]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_6_ ( .D(if_addr_j[8]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[6]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_7_ ( .D(if_addr_j[9]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[7]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_8_ ( .D(if_addr_j[10]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[8]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_9_ ( .D(if_addr_j[11]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[9]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_11_ ( .D(if_addr_j[13]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[0]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_12_ ( .D(if_addr_j[14]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[1]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_13_ ( .D(if_addr_j[15]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[2]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_14_ ( .D(if_addr_j[16]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[3]) );
  DFC1 u_decode_pipe_signext_o_data_immD_reg_15_ ( .D(if_addr_j[17]), .C(clk), 
        .RN(rst_n), .Q(ex_addr_rd[4]) );
  DFC1 u_decode_pipe_con_Wregwrite_reg ( .D(u_decode_control_o_con_regwrite), 
        .C(clk), .RN(rst_n), .Q(ex_con_Wregwrite) );
  DFC1 u_decode_pipe_con_Wmemtoreg_reg ( .D(u_decode_control_o_con_memtoreg), 
        .C(clk), .RN(rst_n), .Q(ex_con_Wmemtoreg) );
  DFC1 u_decode_pipe_con_Mmemwrite_reg ( .D(u_decode_control_o_con_memwrite), 
        .C(clk), .RN(rst_n), .Q(ex_con_Mmemwrite) );
  DFC1 u_decode_pipe_con_Mmemread_reg ( .D(u_decode_control_o_con_memread), 
        .C(clk), .RN(rst_n), .Q(ex_con_Mmemread) );
  DFC1 u_decode_pipe_con_MaluPC4_reg ( .D(u_decode_jbcon_o_con_aluPC4), .C(clk), .RN(rst_n), .Q(ex_con_Malupc8) );
  DFC1 u_decode_pipe_con_Eregdst_reg ( .D(u_decode_control_o_con_regdst), .C(
        clk), .RN(rst_n), .Q(ex_con_Eregdst) );
  DFC1 u_decode_pipe_con_Ealusrc_reg ( .D(u_decode_control_o_con_alusrc), .C(
        clk), .RN(rst_n), .Q(ex_con_Ealusrc) );
  DFC1 u_decode_pipe_con_Ealuop_reg_0_ ( .D(u_decode_control_o_con_aluop_0_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[0]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_1_ ( .D(u_decode_control_o_con_aluop_1_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[1]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_2_ ( .D(u_decode_control_o_con_aluop_2_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[2]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_3_ ( .D(u_decode_control_o_con_aluop_3_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[3]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_4_ ( .D(u_decode_control_o_con_aluop_4_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[4]) );
  DFC1 u_decode_pipe_con_Ealuop_reg_5_ ( .D(u_decode_control_o_con_aluop_5_), 
        .C(clk), .RN(rst_n), .Q(ex_con_Ealuop[5]) );
  DFC1 u_decode_pipe_addr_pc4_reg_2_ ( .D(id_addr_pc4[2]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[2]) );
  DFC1 u_decode_pipe_addr_pc4_reg_3_ ( .D(id_addr_pc4[3]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[3]) );
  DFC1 u_decode_pipe_addr_pc4_reg_4_ ( .D(id_addr_pc4[4]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[4]) );
  DFC1 u_decode_pipe_addr_pc4_reg_5_ ( .D(id_addr_pc4[5]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[5]) );
  DFC1 u_decode_pipe_addr_pc4_reg_6_ ( .D(id_addr_pc4[6]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[6]) );
  DFC1 u_decode_pipe_addr_pc4_reg_7_ ( .D(id_addr_pc4[7]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[7]) );
  DFC1 u_decode_pipe_addr_pc4_reg_8_ ( .D(id_addr_pc4[8]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[8]) );
  DFC1 u_decode_pipe_addr_pc4_reg_9_ ( .D(id_addr_pc4[9]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[9]) );
  DFC1 u_decode_pipe_addr_pc4_reg_10_ ( .D(id_addr_pc4[10]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[10]) );
  DFC1 u_decode_pipe_addr_pc4_reg_11_ ( .D(id_addr_pc4[11]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[11]) );
  DFC1 u_decode_pipe_addr_pc4_reg_12_ ( .D(id_addr_pc4[12]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[12]) );
  DFC1 u_decode_pipe_addr_pc4_reg_13_ ( .D(id_addr_pc4[13]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[13]) );
  DFC1 u_decode_pipe_addr_pc4_reg_14_ ( .D(id_addr_pc4[14]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[14]) );
  DFC1 u_decode_pipe_addr_pc4_reg_15_ ( .D(id_addr_pc4[15]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[15]) );
  DFC1 u_decode_pipe_addr_pc4_reg_16_ ( .D(id_addr_pc4[16]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[16]) );
  DFC1 u_decode_pipe_addr_pc4_reg_17_ ( .D(id_addr_pc4[17]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[17]) );
  DFC1 u_decode_pipe_addr_pc4_reg_18_ ( .D(id_addr_pc4[18]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[18]) );
  DFC1 u_decode_pipe_addr_pc4_reg_19_ ( .D(id_addr_pc4[19]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[19]) );
  DFC1 u_decode_pipe_addr_pc4_reg_20_ ( .D(id_addr_pc4[20]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[20]) );
  DFC1 u_decode_pipe_addr_pc4_reg_21_ ( .D(id_addr_pc4[21]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[21]) );
  DFC1 u_decode_pipe_addr_pc4_reg_22_ ( .D(id_addr_pc4[22]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[22]) );
  DFC1 u_decode_pipe_addr_pc4_reg_23_ ( .D(id_addr_pc4[23]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[23]) );
  DFC1 u_decode_pipe_addr_pc4_reg_24_ ( .D(id_addr_pc4[24]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[24]) );
  DFC1 u_decode_pipe_addr_pc4_reg_25_ ( .D(id_addr_pc4[25]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[25]) );
  DFC1 u_decode_pipe_addr_pc4_reg_26_ ( .D(id_addr_pc4[26]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[26]) );
  DFC1 u_decode_pipe_addr_pc4_reg_27_ ( .D(id_addr_pc4[27]), .C(clk), .RN(
        rst_n), .Q(ex_data_pc4[27]) );
  DFC1 u_decode_pipe_addr_pc4_reg_28_ ( .D(if_addr_j[28]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[28]) );
  DFC1 u_decode_pipe_addr_pc4_reg_29_ ( .D(if_addr_j[29]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[29]) );
  DFC1 u_decode_pipe_addr_pc4_reg_30_ ( .D(if_addr_j[30]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[30]) );
  DFC1 u_decode_pipe_addr_pc4_reg_31_ ( .D(if_addr_j[31]), .C(clk), .RN(rst_n), 
        .Q(ex_data_pc4[31]) );
  DFC1 u_decode_pipe_addr_rt_reg_0_ ( .D(if_addr_j[18]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[0]) );
  DFC1 u_decode_pipe_addr_rt_reg_1_ ( .D(if_addr_j[19]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[1]) );
  DFC1 u_decode_pipe_addr_rt_reg_2_ ( .D(if_addr_j[20]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[2]) );
  DFC1 u_decode_pipe_addr_rt_reg_3_ ( .D(if_addr_j[21]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[3]) );
  DFC1 u_decode_pipe_addr_rt_reg_4_ ( .D(if_addr_j[22]), .C(clk), .RN(rst_n), 
        .Q(ex_addr_rt[4]) );
  DFC1 u_decode_pipe_data_rt_reg_0_ ( .D(u_decode_regbank_o_data_Rt[0]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[0]) );
  DFC1 u_decode_pipe_data_rt_reg_1_ ( .D(u_decode_regbank_o_data_Rt[1]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[1]) );
  DFC1 u_decode_pipe_data_rt_reg_2_ ( .D(u_decode_regbank_o_data_Rt[2]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[2]) );
  DFC1 u_decode_pipe_data_rt_reg_3_ ( .D(u_decode_regbank_o_data_Rt[3]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[3]) );
  DFC1 u_decode_pipe_data_rt_reg_4_ ( .D(u_decode_regbank_o_data_Rt[4]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[4]) );
  DFC1 u_decode_pipe_data_rt_reg_5_ ( .D(u_decode_regbank_o_data_Rt[5]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[5]) );
  DFC1 u_decode_pipe_data_rt_reg_6_ ( .D(u_decode_regbank_o_data_Rt[6]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[6]) );
  DFC1 u_decode_pipe_data_rt_reg_7_ ( .D(u_decode_regbank_o_data_Rt[7]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[7]) );
  DFC1 u_decode_pipe_data_rt_reg_8_ ( .D(u_decode_regbank_o_data_Rt[8]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[8]) );
  DFC1 u_decode_pipe_data_rt_reg_9_ ( .D(u_decode_regbank_o_data_Rt[9]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[9]) );
  DFC1 u_decode_pipe_data_rt_reg_10_ ( .D(u_decode_regbank_o_data_Rt[10]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[10]) );
  DFC1 u_decode_pipe_data_rt_reg_11_ ( .D(u_decode_regbank_o_data_Rt[11]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[11]) );
  DFC1 u_decode_pipe_data_rt_reg_12_ ( .D(u_decode_regbank_o_data_Rt[12]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[12]) );
  DFC1 u_decode_pipe_data_rt_reg_13_ ( .D(u_decode_regbank_o_data_Rt[13]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[13]) );
  DFC1 u_decode_pipe_data_rt_reg_14_ ( .D(u_decode_regbank_o_data_Rt[14]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[14]) );
  DFC1 u_decode_pipe_data_rt_reg_15_ ( .D(u_decode_regbank_o_data_Rt[15]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[15]) );
  DFC1 u_decode_pipe_data_rt_reg_16_ ( .D(u_decode_regbank_o_data_Rt[16]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[16]) );
  DFC1 u_decode_pipe_data_rt_reg_17_ ( .D(u_decode_regbank_o_data_Rt[17]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[17]) );
  DFC1 u_decode_pipe_data_rt_reg_18_ ( .D(u_decode_regbank_o_data_Rt[18]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[18]) );
  DFC1 u_decode_pipe_data_rt_reg_19_ ( .D(u_decode_regbank_o_data_Rt[19]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[19]) );
  DFC1 u_decode_pipe_data_rt_reg_20_ ( .D(u_decode_regbank_o_data_Rt[20]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[20]) );
  DFC1 u_decode_pipe_data_rt_reg_21_ ( .D(u_decode_regbank_o_data_Rt[21]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[21]) );
  DFC1 u_decode_pipe_data_rt_reg_22_ ( .D(u_decode_regbank_o_data_Rt[22]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[22]) );
  DFC1 u_decode_pipe_data_rt_reg_23_ ( .D(u_decode_regbank_o_data_Rt[23]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[23]) );
  DFC1 u_decode_pipe_data_rt_reg_24_ ( .D(u_decode_regbank_o_data_Rt[24]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[24]) );
  DFC1 u_decode_pipe_data_rt_reg_25_ ( .D(u_decode_regbank_o_data_Rt[25]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[25]) );
  DFC1 u_decode_pipe_data_rt_reg_26_ ( .D(u_decode_regbank_o_data_Rt[26]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[26]) );
  DFC1 u_decode_pipe_data_rt_reg_27_ ( .D(u_decode_regbank_o_data_Rt[27]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[27]) );
  DFC1 u_decode_pipe_data_rt_reg_28_ ( .D(u_decode_regbank_o_data_Rt[28]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[28]) );
  DFC1 u_decode_pipe_data_rt_reg_29_ ( .D(u_decode_regbank_o_data_Rt[29]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[29]) );
  DFC1 u_decode_pipe_data_rt_reg_30_ ( .D(u_decode_regbank_o_data_Rt[30]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[30]) );
  DFC1 u_decode_pipe_data_rt_reg_31_ ( .D(u_decode_regbank_o_data_Rt[31]), .C(
        clk), .RN(rst_n), .Q(ex_data_rt[31]) );
  DFC1 u_decode_pipe_data_rs_reg_0_ ( .D(id_data_jr[0]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[0]) );
  DFC1 u_decode_pipe_data_rs_reg_1_ ( .D(id_data_jr[1]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[1]) );
  DFC1 u_decode_pipe_data_rs_reg_2_ ( .D(id_data_jr[2]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[2]) );
  DFC1 u_decode_pipe_data_rs_reg_3_ ( .D(id_data_jr[3]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[3]) );
  DFC1 u_decode_pipe_data_rs_reg_4_ ( .D(id_data_jr[4]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[4]) );
  DFC1 u_decode_pipe_data_rs_reg_5_ ( .D(id_data_jr[5]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[5]) );
  DFC1 u_decode_pipe_data_rs_reg_6_ ( .D(id_data_jr[6]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[6]) );
  DFC1 u_decode_pipe_data_rs_reg_7_ ( .D(id_data_jr[7]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[7]) );
  DFC1 u_decode_pipe_data_rs_reg_8_ ( .D(id_data_jr[8]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[8]) );
  DFC1 u_decode_pipe_data_rs_reg_9_ ( .D(id_data_jr[9]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[9]) );
  DFC1 u_decode_pipe_data_rs_reg_10_ ( .D(id_data_jr[10]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[10]) );
  DFC1 u_decode_pipe_data_rs_reg_11_ ( .D(id_data_jr[11]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[11]) );
  DFC1 u_decode_pipe_data_rs_reg_12_ ( .D(id_data_jr[12]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[12]) );
  DFC1 u_decode_pipe_data_rs_reg_13_ ( .D(id_data_jr[13]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[13]) );
  DFC1 u_decode_pipe_data_rs_reg_14_ ( .D(id_data_jr[14]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[14]) );
  DFC1 u_decode_pipe_data_rs_reg_15_ ( .D(id_data_jr[15]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[15]) );
  DFC1 u_decode_pipe_data_rs_reg_16_ ( .D(id_data_jr[16]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[16]) );
  DFC1 u_decode_pipe_data_rs_reg_17_ ( .D(id_data_jr[17]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[17]) );
  DFC1 u_decode_pipe_data_rs_reg_18_ ( .D(id_data_jr[18]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[18]) );
  DFC1 u_decode_pipe_data_rs_reg_19_ ( .D(id_data_jr[19]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[19]) );
  DFC1 u_decode_pipe_data_rs_reg_20_ ( .D(id_data_jr[20]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[20]) );
  DFC1 u_decode_pipe_data_rs_reg_21_ ( .D(id_data_jr[21]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[21]) );
  DFC1 u_decode_pipe_data_rs_reg_22_ ( .D(id_data_jr[22]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[22]) );
  DFC1 u_decode_pipe_data_rs_reg_23_ ( .D(id_data_jr[23]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[23]) );
  DFC1 u_decode_pipe_data_rs_reg_24_ ( .D(id_data_jr[24]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[24]) );
  DFC1 u_decode_pipe_data_rs_reg_25_ ( .D(id_data_jr[25]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[25]) );
  DFC1 u_decode_pipe_data_rs_reg_26_ ( .D(id_data_jr[26]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[26]) );
  DFC1 u_decode_pipe_data_rs_reg_27_ ( .D(id_data_jr[27]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[27]) );
  DFC1 u_decode_pipe_data_rs_reg_28_ ( .D(id_data_jr[28]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[28]) );
  DFC1 u_decode_pipe_data_rs_reg_29_ ( .D(id_data_jr[29]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[29]) );
  DFC1 u_decode_pipe_data_rs_reg_30_ ( .D(id_data_jr[30]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[30]) );
  DFC1 u_decode_pipe_data_rs_reg_31_ ( .D(id_data_jr[31]), .C(clk), .RN(rst_n), 
        .Q(id_data_rs[31]) );
  DFC1 u_decode_pipe_bop_reg_0_ ( .D(u_decode_jbcon_o_con_bop[0]), .C(clk), 
        .RN(rst_n), .Q(ex_con_bop[0]) );
  DFC1 u_decode_pipe_bop_reg_1_ ( .D(u_decode_jbcon_o_con_bop[1]), .C(clk), 
        .RN(rst_n), .Q(ex_con_bop[1]) );
  DFC1 u_decode_pipe_bop_reg_2_ ( .D(u_decode_n6), .C(clk), .RN(rst_n), .Q(
        ex_con_bop[2]) );
  D_register_bank u_decode_u_regbank ( .i_clk(clk), .i_rst_n(rst_n), 
        .i_addr_Rs(if_addr_j[27:23]), .i_con_RegWr(id_con_Wregwrite), 
        .i_addr_Rd(id_addr_Wregwrite), .i_data_Rd(id_data_Wregwrite), 
        .o_data_Rs(id_data_jr), .o_data_Rt(u_decode_regbank_o_data_Rt), 
        .i_addr_Rt_4_(if_addr_j[22]), .i_addr_Rt_3_(if_addr_j[21]), 
        .i_addr_Rt_2_(if_addr_j[20]), .i_addr_Rt_1_(if_addr_j[19]), 
        .i_addr_Rt_0_(if_addr_j[18]) );
  DFC3 u_fetch_pipe_instr_reg_16_ ( .D(read_instruction[16]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[18]), .QN(n187) );
  DFC3 u_fetch_pipe_instr_reg_17_ ( .D(read_instruction[17]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[19]), .QN(n198) );
  DFC3 u_fetch_pipe_instr_reg_18_ ( .D(read_instruction[18]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[20]), .QN(n197) );
  DFC3 u_fetch_pipe_instr_reg_19_ ( .D(read_instruction[19]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[21]), .QN(n201) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_16_ ( .D(u_decode_n1), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[31]) );
  DFC3 u_decode_pipe_con_Efbmux_reg_1_ ( .D(u_decode_for_o_con_fb[1]), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[1]) );
  DFC3 u_decode_pipe_con_Efbmux_reg_2_ ( .D(u_decode_for_o_con_fb[2]), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[2]) );
  DFC3 u_fetch_u_pc_program_counter_reg_2_ ( .D(n135), .C(clk), .RN(rst_n), 
        .Q(instruction_address[2]), .QN(u_fetch_jmux_i_addr_pc4_2_) );
  DFC3 u_decode_pipe_con_Efbmux_reg_0_ ( .D(u_decode_for_o_con_fb[0]), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efbmux[0]) );
  DFC3 u_fetch_u_pc_program_counter_reg_3_ ( .D(n134), .C(clk), .RN(rst_n), 
        .Q(instruction_address[3]) );
  DFC3 u_decode_pipe_con_Efamux_reg_1_ ( .D(u_decode_for_o_con_fa_1_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[1]) );
  DFC3 u_decode_pipe_con_Efamux_reg_2_ ( .D(u_decode_for_o_con_fa_2_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[2]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_1_ ( .D(if_addr_j[3]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[1]) );
  DFC3 u_decode_pipe_signext_o_data_immD_reg_10_ ( .D(if_addr_j[12]), .C(clk), 
        .RN(rst_n), .Q(ex_data_immext[10]) );
  DFC3 u_mem_pipe_con_Wmemtoreg_reg ( .D(mem_con_Wmemtoreg), .C(clk), .RN(
        rst_n), .Q(wb_con_Wmemtoreg) );
  XNR21 u_decode_add_x_16_U17 ( .A(u_decode_add_x_16_n3), .B(
        u_decode_add_x_16_n39), .Q(u_decode_pcadd_o_addr_pcbranchE[21]) );
  XNR21 u_decode_add_x_16_U31 ( .A(u_decode_add_x_16_n5), .B(
        u_decode_add_x_16_n47), .Q(u_decode_pcadd_o_addr_pcbranchE[19]) );
  XNR21 u_decode_add_x_16_U45 ( .A(u_decode_add_x_16_n7), .B(
        u_decode_add_x_16_n55), .Q(u_decode_pcadd_o_addr_pcbranchE[17]) );
  XNR21 u_decode_add_x_16_U59 ( .A(u_decode_add_x_16_n9), .B(
        u_decode_add_x_16_n63), .Q(u_decode_pcadd_o_addr_pcbranchE[15]) );
  XNR21 u_decode_add_x_16_U73 ( .A(u_decode_add_x_16_n11), .B(
        u_decode_add_x_16_n71), .Q(u_decode_pcadd_o_addr_pcbranchE[13]) );
  XNR21 u_decode_add_x_16_U87 ( .A(u_decode_add_x_16_n13), .B(
        u_decode_add_x_16_n79), .Q(u_decode_pcadd_o_addr_pcbranchE[11]) );
  XNR21 u_decode_add_x_16_U101 ( .A(u_decode_add_x_16_n15), .B(
        u_decode_add_x_16_n90), .Q(u_decode_pcadd_o_addr_pcbranchE[9]) );
  XNR21 u_decode_add_x_16_U126 ( .A(u_decode_add_x_16_n18), .B(
        u_decode_add_x_16_n103), .Q(u_decode_pcadd_o_addr_pcbranchE[6]) );
  XNR21 u_decode_add_x_16_U134 ( .A(u_decode_add_x_16_n19), .B(
        u_decode_add_x_16_n109), .Q(u_decode_pcadd_o_addr_pcbranchE[5]) );
  NOR21 u_decode_add_x_16_U124 ( .A(id_addr_pc4[7]), .B(if_addr_j[7]), .Q(
        u_decode_add_x_16_n96) );
  NOR21 u_decode_add_x_16_U110 ( .A(id_addr_pc4[9]), .B(if_addr_j[9]), .Q(
        u_decode_add_x_16_n88) );
  NOR21 u_decode_add_x_16_U116 ( .A(id_addr_pc4[8]), .B(if_addr_j[8]), .Q(
        u_decode_add_x_16_n91) );
  NOR21 u_decode_add_x_16_U141 ( .A(id_addr_pc4[5]), .B(if_addr_j[5]), .Q(
        u_decode_add_x_16_n107) );
  NOR21 u_decode_add_x_16_U93 ( .A(id_addr_pc4[11]), .B(if_addr_j[11]), .Q(
        u_decode_add_x_16_n77) );
  NOR21 u_decode_add_x_16_U120 ( .A(u_decode_add_x_16_n96), .B(
        u_decode_add_x_16_n101), .Q(u_decode_add_x_16_n94) );
  NOR21 u_decode_add_x_16_U106 ( .A(u_decode_add_x_16_n88), .B(
        u_decode_add_x_16_n91), .Q(u_decode_add_x_16_n86) );
  NAND22 u_decode_add_x_16_U104 ( .A(u_decode_add_x_16_n94), .B(
        u_decode_add_x_16_n86), .Q(u_decode_add_x_16_n84) );
  OAI212 u_decode_add_x_16_U151 ( .A(u_decode_add_x_16_n117), .B(
        u_decode_add_x_16_n114), .C(u_decode_add_x_16_n115), .Q(
        u_decode_add_x_16_n113) );
  NOR21 u_decode_add_x_16_U147 ( .A(id_addr_pc4[4]), .B(if_addr_j[4]), .Q(
        u_decode_add_x_16_n110) );
  NOR21 u_decode_add_x_16_U137 ( .A(u_decode_add_x_16_n107), .B(
        u_decode_add_x_16_n110), .Q(u_decode_add_x_16_n105) );
  AOI211 u_decode_add_x_16_U105 ( .A(u_decode_add_x_16_n95), .B(
        u_decode_add_x_16_n86), .C(u_decode_add_x_16_n87), .Q(
        u_decode_add_x_16_n85) );
  OAI212 u_decode_add_x_16_U103 ( .A(u_decode_add_x_16_n84), .B(
        u_decode_add_x_16_n104), .C(u_decode_add_x_16_n85), .Q(
        u_decode_add_x_16_n83) );
  NOR21 u_decode_add_x_16_U89 ( .A(u_decode_add_x_16_n77), .B(
        u_decode_add_x_16_n80), .Q(u_decode_add_x_16_n75) );
  OAI212 u_decode_add_x_16_U82 ( .A(u_decode_add_x_16_n72), .B(
        u_decode_add_x_16_n74), .C(u_decode_add_x_16_n73), .Q(
        u_decode_add_x_16_n71) );
  OAI212 u_decode_add_x_16_U68 ( .A(u_decode_add_x_16_n64), .B(
        u_decode_add_x_16_n66), .C(u_decode_add_x_16_n65), .Q(
        u_decode_add_x_16_n63) );
  OAI212 u_decode_add_x_16_U54 ( .A(u_decode_add_x_16_n56), .B(
        u_decode_add_x_16_n58), .C(u_decode_add_x_16_n57), .Q(
        u_decode_add_x_16_n55) );
  OAI212 u_decode_add_x_16_U40 ( .A(u_decode_add_x_16_n48), .B(
        u_decode_add_x_16_n50), .C(u_decode_add_x_16_n49), .Q(
        u_decode_add_x_16_n47) );
  OAI212 u_decode_add_x_16_U26 ( .A(u_decode_add_x_16_n40), .B(
        u_decode_add_x_16_n42), .C(u_decode_add_x_16_n41), .Q(
        u_decode_add_x_16_n39) );
  OAI212 u_decode_add_x_16_U12 ( .A(u_decode_add_x_16_n32), .B(
        u_decode_add_x_16_n34), .C(u_decode_add_x_16_n33), .Q(
        u_decode_add_x_16_n31) );
  NOR20 u_decode_add_x_16_U37 ( .A(id_addr_pc4[19]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n45) );
  NOR20 u_decode_add_x_16_U51 ( .A(id_addr_pc4[17]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n53) );
  NAND22 u_decode_add_x_16_U63 ( .A(u_decode_add_x_16_n59), .B(
        u_decode_add_x_16_n62), .Q(u_decode_add_x_16_n9) );
  NAND22 u_decode_add_x_16_U160 ( .A(if_addr_j[2]), .B(id_addr_pc4[2]), .Q(
        u_decode_add_x_16_n117) );
  NAND22 u_decode_add_x_16_U148 ( .A(if_addr_j[4]), .B(id_addr_pc4[4]), .Q(
        u_decode_add_x_16_n111) );
  ADD31 u_decode_add_x_16_U3 ( .A(if_addr_j[17]), .B(if_addr_j[30]), .CI(
        u_decode_add_x_16_n24), .CO(u_decode_add_x_16_n23), .S(
        u_decode_pcadd_o_addr_pcbranchE[30]) );
  ADD31 u_decode_add_x_16_U4 ( .A(if_addr_j[17]), .B(if_addr_j[29]), .CI(
        u_decode_add_x_16_n25), .CO(u_decode_add_x_16_n24), .S(
        u_decode_pcadd_o_addr_pcbranchE[29]) );
  NAND22 u_decode_add_x_16_U133 ( .A(if_addr_j[6]), .B(id_addr_pc4[6]), .Q(
        u_decode_add_x_16_n102) );
  NAND22 u_decode_add_x_16_U117 ( .A(if_addr_j[8]), .B(id_addr_pc4[8]), .Q(
        u_decode_add_x_16_n92) );
  DFC3 u_decode_pipe_con_Efamux_reg_0_ ( .D(u_decode_for_o_con_fa_0_), .C(clk), 
        .RN(rst_n), .Q(for_o_con_Efamux[0]) );
  ADD22 add_x_4_U3 ( .A(add_x_4_n3), .B(instruction_address[29]), .CO(
        add_x_4_n2), .S(u_fetch_jmux_i_addr_pc4_29_) );
  ADD22 add_x_4_U4 ( .A(add_x_4_n4), .B(instruction_address[28]), .CO(
        add_x_4_n3), .S(u_fetch_jmux_i_addr_pc4_28_) );
  DFC3 u_fetch_pipe_instr_reg_20_ ( .D(read_instruction[20]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[22]), .QN(n199) );
  DFC3 u_mem_pipe_addr_regdst_reg_0_ ( .D(mem_addr_regdst[0]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[0]) );
  DFC3 u_mem_pipe_addr_regdst_reg_3_ ( .D(mem_addr_regdst[3]), .C(clk), .RN(
        rst_n), .Q(id_addr_Wregwrite[3]) );
  NOR21 u_decode_add_x_16_U132 ( .A(id_addr_pc4[6]), .B(if_addr_j[6]), .Q(
        u_decode_add_x_16_n101) );
  NAND21 u_decode_add_x_16_U125 ( .A(if_addr_j[7]), .B(id_addr_pc4[7]), .Q(
        u_decode_add_x_16_n97) );
  NAND21 u_decode_add_x_16_U142 ( .A(if_addr_j[5]), .B(id_addr_pc4[5]), .Q(
        u_decode_add_x_16_n108) );
  NOR21 u_decode_add_x_16_U154 ( .A(id_addr_pc4[3]), .B(if_addr_j[3]), .Q(
        u_decode_add_x_16_n114) );
  NAND22 u_decode_add_x_16_U155 ( .A(if_addr_j[3]), .B(id_addr_pc4[3]), .Q(
        u_decode_add_x_16_n115) );
  NOR21 u_decode_add_x_16_U57 ( .A(id_addr_pc4[16]), .B(if_addr_j[16]), .Q(
        u_decode_add_x_16_n56) );
  NAND22 u_decode_add_x_16_U58 ( .A(if_addr_j[16]), .B(id_addr_pc4[16]), .Q(
        u_decode_add_x_16_n57) );
  NAND22 u_decode_add_x_16_U86 ( .A(if_addr_j[12]), .B(id_addr_pc4[12]), .Q(
        u_decode_add_x_16_n73) );
  NOR21 u_decode_add_x_16_U85 ( .A(id_addr_pc4[12]), .B(if_addr_j[12]), .Q(
        u_decode_add_x_16_n72) );
  NAND22 u_decode_add_x_16_U80 ( .A(if_addr_j[13]), .B(id_addr_pc4[13]), .Q(
        u_decode_add_x_16_n70) );
  NOR21 u_decode_add_x_16_U79 ( .A(id_addr_pc4[13]), .B(if_addr_j[13]), .Q(
        u_decode_add_x_16_n69) );
  NOR21 u_decode_add_x_16_U65 ( .A(id_addr_pc4[15]), .B(if_addr_j[15]), .Q(
        u_decode_add_x_16_n61) );
  NAND22 u_decode_add_x_16_U72 ( .A(if_addr_j[14]), .B(id_addr_pc4[14]), .Q(
        u_decode_add_x_16_n65) );
  NOR21 u_decode_add_x_16_U71 ( .A(id_addr_pc4[14]), .B(if_addr_j[14]), .Q(
        u_decode_add_x_16_n64) );
  NAND22 u_decode_add_x_16_U66 ( .A(if_addr_j[15]), .B(id_addr_pc4[15]), .Q(
        u_decode_add_x_16_n62) );
  NAND21 u_decode_add_x_16_U94 ( .A(if_addr_j[11]), .B(id_addr_pc4[11]), .Q(
        u_decode_add_x_16_n78) );
  NOR21 u_decode_add_x_16_U99 ( .A(id_addr_pc4[10]), .B(if_addr_j[10]), .Q(
        u_decode_add_x_16_n80) );
  NAND22 u_decode_add_x_16_U100 ( .A(if_addr_j[10]), .B(id_addr_pc4[10]), .Q(
        u_decode_add_x_16_n81) );
  NAND21 u_decode_add_x_16_U111 ( .A(if_addr_j[9]), .B(id_addr_pc4[9]), .Q(
        u_decode_add_x_16_n89) );
  NAND21 u_decode_add_x_16_U38 ( .A(if_addr_j[17]), .B(id_addr_pc4[19]), .Q(
        u_decode_add_x_16_n46) );
  NOR21 u_decode_add_x_16_U43 ( .A(id_addr_pc4[18]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n48) );
  NAND21 u_decode_add_x_16_U44 ( .A(if_addr_j[17]), .B(id_addr_pc4[18]), .Q(
        u_decode_add_x_16_n49) );
  OAI211 u_decode_add_x_16_U107 ( .A(u_decode_add_x_16_n92), .B(
        u_decode_add_x_16_n88), .C(u_decode_add_x_16_n89), .Q(
        u_decode_add_x_16_n87) );
  OAI211 u_decode_add_x_16_U138 ( .A(u_decode_add_x_16_n111), .B(
        u_decode_add_x_16_n107), .C(u_decode_add_x_16_n108), .Q(
        u_decode_add_x_16_n106) );
  NAND21 u_decode_add_x_16_U30 ( .A(if_addr_j[17]), .B(id_addr_pc4[20]), .Q(
        u_decode_add_x_16_n41) );
  NOR21 u_decode_add_x_16_U29 ( .A(id_addr_pc4[20]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n40) );
  NAND21 u_decode_add_x_16_U52 ( .A(if_addr_j[17]), .B(id_addr_pc4[17]), .Q(
        u_decode_add_x_16_n54) );
  OAI211 u_decode_add_x_16_U90 ( .A(u_decode_add_x_16_n81), .B(
        u_decode_add_x_16_n77), .C(u_decode_add_x_16_n78), .Q(
        u_decode_add_x_16_n76) );
  OAI211 u_decode_add_x_16_U121 ( .A(u_decode_add_x_16_n102), .B(
        u_decode_add_x_16_n96), .C(u_decode_add_x_16_n97), .Q(
        u_decode_add_x_16_n95) );
  NAND22 u_decode_add_x_16_U16 ( .A(if_addr_j[17]), .B(id_addr_pc4[22]), .Q(
        u_decode_add_x_16_n33) );
  NOR21 u_decode_add_x_16_U15 ( .A(id_addr_pc4[22]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n32) );
  NAND22 u_decode_add_x_16_U130 ( .A(u_decode_add_x_16_n99), .B(
        u_decode_add_x_16_n102), .Q(u_decode_add_x_16_n18) );
  NAND22 u_decode_add_x_16_U77 ( .A(u_decode_add_x_16_n67), .B(
        u_decode_add_x_16_n70), .Q(u_decode_add_x_16_n11) );
  AOI211 u_decode_add_x_16_U136 ( .A(u_decode_add_x_16_n113), .B(
        u_decode_add_x_16_n105), .C(u_decode_add_x_16_n106), .Q(
        u_decode_add_x_16_n104) );
  NAND22 u_decode_add_x_16_U108 ( .A(u_decode_add_x_16_n131), .B(
        u_decode_add_x_16_n89), .Q(u_decode_add_x_16_n15) );
  NAND22 u_decode_add_x_16_U91 ( .A(u_decode_add_x_16_n129), .B(
        u_decode_add_x_16_n78), .Q(u_decode_add_x_16_n13) );
  NAND22 u_decode_add_x_16_U139 ( .A(u_decode_add_x_16_n135), .B(
        u_decode_add_x_16_n108), .Q(u_decode_add_x_16_n19) );
  OAI211 u_decode_add_x_16_U144 ( .A(u_decode_add_x_16_n110), .B(
        u_decode_add_x_16_n112), .C(u_decode_add_x_16_n111), .Q(
        u_decode_add_x_16_n109) );
  AOI211 u_decode_add_x_16_U88 ( .A(u_decode_add_x_16_n83), .B(
        u_decode_add_x_16_n75), .C(u_decode_add_x_16_n76), .Q(
        u_decode_add_x_16_n74) );
  AOI211 u_decode_add_x_16_U119 ( .A(u_decode_add_x_16_n103), .B(
        u_decode_add_x_16_n94), .C(u_decode_add_x_16_n95), .Q(
        u_decode_add_x_16_n93) );
  OAI211 u_decode_add_x_16_U96 ( .A(u_decode_add_x_16_n80), .B(
        u_decode_add_x_16_n82), .C(u_decode_add_x_16_n81), .Q(
        u_decode_add_x_16_n79) );
  OAI211 u_decode_add_x_16_U113 ( .A(u_decode_add_x_16_n91), .B(
        u_decode_add_x_16_n93), .C(u_decode_add_x_16_n92), .Q(
        u_decode_add_x_16_n90) );
  AOI211 u_decode_add_x_16_U74 ( .A(u_decode_add_x_16_n71), .B(
        u_decode_add_x_16_n67), .C(u_decode_add_x_16_n68), .Q(
        u_decode_add_x_16_n66) );
  AOI211 u_decode_add_x_16_U60 ( .A(u_decode_add_x_16_n63), .B(
        u_decode_add_x_16_n59), .C(u_decode_add_x_16_n60), .Q(
        u_decode_add_x_16_n58) );
  AOI211 u_decode_add_x_16_U46 ( .A(u_decode_add_x_16_n55), .B(
        u_decode_add_x_16_n51), .C(u_decode_add_x_16_n52), .Q(
        u_decode_add_x_16_n50) );
  AOI211 u_decode_add_x_16_U32 ( .A(u_decode_add_x_16_n47), .B(
        u_decode_add_x_16_n43), .C(u_decode_add_x_16_n44), .Q(
        u_decode_add_x_16_n42) );
  ADD22 add_x_1_U4 ( .A(add_x_1_n4), .B(mem_data_pc4[28]), .CO(add_x_1_n3), 
        .S(u_mem_pc8[28]) );
  NAND22 u_decode_add_x_16_U24 ( .A(if_addr_j[17]), .B(id_addr_pc4[21]), .Q(
        u_decode_add_x_16_n38) );
  NOR21 u_decode_add_x_16_U23 ( .A(id_addr_pc4[21]), .B(if_addr_j[17]), .Q(
        u_decode_add_x_16_n37) );
  NAND21 u_decode_add_x_16_U35 ( .A(u_decode_add_x_16_n43), .B(
        u_decode_add_x_16_n46), .Q(u_decode_add_x_16_n5) );
  NAND21 u_decode_add_x_16_U49 ( .A(u_decode_add_x_16_n51), .B(
        u_decode_add_x_16_n54), .Q(u_decode_add_x_16_n7) );
  NAND21 u_decode_add_x_16_U21 ( .A(u_decode_add_x_16_n35), .B(
        u_decode_add_x_16_n38), .Q(u_decode_add_x_16_n3) );
  ADD32 u_decode_add_x_16_U10 ( .A(if_addr_j[17]), .B(id_addr_pc4[23]), .CI(
        u_decode_add_x_16_n31), .CO(u_decode_add_x_16_n30), .S(
        u_decode_pcadd_o_addr_pcbranchE[23]) );
  ADD32 u_decode_add_x_16_U9 ( .A(if_addr_j[17]), .B(id_addr_pc4[24]), .CI(
        u_decode_add_x_16_n30), .CO(u_decode_add_x_16_n29), .S(
        u_decode_pcadd_o_addr_pcbranchE[24]) );
  ADD32 u_decode_add_x_16_U8 ( .A(if_addr_j[17]), .B(id_addr_pc4[25]), .CI(
        u_decode_add_x_16_n29), .CO(u_decode_add_x_16_n28), .S(
        u_decode_pcadd_o_addr_pcbranchE[25]) );
  ADD32 u_decode_add_x_16_U7 ( .A(if_addr_j[17]), .B(id_addr_pc4[26]), .CI(
        u_decode_add_x_16_n28), .CO(u_decode_add_x_16_n27), .S(
        u_decode_pcadd_o_addr_pcbranchE[26]) );
  ADD32 u_decode_add_x_16_U6 ( .A(if_addr_j[17]), .B(id_addr_pc4[27]), .CI(
        u_decode_add_x_16_n27), .CO(u_decode_add_x_16_n26), .S(
        u_decode_pcadd_o_addr_pcbranchE[27]) );
  ADD32 u_decode_add_x_16_U5 ( .A(if_addr_j[17]), .B(if_addr_j[28]), .CI(
        u_decode_add_x_16_n26), .CO(u_decode_add_x_16_n25), .S(
        u_decode_pcadd_o_addr_pcbranchE[28]) );
  AOI211 u_decode_add_x_16_U18 ( .A(u_decode_add_x_16_n39), .B(
        u_decode_add_x_16_n35), .C(u_decode_add_x_16_n36), .Q(
        u_decode_add_x_16_n34) );
  DFC3 u_fetch_pipe_instr_reg_15_ ( .D(read_instruction[15]), .C(clk), .RN(
        rst_n), .Q(if_addr_j[17]), .QN(n188) );
  OAI2111 U204 ( .A(n405), .B(n404), .C(n403), .D(n402), .Q(n107) );
  BUF2 U205 ( .A(n400), .Q(n169) );
  BUF2 U206 ( .A(n401), .Q(n205) );
  NOR22 U207 ( .A(n171), .B(n173), .Q(n174) );
  NAND22 U208 ( .A(add_x_1_n28), .B(mem_data_pc4[4]), .Q(n175) );
  NAND22 U209 ( .A(add_x_4_n2), .B(instruction_address[30]), .Q(n181) );
  NAND22 U210 ( .A(add_x_4_n12), .B(instruction_address[20]), .Q(n178) );
  OAI220 U211 ( .A(if_con_j[0]), .B(n305), .C(if_con_j[1]), .D(n311), .Q(n140)
         );
  NOR30 U212 ( .A(if_con_b), .B(n398), .C(n140), .Q(n310) );
  CLKIN0 U213 ( .A(u_decode_add_x_16_n49), .Q(n141) );
  NOR20 U214 ( .A(u_decode_add_x_16_n48), .B(n141), .Q(n142) );
  XNR20 U215 ( .A(u_decode_add_x_16_n50), .B(n142), .Q(
        u_decode_pcadd_o_addr_pcbranchE[18]) );
  CLKIN0 U216 ( .A(u_decode_add_x_16_n73), .Q(n143) );
  NOR20 U217 ( .A(u_decode_add_x_16_n72), .B(n143), .Q(n144) );
  XNR20 U218 ( .A(u_decode_add_x_16_n74), .B(n144), .Q(
        u_decode_pcadd_o_addr_pcbranchE[12]) );
  CLKIN0 U219 ( .A(u_decode_add_x_16_n92), .Q(n145) );
  NOR20 U220 ( .A(u_decode_add_x_16_n91), .B(n145), .Q(n146) );
  XNR20 U221 ( .A(u_decode_add_x_16_n93), .B(n146), .Q(
        u_decode_pcadd_o_addr_pcbranchE[8]) );
  CLKIN0 U222 ( .A(u_decode_add_x_16_n115), .Q(n147) );
  NOR20 U223 ( .A(u_decode_add_x_16_n114), .B(n147), .Q(n148) );
  XNR20 U224 ( .A(u_decode_add_x_16_n117), .B(n148), .Q(
        u_decode_pcadd_o_addr_pcbranchE[3]) );
  XOR30 U225 ( .A(if_addr_j[17]), .B(if_addr_j[31]), .C(u_decode_add_x_16_n23), 
        .Q(u_decode_pcadd_o_addr_pcbranchE[31]) );
  CLKIN0 U226 ( .A(u_decode_add_x_16_n33), .Q(n149) );
  NOR20 U227 ( .A(u_decode_add_x_16_n32), .B(n149), .Q(n150) );
  XNR20 U228 ( .A(u_decode_add_x_16_n34), .B(n150), .Q(
        u_decode_pcadd_o_addr_pcbranchE[22]) );
  CLKIN0 U229 ( .A(u_decode_add_x_16_n41), .Q(n151) );
  NOR20 U230 ( .A(u_decode_add_x_16_n40), .B(n151), .Q(n152) );
  XNR20 U231 ( .A(u_decode_add_x_16_n42), .B(n152), .Q(
        u_decode_pcadd_o_addr_pcbranchE[20]) );
  CLKIN0 U232 ( .A(u_decode_add_x_16_n57), .Q(n153) );
  NOR20 U233 ( .A(u_decode_add_x_16_n56), .B(n153), .Q(n154) );
  XNR20 U234 ( .A(u_decode_add_x_16_n58), .B(n154), .Q(
        u_decode_pcadd_o_addr_pcbranchE[16]) );
  CLKIN0 U235 ( .A(u_decode_add_x_16_n65), .Q(n155) );
  NOR20 U236 ( .A(u_decode_add_x_16_n64), .B(n155), .Q(n156) );
  XNR20 U237 ( .A(u_decode_add_x_16_n66), .B(n156), .Q(
        u_decode_pcadd_o_addr_pcbranchE[14]) );
  CLKIN0 U238 ( .A(u_decode_add_x_16_n81), .Q(n157) );
  NOR20 U239 ( .A(u_decode_add_x_16_n80), .B(n157), .Q(n158) );
  XNR20 U240 ( .A(u_decode_add_x_16_n82), .B(n158), .Q(
        u_decode_pcadd_o_addr_pcbranchE[10]) );
  CLKIN0 U241 ( .A(u_decode_add_x_16_n102), .Q(n159) );
  AOI210 U242 ( .A(u_decode_add_x_16_n103), .B(u_decode_add_x_16_n99), .C(n159), .Q(n160) );
  CLKIN0 U243 ( .A(u_decode_add_x_16_n97), .Q(n161) );
  NOR20 U244 ( .A(u_decode_add_x_16_n96), .B(n161), .Q(n162) );
  XNR20 U245 ( .A(n160), .B(n162), .Q(u_decode_pcadd_o_addr_pcbranchE[7]) );
  CLKIN0 U246 ( .A(u_decode_add_x_16_n111), .Q(n163) );
  NOR20 U247 ( .A(u_decode_add_x_16_n110), .B(n163), .Q(n164) );
  XNR20 U248 ( .A(u_decode_add_x_16_n112), .B(n164), .Q(
        u_decode_pcadd_o_addr_pcbranchE[4]) );
  OAI210 U249 ( .A(if_addr_j[2]), .B(id_addr_pc4[2]), .C(
        u_decode_add_x_16_n117), .Q(n165) );
  CLKIN0 U250 ( .A(n165), .Q(u_decode_pcadd_o_addr_pcbranchE[2]) );
  MUX21 U251 ( .A(data_address[31]), .B(u_mem_pc8[31]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[31]) );
  XNR20 U252 ( .A(n171), .B(mem_data_pc4[13]), .Q(n166) );
  MUX21 U253 ( .A(data_address[13]), .B(n166), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[13]) );
  CLKIN0 U254 ( .A(data_address[2]), .Q(n167) );
  IMUX20 U255 ( .A(n167), .B(mem_data_pc4[2]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[2]) );
  XNR20 U256 ( .A(n180), .B(instruction_address[18]), .Q(
        u_fetch_jmux_i_addr_pc4_18_) );
  NAND22 U257 ( .A(add_x_1_n6), .B(mem_data_pc4[26]), .Q(n177) );
  XOR20 U258 ( .A(add_x_1_n6), .B(mem_data_pc4[26]), .Q(u_mem_pc8[26]) );
  INV2 U259 ( .A(u_fetch_jmux_i_addr_pc4_26_), .Q(n388) );
  AOI221 U260 ( .A(n205), .B(id_data_jr[15]), .C(n169), .D(if_addr_j[15]), .Q(
        n353) );
  AOI221 U261 ( .A(n205), .B(id_data_jr[6]), .C(n169), .D(if_addr_j[6]), .Q(
        n326) );
  AOI221 U262 ( .A(n205), .B(id_data_jr[7]), .C(n169), .D(if_addr_j[7]), .Q(
        n329) );
  AOI221 U263 ( .A(n205), .B(id_data_jr[4]), .C(n169), .D(if_addr_j[4]), .Q(
        n320) );
  AOI221 U264 ( .A(n205), .B(id_data_jr[12]), .C(n169), .D(if_addr_j[12]), .Q(
        n344) );
  AOI221 U265 ( .A(n205), .B(id_data_jr[2]), .C(n169), .D(if_addr_j[2]), .Q(
        n315) );
  AOI221 U266 ( .A(n205), .B(id_data_jr[11]), .C(n169), .D(if_addr_j[11]), .Q(
        n341) );
  AOI221 U267 ( .A(n205), .B(id_data_jr[8]), .C(n169), .D(if_addr_j[8]), .Q(
        n332) );
  AOI221 U268 ( .A(n205), .B(id_data_jr[10]), .C(n169), .D(if_addr_j[10]), .Q(
        n338) );
  AOI221 U269 ( .A(n205), .B(id_data_jr[13]), .C(n169), .D(if_addr_j[13]), .Q(
        n347) );
  AOI221 U270 ( .A(n205), .B(id_data_jr[14]), .C(n169), .D(if_addr_j[14]), .Q(
        n350) );
  AOI221 U271 ( .A(n205), .B(id_data_jr[5]), .C(n169), .D(if_addr_j[5]), .Q(
        n323) );
  NOR22 U272 ( .A(n306), .B(n398), .Q(n399) );
  NOR40 U273 ( .A(if_con_b), .B(if_con_j[1]), .C(n398), .D(n311), .Q(n400) );
  INV2 U274 ( .A(u_fetch_jmux_i_addr_pc4_18_), .Q(n364) );
  MUX22 U275 ( .A(data_address[17]), .B(u_mem_pc8[17]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[17]) );
  INV3 U276 ( .A(u_decode_add_x_16_n104), .Q(u_decode_add_x_16_n103) );
  INV3 U277 ( .A(n175), .Q(add_x_1_n27) );
  INV2 U278 ( .A(n294), .Q(n295) );
  CLKIN3 U279 ( .A(mem_data_pc4[13]), .Q(n173) );
  INV2 U280 ( .A(u_fetch_jmux_i_addr_pc4_27_), .Q(n391) );
  NAND24 U281 ( .A(add_x_1_n9), .B(mem_data_pc4[23]), .Q(n170) );
  INV3 U282 ( .A(n310), .Q(n405) );
  NAND24 U283 ( .A(add_x_1_n20), .B(mem_data_pc4[12]), .Q(n171) );
  AOI210 U284 ( .A(n293), .B(n294), .C(u_decode_control_o_con_aluop_1_), .Q(
        n292) );
  INV3 U285 ( .A(u_decode_add_x_16_n37), .Q(u_decode_add_x_16_n35) );
  INV3 U286 ( .A(u_decode_add_x_16_n38), .Q(u_decode_add_x_16_n36) );
  MUX22 U287 ( .A(data_address[30]), .B(u_mem_pc8[30]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[30]) );
  XOR21 U288 ( .A(add_x_1_n1), .B(mem_data_pc4[31]), .Q(u_mem_pc8[31]) );
  MUX22 U289 ( .A(data_address[29]), .B(u_mem_pc8[29]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[29]) );
  MUX22 U290 ( .A(data_address[28]), .B(u_mem_pc8[28]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[28]) );
  MUX22 U291 ( .A(data_address[27]), .B(u_mem_pc8[27]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[27]) );
  INV2 U292 ( .A(u_fetch_jmux_i_addr_pc4_29_), .Q(n397) );
  INV2 U293 ( .A(u_fetch_jmux_i_addr_pc4_28_), .Q(n394) );
  MUX22 U294 ( .A(data_address[26]), .B(u_mem_pc8[26]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[26]) );
  MUX22 U295 ( .A(data_address[25]), .B(u_mem_pc8[25]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[25]) );
  MUX22 U296 ( .A(data_address[24]), .B(u_mem_pc8[24]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[24]) );
  INV10 U297 ( .A(n184), .Q(add_x_4_n5) );
  OAI211 U298 ( .A(n309), .B(n202), .C(n307), .Q(n137) );
  INV2 U299 ( .A(u_fetch_jmux_i_addr_pc4_25_), .Q(n385) );
  OAI211 U300 ( .A(n309), .B(n203), .C(n308), .Q(n136) );
  INV2 U301 ( .A(u_fetch_jmux_i_addr_pc4_24_), .Q(n382) );
  AOI221 U302 ( .A(n205), .B(id_data_jr[16]), .C(n169), .D(if_addr_j[16]), .Q(
        n356) );
  INV2 U303 ( .A(u_fetch_jmux_i_addr_pc4_23_), .Q(n379) );
  AOI221 U304 ( .A(n205), .B(id_data_jr[30]), .C(n169), .D(if_addr_j[30]), .Q(
        n402) );
  AOI221 U305 ( .A(n205), .B(id_data_jr[31]), .C(n169), .D(if_addr_j[31]), .Q(
        n312) );
  AOI221 U306 ( .A(n205), .B(id_data_jr[3]), .C(n169), .D(if_addr_j[3]), .Q(
        n317) );
  AOI221 U307 ( .A(n205), .B(id_data_jr[29]), .C(n169), .D(if_addr_j[29]), .Q(
        n395) );
  NAND23 U308 ( .A(add_x_1_n10), .B(mem_data_pc4[22]), .Q(n172) );
  MUX22 U309 ( .A(data_address[21]), .B(u_mem_pc8[21]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[21]) );
  INV2 U310 ( .A(u_fetch_jmux_i_addr_pc4_22_), .Q(n376) );
  NOR40 U311 ( .A(if_con_b), .B(if_con_j[0]), .C(n398), .D(n305), .Q(n401) );
  MUX22 U312 ( .A(data_address[20]), .B(u_mem_pc8[20]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[20]) );
  INV2 U313 ( .A(u_fetch_jmux_i_addr_pc4_21_), .Q(n373) );
  MUX22 U314 ( .A(data_address[19]), .B(u_mem_pc8[19]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[19]) );
  INV1 U315 ( .A(u_fetch_jmux_i_addr_pc4_20_), .Q(n370) );
  INV2 U316 ( .A(u_fetch_jmux_i_addr_pc4_19_), .Q(n367) );
  INV1 U317 ( .A(u_fetch_jmux_i_addr_pc4_17_), .Q(n361) );
  INV2 U318 ( .A(u_fetch_jmux_i_addr_pc4_16_), .Q(n358) );
  INV2 U319 ( .A(u_fetch_jmux_i_addr_pc4_15_), .Q(n355) );
  INV2 U320 ( .A(u_fetch_jmux_i_addr_pc4_14_), .Q(n352) );
  INV2 U321 ( .A(u_fetch_jmux_i_addr_pc4_13_), .Q(n349) );
  INV2 U322 ( .A(u_fetch_jmux_i_addr_pc4_12_), .Q(n346) );
  INV2 U323 ( .A(u_fetch_jmux_i_addr_pc4_11_), .Q(n343) );
  INV2 U324 ( .A(u_fetch_jmux_i_addr_pc4_10_), .Q(n340) );
  OAI2111 U325 ( .A(mem_addr_regdst[1]), .B(n269), .C(n270), .D(n271), .Q(n260) );
  INV2 U326 ( .A(u_fetch_jmux_i_addr_pc4_9_), .Q(n337) );
  AOI211 U327 ( .A(n208), .B(n209), .C(n188), .Q(u_decode_n1) );
  INV2 U328 ( .A(u_fetch_jmux_i_addr_pc4_8_), .Q(n334) );
  INV2 U329 ( .A(n256), .Q(n255) );
  OAI210 U330 ( .A(n300), .B(n301), .C(n209), .Q(
        u_decode_control_o_con_aluop_3_) );
  INV2 U331 ( .A(u_decode_control_o_con_aluop_4_), .Q(n209) );
  INV2 U332 ( .A(u_fetch_jmux_i_addr_pc4_7_), .Q(n331) );
  OAI211 U333 ( .A(n222), .B(n223), .C(n224), .Q(u_decode_for_o_con_fb[2]) );
  NAND31 U334 ( .A(ex_con_Wregwrite), .B(n239), .C(n240), .Q(n226) );
  INV2 U335 ( .A(n259), .Q(n257) );
  INV2 U336 ( .A(u_fetch_jmux_i_addr_pc4_6_), .Q(n328) );
  OAI2111 U337 ( .A(for_o_addr_Erd[2]), .B(n190), .C(n277), .D(n278), .Q(n276)
         );
  INV3 U338 ( .A(u_decode_add_x_16_n83), .Q(u_decode_add_x_16_n82) );
  INV2 U339 ( .A(n292), .Q(u_decode_control_o_con_regwrite) );
  OAI210 U340 ( .A(n218), .B(n301), .C(n302), .Q(
        u_decode_control_o_con_aluop_2_) );
  AOI211 U341 ( .A(n304), .B(n298), .C(n192), .Q(
        u_decode_control_o_con_aluop_4_) );
  OAI212 U342 ( .A(id_data_instr[28]), .B(n215), .C(n213), .Q(if_con_j[0]) );
  NAND21 U343 ( .A(ex_con_Wregwrite), .B(n280), .Q(n275) );
  INV1 U344 ( .A(u_decode_control_o_con_aluop_5_), .Q(n302) );
  INV2 U345 ( .A(n223), .Q(n225) );
  INV2 U346 ( .A(u_fetch_jmux_i_addr_pc4_5_), .Q(n325) );
  NOR20 U347 ( .A(n296), .B(n214), .Q(u_decode_control_o_con_regdst) );
  INV2 U348 ( .A(n268), .Q(n261) );
  NOR21 U349 ( .A(n200), .B(n297), .Q(u_decode_control_o_con_memwrite) );
  NAND41 U350 ( .A(for_FWmemread), .B(n285), .C(n286), .D(n268), .Q(n258) );
  OAI211 U351 ( .A(n192), .B(n298), .C(n299), .Q(
        u_decode_control_o_con_memread) );
  NOR21 U352 ( .A(id_data_instr[27]), .B(n216), .Q(n215) );
  NAND31 U353 ( .A(for_FWmemread), .B(n249), .C(n250), .Q(n223) );
  NAND41 U354 ( .A(mem_read), .B(n229), .C(n228), .D(n230), .Q(n224) );
  INV2 U355 ( .A(u_fetch_jmux_i_addr_pc4_4_), .Q(n322) );
  INV2 U356 ( .A(u_decode_add_x_16_n46), .Q(u_decode_add_x_16_n44) );
  INV3 U357 ( .A(u_decode_add_x_16_n113), .Q(u_decode_add_x_16_n112) );
  INV2 U358 ( .A(u_decode_add_x_16_n45), .Q(u_decode_add_x_16_n43) );
  INV2 U359 ( .A(u_decode_add_x_16_n54), .Q(u_decode_add_x_16_n52) );
  INV2 U360 ( .A(u_decode_add_x_16_n53), .Q(u_decode_add_x_16_n51) );
  INV2 U361 ( .A(u_fetch_jmux_i_addr_pc4_3_), .Q(n319) );
  INV1 U362 ( .A(n213), .Q(n296) );
  NAND41 U363 ( .A(mem_read), .B(n265), .C(n266), .D(n267), .Q(n264) );
  INV2 U364 ( .A(u_decode_add_x_16_n77), .Q(u_decode_add_x_16_n129) );
  NAND21 U365 ( .A(id_data_instr[26]), .B(n303), .Q(n298) );
  INV2 U366 ( .A(n303), .Q(n301) );
  NAND22 U367 ( .A(n287), .B(n194), .Q(n268) );
  INV2 U368 ( .A(u_decode_add_x_16_n101), .Q(u_decode_add_x_16_n99) );
  INV1 U369 ( .A(u_decode_add_x_16_n107), .Q(u_decode_add_x_16_n135) );
  INV2 U370 ( .A(u_decode_add_x_16_n88), .Q(u_decode_add_x_16_n131) );
  NAND22 U371 ( .A(n235), .B(n199), .Q(n228) );
  OAI212 U372 ( .A(id_data_instr[28]), .B(n218), .C(n213), .Q(if_con_ifstall)
         );
  AOI311 U373 ( .A(if_addr_j[5]), .B(n217), .C(n196), .D(id_data_instr[26]), 
        .Q(n216) );
  NAND22 U374 ( .A(n300), .B(n189), .Q(n214) );
  MUX22 U375 ( .A(mem_data_alures[8]), .B(wb_data_memout[8]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[8]) );
  MUX22 U376 ( .A(mem_data_alures[25]), .B(wb_data_memout[25]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[25]) );
  MUX22 U377 ( .A(mem_data_alures[26]), .B(wb_data_memout[26]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[26]) );
  MUX22 U378 ( .A(mem_data_alures[19]), .B(wb_data_memout[19]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[19]) );
  MUX22 U379 ( .A(mem_data_alures[20]), .B(wb_data_memout[20]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[20]) );
  INV1 U380 ( .A(mem_con_Wregwrite), .Q(n248) );
  MUX22 U381 ( .A(mem_data_alures[9]), .B(wb_data_memout[9]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[9]) );
  MUX22 U382 ( .A(mem_data_alures[23]), .B(wb_data_memout[23]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[23]) );
  MUX22 U383 ( .A(mem_data_alures[28]), .B(wb_data_memout[28]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[28]) );
  MUX22 U384 ( .A(mem_data_alures[21]), .B(wb_data_memout[21]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[21]) );
  MUX22 U385 ( .A(mem_data_alures[27]), .B(wb_data_memout[27]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[27]) );
  MUX22 U386 ( .A(mem_data_alures[1]), .B(wb_data_memout[1]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[1]) );
  MUX22 U387 ( .A(mem_data_alures[18]), .B(wb_data_memout[18]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[18]) );
  MUX22 U388 ( .A(mem_data_alures[16]), .B(wb_data_memout[16]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[16]) );
  MUX22 U389 ( .A(mem_data_alures[4]), .B(wb_data_memout[4]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[4]) );
  MUX22 U390 ( .A(mem_data_alures[17]), .B(wb_data_memout[17]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[17]) );
  MUX22 U391 ( .A(mem_data_alures[3]), .B(wb_data_memout[3]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[3]) );
  MUX22 U392 ( .A(mem_data_alures[22]), .B(wb_data_memout[22]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[22]) );
  NOR21 U393 ( .A(n186), .B(id_data_instr[30]), .Q(n210) );
  MUX22 U394 ( .A(mem_data_alures[30]), .B(wb_data_memout[30]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[30]) );
  MUX22 U395 ( .A(mem_data_alures[14]), .B(wb_data_memout[14]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[14]) );
  MUX22 U396 ( .A(mem_data_alures[12]), .B(wb_data_memout[12]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[12]) );
  MUX22 U397 ( .A(mem_data_alures[15]), .B(wb_data_memout[15]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[15]) );
  NOR21 U398 ( .A(id_data_instr[27]), .B(n185), .Q(n218) );
  MUX22 U399 ( .A(mem_data_alures[5]), .B(wb_data_memout[5]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[5]) );
  NOR21 U400 ( .A(id_data_instr[26]), .B(id_data_instr[27]), .Q(n300) );
  MUX22 U401 ( .A(mem_data_alures[2]), .B(wb_data_memout[2]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[2]) );
  MUX22 U402 ( .A(mem_data_alures[6]), .B(wb_data_memout[6]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[6]) );
  MUX22 U403 ( .A(mem_data_alures[13]), .B(wb_data_memout[13]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[13]) );
  MUX22 U404 ( .A(mem_data_alures[7]), .B(wb_data_memout[7]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[7]) );
  MUX22 U405 ( .A(mem_data_alures[10]), .B(wb_data_memout[10]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[10]) );
  MUX22 U406 ( .A(mem_data_alures[0]), .B(wb_data_memout[0]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[0]) );
  MUX22 U407 ( .A(mem_data_alures[11]), .B(wb_data_memout[11]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[11]) );
  MUX22 U408 ( .A(mem_data_alures[24]), .B(wb_data_memout[24]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[24]) );
  MUX22 U409 ( .A(mem_data_alures[29]), .B(wb_data_memout[29]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[29]) );
  NOR31 U410 ( .A(id_data_instr[30]), .B(id_data_instr[29]), .C(
        id_data_instr[31]), .Q(n213) );
  MUX22 U411 ( .A(mem_data_alures[31]), .B(wb_data_memout[31]), .S(
        wb_con_Wmemtoreg), .Q(id_data_Wregwrite[31]) );
  INV3 U412 ( .A(n176), .Q(add_x_1_n13) );
  XOR20 U413 ( .A(add_x_1_n9), .B(mem_data_pc4[23]), .Q(u_mem_pc8[23]) );
  XOR20 U414 ( .A(add_x_1_n10), .B(mem_data_pc4[22]), .Q(u_mem_pc8[22]) );
  XOR20 U415 ( .A(add_x_1_n14), .B(mem_data_pc4[18]), .Q(u_mem_pc8[18]) );
  XOR20 U416 ( .A(add_x_1_n20), .B(mem_data_pc4[12]), .Q(u_mem_pc8[12]) );
  XOR20 U417 ( .A(add_x_1_n28), .B(mem_data_pc4[4]), .Q(u_mem_pc8[4]) );
  ADD22 U418 ( .A(add_x_1_n16), .B(mem_data_pc4[16]), .CO(add_x_1_n15), .S(
        u_mem_pc8[16]) );
  ADD22 U419 ( .A(add_x_1_n15), .B(mem_data_pc4[17]), .CO(add_x_1_n14), .S(
        u_mem_pc8[17]) );
  ADD22 U420 ( .A(add_x_1_n12), .B(mem_data_pc4[20]), .CO(add_x_1_n11), .S(
        u_mem_pc8[20]) );
  ADD22 U421 ( .A(add_x_1_n11), .B(mem_data_pc4[21]), .CO(add_x_1_n10), .S(
        u_mem_pc8[21]) );
  ADD22 U422 ( .A(add_x_1_n8), .B(mem_data_pc4[24]), .CO(add_x_1_n7), .S(
        u_mem_pc8[24]) );
  ADD22 U423 ( .A(add_x_1_n3), .B(mem_data_pc4[29]), .CO(add_x_1_n2), .S(
        u_mem_pc8[29]) );
  ADD22 U424 ( .A(add_x_1_n2), .B(mem_data_pc4[30]), .CO(add_x_1_n1), .S(
        u_mem_pc8[30]) );
  ADD22 U425 ( .A(add_x_1_n22), .B(mem_data_pc4[10]), .CO(add_x_1_n21), .S(
        u_mem_pc8[10]) );
  ADD22 U426 ( .A(add_x_1_n21), .B(mem_data_pc4[11]), .CO(add_x_1_n20), .S(
        u_mem_pc8[11]) );
  ADD22 U427 ( .A(n174), .B(mem_data_pc4[14]), .CO(add_x_1_n17), .S(
        u_mem_pc8[14]) );
  ADD22 U428 ( .A(add_x_1_n17), .B(mem_data_pc4[15]), .CO(add_x_1_n16), .S(
        u_mem_pc8[15]) );
  ADD22 U429 ( .A(add_x_1_n13), .B(mem_data_pc4[19]), .CO(add_x_1_n12), .S(
        u_mem_pc8[19]) );
  ADD22 U430 ( .A(mem_data_pc4[2]), .B(mem_data_pc4[3]), .CO(add_x_1_n28), .S(
        u_mem_pc8[3]) );
  NAND23 U431 ( .A(add_x_1_n14), .B(mem_data_pc4[18]), .Q(n176) );
  ADD22 U432 ( .A(add_x_1_n23), .B(mem_data_pc4[9]), .CO(add_x_1_n22), .S(
        u_mem_pc8[9]) );
  ADD22 U433 ( .A(add_x_1_n25), .B(mem_data_pc4[7]), .CO(add_x_1_n24), .S(
        u_mem_pc8[7]) );
  ADD22 U434 ( .A(add_x_1_n24), .B(mem_data_pc4[8]), .CO(add_x_1_n23), .S(
        u_mem_pc8[8]) );
  ADD22 U435 ( .A(add_x_1_n5), .B(mem_data_pc4[27]), .CO(add_x_1_n4), .S(
        u_mem_pc8[27]) );
  ADD22 U436 ( .A(add_x_1_n27), .B(mem_data_pc4[5]), .CO(add_x_1_n26), .S(
        u_mem_pc8[5]) );
  ADD22 U437 ( .A(add_x_1_n26), .B(mem_data_pc4[6]), .CO(add_x_1_n25), .S(
        u_mem_pc8[6]) );
  ADD22 U438 ( .A(add_x_1_n7), .B(mem_data_pc4[25]), .CO(add_x_1_n6), .S(
        u_mem_pc8[25]) );
  INV6 U439 ( .A(n170), .Q(add_x_1_n8) );
  INV3 U440 ( .A(n172), .Q(add_x_1_n9) );
  INV3 U441 ( .A(n177), .Q(add_x_1_n5) );
  INV3 U442 ( .A(n181), .Q(add_x_4_n1) );
  XOR21 U443 ( .A(add_x_4_n2), .B(instruction_address[30]), .Q(
        u_fetch_jmux_i_addr_pc4_30_) );
  XOR21 U444 ( .A(add_x_4_n5), .B(instruction_address[27]), .Q(
        u_fetch_jmux_i_addr_pc4_27_) );
  XOR21 U445 ( .A(add_x_4_n6), .B(instruction_address[26]), .Q(
        u_fetch_jmux_i_addr_pc4_26_) );
  XOR20 U446 ( .A(add_x_4_n12), .B(instruction_address[20]), .Q(
        u_fetch_jmux_i_addr_pc4_20_) );
  XOR20 U447 ( .A(add_x_4_n15), .B(instruction_address[17]), .Q(
        u_fetch_jmux_i_addr_pc4_17_) );
  NOR24 U448 ( .A(n180), .B(n168), .Q(n182) );
  ADD22 U449 ( .A(add_x_4_n17), .B(instruction_address[15]), .CO(add_x_4_n16), 
        .S(u_fetch_jmux_i_addr_pc4_15_) );
  ADD22 U450 ( .A(add_x_4_n16), .B(instruction_address[16]), .CO(add_x_4_n15), 
        .S(u_fetch_jmux_i_addr_pc4_16_) );
  ADD22 U451 ( .A(add_x_4_n8), .B(instruction_address[24]), .CO(add_x_4_n7), 
        .S(u_fetch_jmux_i_addr_pc4_24_) );
  ADD22 U452 ( .A(add_x_4_n7), .B(instruction_address[25]), .CO(add_x_4_n6), 
        .S(u_fetch_jmux_i_addr_pc4_25_) );
  XNR22 U453 ( .A(n179), .B(add_x_4_n1), .Q(u_fetch_jmux_i_addr_pc4_31_) );
  ADD22 U454 ( .A(n182), .B(instruction_address[19]), .CO(add_x_4_n12), .S(
        u_fetch_jmux_i_addr_pc4_19_) );
  ADD22 U455 ( .A(add_x_4_n19), .B(instruction_address[13]), .CO(add_x_4_n18), 
        .S(u_fetch_jmux_i_addr_pc4_13_) );
  ADD22 U456 ( .A(add_x_4_n18), .B(instruction_address[14]), .CO(add_x_4_n17), 
        .S(u_fetch_jmux_i_addr_pc4_14_) );
  ADD22 U457 ( .A(add_x_4_n10), .B(instruction_address[22]), .CO(add_x_4_n9), 
        .S(u_fetch_jmux_i_addr_pc4_22_) );
  ADD22 U458 ( .A(add_x_4_n9), .B(instruction_address[23]), .CO(add_x_4_n8), 
        .S(u_fetch_jmux_i_addr_pc4_23_) );
  ADD22 U459 ( .A(add_x_4_n20), .B(instruction_address[12]), .CO(add_x_4_n19), 
        .S(u_fetch_jmux_i_addr_pc4_12_) );
  ADD22 U460 ( .A(add_x_4_n11), .B(instruction_address[21]), .CO(add_x_4_n10), 
        .S(u_fetch_jmux_i_addr_pc4_21_) );
  NAND26 U461 ( .A(add_x_4_n15), .B(instruction_address[17]), .Q(n180) );
  ADD22 U462 ( .A(instruction_address[2]), .B(instruction_address[3]), .CO(
        add_x_4_n28), .S(u_fetch_jmux_i_addr_pc4_3_) );
  INV3 U463 ( .A(n178), .Q(add_x_4_n11) );
  ADD22 U464 ( .A(add_x_4_n22), .B(instruction_address[10]), .CO(add_x_4_n21), 
        .S(u_fetch_jmux_i_addr_pc4_10_) );
  ADD22 U465 ( .A(add_x_4_n21), .B(instruction_address[11]), .CO(add_x_4_n20), 
        .S(u_fetch_jmux_i_addr_pc4_11_) );
  ADD22 U466 ( .A(add_x_4_n24), .B(instruction_address[8]), .CO(add_x_4_n23), 
        .S(u_fetch_jmux_i_addr_pc4_8_) );
  ADD22 U467 ( .A(add_x_4_n23), .B(instruction_address[9]), .CO(add_x_4_n22), 
        .S(u_fetch_jmux_i_addr_pc4_9_) );
  ADD22 U468 ( .A(add_x_4_n26), .B(instruction_address[6]), .CO(add_x_4_n25), 
        .S(u_fetch_jmux_i_addr_pc4_6_) );
  ADD22 U469 ( .A(add_x_4_n25), .B(instruction_address[7]), .CO(add_x_4_n24), 
        .S(u_fetch_jmux_i_addr_pc4_7_) );
  NAND26 U470 ( .A(add_x_4_n6), .B(instruction_address[26]), .Q(n184) );
  NAND28 U471 ( .A(add_x_4_n5), .B(instruction_address[27]), .Q(n183) );
  INV6 U472 ( .A(n183), .Q(add_x_4_n4) );
  ADD22 U473 ( .A(add_x_4_n28), .B(instruction_address[4]), .CO(add_x_4_n27), 
        .S(u_fetch_jmux_i_addr_pc4_4_) );
  ADD22 U474 ( .A(add_x_4_n27), .B(instruction_address[5]), .CO(add_x_4_n26), 
        .S(u_fetch_jmux_i_addr_pc4_5_) );
  OAI2110 U475 ( .A(instruction_address[2]), .B(n405), .C(n316), .D(n315), .Q(
        n135) );
  OAI2112 U476 ( .A(n405), .B(n314), .C(n313), .D(n312), .Q(n138) );
  NAND20 U477 ( .A(n213), .B(n218), .Q(n220) );
  AOI221 U478 ( .A(n205), .B(id_data_jr[1]), .C(n399), .D(ex_data_pc4[1]), .Q(
        n308) );
  AOI221 U479 ( .A(n205), .B(id_data_jr[0]), .C(n399), .D(ex_data_pc4[0]), .Q(
        n307) );
  NOR21 U480 ( .A(n310), .B(n398), .Q(n309) );
  AOI221 U481 ( .A(n205), .B(id_data_jr[28]), .C(n169), .D(if_addr_j[28]), .Q(
        n392) );
  BUF6 U482 ( .A(ex_data_immext[6]), .Q(n206) );
  AOI220 U483 ( .A(if_addr_b[3]), .B(n399), .C(instruction_address[3]), .D(
        n398), .Q(n318) );
  INV3 U484 ( .A(if_con_ifstall), .Q(n398) );
  INV3 U485 ( .A(u_fetch_jmux_i_addr_pc4_30_), .Q(n404) );
  INV3 U486 ( .A(u_fetch_jmux_i_addr_pc4_31_), .Q(n314) );
  NOR40 U487 ( .A(n261), .B(n262), .C(n263), .D(n264), .Q(n259) );
  NAND30 U488 ( .A(id_data_instr[28]), .B(n213), .C(n185), .Q(n221) );
  NOR20 U489 ( .A(id_data_instr[31]), .B(n297), .Q(
        u_decode_control_o_con_aluop_0_) );
  NOR30 U490 ( .A(n185), .B(n192), .C(id_data_instr[28]), .Q(n294) );
  MUX21 U491 ( .A(data_address[6]), .B(u_mem_pc8[6]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[6]) );
  MUX21 U492 ( .A(data_address[1]), .B(u_mem_pc8[1]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[1]) );
  MUX21 U493 ( .A(data_address[4]), .B(u_mem_pc8[4]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[4]) );
  MUX21 U494 ( .A(data_address[5]), .B(u_mem_pc8[5]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[5]) );
  MUX21 U495 ( .A(data_address[0]), .B(u_mem_pc8[0]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[0]) );
  MUX21 U496 ( .A(data_address[3]), .B(u_mem_pc8[3]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[3]) );
  MUX21 U497 ( .A(data_address[7]), .B(u_mem_pc8[7]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[7]) );
  MUX21 U498 ( .A(data_address[8]), .B(u_mem_pc8[8]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[8]) );
  NOR21 U499 ( .A(n295), .B(n296), .Q(u_decode_jbcon_o_con_aluPC4) );
  MUX21 U500 ( .A(data_address[9]), .B(u_mem_pc8[9]), .S(mem_con_Malupc8), .Q(
        u_mem_resmux_o_data_alu[9]) );
  MUX21 U501 ( .A(data_address[10]), .B(u_mem_pc8[10]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[10]) );
  MUX21 U502 ( .A(data_address[11]), .B(u_mem_pc8[11]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[11]) );
  NOR31 U503 ( .A(n225), .B(n222), .C(n226), .Q(u_decode_for_o_con_fb[1]) );
  MUX21 U504 ( .A(data_address[12]), .B(u_mem_pc8[12]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[12]) );
  AOI211 U505 ( .A(n223), .B(n227), .C(n222), .Q(u_decode_for_o_con_fb[0]) );
  NAND41 U506 ( .A(n236), .B(n226), .C(n237), .D(n238), .Q(n227) );
  IMUX20 U507 ( .A(if_addr_j[20]), .B(n197), .S(for_o_addr_Erd[2]), .Q(n240)
         );
  IMUX20 U508 ( .A(n187), .B(if_addr_j[18]), .S(for_o_addr_Erd[0]), .Q(n244)
         );
  IMUX20 U509 ( .A(n201), .B(if_addr_j[21]), .S(for_o_addr_Erd[3]), .Q(n243)
         );
  IMUX20 U510 ( .A(n198), .B(if_addr_j[19]), .S(for_o_addr_Erd[1]), .Q(n242)
         );
  MUX21 U511 ( .A(data_address[14]), .B(u_mem_pc8[14]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[14]) );
  NOR21 U512 ( .A(n255), .B(u_decode_for_o_con_fa_2_), .Q(
        u_decode_for_o_con_fa_1_) );
  NAND22 U513 ( .A(n257), .B(n258), .Q(u_decode_for_o_con_fa_2_) );
  MUX21 U514 ( .A(data_address[15]), .B(u_mem_pc8[15]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[15]) );
  MUX21 U515 ( .A(data_address[16]), .B(u_mem_pc8[16]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[16]) );
  AOI211 U516 ( .A(n258), .B(n260), .C(n259), .Q(u_decode_for_o_con_fa_0_) );
  IMUX20 U517 ( .A(if_addr_j[23]), .B(n193), .S(for_o_addr_Erd[0]), .Q(n277)
         );
  MUX21 U518 ( .A(data_address[18]), .B(u_mem_pc8[18]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[18]) );
  MUX21 U519 ( .A(data_address[22]), .B(u_mem_pc8[22]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[22]) );
  MUX21 U520 ( .A(data_address[23]), .B(u_mem_pc8[23]), .S(mem_con_Malupc8), 
        .Q(u_mem_resmux_o_data_alu[23]) );
  INV3 U521 ( .A(u_decode_add_x_16_n62), .Q(u_decode_add_x_16_n60) );
  INV3 U522 ( .A(u_decode_add_x_16_n70), .Q(u_decode_add_x_16_n68) );
  OAI2111 U523 ( .A(n405), .B(n337), .C(n336), .D(n335), .Q(n128) );
  OAI2111 U524 ( .A(n405), .B(n373), .C(n372), .D(n371), .Q(n116) );
  OAI2111 U525 ( .A(n405), .B(n388), .C(n387), .D(n386), .Q(n111) );
  OAI2111 U526 ( .A(n405), .B(n346), .C(n345), .D(n344), .Q(n125) );
  OAI2111 U527 ( .A(n405), .B(n397), .C(n396), .D(n395), .Q(n108) );
  OAI2111 U528 ( .A(n405), .B(n331), .C(n330), .D(n329), .Q(n130) );
  OAI2111 U529 ( .A(n405), .B(n376), .C(n375), .D(n374), .Q(n115) );
  OAI2111 U530 ( .A(n405), .B(n349), .C(n348), .D(n347), .Q(n124) );
  OAI2111 U531 ( .A(n405), .B(n391), .C(n390), .D(n389), .Q(n110) );
  OAI2111 U532 ( .A(n405), .B(n367), .C(n366), .D(n365), .Q(n118) );
  OAI2111 U533 ( .A(n405), .B(n394), .C(n393), .D(n392), .Q(n109) );
  OAI2111 U534 ( .A(n405), .B(n364), .C(n363), .D(n362), .Q(n119) );
  OAI2111 U535 ( .A(n405), .B(n322), .C(n321), .D(n320), .Q(n133) );
  OAI2111 U536 ( .A(n405), .B(n361), .C(n360), .D(n359), .Q(n120) );
  OAI2111 U537 ( .A(n405), .B(n352), .C(n351), .D(n350), .Q(n123) );
  OAI2111 U538 ( .A(n405), .B(n382), .C(n381), .D(n380), .Q(n113) );
  OAI2111 U539 ( .A(n405), .B(n379), .C(n378), .D(n377), .Q(n114) );
  OAI2111 U540 ( .A(n405), .B(n343), .C(n342), .D(n341), .Q(n126) );
  OAI2111 U541 ( .A(n405), .B(n319), .C(n318), .D(n317), .Q(n134) );
  OAI2111 U542 ( .A(n405), .B(n325), .C(n324), .D(n323), .Q(n132) );
  OAI2111 U543 ( .A(n405), .B(n358), .C(n357), .D(n356), .Q(n121) );
  OAI2111 U544 ( .A(n405), .B(n355), .C(n354), .D(n353), .Q(n122) );
  OAI2111 U545 ( .A(n405), .B(n370), .C(n369), .D(n368), .Q(n117) );
  OAI2111 U546 ( .A(n405), .B(n385), .C(n384), .D(n383), .Q(n112) );
  OAI2111 U547 ( .A(n405), .B(n340), .C(n339), .D(n338), .Q(n127) );
  OAI2111 U548 ( .A(n405), .B(n334), .C(n333), .D(n332), .Q(n129) );
  OAI2111 U549 ( .A(n405), .B(n328), .C(n327), .D(n326), .Q(n131) );
  INV3 U550 ( .A(if_con_b), .Q(n306) );
  BUF6 U551 ( .A(ex_data_immext[8]), .Q(n207) );
  INV3 U552 ( .A(n210), .Q(n297) );
  NAND22 U553 ( .A(n228), .B(n224), .Q(n222) );
  INV3 U554 ( .A(u_decode_add_x_16_n61), .Q(u_decode_add_x_16_n59) );
  INV3 U555 ( .A(u_decode_add_x_16_n69), .Q(u_decode_add_x_16_n67) );
  INV3 U556 ( .A(if_con_j[0]), .Q(n311) );
  INV3 U557 ( .A(if_con_j[1]), .Q(n305) );
  NAND22 U558 ( .A(n213), .B(n214), .Q(if_con_j[1]) );
  LOGIC0 U559 ( .Q(n204) );
  AOI310 U560 ( .A(n210), .B(n189), .C(n211), .D(
        u_decode_control_o_con_memtoreg), .Q(n208) );
  AOI210 U561 ( .A(n189), .B(id_data_instr[27]), .C(n212), .Q(u_decode_n6) );
  OAI2110 U562 ( .A(n189), .B(id_data_instr[27]), .C(n213), .D(
        id_data_instr[26]), .Q(n212) );
  NOR40 U563 ( .A(if_addr_j[2]), .B(if_addr_j[3]), .C(if_addr_j[4]), .D(
        if_addr_j[6]), .Q(n217) );
  OAI220 U564 ( .A(n219), .B(n220), .C(n192), .D(n221), .Q(
        u_decode_jbcon_o_con_bop[1]) );
  NOR20 U565 ( .A(if_addr_j[18]), .B(id_data_instr[28]), .Q(n219) );
  OAI310 U566 ( .A(if_addr_j[18]), .B(id_data_instr[28]), .C(n220), .D(n221), 
        .Q(u_decode_jbcon_o_con_bop[0]) );
  IMUX20 U567 ( .A(if_addr_j[20]), .B(n197), .S(for_addr_rtM[2]), .Q(n230) );
  NOR40 U568 ( .A(n231), .B(n232), .C(n233), .D(n234), .Q(n229) );
  IMUX20 U569 ( .A(n201), .B(if_addr_j[21]), .S(for_addr_rtM[3]), .Q(n234) );
  IMUX20 U570 ( .A(n198), .B(if_addr_j[19]), .S(for_addr_rtM[1]), .Q(n233) );
  IMUX20 U571 ( .A(n199), .B(if_addr_j[22]), .S(for_addr_rtM[4]), .Q(n232) );
  IMUX20 U572 ( .A(n187), .B(if_addr_j[18]), .S(for_addr_rtM[0]), .Q(n231) );
  NOR40 U573 ( .A(if_addr_j[19]), .B(if_addr_j[21]), .C(if_addr_j[18]), .D(
        if_addr_j[20]), .Q(n235) );
  IMUX20 U574 ( .A(if_addr_j[18]), .B(n187), .S(mem_addr_regdst[0]), .Q(n238)
         );
  IMUX20 U575 ( .A(if_addr_j[19]), .B(n198), .S(mem_addr_regdst[1]), .Q(n237)
         );
  NOR40 U576 ( .A(n241), .B(n242), .C(n243), .D(n244), .Q(n239) );
  IMUX20 U577 ( .A(n199), .B(if_addr_j[22]), .S(for_o_addr_Erd[4]), .Q(n241)
         );
  NOR40 U578 ( .A(n245), .B(n246), .C(n247), .D(n248), .Q(n236) );
  IMUX20 U579 ( .A(n201), .B(if_addr_j[21]), .S(mem_addr_regdst[3]), .Q(n247)
         );
  IMUX20 U580 ( .A(n197), .B(if_addr_j[20]), .S(mem_addr_regdst[2]), .Q(n246)
         );
  IMUX20 U581 ( .A(n199), .B(if_addr_j[22]), .S(mem_addr_regdst[4]), .Q(n245)
         );
  IMUX20 U582 ( .A(if_addr_j[22]), .B(n199), .S(for_addr_rtW[4]), .Q(n250) );
  NOR40 U583 ( .A(n251), .B(n252), .C(n253), .D(n254), .Q(n249) );
  IMUX20 U584 ( .A(n187), .B(if_addr_j[18]), .S(for_addr_rtW[0]), .Q(n254) );
  IMUX20 U585 ( .A(n198), .B(if_addr_j[19]), .S(for_addr_rtW[1]), .Q(n253) );
  IMUX20 U586 ( .A(n197), .B(if_addr_j[20]), .S(for_addr_rtW[2]), .Q(n252) );
  IMUX20 U587 ( .A(n201), .B(if_addr_j[21]), .S(for_addr_rtW[3]), .Q(n251) );
  IMUX20 U588 ( .A(if_addr_j[25]), .B(n190), .S(for_addr_rtM[2]), .Q(n267) );
  IMUX20 U589 ( .A(if_addr_j[26]), .B(n195), .S(for_addr_rtM[3]), .Q(n266) );
  IMUX20 U590 ( .A(if_addr_j[27]), .B(n194), .S(for_addr_rtM[4]), .Q(n265) );
  IMUX20 U591 ( .A(n193), .B(if_addr_j[23]), .S(for_addr_rtM[0]), .Q(n263) );
  IMUX20 U592 ( .A(n191), .B(if_addr_j[24]), .S(for_addr_rtM[1]), .Q(n262) );
  AOI2110 U593 ( .A(mem_addr_regdst[1]), .B(n191), .C(n256), .D(n272), .Q(n271) );
  IMUX20 U594 ( .A(n190), .B(if_addr_j[25]), .S(mem_addr_regdst[2]), .Q(n272)
         );
  NOR40 U595 ( .A(n273), .B(n274), .C(n275), .D(n276), .Q(n256) );
  OAI210 U596 ( .A(for_o_addr_Erd[2]), .B(n279), .C(n190), .Q(n278) );
  NOR40 U597 ( .A(for_o_addr_Erd[1]), .B(for_o_addr_Erd[3]), .C(
        for_o_addr_Erd[0]), .D(if_addr_j[27]), .Q(n279) );
  IMUX20 U598 ( .A(if_addr_j[27]), .B(n194), .S(for_o_addr_Erd[4]), .Q(n280)
         );
  IMUX20 U599 ( .A(n195), .B(if_addr_j[26]), .S(for_o_addr_Erd[3]), .Q(n274)
         );
  IMUX20 U600 ( .A(n191), .B(if_addr_j[24]), .S(for_o_addr_Erd[1]), .Q(n273)
         );
  NOR40 U601 ( .A(n281), .B(n282), .C(n283), .D(n248), .Q(n270) );
  IMUX20 U602 ( .A(n194), .B(if_addr_j[27]), .S(mem_addr_regdst[4]), .Q(n283)
         );
  IMUX20 U603 ( .A(n195), .B(if_addr_j[26]), .S(mem_addr_regdst[3]), .Q(n282)
         );
  IMUX20 U604 ( .A(n193), .B(if_addr_j[23]), .S(mem_addr_regdst[0]), .Q(n281)
         );
  NOR20 U605 ( .A(if_addr_j[24]), .B(n284), .Q(n269) );
  NOR40 U606 ( .A(mem_addr_regdst[0]), .B(mem_addr_regdst[4]), .C(
        mem_addr_regdst[2]), .D(mem_addr_regdst[3]), .Q(n284) );
  NOR40 U607 ( .A(if_addr_j[23]), .B(if_addr_j[25]), .C(if_addr_j[26]), .D(
        if_addr_j[24]), .Q(n287) );
  IMUX20 U608 ( .A(if_addr_j[26]), .B(n195), .S(for_addr_rtW[3]), .Q(n286) );
  NOR40 U609 ( .A(n288), .B(n289), .C(n290), .D(n291), .Q(n285) );
  IMUX20 U610 ( .A(n190), .B(if_addr_j[25]), .S(for_addr_rtW[2]), .Q(n291) );
  IMUX20 U611 ( .A(n194), .B(if_addr_j[27]), .S(for_addr_rtW[4]), .Q(n290) );
  IMUX20 U612 ( .A(n193), .B(if_addr_j[23]), .S(for_addr_rtW[0]), .Q(n289) );
  IMUX20 U613 ( .A(n191), .B(if_addr_j[24]), .S(for_addr_rtW[1]), .Q(n288) );
  AOI2110 U614 ( .A(n186), .B(n295), .C(id_data_instr[30]), .D(n200), .Q(
        u_decode_control_o_con_memtoreg) );
  NAND30 U615 ( .A(n293), .B(n294), .C(id_data_instr[31]), .Q(n299) );
  NOR20 U616 ( .A(id_data_instr[30]), .B(id_data_instr[29]), .Q(n293) );
  OAI310 U617 ( .A(id_data_instr[30]), .B(n295), .C(n200), .D(n297), .Q(
        u_decode_control_o_con_alusrc) );
  AOI2110 U618 ( .A(n186), .B(n214), .C(id_data_instr[30]), .D(
        id_data_instr[31]), .Q(u_decode_control_o_con_aluop_1_) );
  NOR40 U619 ( .A(id_data_instr[28]), .B(id_data_instr[31]), .C(n211), .D(n297), .Q(u_decode_control_o_con_aluop_5_) );
  NAND20 U620 ( .A(id_data_instr[26]), .B(id_data_instr[27]), .Q(n211) );
  NOR40 U621 ( .A(id_data_instr[30]), .B(id_data_instr[31]), .C(n186), .D(n189), .Q(n303) );
  NAND30 U622 ( .A(u_decode_control_o_con_aluop_0_), .B(n189), .C(n185), .Q(
        n304) );
  AOI220 U623 ( .A(if_addr_b[31]), .B(n399), .C(instruction_address[31]), .D(
        n398), .Q(n313) );
  AOI220 U624 ( .A(if_addr_b[2]), .B(n399), .C(instruction_address[2]), .D(
        n398), .Q(n316) );
  AOI220 U625 ( .A(if_addr_b[4]), .B(n399), .C(instruction_address[4]), .D(
        n398), .Q(n321) );
  AOI220 U626 ( .A(if_addr_b[5]), .B(n399), .C(instruction_address[5]), .D(
        n398), .Q(n324) );
  AOI220 U627 ( .A(if_addr_b[6]), .B(n399), .C(instruction_address[6]), .D(
        n398), .Q(n327) );
  AOI220 U628 ( .A(if_addr_b[7]), .B(n399), .C(instruction_address[7]), .D(
        n398), .Q(n330) );
  AOI220 U629 ( .A(if_addr_b[8]), .B(n399), .C(instruction_address[8]), .D(
        n398), .Q(n333) );
  AOI220 U630 ( .A(if_addr_b[9]), .B(n399), .C(instruction_address[9]), .D(
        n398), .Q(n336) );
  AOI220 U631 ( .A(n401), .B(id_data_jr[9]), .C(n169), .D(if_addr_j[9]), .Q(
        n335) );
  AOI220 U632 ( .A(if_addr_b[10]), .B(n399), .C(instruction_address[10]), .D(
        n398), .Q(n339) );
  AOI220 U633 ( .A(if_addr_b[11]), .B(n399), .C(instruction_address[11]), .D(
        n398), .Q(n342) );
  AOI220 U634 ( .A(if_addr_b[12]), .B(n399), .C(instruction_address[12]), .D(
        n398), .Q(n345) );
  AOI220 U635 ( .A(if_addr_b[13]), .B(n399), .C(instruction_address[13]), .D(
        n398), .Q(n348) );
  AOI220 U636 ( .A(if_addr_b[14]), .B(n399), .C(instruction_address[14]), .D(
        n398), .Q(n351) );
  AOI220 U637 ( .A(if_addr_b[15]), .B(n399), .C(instruction_address[15]), .D(
        n398), .Q(n354) );
  AOI220 U638 ( .A(if_addr_b[16]), .B(n399), .C(instruction_address[16]), .D(
        n398), .Q(n357) );
  AOI220 U639 ( .A(if_addr_b[17]), .B(n399), .C(instruction_address[17]), .D(
        n398), .Q(n360) );
  AOI220 U640 ( .A(n205), .B(id_data_jr[17]), .C(n169), .D(if_addr_j[17]), .Q(
        n359) );
  AOI220 U641 ( .A(if_addr_b[18]), .B(n399), .C(instruction_address[18]), .D(
        n398), .Q(n363) );
  AOI220 U642 ( .A(n205), .B(id_data_jr[18]), .C(n169), .D(if_addr_j[18]), .Q(
        n362) );
  AOI220 U643 ( .A(if_addr_b[19]), .B(n399), .C(instruction_address[19]), .D(
        n398), .Q(n366) );
  AOI220 U644 ( .A(n205), .B(id_data_jr[19]), .C(n169), .D(if_addr_j[19]), .Q(
        n365) );
  AOI220 U645 ( .A(if_addr_b[20]), .B(n399), .C(instruction_address[20]), .D(
        n398), .Q(n369) );
  AOI220 U646 ( .A(n205), .B(id_data_jr[20]), .C(n169), .D(if_addr_j[20]), .Q(
        n368) );
  AOI220 U647 ( .A(if_addr_b[21]), .B(n399), .C(instruction_address[21]), .D(
        n398), .Q(n372) );
  AOI220 U648 ( .A(n205), .B(id_data_jr[21]), .C(n169), .D(if_addr_j[21]), .Q(
        n371) );
  AOI220 U649 ( .A(if_addr_b[22]), .B(n399), .C(instruction_address[22]), .D(
        n398), .Q(n375) );
  AOI220 U650 ( .A(n205), .B(id_data_jr[22]), .C(n169), .D(if_addr_j[22]), .Q(
        n374) );
  AOI220 U651 ( .A(if_addr_b[23]), .B(n399), .C(instruction_address[23]), .D(
        n398), .Q(n378) );
  AOI220 U652 ( .A(n205), .B(id_data_jr[23]), .C(n169), .D(if_addr_j[23]), .Q(
        n377) );
  AOI220 U653 ( .A(if_addr_b[24]), .B(n399), .C(instruction_address[24]), .D(
        n398), .Q(n381) );
  AOI220 U654 ( .A(n205), .B(id_data_jr[24]), .C(n169), .D(if_addr_j[24]), .Q(
        n380) );
  AOI220 U655 ( .A(if_addr_b[25]), .B(n399), .C(instruction_address[25]), .D(
        n398), .Q(n384) );
  AOI220 U656 ( .A(n205), .B(id_data_jr[25]), .C(n169), .D(if_addr_j[25]), .Q(
        n383) );
  AOI220 U657 ( .A(if_addr_b[26]), .B(n399), .C(instruction_address[26]), .D(
        n398), .Q(n387) );
  AOI220 U658 ( .A(n205), .B(id_data_jr[26]), .C(n169), .D(if_addr_j[26]), .Q(
        n386) );
  AOI220 U659 ( .A(if_addr_b[27]), .B(n399), .C(instruction_address[27]), .D(
        n398), .Q(n390) );
  AOI220 U660 ( .A(n205), .B(id_data_jr[27]), .C(n169), .D(if_addr_j[27]), .Q(
        n389) );
  AOI220 U661 ( .A(if_addr_b[28]), .B(n399), .C(instruction_address[28]), .D(
        n398), .Q(n393) );
  AOI220 U662 ( .A(if_addr_b[29]), .B(n399), .C(instruction_address[29]), .D(
        n398), .Q(n396) );
  AOI220 U663 ( .A(if_addr_b[30]), .B(n399), .C(instruction_address[30]), .D(
        n398), .Q(n403) );
endmodule

